module fake_netlist_6_3814_n_1732 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1732);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1732;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_913;
wire n_407;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_850;
wire n_690;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1669;
wire n_1403;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1702;
wire n_1570;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_228;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_106),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_136),
.Y(n_157)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_57),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_18),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_13),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_50),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_109),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_58),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_1),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_62),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_37),
.Y(n_166)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_73),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_29),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_101),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_115),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_102),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_10),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_151),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_36),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_0),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_88),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_113),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_44),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_47),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_64),
.Y(n_180)
);

BUFx10_ASAP7_75t_L g181 ( 
.A(n_29),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_146),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_46),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_87),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_11),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_104),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_10),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_141),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_110),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_60),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_93),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_33),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_59),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_50),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_8),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_0),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_150),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_37),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_13),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_84),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_39),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_145),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_107),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_147),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_121),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_1),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_17),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_59),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_15),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_116),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_26),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_58),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_14),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_66),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_81),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_80),
.Y(n_216)
);

INVx2_ASAP7_75t_SL g217 ( 
.A(n_52),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_48),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_20),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_2),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_57),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_74),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_8),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_149),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_72),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_4),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_18),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_54),
.Y(n_228)
);

BUFx10_ASAP7_75t_L g229 ( 
.A(n_17),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_5),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_127),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_77),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_4),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_86),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_28),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_111),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_134),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_52),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_95),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_100),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_68),
.Y(n_241)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_6),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_82),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_56),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_139),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_90),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_19),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_38),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_126),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_137),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_32),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_26),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_142),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_97),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_132),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_118),
.Y(n_256)
);

BUFx5_ASAP7_75t_L g257 ( 
.A(n_43),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_31),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_53),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_42),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_56),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_131),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_21),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_14),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_30),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_51),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_2),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_33),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_144),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_55),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_89),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_41),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_24),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_94),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_129),
.Y(n_275)
);

INVx2_ASAP7_75t_SL g276 ( 
.A(n_71),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_25),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_16),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_69),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_27),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_16),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_96),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_36),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_105),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_6),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_63),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_27),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_47),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_98),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_70),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_79),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_123),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_38),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_91),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_23),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_20),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_148),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_83),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_53),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_108),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_112),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_49),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_43),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_55),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_120),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_124),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_19),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_9),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_15),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_257),
.Y(n_310)
);

NOR2xp67_ASAP7_75t_L g311 ( 
.A(n_290),
.B(n_3),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g312 ( 
.A(n_158),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_257),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_156),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_157),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_162),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_169),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_257),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_257),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_257),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_257),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_170),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_158),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_257),
.Y(n_324)
);

BUFx10_ASAP7_75t_L g325 ( 
.A(n_165),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_286),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_257),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_292),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_257),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_180),
.Y(n_330)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_293),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_183),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_293),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_293),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_R g335 ( 
.A(n_231),
.B(n_119),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_293),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_176),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_183),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_177),
.Y(n_339)
);

NOR2xp67_ASAP7_75t_L g340 ( 
.A(n_290),
.B(n_3),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_186),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_188),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_293),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_293),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_196),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_167),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g347 ( 
.A(n_167),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_231),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_196),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_196),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_191),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_197),
.Y(n_352)
);

NOR2xp67_ASAP7_75t_L g353 ( 
.A(n_290),
.B(n_5),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_196),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_242),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_196),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_272),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_289),
.B(n_7),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_211),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_289),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_200),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_272),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_211),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_202),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_223),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_203),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_204),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_223),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_205),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_210),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_215),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_227),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_216),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_227),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_222),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_225),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_247),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_247),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_263),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_232),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_263),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_181),
.Y(n_382)
);

INVxp67_ASAP7_75t_SL g383 ( 
.A(n_290),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_236),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_264),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_334),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_321),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_330),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_330),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_330),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_321),
.Y(n_391)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_330),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_310),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_332),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_310),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_334),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_336),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_336),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_383),
.B(n_173),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_345),
.B(n_165),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_343),
.Y(n_401)
);

BUFx8_ASAP7_75t_L g402 ( 
.A(n_360),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_330),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_343),
.Y(n_404)
);

AND2x4_ASAP7_75t_L g405 ( 
.A(n_311),
.B(n_276),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_313),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_344),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_344),
.Y(n_408)
);

AND2x4_ASAP7_75t_L g409 ( 
.A(n_340),
.B(n_276),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_313),
.Y(n_410)
);

NOR2x1_ASAP7_75t_L g411 ( 
.A(n_353),
.B(n_171),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_318),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_318),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_331),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_331),
.B(n_173),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_351),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_331),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_333),
.B(n_182),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_333),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_345),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_319),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_349),
.B(n_241),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_319),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_349),
.B(n_243),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_320),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_320),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_324),
.Y(n_427)
);

AND2x4_ASAP7_75t_L g428 ( 
.A(n_350),
.B(n_171),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_324),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_350),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_354),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_354),
.Y(n_432)
);

AND2x4_ASAP7_75t_L g433 ( 
.A(n_356),
.B(n_189),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_358),
.B(n_181),
.Y(n_434)
);

BUFx2_ASAP7_75t_L g435 ( 
.A(n_348),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_356),
.B(n_189),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_327),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_327),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_329),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_329),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_374),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_374),
.B(n_182),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_359),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_346),
.B(n_245),
.Y(n_444)
);

NAND2xp33_ASAP7_75t_L g445 ( 
.A(n_335),
.B(n_217),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_359),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_347),
.B(n_273),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_363),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_363),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_365),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_365),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g452 ( 
.A(n_357),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_368),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_368),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_372),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_372),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_377),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_387),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_388),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_388),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_418),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_405),
.B(n_314),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_434),
.B(n_316),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_388),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_388),
.Y(n_465)
);

AND2x6_ASAP7_75t_L g466 ( 
.A(n_399),
.B(n_262),
.Y(n_466)
);

OR2x2_ASAP7_75t_L g467 ( 
.A(n_394),
.B(n_323),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_387),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_399),
.B(n_360),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_437),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_437),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_437),
.Y(n_472)
);

INVx5_ASAP7_75t_L g473 ( 
.A(n_412),
.Y(n_473)
);

INVx2_ASAP7_75t_SL g474 ( 
.A(n_447),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_416),
.Y(n_475)
);

INVx1_ASAP7_75t_SL g476 ( 
.A(n_416),
.Y(n_476)
);

BUFx4f_ASAP7_75t_L g477 ( 
.A(n_412),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_387),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_418),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_387),
.Y(n_480)
);

OR2x2_ASAP7_75t_L g481 ( 
.A(n_394),
.B(n_338),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_434),
.B(n_317),
.Y(n_482)
);

OR2x6_ASAP7_75t_L g483 ( 
.A(n_444),
.B(n_184),
.Y(n_483)
);

OR2x2_ASAP7_75t_L g484 ( 
.A(n_452),
.B(n_338),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_391),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_439),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_391),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_444),
.B(n_322),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_439),
.Y(n_489)
);

AND2x4_ASAP7_75t_L g490 ( 
.A(n_418),
.B(n_184),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_439),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_391),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_440),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_440),
.Y(n_494)
);

INVx4_ASAP7_75t_L g495 ( 
.A(n_412),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_440),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_399),
.B(n_337),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_405),
.B(n_339),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_418),
.Y(n_499)
);

AO21x2_ASAP7_75t_L g500 ( 
.A1(n_422),
.A2(n_234),
.B(n_224),
.Y(n_500)
);

INVx5_ASAP7_75t_L g501 ( 
.A(n_412),
.Y(n_501)
);

OR2x2_ASAP7_75t_L g502 ( 
.A(n_452),
.B(n_362),
.Y(n_502)
);

INVx4_ASAP7_75t_L g503 ( 
.A(n_412),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_405),
.B(n_341),
.Y(n_504)
);

AOI22xp33_ASAP7_75t_L g505 ( 
.A1(n_399),
.A2(n_312),
.B1(n_260),
.B2(n_217),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_421),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_442),
.B(n_385),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_405),
.A2(n_369),
.B1(n_384),
.B2(n_352),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_421),
.Y(n_509)
);

AND2x4_ASAP7_75t_L g510 ( 
.A(n_442),
.B(n_224),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_442),
.B(n_385),
.Y(n_511)
);

BUFx4f_ASAP7_75t_L g512 ( 
.A(n_412),
.Y(n_512)
);

INVx5_ASAP7_75t_L g513 ( 
.A(n_412),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_421),
.Y(n_514)
);

BUFx4f_ASAP7_75t_L g515 ( 
.A(n_412),
.Y(n_515)
);

INVx5_ASAP7_75t_L g516 ( 
.A(n_412),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_421),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_402),
.B(n_342),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_391),
.Y(n_519)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_442),
.B(n_377),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_393),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_393),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_421),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_SL g524 ( 
.A1(n_402),
.A2(n_362),
.B1(n_382),
.B2(n_206),
.Y(n_524)
);

BUFx3_ASAP7_75t_L g525 ( 
.A(n_415),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_402),
.B(n_361),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_L g527 ( 
.A1(n_405),
.A2(n_260),
.B1(n_264),
.B2(n_355),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_393),
.Y(n_528)
);

AND2x2_ASAP7_75t_SL g529 ( 
.A(n_405),
.B(n_262),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_409),
.B(n_422),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_388),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_393),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_421),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_427),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_395),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_415),
.Y(n_536)
);

INVx1_ASAP7_75t_SL g537 ( 
.A(n_435),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_409),
.B(n_370),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_427),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_388),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_388),
.Y(n_541)
);

AND2x4_ASAP7_75t_L g542 ( 
.A(n_415),
.B(n_234),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_452),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_395),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_402),
.B(n_371),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_409),
.B(n_325),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_SL g547 ( 
.A(n_402),
.B(n_364),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_395),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_402),
.B(n_382),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_427),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_395),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_447),
.B(n_366),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_427),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_447),
.B(n_367),
.Y(n_554)
);

NAND2xp33_ASAP7_75t_L g555 ( 
.A(n_411),
.B(n_180),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_406),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_427),
.Y(n_557)
);

BUFx3_ASAP7_75t_L g558 ( 
.A(n_415),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_409),
.B(n_325),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_406),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_427),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_388),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_388),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_424),
.B(n_373),
.Y(n_564)
);

NAND2xp33_ASAP7_75t_L g565 ( 
.A(n_411),
.B(n_180),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_406),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_410),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_409),
.B(n_375),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_410),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_410),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_413),
.Y(n_571)
);

BUFx6f_ASAP7_75t_SL g572 ( 
.A(n_409),
.Y(n_572)
);

AND2x4_ASAP7_75t_L g573 ( 
.A(n_411),
.B(n_237),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_390),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_424),
.B(n_376),
.Y(n_575)
);

BUFx4f_ASAP7_75t_L g576 ( 
.A(n_423),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_413),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_390),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_413),
.Y(n_579)
);

INVx2_ASAP7_75t_SL g580 ( 
.A(n_428),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_428),
.B(n_380),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_413),
.B(n_325),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_446),
.B(n_378),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_435),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_425),
.B(n_325),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_425),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_425),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_425),
.B(n_214),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_426),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_426),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_426),
.Y(n_591)
);

AND2x6_ASAP7_75t_L g592 ( 
.A(n_426),
.B(n_294),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_428),
.Y(n_593)
);

NOR2x1p5_ASAP7_75t_L g594 ( 
.A(n_446),
.B(n_273),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_429),
.Y(n_595)
);

OAI21xp5_ASAP7_75t_L g596 ( 
.A1(n_429),
.A2(n_239),
.B(n_237),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_429),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_429),
.Y(n_598)
);

OAI22xp33_ASAP7_75t_L g599 ( 
.A1(n_400),
.A2(n_304),
.B1(n_238),
.B2(n_278),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_414),
.B(n_250),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_390),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_428),
.B(n_253),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_390),
.Y(n_603)
);

OR2x2_ASAP7_75t_L g604 ( 
.A(n_435),
.B(n_281),
.Y(n_604)
);

INVx1_ASAP7_75t_SL g605 ( 
.A(n_445),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_386),
.Y(n_606)
);

OAI22xp33_ASAP7_75t_L g607 ( 
.A1(n_483),
.A2(n_246),
.B1(n_240),
.B2(n_298),
.Y(n_607)
);

BUFx2_ASAP7_75t_L g608 ( 
.A(n_543),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_488),
.B(n_445),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_474),
.B(n_315),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_461),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_497),
.B(n_187),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_474),
.B(n_326),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_529),
.B(n_423),
.Y(n_614)
);

INVx1_ASAP7_75t_SL g615 ( 
.A(n_467),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_529),
.B(n_423),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_479),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_479),
.Y(n_618)
);

OAI22xp33_ASAP7_75t_L g619 ( 
.A1(n_483),
.A2(n_239),
.B1(n_240),
.B2(n_298),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_499),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_530),
.B(n_499),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_499),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_470),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_525),
.B(n_423),
.Y(n_624)
);

INVx4_ASAP7_75t_SL g625 ( 
.A(n_466),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_525),
.B(n_423),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_470),
.Y(n_627)
);

O2A1O1Ixp33_ASAP7_75t_L g628 ( 
.A1(n_596),
.A2(n_469),
.B(n_472),
.C(n_471),
.Y(n_628)
);

OAI22xp33_ASAP7_75t_L g629 ( 
.A1(n_483),
.A2(n_246),
.B1(n_256),
.B2(n_284),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_507),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_507),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_605),
.B(n_160),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_511),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_525),
.B(n_423),
.Y(n_634)
);

NOR2x1p5_ASAP7_75t_SL g635 ( 
.A(n_521),
.B(n_414),
.Y(n_635)
);

INVx4_ASAP7_75t_L g636 ( 
.A(n_536),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_511),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_471),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_564),
.B(n_161),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_462),
.B(n_163),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_520),
.Y(n_641)
);

INVx8_ASAP7_75t_L g642 ( 
.A(n_572),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_536),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_L g644 ( 
.A1(n_466),
.A2(n_159),
.B1(n_164),
.B2(n_168),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_466),
.A2(n_328),
.B1(n_255),
.B2(n_306),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_472),
.Y(n_646)
);

AND2x4_ASAP7_75t_L g647 ( 
.A(n_520),
.B(n_281),
.Y(n_647)
);

BUFx2_ASAP7_75t_SL g648 ( 
.A(n_572),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_498),
.B(n_166),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_552),
.B(n_181),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_469),
.B(n_181),
.Y(n_651)
);

AOI22xp5_ASAP7_75t_L g652 ( 
.A1(n_466),
.A2(n_291),
.B1(n_297),
.B2(n_300),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_580),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_536),
.B(n_423),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_467),
.B(n_229),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_475),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_486),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_558),
.B(n_423),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_580),
.Y(n_659)
);

BUFx2_ASAP7_75t_L g660 ( 
.A(n_543),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_558),
.B(n_438),
.Y(n_661)
);

NOR3xp33_ASAP7_75t_L g662 ( 
.A(n_508),
.B(n_185),
.C(n_174),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_558),
.B(n_486),
.Y(n_663)
);

NAND2xp33_ASAP7_75t_L g664 ( 
.A(n_466),
.B(n_504),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_604),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_489),
.B(n_438),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_583),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_489),
.B(n_438),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_583),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_538),
.B(n_192),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_491),
.B(n_438),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_575),
.B(n_193),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_491),
.Y(n_673)
);

INVx2_ASAP7_75t_SL g674 ( 
.A(n_604),
.Y(n_674)
);

INVx4_ASAP7_75t_L g675 ( 
.A(n_572),
.Y(n_675)
);

OAI21xp33_ASAP7_75t_L g676 ( 
.A1(n_505),
.A2(n_164),
.B(n_159),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_493),
.B(n_438),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_593),
.B(n_542),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_493),
.B(n_494),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_593),
.B(n_542),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_483),
.B(n_463),
.Y(n_681)
);

BUFx12f_ASAP7_75t_SL g682 ( 
.A(n_483),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_494),
.B(n_438),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_606),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_496),
.B(n_438),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_460),
.Y(n_686)
);

INVxp33_ASAP7_75t_SL g687 ( 
.A(n_547),
.Y(n_687)
);

BUFx8_ASAP7_75t_L g688 ( 
.A(n_484),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_594),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_496),
.B(n_438),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_542),
.B(n_438),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_542),
.B(n_180),
.Y(n_692)
);

INVx2_ASAP7_75t_SL g693 ( 
.A(n_594),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_606),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_573),
.B(n_490),
.Y(n_695)
);

AOI22xp5_ASAP7_75t_L g696 ( 
.A1(n_482),
.A2(n_271),
.B1(n_275),
.B2(n_274),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_581),
.B(n_554),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_476),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_484),
.B(n_229),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_573),
.B(n_180),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_458),
.Y(n_701)
);

XNOR2xp5_ASAP7_75t_L g702 ( 
.A(n_524),
.B(n_244),
.Y(n_702)
);

INVx8_ASAP7_75t_L g703 ( 
.A(n_584),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_588),
.B(n_428),
.Y(n_704)
);

INVxp67_ASAP7_75t_L g705 ( 
.A(n_502),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_546),
.B(n_194),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_510),
.B(n_506),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_573),
.B(n_294),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_573),
.B(n_301),
.Y(n_709)
);

A2O1A1Ixp33_ASAP7_75t_L g710 ( 
.A1(n_490),
.A2(n_301),
.B(n_436),
.C(n_433),
.Y(n_710)
);

CKINVDCx8_ASAP7_75t_R g711 ( 
.A(n_510),
.Y(n_711)
);

INVxp67_ASAP7_75t_L g712 ( 
.A(n_502),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_510),
.B(n_506),
.Y(n_713)
);

OR2x2_ASAP7_75t_L g714 ( 
.A(n_481),
.B(n_198),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_458),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_559),
.B(n_269),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_509),
.B(n_433),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_568),
.B(n_199),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_490),
.B(n_509),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_514),
.B(n_433),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_478),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_517),
.Y(n_722)
);

NOR2xp67_ASAP7_75t_L g723 ( 
.A(n_518),
.B(n_400),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_490),
.B(n_433),
.Y(n_724)
);

OAI21xp33_ASAP7_75t_L g725 ( 
.A1(n_527),
.A2(n_172),
.B(n_168),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_517),
.Y(n_726)
);

NAND2x1_ASAP7_75t_L g727 ( 
.A(n_459),
.B(n_389),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_523),
.B(n_433),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_523),
.B(n_533),
.Y(n_729)
);

INVx2_ASAP7_75t_SL g730 ( 
.A(n_481),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_533),
.B(n_436),
.Y(n_731)
);

OR2x2_ASAP7_75t_L g732 ( 
.A(n_537),
.B(n_207),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_500),
.A2(n_268),
.B1(n_175),
.B2(n_178),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_478),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_526),
.A2(n_305),
.B1(n_436),
.B2(n_256),
.Y(n_735)
);

NOR2xp67_ASAP7_75t_L g736 ( 
.A(n_545),
.B(n_446),
.Y(n_736)
);

BUFx6f_ASAP7_75t_SL g737 ( 
.A(n_592),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_534),
.B(n_436),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_480),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_539),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_550),
.B(n_436),
.Y(n_741)
);

BUFx3_ASAP7_75t_L g742 ( 
.A(n_553),
.Y(n_742)
);

BUFx3_ASAP7_75t_L g743 ( 
.A(n_553),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_557),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_557),
.B(n_443),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_600),
.B(n_208),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_561),
.B(n_414),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_561),
.B(n_443),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_582),
.B(n_417),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_480),
.Y(n_750)
);

OR2x6_ASAP7_75t_L g751 ( 
.A(n_549),
.B(n_172),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_585),
.B(n_417),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_460),
.B(n_443),
.Y(n_753)
);

NOR3xp33_ASAP7_75t_L g754 ( 
.A(n_599),
.B(n_602),
.C(n_212),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_500),
.B(n_417),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_460),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_500),
.B(n_386),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_485),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_592),
.A2(n_175),
.B1(n_302),
.B2(n_178),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_459),
.B(n_386),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_485),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_460),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_566),
.Y(n_763)
);

INVxp67_ASAP7_75t_L g764 ( 
.A(n_555),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_459),
.B(n_396),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_667),
.B(n_566),
.Y(n_766)
);

A2O1A1Ixp33_ASAP7_75t_L g767 ( 
.A1(n_612),
.A2(n_249),
.B(n_254),
.C(n_279),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_667),
.B(n_669),
.Y(n_768)
);

OAI21xp5_ASAP7_75t_L g769 ( 
.A1(n_614),
.A2(n_512),
.B(n_477),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_643),
.B(n_460),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_621),
.A2(n_512),
.B(n_477),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_695),
.A2(n_512),
.B(n_477),
.Y(n_772)
);

INVx4_ASAP7_75t_L g773 ( 
.A(n_643),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_615),
.B(n_229),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_695),
.A2(n_576),
.B(n_515),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_616),
.A2(n_576),
.B(n_515),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_678),
.A2(n_503),
.B(n_495),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_643),
.Y(n_778)
);

A2O1A1Ixp33_ASAP7_75t_L g779 ( 
.A1(n_612),
.A2(n_285),
.B(n_190),
.C(n_195),
.Y(n_779)
);

A2O1A1Ixp33_ASAP7_75t_L g780 ( 
.A1(n_639),
.A2(n_249),
.B(n_254),
.C(n_279),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_678),
.A2(n_503),
.B(n_495),
.Y(n_781)
);

INVx2_ASAP7_75t_SL g782 ( 
.A(n_608),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_643),
.B(n_460),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_733),
.A2(n_190),
.B1(n_252),
.B2(n_285),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_655),
.B(n_229),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_611),
.B(n_567),
.Y(n_786)
);

INVx4_ASAP7_75t_L g787 ( 
.A(n_642),
.Y(n_787)
);

BUFx6f_ASAP7_75t_L g788 ( 
.A(n_756),
.Y(n_788)
);

INVx3_ASAP7_75t_L g789 ( 
.A(n_636),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_680),
.A2(n_503),
.B(n_495),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_609),
.B(n_639),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_618),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_618),
.B(n_746),
.Y(n_793)
);

AOI21xp33_ASAP7_75t_L g794 ( 
.A1(n_672),
.A2(n_565),
.B(n_284),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_650),
.B(n_378),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_680),
.A2(n_503),
.B(n_495),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_623),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_724),
.A2(n_531),
.B(n_464),
.Y(n_798)
);

AOI21xp33_ASAP7_75t_L g799 ( 
.A1(n_672),
.A2(n_282),
.B(n_213),
.Y(n_799)
);

AOI21x1_ASAP7_75t_L g800 ( 
.A1(n_658),
.A2(n_570),
.B(n_567),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_746),
.B(n_570),
.Y(n_801)
);

AND2x4_ASAP7_75t_L g802 ( 
.A(n_641),
.B(n_449),
.Y(n_802)
);

NOR3xp33_ASAP7_75t_L g803 ( 
.A(n_610),
.B(n_282),
.C(n_219),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_724),
.A2(n_531),
.B(n_464),
.Y(n_804)
);

BUFx2_ASAP7_75t_L g805 ( 
.A(n_660),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_617),
.B(n_571),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_704),
.A2(n_531),
.B(n_464),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_620),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_705),
.B(n_287),
.Y(n_809)
);

AOI21xp5_ASAP7_75t_L g810 ( 
.A1(n_664),
.A2(n_531),
.B(n_464),
.Y(n_810)
);

AOI21x1_ASAP7_75t_L g811 ( 
.A1(n_658),
.A2(n_579),
.B(n_577),
.Y(n_811)
);

A2O1A1Ixp33_ASAP7_75t_L g812 ( 
.A1(n_681),
.A2(n_296),
.B(n_179),
.C(n_195),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_624),
.A2(n_531),
.B(n_464),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_622),
.B(n_641),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_706),
.B(n_577),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_626),
.A2(n_601),
.B(n_501),
.Y(n_816)
);

OAI22xp5_ASAP7_75t_L g817 ( 
.A1(n_681),
.A2(n_299),
.B1(n_579),
.B2(n_591),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_634),
.A2(n_601),
.B(n_501),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_706),
.B(n_591),
.Y(n_819)
);

BUFx2_ASAP7_75t_L g820 ( 
.A(n_698),
.Y(n_820)
);

BUFx3_ASAP7_75t_L g821 ( 
.A(n_703),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_654),
.A2(n_601),
.B(n_501),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_623),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_627),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_691),
.A2(n_762),
.B(n_756),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_636),
.B(n_595),
.Y(n_826)
);

OAI21xp5_ASAP7_75t_L g827 ( 
.A1(n_707),
.A2(n_595),
.B(n_535),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_632),
.B(n_532),
.Y(n_828)
);

A2O1A1Ixp33_ASAP7_75t_L g829 ( 
.A1(n_697),
.A2(n_544),
.B(n_598),
.C(n_548),
.Y(n_829)
);

A2O1A1Ixp33_ASAP7_75t_L g830 ( 
.A1(n_697),
.A2(n_544),
.B(n_598),
.C(n_551),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_651),
.B(n_379),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_691),
.A2(n_601),
.B(n_501),
.Y(n_832)
);

A2O1A1Ixp33_ASAP7_75t_L g833 ( 
.A1(n_628),
.A2(n_551),
.B(n_556),
.C(n_590),
.Y(n_833)
);

OAI21xp5_ASAP7_75t_L g834 ( 
.A1(n_713),
.A2(n_548),
.B(n_535),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_756),
.Y(n_835)
);

OAI21xp5_ASAP7_75t_L g836 ( 
.A1(n_719),
.A2(n_560),
.B(n_556),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_756),
.A2(n_601),
.B(n_501),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_638),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_625),
.B(n_601),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_625),
.B(n_465),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_762),
.A2(n_501),
.B(n_473),
.Y(n_841)
);

OAI21xp5_ASAP7_75t_L g842 ( 
.A1(n_719),
.A2(n_586),
.B(n_560),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_638),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_762),
.A2(n_513),
.B(n_473),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_646),
.Y(n_845)
);

OAI21xp5_ASAP7_75t_L g846 ( 
.A1(n_661),
.A2(n_589),
.B(n_587),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_762),
.A2(n_513),
.B(n_473),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_663),
.A2(n_513),
.B(n_473),
.Y(n_848)
);

HB1xp67_ASAP7_75t_L g849 ( 
.A(n_665),
.Y(n_849)
);

BUFx6f_ASAP7_75t_L g850 ( 
.A(n_742),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_640),
.B(n_589),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_640),
.B(n_590),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_674),
.B(n_699),
.Y(n_853)
);

NOR2x1_ASAP7_75t_L g854 ( 
.A(n_675),
.B(n_465),
.Y(n_854)
);

OAI321xp33_ASAP7_75t_L g855 ( 
.A1(n_607),
.A2(n_235),
.A3(n_233),
.B1(n_228),
.B2(n_218),
.C(n_201),
.Y(n_855)
);

HB1xp67_ASAP7_75t_L g856 ( 
.A(n_730),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_679),
.A2(n_513),
.B(n_473),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_717),
.A2(n_516),
.B(n_513),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_712),
.B(n_521),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_720),
.A2(n_516),
.B(n_465),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_649),
.B(n_521),
.Y(n_861)
);

NOR2xp67_ASAP7_75t_L g862 ( 
.A(n_656),
.B(n_449),
.Y(n_862)
);

AO21x1_ASAP7_75t_L g863 ( 
.A1(n_757),
.A2(n_201),
.B(n_179),
.Y(n_863)
);

OR2x6_ASAP7_75t_L g864 ( 
.A(n_703),
.B(n_218),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_625),
.B(n_540),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_728),
.A2(n_516),
.B(n_603),
.Y(n_866)
);

CKINVDCx6p67_ASAP7_75t_R g867 ( 
.A(n_703),
.Y(n_867)
);

OAI21xp5_ASAP7_75t_L g868 ( 
.A1(n_755),
.A2(n_528),
.B(n_522),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_731),
.A2(n_516),
.B(n_603),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_630),
.B(n_379),
.Y(n_870)
);

AO21x1_ASAP7_75t_L g871 ( 
.A1(n_619),
.A2(n_233),
.B(n_228),
.Y(n_871)
);

AND2x4_ASAP7_75t_L g872 ( 
.A(n_631),
.B(n_449),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_723),
.B(n_540),
.Y(n_873)
);

AOI22xp5_ASAP7_75t_L g874 ( 
.A1(n_649),
.A2(n_592),
.B1(n_597),
.B2(n_522),
.Y(n_874)
);

NOR3xp33_ASAP7_75t_L g875 ( 
.A(n_613),
.B(n_259),
.C(n_209),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_741),
.A2(n_603),
.B(n_540),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_657),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_714),
.B(n_522),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_670),
.B(n_528),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_749),
.A2(n_540),
.B(n_541),
.Y(n_880)
);

AO21x1_ASAP7_75t_L g881 ( 
.A1(n_629),
.A2(n_252),
.B(n_302),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_742),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_752),
.A2(n_562),
.B(n_541),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_729),
.A2(n_562),
.B(n_541),
.Y(n_884)
);

AOI33xp33_ASAP7_75t_L g885 ( 
.A1(n_633),
.A2(n_235),
.A3(n_296),
.B1(n_295),
.B2(n_280),
.B3(n_268),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_729),
.A2(n_541),
.B(n_562),
.Y(n_886)
);

AND2x4_ASAP7_75t_L g887 ( 
.A(n_637),
.B(n_450),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_673),
.Y(n_888)
);

NOR3xp33_ASAP7_75t_L g889 ( 
.A(n_662),
.B(n_230),
.C(n_221),
.Y(n_889)
);

O2A1O1Ixp33_ASAP7_75t_L g890 ( 
.A1(n_708),
.A2(n_597),
.B(n_569),
.C(n_468),
.Y(n_890)
);

A2O1A1Ixp33_ASAP7_75t_L g891 ( 
.A1(n_718),
.A2(n_736),
.B(n_659),
.C(n_653),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_738),
.A2(n_563),
.B(n_578),
.Y(n_892)
);

A2O1A1Ixp33_ASAP7_75t_L g893 ( 
.A1(n_718),
.A2(n_597),
.B(n_569),
.C(n_574),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_684),
.B(n_569),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_673),
.B(n_694),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_647),
.B(n_381),
.Y(n_896)
);

AND2x4_ASAP7_75t_L g897 ( 
.A(n_689),
.B(n_450),
.Y(n_897)
);

O2A1O1Ixp5_ASAP7_75t_L g898 ( 
.A1(n_708),
.A2(n_492),
.B(n_519),
.C(n_487),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_694),
.B(n_563),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_722),
.Y(n_900)
);

A2O1A1Ixp33_ASAP7_75t_L g901 ( 
.A1(n_735),
.A2(n_578),
.B(n_574),
.C(n_563),
.Y(n_901)
);

AND2x4_ASAP7_75t_L g902 ( 
.A(n_693),
.B(n_450),
.Y(n_902)
);

AND2x2_ASAP7_75t_SL g903 ( 
.A(n_733),
.B(n_280),
.Y(n_903)
);

OAI21xp5_ASAP7_75t_L g904 ( 
.A1(n_666),
.A2(n_519),
.B(n_492),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_738),
.A2(n_574),
.B(n_487),
.Y(n_905)
);

AND2x2_ASAP7_75t_SL g906 ( 
.A(n_644),
.B(n_295),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_743),
.B(n_574),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_687),
.B(n_220),
.Y(n_908)
);

AOI22xp33_ASAP7_75t_L g909 ( 
.A1(n_644),
.A2(n_592),
.B1(n_468),
.B2(n_226),
.Y(n_909)
);

AOI22xp33_ASAP7_75t_L g910 ( 
.A1(n_709),
.A2(n_592),
.B1(n_468),
.B2(n_248),
.Y(n_910)
);

BUFx6f_ASAP7_75t_L g911 ( 
.A(n_743),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_682),
.B(n_251),
.Y(n_912)
);

HB1xp67_ASAP7_75t_L g913 ( 
.A(n_647),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_732),
.B(n_381),
.Y(n_914)
);

NOR2x1p5_ASAP7_75t_L g915 ( 
.A(n_675),
.B(n_258),
.Y(n_915)
);

BUFx4f_ASAP7_75t_L g916 ( 
.A(n_642),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_754),
.A2(n_453),
.B(n_457),
.C(n_455),
.Y(n_917)
);

NAND3xp33_ASAP7_75t_L g918 ( 
.A(n_702),
.B(n_261),
.C(n_308),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_686),
.A2(n_390),
.B(n_403),
.Y(n_919)
);

A2O1A1Ixp33_ASAP7_75t_L g920 ( 
.A1(n_635),
.A2(n_453),
.B(n_457),
.C(n_455),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_701),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_642),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_686),
.A2(n_390),
.B(n_403),
.Y(n_923)
);

INVx3_ASAP7_75t_L g924 ( 
.A(n_711),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_668),
.A2(n_390),
.B(n_403),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_671),
.A2(n_390),
.B(n_403),
.Y(n_926)
);

AOI33xp33_ASAP7_75t_L g927 ( 
.A1(n_759),
.A2(n_457),
.A3(n_455),
.B1(n_453),
.B2(n_441),
.B3(n_420),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_677),
.A2(n_390),
.B(n_392),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_SL g929 ( 
.A(n_645),
.B(n_443),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_683),
.A2(n_392),
.B(n_389),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_726),
.Y(n_931)
);

OAI321xp33_ASAP7_75t_L g932 ( 
.A1(n_676),
.A2(n_420),
.A3(n_432),
.B1(n_431),
.B2(n_430),
.C(n_441),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_740),
.B(n_443),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_SL g934 ( 
.A(n_648),
.B(n_265),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_744),
.Y(n_935)
);

AOI21xp33_ASAP7_75t_L g936 ( 
.A1(n_751),
.A2(n_266),
.B(n_267),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_R g937 ( 
.A(n_916),
.B(n_688),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_823),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_791),
.B(n_751),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_SL g940 ( 
.A(n_820),
.B(n_688),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_793),
.A2(n_709),
.B(n_685),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_795),
.B(n_764),
.Y(n_942)
);

OR2x6_ASAP7_75t_SL g943 ( 
.A(n_918),
.B(n_270),
.Y(n_943)
);

BUFx2_ASAP7_75t_L g944 ( 
.A(n_805),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_R g945 ( 
.A(n_916),
.B(n_737),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_850),
.B(n_696),
.Y(n_946)
);

BUFx4f_ASAP7_75t_L g947 ( 
.A(n_922),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_769),
.A2(n_690),
.B(n_710),
.Y(n_948)
);

A2O1A1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_799),
.A2(n_700),
.B(n_692),
.C(n_716),
.Y(n_949)
);

O2A1O1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_767),
.A2(n_700),
.B(n_692),
.C(n_725),
.Y(n_950)
);

O2A1O1Ixp5_ASAP7_75t_L g951 ( 
.A1(n_794),
.A2(n_929),
.B(n_863),
.C(n_771),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_831),
.B(n_763),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_908),
.B(n_652),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_787),
.B(n_701),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_772),
.A2(n_753),
.B(n_760),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_908),
.B(n_747),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_850),
.B(n_715),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_775),
.A2(n_765),
.B(n_727),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_878),
.B(n_859),
.Y(n_959)
);

OAI22xp5_ASAP7_75t_L g960 ( 
.A1(n_801),
.A2(n_759),
.B1(n_721),
.B2(n_758),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_877),
.Y(n_961)
);

A2O1A1Ixp33_ASAP7_75t_SL g962 ( 
.A1(n_889),
.A2(n_761),
.B(n_758),
.C(n_750),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_R g963 ( 
.A(n_924),
.B(n_737),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_888),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_911),
.B(n_862),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_859),
.B(n_721),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_L g967 ( 
.A(n_809),
.B(n_734),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_R g968 ( 
.A(n_924),
.B(n_739),
.Y(n_968)
);

BUFx12f_ASAP7_75t_L g969 ( 
.A(n_782),
.Y(n_969)
);

INVx3_ASAP7_75t_L g970 ( 
.A(n_778),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_914),
.B(n_761),
.Y(n_971)
);

AND2x4_ASAP7_75t_L g972 ( 
.A(n_787),
.B(n_745),
.Y(n_972)
);

NOR2xp67_ASAP7_75t_L g973 ( 
.A(n_853),
.B(n_61),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_792),
.Y(n_974)
);

O2A1O1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_812),
.A2(n_748),
.B(n_745),
.C(n_420),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_807),
.A2(n_748),
.B(n_389),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_802),
.B(n_397),
.Y(n_977)
);

A2O1A1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_891),
.A2(n_277),
.B(n_307),
.C(n_283),
.Y(n_978)
);

INVx3_ASAP7_75t_L g979 ( 
.A(n_778),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_797),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_785),
.B(n_288),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_809),
.B(n_303),
.Y(n_982)
);

A2O1A1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_768),
.A2(n_309),
.B(n_456),
.C(n_448),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_861),
.A2(n_389),
.B(n_392),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_824),
.Y(n_985)
);

BUFx3_ASAP7_75t_L g986 ( 
.A(n_821),
.Y(n_986)
);

INVx6_ASAP7_75t_L g987 ( 
.A(n_922),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_922),
.Y(n_988)
);

NOR2x1_ASAP7_75t_L g989 ( 
.A(n_773),
.B(n_882),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_922),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_911),
.B(n_448),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_911),
.B(n_778),
.Y(n_992)
);

NOR3xp33_ASAP7_75t_SL g993 ( 
.A(n_912),
.B(n_432),
.C(n_431),
.Y(n_993)
);

CKINVDCx16_ASAP7_75t_R g994 ( 
.A(n_934),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_879),
.A2(n_389),
.B(n_392),
.Y(n_995)
);

BUFx2_ASAP7_75t_L g996 ( 
.A(n_856),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_929),
.A2(n_392),
.B(n_403),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_856),
.B(n_7),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_849),
.B(n_9),
.Y(n_999)
);

O2A1O1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_812),
.A2(n_431),
.B(n_430),
.C(n_432),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_802),
.B(n_397),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_849),
.B(n_11),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_815),
.A2(n_397),
.B1(n_408),
.B2(n_398),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_913),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_776),
.A2(n_403),
.B(n_401),
.Y(n_1005)
);

INVx3_ASAP7_75t_L g1006 ( 
.A(n_778),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_911),
.B(n_456),
.Y(n_1007)
);

NOR3xp33_ASAP7_75t_SL g1008 ( 
.A(n_912),
.B(n_430),
.C(n_441),
.Y(n_1008)
);

O2A1O1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_779),
.A2(n_398),
.B(n_401),
.C(n_404),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_851),
.A2(n_404),
.B(n_407),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_814),
.B(n_404),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_913),
.B(n_12),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_852),
.A2(n_407),
.B(n_408),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_872),
.B(n_407),
.Y(n_1014)
);

BUFx3_ASAP7_75t_L g1015 ( 
.A(n_867),
.Y(n_1015)
);

O2A1O1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_779),
.A2(n_780),
.B(n_936),
.C(n_803),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_813),
.A2(n_819),
.B(n_810),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_872),
.B(n_408),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_838),
.Y(n_1019)
);

NAND2x1p5_ASAP7_75t_L g1020 ( 
.A(n_773),
.B(n_419),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_774),
.B(n_448),
.Y(n_1021)
);

BUFx3_ASAP7_75t_L g1022 ( 
.A(n_896),
.Y(n_1022)
);

A2O1A1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_803),
.A2(n_456),
.B(n_448),
.C(n_419),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_828),
.A2(n_419),
.B(n_454),
.C(n_451),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_843),
.Y(n_1025)
);

NOR3xp33_ASAP7_75t_SL g1026 ( 
.A(n_855),
.B(n_21),
.C(n_22),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_864),
.Y(n_1027)
);

O2A1O1Ixp5_ASAP7_75t_L g1028 ( 
.A1(n_917),
.A2(n_592),
.B(n_76),
.C(n_78),
.Y(n_1028)
);

O2A1O1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_817),
.A2(n_22),
.B(n_23),
.C(n_24),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_887),
.B(n_903),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_868),
.A2(n_454),
.B(n_451),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_887),
.B(n_454),
.Y(n_1032)
);

AND2x2_ASAP7_75t_L g1033 ( 
.A(n_870),
.B(n_443),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_897),
.B(n_85),
.Y(n_1034)
);

OAI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_789),
.A2(n_454),
.B1(n_451),
.B2(n_443),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_808),
.B(n_25),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_895),
.A2(n_454),
.B(n_451),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_827),
.A2(n_454),
.B(n_451),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_897),
.B(n_28),
.Y(n_1039)
);

O2A1O1Ixp5_ASAP7_75t_L g1040 ( 
.A1(n_873),
.A2(n_592),
.B(n_99),
.C(n_103),
.Y(n_1040)
);

INVxp67_ASAP7_75t_L g1041 ( 
.A(n_864),
.Y(n_1041)
);

OAI22xp33_ASAP7_75t_SL g1042 ( 
.A1(n_864),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_902),
.B(n_34),
.Y(n_1043)
);

NOR3xp33_ASAP7_75t_L g1044 ( 
.A(n_875),
.B(n_34),
.C(n_35),
.Y(n_1044)
);

OAI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_789),
.A2(n_454),
.B1(n_451),
.B2(n_443),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_R g1046 ( 
.A(n_900),
.B(n_114),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_826),
.A2(n_454),
.B(n_451),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_798),
.A2(n_451),
.B(n_443),
.Y(n_1048)
);

INVx1_ASAP7_75t_SL g1049 ( 
.A(n_902),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_804),
.A2(n_75),
.B(n_154),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_889),
.B(n_931),
.Y(n_1051)
);

NAND2x1p5_ASAP7_75t_L g1052 ( 
.A(n_788),
.B(n_67),
.Y(n_1052)
);

O2A1O1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_920),
.A2(n_35),
.B(n_39),
.C(n_40),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_901),
.A2(n_117),
.B(n_153),
.Y(n_1054)
);

AND2x2_ASAP7_75t_L g1055 ( 
.A(n_903),
.B(n_40),
.Y(n_1055)
);

A2O1A1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_935),
.A2(n_41),
.B(n_44),
.C(n_45),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_777),
.A2(n_122),
.B(n_152),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_915),
.B(n_92),
.Y(n_1058)
);

AND2x2_ASAP7_75t_SL g1059 ( 
.A(n_906),
.B(n_45),
.Y(n_1059)
);

A2O1A1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_784),
.A2(n_46),
.B(n_48),
.C(n_49),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_781),
.A2(n_130),
.B(n_143),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_790),
.A2(n_128),
.B(n_140),
.Y(n_1062)
);

OR2x2_ASAP7_75t_L g1063 ( 
.A(n_845),
.B(n_766),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_788),
.B(n_125),
.Y(n_1064)
);

INVx4_ASAP7_75t_L g1065 ( 
.A(n_788),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_921),
.Y(n_1066)
);

HB1xp67_ASAP7_75t_L g1067 ( 
.A(n_788),
.Y(n_1067)
);

BUFx6f_ASAP7_75t_SL g1068 ( 
.A(n_906),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_784),
.B(n_885),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_907),
.B(n_60),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_874),
.A2(n_876),
.B(n_890),
.C(n_796),
.Y(n_1071)
);

OAI21x1_ASAP7_75t_L g1072 ( 
.A1(n_1005),
.A2(n_800),
.B(n_811),
.Y(n_1072)
);

OR2x6_ASAP7_75t_L g1073 ( 
.A(n_1034),
.B(n_835),
.Y(n_1073)
);

O2A1O1Ixp33_ASAP7_75t_SL g1074 ( 
.A1(n_949),
.A2(n_839),
.B(n_840),
.C(n_865),
.Y(n_1074)
);

AOI221xp5_ASAP7_75t_L g1075 ( 
.A1(n_982),
.A2(n_871),
.B1(n_881),
.B2(n_932),
.C(n_910),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_938),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_1066),
.Y(n_1077)
);

NOR2xp67_ASAP7_75t_L g1078 ( 
.A(n_942),
.B(n_806),
.Y(n_1078)
);

OAI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_956),
.A2(n_905),
.B(n_892),
.Y(n_1079)
);

O2A1O1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_1051),
.A2(n_893),
.B(n_830),
.C(n_829),
.Y(n_1080)
);

HB1xp67_ASAP7_75t_L g1081 ( 
.A(n_996),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_L g1082 ( 
.A1(n_1005),
.A2(n_898),
.B(n_818),
.Y(n_1082)
);

AND2x4_ASAP7_75t_L g1083 ( 
.A(n_1022),
.B(n_854),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_959),
.A2(n_839),
.B(n_825),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_939),
.B(n_783),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_1071),
.A2(n_770),
.B(n_880),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_961),
.Y(n_1087)
);

NOR2xp67_ASAP7_75t_L g1088 ( 
.A(n_1021),
.B(n_952),
.Y(n_1088)
);

OAI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_953),
.A2(n_786),
.B1(n_835),
.B2(n_910),
.Y(n_1089)
);

OAI21x1_ASAP7_75t_L g1090 ( 
.A1(n_976),
.A2(n_898),
.B(n_822),
.Y(n_1090)
);

AOI221xp5_ASAP7_75t_SL g1091 ( 
.A1(n_1029),
.A2(n_909),
.B1(n_883),
.B2(n_894),
.C(n_933),
.Y(n_1091)
);

AOI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_1059),
.A2(n_909),
.B1(n_899),
.B2(n_836),
.Y(n_1092)
);

OAI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_951),
.A2(n_884),
.B(n_886),
.Y(n_1093)
);

O2A1O1Ixp33_ASAP7_75t_L g1094 ( 
.A1(n_1044),
.A2(n_833),
.B(n_865),
.C(n_840),
.Y(n_1094)
);

NOR2xp67_ASAP7_75t_SL g1095 ( 
.A(n_994),
.B(n_835),
.Y(n_1095)
);

AND2x4_ASAP7_75t_L g1096 ( 
.A(n_1049),
.B(n_835),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_948),
.A2(n_816),
.B(n_834),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_976),
.A2(n_958),
.B(n_997),
.Y(n_1098)
);

OA21x2_ASAP7_75t_L g1099 ( 
.A1(n_1031),
.A2(n_904),
.B(n_846),
.Y(n_1099)
);

BUFx12f_ASAP7_75t_L g1100 ( 
.A(n_969),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_1016),
.A2(n_927),
.B(n_930),
.C(n_860),
.Y(n_1101)
);

AND2x4_ASAP7_75t_L g1102 ( 
.A(n_986),
.B(n_842),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_941),
.A2(n_869),
.B(n_866),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_941),
.A2(n_848),
.B(n_857),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_L g1105 ( 
.A1(n_997),
.A2(n_928),
.B(n_926),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_955),
.A2(n_925),
.B(n_923),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_1030),
.A2(n_832),
.B1(n_858),
.B2(n_837),
.Y(n_1107)
);

INVx4_ASAP7_75t_L g1108 ( 
.A(n_947),
.Y(n_1108)
);

AO31x2_ASAP7_75t_L g1109 ( 
.A1(n_1024),
.A2(n_919),
.A3(n_847),
.B(n_844),
.Y(n_1109)
);

AO31x2_ASAP7_75t_L g1110 ( 
.A1(n_983),
.A2(n_841),
.A3(n_133),
.B(n_135),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_SL g1111 ( 
.A1(n_1068),
.A2(n_65),
.B(n_138),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_L g1112 ( 
.A1(n_984),
.A2(n_155),
.B(n_995),
.Y(n_1112)
);

AO31x2_ASAP7_75t_L g1113 ( 
.A1(n_1054),
.A2(n_978),
.A3(n_1023),
.B(n_1038),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_1068),
.A2(n_971),
.B1(n_967),
.B2(n_1069),
.Y(n_1114)
);

A2O1A1Ixp33_ASAP7_75t_L g1115 ( 
.A1(n_950),
.A2(n_1070),
.B(n_973),
.C(n_1008),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1063),
.B(n_981),
.Y(n_1116)
);

INVx2_ASAP7_75t_SL g1117 ( 
.A(n_947),
.Y(n_1117)
);

AOI221xp5_ASAP7_75t_L g1118 ( 
.A1(n_1055),
.A2(n_998),
.B1(n_999),
.B2(n_1002),
.C(n_1053),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_964),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_946),
.A2(n_966),
.B(n_960),
.Y(n_1120)
);

BUFx3_ASAP7_75t_L g1121 ( 
.A(n_1015),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_1054),
.A2(n_1033),
.B(n_1061),
.Y(n_1122)
);

AOI31xp67_ASAP7_75t_L g1123 ( 
.A1(n_1064),
.A2(n_957),
.A3(n_1011),
.B(n_991),
.Y(n_1123)
);

OAI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_1034),
.A2(n_974),
.B1(n_985),
.B2(n_1025),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_SL g1125 ( 
.A1(n_1057),
.A2(n_1050),
.B(n_1062),
.Y(n_1125)
);

INVx4_ASAP7_75t_L g1126 ( 
.A(n_988),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_980),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1057),
.A2(n_962),
.B(n_965),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1019),
.Y(n_1129)
);

BUFx2_ASAP7_75t_L g1130 ( 
.A(n_1004),
.Y(n_1130)
);

HB1xp67_ASAP7_75t_L g1131 ( 
.A(n_968),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_977),
.B(n_1001),
.Y(n_1132)
);

OA21x2_ASAP7_75t_L g1133 ( 
.A1(n_1048),
.A2(n_1047),
.B(n_1028),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_937),
.Y(n_1134)
);

OR2x2_ASAP7_75t_L g1135 ( 
.A(n_1014),
.B(n_1018),
.Y(n_1135)
);

AO31x2_ASAP7_75t_L g1136 ( 
.A1(n_1003),
.A2(n_1047),
.A3(n_1013),
.B(n_1010),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1039),
.B(n_1043),
.Y(n_1137)
);

A2O1A1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_993),
.A2(n_1026),
.B(n_1036),
.C(n_975),
.Y(n_1138)
);

O2A1O1Ixp33_ASAP7_75t_SL g1139 ( 
.A1(n_1060),
.A2(n_1056),
.B(n_992),
.C(n_1032),
.Y(n_1139)
);

HB1xp67_ASAP7_75t_L g1140 ( 
.A(n_1067),
.Y(n_1140)
);

BUFx10_ASAP7_75t_L g1141 ( 
.A(n_1012),
.Y(n_1141)
);

BUFx3_ASAP7_75t_L g1142 ( 
.A(n_988),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_1037),
.A2(n_1050),
.B(n_1020),
.Y(n_1143)
);

OA21x2_ASAP7_75t_L g1144 ( 
.A1(n_1037),
.A2(n_1040),
.B(n_1007),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_943),
.B(n_1041),
.Y(n_1145)
);

INVx6_ASAP7_75t_L g1146 ( 
.A(n_990),
.Y(n_1146)
);

CKINVDCx11_ASAP7_75t_R g1147 ( 
.A(n_990),
.Y(n_1147)
);

O2A1O1Ixp5_ASAP7_75t_SL g1148 ( 
.A1(n_970),
.A2(n_979),
.B(n_1006),
.C(n_1035),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_1020),
.A2(n_1045),
.B(n_989),
.Y(n_1149)
);

O2A1O1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_1042),
.A2(n_1058),
.B(n_1000),
.C(n_1009),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_954),
.A2(n_972),
.B(n_1065),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_954),
.A2(n_972),
.B(n_979),
.Y(n_1152)
);

NAND3xp33_ASAP7_75t_L g1153 ( 
.A(n_940),
.B(n_1058),
.C(n_1027),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_963),
.B(n_1046),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1052),
.A2(n_945),
.B(n_987),
.Y(n_1155)
);

AOI22xp33_ASAP7_75t_L g1156 ( 
.A1(n_987),
.A2(n_953),
.B1(n_1059),
.B2(n_639),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_987),
.B(n_1052),
.Y(n_1157)
);

AOI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_1059),
.A2(n_953),
.B1(n_612),
.B2(n_639),
.Y(n_1158)
);

BUFx2_ASAP7_75t_L g1159 ( 
.A(n_944),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1017),
.A2(n_791),
.B(n_621),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_938),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_956),
.B(n_994),
.Y(n_1162)
);

AND2x4_ASAP7_75t_L g1163 ( 
.A(n_1022),
.B(n_922),
.Y(n_1163)
);

AO31x2_ASAP7_75t_L g1164 ( 
.A1(n_1071),
.A2(n_863),
.A3(n_1024),
.B(n_1017),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_956),
.B(n_959),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_1017),
.A2(n_791),
.B(n_621),
.Y(n_1166)
);

A2O1A1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_953),
.A2(n_681),
.B(n_639),
.C(n_1016),
.Y(n_1167)
);

OR2x6_ASAP7_75t_L g1168 ( 
.A(n_1034),
.B(n_922),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1017),
.A2(n_791),
.B(n_621),
.Y(n_1169)
);

INVxp67_ASAP7_75t_L g1170 ( 
.A(n_996),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1017),
.A2(n_791),
.B(n_621),
.Y(n_1171)
);

AO21x2_ASAP7_75t_L g1172 ( 
.A1(n_1017),
.A2(n_948),
.B(n_1071),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1017),
.A2(n_791),
.B(n_621),
.Y(n_1173)
);

O2A1O1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_982),
.A2(n_799),
.B(n_639),
.C(n_612),
.Y(n_1174)
);

O2A1O1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_982),
.A2(n_799),
.B(n_639),
.C(n_612),
.Y(n_1175)
);

AND2x2_ASAP7_75t_L g1176 ( 
.A(n_981),
.B(n_615),
.Y(n_1176)
);

CKINVDCx20_ASAP7_75t_R g1177 ( 
.A(n_994),
.Y(n_1177)
);

INVx3_ASAP7_75t_L g1178 ( 
.A(n_954),
.Y(n_1178)
);

A2O1A1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_953),
.A2(n_681),
.B(n_639),
.C(n_1016),
.Y(n_1179)
);

O2A1O1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_982),
.A2(n_799),
.B(n_639),
.C(n_612),
.Y(n_1180)
);

OAI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_956),
.A2(n_791),
.B(n_939),
.Y(n_1181)
);

AOI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1059),
.A2(n_953),
.B1(n_612),
.B2(n_639),
.Y(n_1182)
);

NOR2xp67_ASAP7_75t_SL g1183 ( 
.A(n_994),
.B(n_656),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_938),
.Y(n_1184)
);

A2O1A1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_953),
.A2(n_681),
.B(n_639),
.C(n_1016),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_L g1186 ( 
.A(n_956),
.B(n_959),
.Y(n_1186)
);

AOI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1059),
.A2(n_953),
.B1(n_612),
.B2(n_639),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1017),
.A2(n_791),
.B(n_621),
.Y(n_1188)
);

AOI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1059),
.A2(n_953),
.B1(n_612),
.B2(n_639),
.Y(n_1189)
);

CKINVDCx11_ASAP7_75t_R g1190 ( 
.A(n_969),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_956),
.B(n_959),
.Y(n_1191)
);

O2A1O1Ixp33_ASAP7_75t_SL g1192 ( 
.A1(n_949),
.A2(n_978),
.B(n_791),
.C(n_780),
.Y(n_1192)
);

NOR3xp33_ASAP7_75t_L g1193 ( 
.A(n_953),
.B(n_639),
.C(n_799),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_L g1194 ( 
.A(n_956),
.B(n_315),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1017),
.A2(n_791),
.B(n_621),
.Y(n_1195)
);

BUFx3_ASAP7_75t_L g1196 ( 
.A(n_969),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_953),
.A2(n_1059),
.B1(n_639),
.B2(n_799),
.Y(n_1197)
);

NAND2xp33_ASAP7_75t_L g1198 ( 
.A(n_945),
.B(n_922),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1005),
.A2(n_976),
.B(n_958),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1017),
.A2(n_791),
.B(n_621),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_L g1201 ( 
.A(n_956),
.B(n_315),
.Y(n_1201)
);

AO31x2_ASAP7_75t_L g1202 ( 
.A1(n_1071),
.A2(n_863),
.A3(n_1024),
.B(n_1017),
.Y(n_1202)
);

O2A1O1Ixp33_ASAP7_75t_SL g1203 ( 
.A1(n_949),
.A2(n_978),
.B(n_791),
.C(n_780),
.Y(n_1203)
);

AO31x2_ASAP7_75t_L g1204 ( 
.A1(n_1071),
.A2(n_863),
.A3(n_1024),
.B(n_1017),
.Y(n_1204)
);

O2A1O1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_982),
.A2(n_799),
.B(n_639),
.C(n_612),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1005),
.A2(n_976),
.B(n_958),
.Y(n_1206)
);

AO31x2_ASAP7_75t_L g1207 ( 
.A1(n_1071),
.A2(n_863),
.A3(n_1024),
.B(n_1017),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1005),
.A2(n_976),
.B(n_958),
.Y(n_1208)
);

INVx1_ASAP7_75t_SL g1209 ( 
.A(n_1159),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_SL g1210 ( 
.A1(n_1194),
.A2(n_1201),
.B1(n_1141),
.B2(n_1165),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1076),
.Y(n_1211)
);

BUFx8_ASAP7_75t_L g1212 ( 
.A(n_1100),
.Y(n_1212)
);

BUFx6f_ASAP7_75t_L g1213 ( 
.A(n_1147),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1186),
.B(n_1191),
.Y(n_1214)
);

INVx4_ASAP7_75t_L g1215 ( 
.A(n_1108),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_SL g1216 ( 
.A1(n_1141),
.A2(n_1153),
.B1(n_1137),
.B2(n_1189),
.Y(n_1216)
);

BUFx6f_ASAP7_75t_L g1217 ( 
.A(n_1168),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1193),
.A2(n_1182),
.B1(n_1187),
.B2(n_1158),
.Y(n_1218)
);

CKINVDCx11_ASAP7_75t_R g1219 ( 
.A(n_1190),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_SL g1220 ( 
.A1(n_1158),
.A2(n_1189),
.B1(n_1187),
.B2(n_1182),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1087),
.Y(n_1221)
);

CKINVDCx11_ASAP7_75t_R g1222 ( 
.A(n_1177),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1197),
.A2(n_1118),
.B1(n_1156),
.B2(n_1181),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1176),
.B(n_1116),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1075),
.A2(n_1114),
.B1(n_1078),
.B2(n_1162),
.Y(n_1225)
);

OAI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1167),
.A2(n_1179),
.B1(n_1185),
.B2(n_1180),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_L g1227 ( 
.A1(n_1078),
.A2(n_1135),
.B1(n_1085),
.B2(n_1132),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_1134),
.Y(n_1228)
);

CKINVDCx20_ASAP7_75t_R g1229 ( 
.A(n_1196),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1119),
.Y(n_1230)
);

AOI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1145),
.A2(n_1088),
.B1(n_1120),
.B2(n_1205),
.Y(n_1231)
);

INVx3_ASAP7_75t_SL g1232 ( 
.A(n_1163),
.Y(n_1232)
);

AOI22xp33_ASAP7_75t_L g1233 ( 
.A1(n_1088),
.A2(n_1175),
.B1(n_1174),
.B2(n_1129),
.Y(n_1233)
);

CKINVDCx20_ASAP7_75t_R g1234 ( 
.A(n_1154),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1073),
.A2(n_1168),
.B1(n_1131),
.B2(n_1138),
.Y(n_1235)
);

INVx1_ASAP7_75t_SL g1236 ( 
.A(n_1130),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1073),
.A2(n_1168),
.B1(n_1124),
.B2(n_1115),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1161),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1127),
.A2(n_1172),
.B1(n_1102),
.B2(n_1184),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_SL g1240 ( 
.A1(n_1089),
.A2(n_1102),
.B1(n_1125),
.B2(n_1083),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1183),
.B(n_1081),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1172),
.A2(n_1092),
.B1(n_1077),
.B2(n_1079),
.Y(n_1242)
);

BUFx2_ASAP7_75t_L g1243 ( 
.A(n_1170),
.Y(n_1243)
);

BUFx3_ASAP7_75t_L g1244 ( 
.A(n_1121),
.Y(n_1244)
);

INVx4_ASAP7_75t_L g1245 ( 
.A(n_1146),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1095),
.B(n_1140),
.Y(n_1246)
);

BUFx3_ASAP7_75t_L g1247 ( 
.A(n_1142),
.Y(n_1247)
);

BUFx8_ASAP7_75t_SL g1248 ( 
.A(n_1073),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1096),
.B(n_1178),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_1146),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1160),
.A2(n_1171),
.B1(n_1200),
.B2(n_1169),
.Y(n_1251)
);

CKINVDCx6p67_ASAP7_75t_R g1252 ( 
.A(n_1126),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1157),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_1117),
.Y(n_1254)
);

OAI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1151),
.A2(n_1150),
.B1(n_1152),
.B2(n_1155),
.Y(n_1255)
);

INVx6_ASAP7_75t_L g1256 ( 
.A(n_1126),
.Y(n_1256)
);

AOI22xp5_ASAP7_75t_SL g1257 ( 
.A1(n_1111),
.A2(n_1128),
.B1(n_1084),
.B2(n_1107),
.Y(n_1257)
);

CKINVDCx11_ASAP7_75t_R g1258 ( 
.A(n_1198),
.Y(n_1258)
);

INVx5_ASAP7_75t_L g1259 ( 
.A(n_1139),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1094),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_SL g1261 ( 
.A1(n_1122),
.A2(n_1093),
.B1(n_1097),
.B2(n_1188),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1166),
.A2(n_1195),
.B1(n_1173),
.B2(n_1099),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1192),
.B(n_1203),
.Y(n_1263)
);

OAI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1101),
.A2(n_1086),
.B1(n_1080),
.B2(n_1099),
.Y(n_1264)
);

BUFx2_ASAP7_75t_R g1265 ( 
.A(n_1148),
.Y(n_1265)
);

OAI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1144),
.A2(n_1103),
.B1(n_1104),
.B2(n_1133),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1074),
.Y(n_1267)
);

BUFx3_ASAP7_75t_L g1268 ( 
.A(n_1112),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1133),
.A2(n_1072),
.B1(n_1143),
.B2(n_1098),
.Y(n_1269)
);

OAI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1123),
.A2(n_1091),
.B1(n_1113),
.B2(n_1204),
.Y(n_1270)
);

CKINVDCx11_ASAP7_75t_R g1271 ( 
.A(n_1110),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_1110),
.Y(n_1272)
);

OAI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1113),
.A2(n_1164),
.B1(n_1207),
.B2(n_1204),
.Y(n_1273)
);

INVx6_ASAP7_75t_L g1274 ( 
.A(n_1110),
.Y(n_1274)
);

CKINVDCx6p67_ASAP7_75t_R g1275 ( 
.A(n_1149),
.Y(n_1275)
);

CKINVDCx6p67_ASAP7_75t_R g1276 ( 
.A(n_1164),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_SL g1277 ( 
.A1(n_1199),
.A2(n_1208),
.B1(n_1206),
.B2(n_1106),
.Y(n_1277)
);

BUFx12f_ASAP7_75t_L g1278 ( 
.A(n_1164),
.Y(n_1278)
);

BUFx3_ASAP7_75t_L g1279 ( 
.A(n_1202),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1105),
.A2(n_1090),
.B1(n_1082),
.B2(n_1207),
.Y(n_1280)
);

OAI22x1_ASAP7_75t_L g1281 ( 
.A1(n_1202),
.A2(n_1204),
.B1(n_1207),
.B2(n_1136),
.Y(n_1281)
);

OAI22xp33_ASAP7_75t_L g1282 ( 
.A1(n_1136),
.A2(n_1158),
.B1(n_1187),
.B2(n_1182),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1109),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1193),
.A2(n_1158),
.B1(n_1187),
.B2(n_1182),
.Y(n_1284)
);

INVx5_ASAP7_75t_L g1285 ( 
.A(n_1108),
.Y(n_1285)
);

CKINVDCx6p67_ASAP7_75t_R g1286 ( 
.A(n_1190),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1193),
.A2(n_1158),
.B1(n_1187),
.B2(n_1182),
.Y(n_1287)
);

BUFx3_ASAP7_75t_L g1288 ( 
.A(n_1159),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_SL g1289 ( 
.A1(n_1194),
.A2(n_1059),
.B1(n_1068),
.B2(n_1201),
.Y(n_1289)
);

BUFx2_ASAP7_75t_L g1290 ( 
.A(n_1159),
.Y(n_1290)
);

CKINVDCx11_ASAP7_75t_R g1291 ( 
.A(n_1190),
.Y(n_1291)
);

AND2x2_ASAP7_75t_L g1292 ( 
.A(n_1176),
.B(n_1137),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1193),
.A2(n_1158),
.B1(n_1187),
.B2(n_1182),
.Y(n_1293)
);

OAI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1158),
.A2(n_1182),
.B1(n_1189),
.B2(n_1187),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_SL g1295 ( 
.A1(n_1194),
.A2(n_1059),
.B1(n_1068),
.B2(n_1201),
.Y(n_1295)
);

INVx2_ASAP7_75t_SL g1296 ( 
.A(n_1121),
.Y(n_1296)
);

BUFx4f_ASAP7_75t_SL g1297 ( 
.A(n_1100),
.Y(n_1297)
);

NAND2x1p5_ASAP7_75t_L g1298 ( 
.A(n_1095),
.B(n_1108),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1193),
.A2(n_1158),
.B1(n_1187),
.B2(n_1182),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1076),
.Y(n_1300)
);

BUFx2_ASAP7_75t_L g1301 ( 
.A(n_1159),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1193),
.A2(n_1158),
.B1(n_1187),
.B2(n_1182),
.Y(n_1302)
);

CKINVDCx20_ASAP7_75t_R g1303 ( 
.A(n_1177),
.Y(n_1303)
);

INVx4_ASAP7_75t_L g1304 ( 
.A(n_1108),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_SL g1305 ( 
.A1(n_1194),
.A2(n_1059),
.B1(n_1068),
.B2(n_1201),
.Y(n_1305)
);

INVx2_ASAP7_75t_SL g1306 ( 
.A(n_1121),
.Y(n_1306)
);

BUFx2_ASAP7_75t_SL g1307 ( 
.A(n_1108),
.Y(n_1307)
);

BUFx6f_ASAP7_75t_L g1308 ( 
.A(n_1147),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1193),
.A2(n_1158),
.B1(n_1187),
.B2(n_1182),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1158),
.A2(n_1187),
.B1(n_1189),
.B2(n_1182),
.Y(n_1310)
);

CKINVDCx11_ASAP7_75t_R g1311 ( 
.A(n_1190),
.Y(n_1311)
);

BUFx2_ASAP7_75t_L g1312 ( 
.A(n_1159),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1193),
.A2(n_1158),
.B1(n_1187),
.B2(n_1182),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1193),
.A2(n_1158),
.B1(n_1187),
.B2(n_1182),
.Y(n_1314)
);

BUFx8_ASAP7_75t_L g1315 ( 
.A(n_1100),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1158),
.A2(n_1187),
.B1(n_1189),
.B2(n_1182),
.Y(n_1316)
);

BUFx8_ASAP7_75t_SL g1317 ( 
.A(n_1100),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1158),
.A2(n_1187),
.B1(n_1189),
.B2(n_1182),
.Y(n_1318)
);

NAND2x1p5_ASAP7_75t_L g1319 ( 
.A(n_1095),
.B(n_1108),
.Y(n_1319)
);

INVx11_ASAP7_75t_L g1320 ( 
.A(n_1100),
.Y(n_1320)
);

BUFx2_ASAP7_75t_L g1321 ( 
.A(n_1159),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1076),
.Y(n_1322)
);

INVx6_ASAP7_75t_L g1323 ( 
.A(n_1108),
.Y(n_1323)
);

CKINVDCx20_ASAP7_75t_R g1324 ( 
.A(n_1177),
.Y(n_1324)
);

HB1xp67_ASAP7_75t_L g1325 ( 
.A(n_1283),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1218),
.B(n_1284),
.Y(n_1326)
);

INVx2_ASAP7_75t_SL g1327 ( 
.A(n_1274),
.Y(n_1327)
);

AOI21xp33_ASAP7_75t_L g1328 ( 
.A1(n_1226),
.A2(n_1223),
.B(n_1294),
.Y(n_1328)
);

HB1xp67_ASAP7_75t_SL g1329 ( 
.A(n_1213),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1279),
.Y(n_1330)
);

INVx3_ASAP7_75t_L g1331 ( 
.A(n_1278),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1214),
.B(n_1227),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1269),
.A2(n_1251),
.B(n_1262),
.Y(n_1333)
);

BUFx2_ASAP7_75t_L g1334 ( 
.A(n_1278),
.Y(n_1334)
);

OAI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1223),
.A2(n_1287),
.B(n_1284),
.Y(n_1335)
);

HB1xp67_ASAP7_75t_L g1336 ( 
.A(n_1281),
.Y(n_1336)
);

HB1xp67_ASAP7_75t_L g1337 ( 
.A(n_1273),
.Y(n_1337)
);

BUFx2_ASAP7_75t_L g1338 ( 
.A(n_1272),
.Y(n_1338)
);

INVx3_ASAP7_75t_L g1339 ( 
.A(n_1268),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1287),
.B(n_1293),
.Y(n_1340)
);

OAI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1310),
.A2(n_1318),
.B1(n_1316),
.B2(n_1259),
.Y(n_1341)
);

BUFx3_ASAP7_75t_L g1342 ( 
.A(n_1217),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1220),
.A2(n_1313),
.B1(n_1309),
.B2(n_1293),
.Y(n_1343)
);

BUFx2_ASAP7_75t_L g1344 ( 
.A(n_1276),
.Y(n_1344)
);

INVx4_ASAP7_75t_L g1345 ( 
.A(n_1259),
.Y(n_1345)
);

INVx4_ASAP7_75t_L g1346 ( 
.A(n_1259),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1267),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1260),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1299),
.B(n_1302),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1280),
.A2(n_1270),
.B(n_1264),
.Y(n_1350)
);

NAND3xp33_ASAP7_75t_L g1351 ( 
.A(n_1299),
.B(n_1313),
.C(n_1314),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1302),
.A2(n_1309),
.B1(n_1314),
.B2(n_1282),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1211),
.Y(n_1353)
);

OR2x2_ASAP7_75t_L g1354 ( 
.A(n_1242),
.B(n_1239),
.Y(n_1354)
);

NOR2xp33_ASAP7_75t_L g1355 ( 
.A(n_1292),
.B(n_1210),
.Y(n_1355)
);

AO21x2_ASAP7_75t_L g1356 ( 
.A1(n_1266),
.A2(n_1263),
.B(n_1255),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1221),
.Y(n_1357)
);

OR2x2_ASAP7_75t_L g1358 ( 
.A(n_1227),
.B(n_1233),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1233),
.B(n_1231),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1230),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1238),
.Y(n_1361)
);

INVx3_ASAP7_75t_L g1362 ( 
.A(n_1275),
.Y(n_1362)
);

BUFx6f_ASAP7_75t_L g1363 ( 
.A(n_1259),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1300),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1322),
.Y(n_1365)
);

NAND2x1_ASAP7_75t_L g1366 ( 
.A(n_1231),
.B(n_1253),
.Y(n_1366)
);

INVx2_ASAP7_75t_SL g1367 ( 
.A(n_1285),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1240),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1271),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1271),
.Y(n_1370)
);

AOI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1216),
.A2(n_1289),
.B1(n_1295),
.B2(n_1305),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1261),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1225),
.B(n_1224),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1277),
.Y(n_1374)
);

NOR2xp33_ASAP7_75t_L g1375 ( 
.A(n_1234),
.B(n_1209),
.Y(n_1375)
);

HB1xp67_ASAP7_75t_SL g1376 ( 
.A(n_1213),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1237),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1225),
.B(n_1257),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1235),
.A2(n_1298),
.B(n_1319),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1265),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1249),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1246),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1298),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1319),
.Y(n_1384)
);

HB1xp67_ASAP7_75t_L g1385 ( 
.A(n_1290),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1301),
.Y(n_1386)
);

BUFx3_ASAP7_75t_L g1387 ( 
.A(n_1248),
.Y(n_1387)
);

INVxp67_ASAP7_75t_L g1388 ( 
.A(n_1312),
.Y(n_1388)
);

AND2x2_ASAP7_75t_L g1389 ( 
.A(n_1232),
.B(n_1288),
.Y(n_1389)
);

BUFx3_ASAP7_75t_L g1390 ( 
.A(n_1248),
.Y(n_1390)
);

HB1xp67_ASAP7_75t_L g1391 ( 
.A(n_1321),
.Y(n_1391)
);

CKINVDCx11_ASAP7_75t_R g1392 ( 
.A(n_1387),
.Y(n_1392)
);

OAI21xp33_ASAP7_75t_SL g1393 ( 
.A1(n_1371),
.A2(n_1241),
.B(n_1215),
.Y(n_1393)
);

AOI221xp5_ASAP7_75t_L g1394 ( 
.A1(n_1328),
.A2(n_1236),
.B1(n_1243),
.B2(n_1288),
.C(n_1306),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1360),
.Y(n_1395)
);

OR2x2_ASAP7_75t_L g1396 ( 
.A(n_1382),
.B(n_1213),
.Y(n_1396)
);

BUFx6f_ASAP7_75t_L g1397 ( 
.A(n_1387),
.Y(n_1397)
);

O2A1O1Ixp33_ASAP7_75t_L g1398 ( 
.A1(n_1328),
.A2(n_1296),
.B(n_1244),
.C(n_1247),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_1329),
.Y(n_1399)
);

AO21x2_ASAP7_75t_L g1400 ( 
.A1(n_1333),
.A2(n_1258),
.B(n_1307),
.Y(n_1400)
);

NAND2x1p5_ASAP7_75t_L g1401 ( 
.A(n_1363),
.B(n_1215),
.Y(n_1401)
);

AND2x4_ASAP7_75t_L g1402 ( 
.A(n_1331),
.B(n_1213),
.Y(n_1402)
);

AND2x4_ASAP7_75t_L g1403 ( 
.A(n_1331),
.B(n_1308),
.Y(n_1403)
);

OAI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1351),
.A2(n_1335),
.B(n_1343),
.Y(n_1404)
);

OAI22xp5_ASAP7_75t_L g1405 ( 
.A1(n_1371),
.A2(n_1308),
.B1(n_1254),
.B2(n_1323),
.Y(n_1405)
);

OAI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1335),
.A2(n_1304),
.B(n_1303),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1353),
.Y(n_1407)
);

A2O1A1Ixp33_ASAP7_75t_L g1408 ( 
.A1(n_1378),
.A2(n_1308),
.B(n_1258),
.C(n_1244),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1369),
.B(n_1308),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1369),
.B(n_1222),
.Y(n_1410)
);

OR2x2_ASAP7_75t_L g1411 ( 
.A(n_1382),
.B(n_1381),
.Y(n_1411)
);

AOI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1366),
.A2(n_1252),
.B(n_1323),
.Y(n_1412)
);

AOI21xp33_ASAP7_75t_L g1413 ( 
.A1(n_1359),
.A2(n_1304),
.B(n_1324),
.Y(n_1413)
);

AO32x2_ASAP7_75t_L g1414 ( 
.A1(n_1327),
.A2(n_1245),
.A3(n_1222),
.B1(n_1323),
.B2(n_1256),
.Y(n_1414)
);

HB1xp67_ASAP7_75t_L g1415 ( 
.A(n_1325),
.Y(n_1415)
);

OA21x2_ASAP7_75t_L g1416 ( 
.A1(n_1350),
.A2(n_1250),
.B(n_1228),
.Y(n_1416)
);

OR2x6_ASAP7_75t_L g1417 ( 
.A(n_1379),
.B(n_1256),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_1329),
.Y(n_1418)
);

OAI211xp5_ASAP7_75t_SL g1419 ( 
.A1(n_1352),
.A2(n_1332),
.B(n_1359),
.C(n_1388),
.Y(n_1419)
);

AOI221xp5_ASAP7_75t_L g1420 ( 
.A1(n_1341),
.A2(n_1326),
.B1(n_1349),
.B2(n_1340),
.C(n_1378),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1326),
.A2(n_1291),
.B1(n_1219),
.B2(n_1311),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_1376),
.Y(n_1422)
);

NOR2x1_ASAP7_75t_SL g1423 ( 
.A(n_1363),
.B(n_1219),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1370),
.B(n_1229),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1332),
.B(n_1286),
.Y(n_1425)
);

OAI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1378),
.A2(n_1212),
.B(n_1315),
.Y(n_1426)
);

AOI21xp5_ASAP7_75t_SL g1427 ( 
.A1(n_1363),
.A2(n_1291),
.B(n_1311),
.Y(n_1427)
);

INVxp67_ASAP7_75t_SL g1428 ( 
.A(n_1325),
.Y(n_1428)
);

CKINVDCx14_ASAP7_75t_R g1429 ( 
.A(n_1387),
.Y(n_1429)
);

A2O1A1Ixp33_ASAP7_75t_L g1430 ( 
.A1(n_1340),
.A2(n_1349),
.B(n_1366),
.C(n_1358),
.Y(n_1430)
);

NAND2x1_ASAP7_75t_L g1431 ( 
.A(n_1362),
.B(n_1345),
.Y(n_1431)
);

A2O1A1Ixp33_ASAP7_75t_L g1432 ( 
.A1(n_1358),
.A2(n_1368),
.B(n_1377),
.C(n_1372),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1370),
.B(n_1320),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1348),
.B(n_1212),
.Y(n_1434)
);

A2O1A1Ixp33_ASAP7_75t_L g1435 ( 
.A1(n_1355),
.A2(n_1212),
.B(n_1315),
.C(n_1297),
.Y(n_1435)
);

AND2x4_ASAP7_75t_L g1436 ( 
.A(n_1331),
.B(n_1315),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1370),
.B(n_1317),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1348),
.B(n_1317),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1353),
.Y(n_1439)
);

A2O1A1Ixp33_ASAP7_75t_L g1440 ( 
.A1(n_1377),
.A2(n_1368),
.B(n_1338),
.C(n_1379),
.Y(n_1440)
);

O2A1O1Ixp33_ASAP7_75t_L g1441 ( 
.A1(n_1341),
.A2(n_1377),
.B(n_1380),
.C(n_1372),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1376),
.A2(n_1380),
.B1(n_1338),
.B2(n_1373),
.Y(n_1442)
);

OR2x6_ASAP7_75t_L g1443 ( 
.A(n_1379),
.B(n_1344),
.Y(n_1443)
);

AND2x4_ASAP7_75t_L g1444 ( 
.A(n_1331),
.B(n_1342),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1381),
.B(n_1389),
.Y(n_1445)
);

AO32x1_ASAP7_75t_L g1446 ( 
.A1(n_1345),
.A2(n_1346),
.A3(n_1347),
.B1(n_1373),
.B2(n_1330),
.Y(n_1446)
);

OR2x2_ASAP7_75t_L g1447 ( 
.A(n_1364),
.B(n_1365),
.Y(n_1447)
);

OR2x2_ASAP7_75t_SL g1448 ( 
.A(n_1391),
.B(n_1385),
.Y(n_1448)
);

A2O1A1Ixp33_ASAP7_75t_L g1449 ( 
.A1(n_1354),
.A2(n_1337),
.B(n_1333),
.C(n_1350),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1386),
.B(n_1391),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_SL g1451 ( 
.A1(n_1390),
.A2(n_1375),
.B1(n_1334),
.B2(n_1344),
.Y(n_1451)
);

AOI21xp33_ASAP7_75t_SL g1452 ( 
.A1(n_1405),
.A2(n_1388),
.B(n_1386),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1407),
.Y(n_1453)
);

INVx2_ASAP7_75t_SL g1454 ( 
.A(n_1444),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1395),
.Y(n_1455)
);

OA22x2_ASAP7_75t_L g1456 ( 
.A1(n_1404),
.A2(n_1334),
.B1(n_1383),
.B2(n_1384),
.Y(n_1456)
);

HB1xp67_ASAP7_75t_L g1457 ( 
.A(n_1415),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1439),
.Y(n_1458)
);

CKINVDCx14_ASAP7_75t_R g1459 ( 
.A(n_1429),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1411),
.B(n_1337),
.Y(n_1460)
);

INVx1_ASAP7_75t_SL g1461 ( 
.A(n_1396),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_SL g1462 ( 
.A(n_1393),
.B(n_1383),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1445),
.B(n_1336),
.Y(n_1463)
);

INVx1_ASAP7_75t_SL g1464 ( 
.A(n_1450),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1447),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1448),
.B(n_1449),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1428),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1428),
.Y(n_1468)
);

HB1xp67_ASAP7_75t_L g1469 ( 
.A(n_1443),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1417),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1449),
.B(n_1443),
.Y(n_1471)
);

AND2x4_ASAP7_75t_L g1472 ( 
.A(n_1417),
.B(n_1444),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1446),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1430),
.B(n_1357),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1430),
.B(n_1357),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1446),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1440),
.B(n_1361),
.Y(n_1477)
);

INVx2_ASAP7_75t_SL g1478 ( 
.A(n_1431),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1446),
.Y(n_1479)
);

AND2x4_ASAP7_75t_L g1480 ( 
.A(n_1400),
.B(n_1339),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1416),
.Y(n_1481)
);

INVxp67_ASAP7_75t_SL g1482 ( 
.A(n_1398),
.Y(n_1482)
);

NOR2xp33_ASAP7_75t_L g1483 ( 
.A(n_1425),
.B(n_1438),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1414),
.Y(n_1484)
);

AOI221xp5_ASAP7_75t_L g1485 ( 
.A1(n_1482),
.A2(n_1419),
.B1(n_1420),
.B2(n_1432),
.C(n_1441),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1464),
.B(n_1463),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1467),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1468),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1464),
.B(n_1400),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1463),
.B(n_1409),
.Y(n_1490)
);

INVx2_ASAP7_75t_SL g1491 ( 
.A(n_1454),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1455),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1483),
.A2(n_1425),
.B1(n_1413),
.B2(n_1419),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1453),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1455),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1453),
.Y(n_1496)
);

INVx4_ASAP7_75t_L g1497 ( 
.A(n_1472),
.Y(n_1497)
);

NAND2xp33_ASAP7_75t_R g1498 ( 
.A(n_1466),
.B(n_1399),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1471),
.B(n_1414),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1471),
.B(n_1414),
.Y(n_1500)
);

INVxp67_ASAP7_75t_L g1501 ( 
.A(n_1477),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1458),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1458),
.Y(n_1503)
);

BUFx2_ASAP7_75t_L g1504 ( 
.A(n_1469),
.Y(n_1504)
);

AOI221xp5_ASAP7_75t_L g1505 ( 
.A1(n_1452),
.A2(n_1420),
.B1(n_1441),
.B2(n_1394),
.C(n_1421),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1457),
.B(n_1356),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1461),
.B(n_1414),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1466),
.A2(n_1413),
.B1(n_1406),
.B2(n_1394),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1461),
.B(n_1410),
.Y(n_1509)
);

AO21x2_ASAP7_75t_L g1510 ( 
.A1(n_1481),
.A2(n_1476),
.B(n_1473),
.Y(n_1510)
);

NAND3xp33_ASAP7_75t_L g1511 ( 
.A(n_1452),
.B(n_1398),
.C(n_1408),
.Y(n_1511)
);

OAI211xp5_ASAP7_75t_L g1512 ( 
.A1(n_1474),
.A2(n_1421),
.B(n_1408),
.C(n_1427),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1472),
.B(n_1374),
.Y(n_1513)
);

OAI221xp5_ASAP7_75t_L g1514 ( 
.A1(n_1474),
.A2(n_1435),
.B1(n_1426),
.B2(n_1434),
.C(n_1438),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1460),
.B(n_1356),
.Y(n_1515)
);

NOR2xp67_ASAP7_75t_L g1516 ( 
.A(n_1478),
.B(n_1434),
.Y(n_1516)
);

NAND2x1p5_ASAP7_75t_L g1517 ( 
.A(n_1462),
.B(n_1412),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1499),
.B(n_1456),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1499),
.B(n_1456),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1501),
.B(n_1465),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1494),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1494),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1500),
.B(n_1456),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1500),
.B(n_1479),
.Y(n_1524)
);

INVx1_ASAP7_75t_SL g1525 ( 
.A(n_1504),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1507),
.B(n_1479),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1496),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1501),
.B(n_1465),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1492),
.Y(n_1529)
);

INVxp67_ASAP7_75t_SL g1530 ( 
.A(n_1506),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1492),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1496),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1492),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1502),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1510),
.B(n_1479),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1507),
.B(n_1484),
.Y(n_1536)
);

OAI21xp5_ASAP7_75t_SL g1537 ( 
.A1(n_1512),
.A2(n_1459),
.B(n_1436),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_SL g1538 ( 
.A(n_1511),
.B(n_1485),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1502),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1497),
.B(n_1504),
.Y(n_1540)
);

AND2x4_ASAP7_75t_L g1541 ( 
.A(n_1497),
.B(n_1480),
.Y(n_1541)
);

OR2x6_ASAP7_75t_L g1542 ( 
.A(n_1517),
.B(n_1480),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1510),
.B(n_1473),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1495),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1503),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1497),
.B(n_1484),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1497),
.B(n_1476),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1486),
.B(n_1470),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1495),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1487),
.B(n_1475),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1495),
.Y(n_1551)
);

OAI211xp5_ASAP7_75t_SL g1552 ( 
.A1(n_1505),
.A2(n_1392),
.B(n_1475),
.C(n_1477),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1486),
.B(n_1470),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1521),
.Y(n_1554)
);

BUFx2_ASAP7_75t_L g1555 ( 
.A(n_1542),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1538),
.A2(n_1505),
.B1(n_1485),
.B2(n_1508),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1518),
.B(n_1513),
.Y(n_1557)
);

INVx4_ASAP7_75t_L g1558 ( 
.A(n_1542),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1521),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1518),
.B(n_1513),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1550),
.B(n_1510),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1550),
.B(n_1510),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1530),
.B(n_1487),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1531),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1522),
.Y(n_1565)
);

AND2x4_ASAP7_75t_L g1566 ( 
.A(n_1541),
.B(n_1516),
.Y(n_1566)
);

NAND4xp25_ASAP7_75t_L g1567 ( 
.A(n_1538),
.B(n_1511),
.C(n_1512),
.D(n_1493),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1531),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1522),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1527),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1518),
.B(n_1491),
.Y(n_1571)
);

HB1xp67_ASAP7_75t_L g1572 ( 
.A(n_1527),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1531),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1531),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1530),
.B(n_1488),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1532),
.Y(n_1576)
);

AOI22xp5_ASAP7_75t_L g1577 ( 
.A1(n_1552),
.A2(n_1498),
.B1(n_1514),
.B2(n_1451),
.Y(n_1577)
);

INVxp67_ASAP7_75t_L g1578 ( 
.A(n_1525),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1520),
.B(n_1528),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1520),
.B(n_1488),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1519),
.B(n_1523),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1532),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1519),
.B(n_1523),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1528),
.B(n_1515),
.Y(n_1584)
);

INVx2_ASAP7_75t_SL g1585 ( 
.A(n_1540),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1519),
.B(n_1491),
.Y(n_1586)
);

INVx2_ASAP7_75t_SL g1587 ( 
.A(n_1540),
.Y(n_1587)
);

OAI22xp33_ASAP7_75t_SL g1588 ( 
.A1(n_1542),
.A2(n_1514),
.B1(n_1517),
.B2(n_1489),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1523),
.B(n_1516),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1534),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1552),
.B(n_1437),
.Y(n_1591)
);

HB1xp67_ASAP7_75t_L g1592 ( 
.A(n_1525),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1533),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1524),
.B(n_1490),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1534),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1539),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1581),
.B(n_1540),
.Y(n_1597)
);

INVxp67_ASAP7_75t_L g1598 ( 
.A(n_1592),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1556),
.B(n_1548),
.Y(n_1599)
);

OAI21xp5_ASAP7_75t_L g1600 ( 
.A1(n_1567),
.A2(n_1537),
.B(n_1517),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1572),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1572),
.Y(n_1602)
);

INVx1_ASAP7_75t_SL g1603 ( 
.A(n_1589),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1579),
.B(n_1578),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1554),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1571),
.Y(n_1606)
);

AOI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1567),
.A2(n_1537),
.B1(n_1542),
.B2(n_1541),
.Y(n_1607)
);

AND2x4_ASAP7_75t_L g1608 ( 
.A(n_1578),
.B(n_1542),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1554),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1559),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1581),
.B(n_1547),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1571),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1557),
.B(n_1548),
.Y(n_1613)
);

NAND3xp33_ASAP7_75t_L g1614 ( 
.A(n_1577),
.B(n_1543),
.C(n_1542),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1557),
.B(n_1548),
.Y(n_1615)
);

INVxp67_ASAP7_75t_SL g1616 ( 
.A(n_1588),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1583),
.B(n_1594),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1583),
.B(n_1547),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1579),
.B(n_1584),
.Y(n_1619)
);

XNOR2xp5_ASAP7_75t_L g1620 ( 
.A(n_1577),
.B(n_1436),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1584),
.B(n_1543),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1580),
.B(n_1543),
.Y(n_1622)
);

HB1xp67_ASAP7_75t_L g1623 ( 
.A(n_1585),
.Y(n_1623)
);

INVxp67_ASAP7_75t_L g1624 ( 
.A(n_1591),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1596),
.Y(n_1625)
);

NAND2xp33_ASAP7_75t_L g1626 ( 
.A(n_1585),
.B(n_1418),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1594),
.B(n_1547),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1589),
.B(n_1524),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1559),
.Y(n_1629)
);

AOI22xp33_ASAP7_75t_L g1630 ( 
.A1(n_1588),
.A2(n_1542),
.B1(n_1541),
.B2(n_1509),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1580),
.B(n_1515),
.Y(n_1631)
);

INVxp67_ASAP7_75t_L g1632 ( 
.A(n_1585),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1617),
.B(n_1587),
.Y(n_1633)
);

INVx3_ASAP7_75t_SL g1634 ( 
.A(n_1604),
.Y(n_1634)
);

AOI21xp33_ASAP7_75t_SL g1635 ( 
.A1(n_1620),
.A2(n_1587),
.B(n_1566),
.Y(n_1635)
);

AOI32xp33_ASAP7_75t_L g1636 ( 
.A1(n_1616),
.A2(n_1555),
.A3(n_1566),
.B1(n_1558),
.B2(n_1586),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1617),
.Y(n_1637)
);

NOR2xp33_ASAP7_75t_L g1638 ( 
.A(n_1624),
.B(n_1390),
.Y(n_1638)
);

NAND3xp33_ASAP7_75t_L g1639 ( 
.A(n_1614),
.B(n_1587),
.C(n_1558),
.Y(n_1639)
);

OAI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1600),
.A2(n_1555),
.B(n_1558),
.Y(n_1640)
);

OAI32xp33_ASAP7_75t_L g1641 ( 
.A1(n_1599),
.A2(n_1535),
.A3(n_1558),
.B1(n_1562),
.B2(n_1561),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1611),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1605),
.Y(n_1643)
);

NAND3xp33_ASAP7_75t_L g1644 ( 
.A(n_1598),
.B(n_1562),
.C(n_1561),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1597),
.B(n_1560),
.Y(n_1645)
);

AOI21xp33_ASAP7_75t_L g1646 ( 
.A1(n_1604),
.A2(n_1575),
.B(n_1563),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1619),
.B(n_1563),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1605),
.Y(n_1648)
);

NAND2x1_ASAP7_75t_L g1649 ( 
.A(n_1608),
.B(n_1566),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1597),
.B(n_1560),
.Y(n_1650)
);

AOI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1626),
.A2(n_1575),
.B(n_1566),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1610),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1610),
.Y(n_1653)
);

NOR2x1_ASAP7_75t_L g1654 ( 
.A(n_1626),
.B(n_1601),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1619),
.B(n_1606),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1611),
.B(n_1586),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1618),
.B(n_1541),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1629),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1655),
.Y(n_1659)
);

O2A1O1Ixp5_ASAP7_75t_L g1660 ( 
.A1(n_1641),
.A2(n_1602),
.B(n_1608),
.C(n_1612),
.Y(n_1660)
);

NOR2xp67_ASAP7_75t_L g1661 ( 
.A(n_1635),
.B(n_1607),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1655),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1637),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1637),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1643),
.Y(n_1665)
);

NAND4xp25_ASAP7_75t_L g1666 ( 
.A(n_1639),
.B(n_1630),
.C(n_1603),
.D(n_1632),
.Y(n_1666)
);

NOR2xp33_ASAP7_75t_SL g1667 ( 
.A(n_1654),
.B(n_1608),
.Y(n_1667)
);

OAI22xp33_ASAP7_75t_L g1668 ( 
.A1(n_1634),
.A2(n_1612),
.B1(n_1606),
.B2(n_1623),
.Y(n_1668)
);

OAI22xp5_ASAP7_75t_L g1669 ( 
.A1(n_1634),
.A2(n_1620),
.B1(n_1613),
.B2(n_1615),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1648),
.Y(n_1670)
);

INVx1_ASAP7_75t_SL g1671 ( 
.A(n_1633),
.Y(n_1671)
);

AOI211xp5_ASAP7_75t_L g1672 ( 
.A1(n_1640),
.A2(n_1625),
.B(n_1609),
.C(n_1618),
.Y(n_1672)
);

OAI21xp5_ASAP7_75t_SL g1673 ( 
.A1(n_1636),
.A2(n_1628),
.B(n_1627),
.Y(n_1673)
);

OAI21xp5_ASAP7_75t_SL g1674 ( 
.A1(n_1651),
.A2(n_1638),
.B(n_1646),
.Y(n_1674)
);

AOI222xp33_ASAP7_75t_L g1675 ( 
.A1(n_1644),
.A2(n_1628),
.B1(n_1627),
.B2(n_1629),
.C1(n_1526),
.C2(n_1524),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1652),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1633),
.Y(n_1677)
);

AOI211xp5_ASAP7_75t_L g1678 ( 
.A1(n_1667),
.A2(n_1661),
.B(n_1668),
.C(n_1674),
.Y(n_1678)
);

AOI32xp33_ASAP7_75t_L g1679 ( 
.A1(n_1669),
.A2(n_1668),
.A3(n_1672),
.B1(n_1671),
.B2(n_1677),
.Y(n_1679)
);

OAI22xp33_ASAP7_75t_SL g1680 ( 
.A1(n_1659),
.A2(n_1649),
.B1(n_1653),
.B2(n_1658),
.Y(n_1680)
);

AOI21xp33_ASAP7_75t_SL g1681 ( 
.A1(n_1662),
.A2(n_1638),
.B(n_1677),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1663),
.B(n_1656),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1664),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1665),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1673),
.B(n_1656),
.Y(n_1685)
);

INVxp67_ASAP7_75t_L g1686 ( 
.A(n_1666),
.Y(n_1686)
);

XOR2xp5_ASAP7_75t_L g1687 ( 
.A(n_1670),
.B(n_1423),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1676),
.Y(n_1688)
);

AOI211xp5_ASAP7_75t_L g1689 ( 
.A1(n_1680),
.A2(n_1647),
.B(n_1660),
.C(n_1642),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1682),
.Y(n_1690)
);

AOI221xp5_ASAP7_75t_L g1691 ( 
.A1(n_1679),
.A2(n_1686),
.B1(n_1678),
.B2(n_1680),
.C(n_1660),
.Y(n_1691)
);

O2A1O1Ixp33_ASAP7_75t_SL g1692 ( 
.A1(n_1685),
.A2(n_1647),
.B(n_1642),
.C(n_1650),
.Y(n_1692)
);

NOR3xp33_ASAP7_75t_SL g1693 ( 
.A(n_1684),
.B(n_1422),
.C(n_1675),
.Y(n_1693)
);

NOR3x1_ASAP7_75t_L g1694 ( 
.A(n_1688),
.B(n_1621),
.C(n_1622),
.Y(n_1694)
);

NAND4xp25_ASAP7_75t_L g1695 ( 
.A(n_1681),
.B(n_1683),
.C(n_1645),
.D(n_1657),
.Y(n_1695)
);

NOR2xp33_ASAP7_75t_L g1696 ( 
.A(n_1687),
.B(n_1645),
.Y(n_1696)
);

NAND3xp33_ASAP7_75t_L g1697 ( 
.A(n_1678),
.B(n_1622),
.C(n_1621),
.Y(n_1697)
);

NAND4xp25_ASAP7_75t_L g1698 ( 
.A(n_1678),
.B(n_1657),
.C(n_1390),
.D(n_1433),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1682),
.B(n_1541),
.Y(n_1699)
);

AOI221xp5_ASAP7_75t_L g1700 ( 
.A1(n_1691),
.A2(n_1564),
.B1(n_1568),
.B2(n_1573),
.C(n_1593),
.Y(n_1700)
);

A2O1A1Ixp33_ASAP7_75t_L g1701 ( 
.A1(n_1689),
.A2(n_1535),
.B(n_1631),
.C(n_1595),
.Y(n_1701)
);

AOI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1692),
.A2(n_1535),
.B(n_1565),
.Y(n_1702)
);

NAND4xp25_ASAP7_75t_L g1703 ( 
.A(n_1698),
.B(n_1402),
.C(n_1403),
.D(n_1424),
.Y(n_1703)
);

NAND4xp75_ASAP7_75t_L g1704 ( 
.A(n_1694),
.B(n_1690),
.C(n_1693),
.D(n_1696),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1695),
.B(n_1631),
.Y(n_1705)
);

AOI221x1_ASAP7_75t_L g1706 ( 
.A1(n_1701),
.A2(n_1697),
.B1(n_1699),
.B2(n_1565),
.C(n_1576),
.Y(n_1706)
);

OAI321xp33_ASAP7_75t_L g1707 ( 
.A1(n_1705),
.A2(n_1397),
.A3(n_1442),
.B1(n_1574),
.B2(n_1573),
.C(n_1568),
.Y(n_1707)
);

O2A1O1Ixp33_ASAP7_75t_L g1708 ( 
.A1(n_1700),
.A2(n_1596),
.B(n_1595),
.C(n_1569),
.Y(n_1708)
);

AOI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1704),
.A2(n_1403),
.B1(n_1397),
.B2(n_1582),
.Y(n_1709)
);

NOR2xp67_ASAP7_75t_L g1710 ( 
.A(n_1702),
.B(n_1569),
.Y(n_1710)
);

AOI21xp33_ASAP7_75t_SL g1711 ( 
.A1(n_1703),
.A2(n_1576),
.B(n_1570),
.Y(n_1711)
);

NOR3xp33_ASAP7_75t_L g1712 ( 
.A(n_1707),
.B(n_1568),
.C(n_1564),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1710),
.Y(n_1713)
);

AOI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1709),
.A2(n_1397),
.B1(n_1590),
.B2(n_1582),
.Y(n_1714)
);

AND3x4_ASAP7_75t_L g1715 ( 
.A(n_1706),
.B(n_1573),
.C(n_1564),
.Y(n_1715)
);

AOI22xp5_ASAP7_75t_L g1716 ( 
.A1(n_1711),
.A2(n_1590),
.B1(n_1570),
.B2(n_1526),
.Y(n_1716)
);

OAI31xp33_ASAP7_75t_L g1717 ( 
.A1(n_1713),
.A2(n_1708),
.A3(n_1593),
.B(n_1574),
.Y(n_1717)
);

NAND4xp75_ASAP7_75t_L g1718 ( 
.A(n_1714),
.B(n_1593),
.C(n_1574),
.D(n_1526),
.Y(n_1718)
);

AND2x4_ASAP7_75t_L g1719 ( 
.A(n_1716),
.B(n_1509),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1719),
.Y(n_1720)
);

OA22x2_ASAP7_75t_L g1721 ( 
.A1(n_1720),
.A2(n_1715),
.B1(n_1717),
.B2(n_1718),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1721),
.B(n_1712),
.Y(n_1722)
);

INVxp67_ASAP7_75t_L g1723 ( 
.A(n_1721),
.Y(n_1723)
);

AOI22x1_ASAP7_75t_L g1724 ( 
.A1(n_1722),
.A2(n_1544),
.B1(n_1551),
.B2(n_1549),
.Y(n_1724)
);

AOI22xp5_ASAP7_75t_L g1725 ( 
.A1(n_1723),
.A2(n_1546),
.B1(n_1536),
.B2(n_1553),
.Y(n_1725)
);

AO21x2_ASAP7_75t_L g1726 ( 
.A1(n_1725),
.A2(n_1551),
.B(n_1549),
.Y(n_1726)
);

OAI21xp5_ASAP7_75t_L g1727 ( 
.A1(n_1724),
.A2(n_1536),
.B(n_1546),
.Y(n_1727)
);

XNOR2x1_ASAP7_75t_L g1728 ( 
.A(n_1727),
.B(n_1401),
.Y(n_1728)
);

OR2x6_ASAP7_75t_L g1729 ( 
.A(n_1728),
.B(n_1726),
.Y(n_1729)
);

XNOR2xp5_ASAP7_75t_L g1730 ( 
.A(n_1729),
.B(n_1401),
.Y(n_1730)
);

OAI221xp5_ASAP7_75t_R g1731 ( 
.A1(n_1730),
.A2(n_1536),
.B1(n_1546),
.B2(n_1549),
.C(n_1551),
.Y(n_1731)
);

AOI211xp5_ASAP7_75t_L g1732 ( 
.A1(n_1731),
.A2(n_1367),
.B(n_1529),
.C(n_1545),
.Y(n_1732)
);


endmodule