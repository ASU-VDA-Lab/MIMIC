module fake_ariane_2016_n_111 (n_8, n_7, n_1, n_6, n_13, n_17, n_4, n_2, n_18, n_9, n_11, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_10, n_111);

input n_8;
input n_7;
input n_1;
input n_6;
input n_13;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_10;

output n_111;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_90;
wire n_38;
wire n_47;
wire n_110;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_34;
wire n_69;
wire n_95;
wire n_92;
wire n_98;
wire n_74;
wire n_33;
wire n_40;
wire n_106;
wire n_53;
wire n_21;
wire n_66;
wire n_71;
wire n_24;
wire n_109;
wire n_96;
wire n_49;
wire n_20;
wire n_100;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_103;
wire n_79;
wire n_26;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_107;
wire n_72;
wire n_105;
wire n_44;
wire n_30;
wire n_82;
wire n_31;
wire n_42;
wire n_57;
wire n_70;
wire n_85;
wire n_48;
wire n_94;
wire n_101;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_93;
wire n_23;
wire n_61;
wire n_108;
wire n_102;
wire n_22;
wire n_81;
wire n_87;
wire n_43;
wire n_27;
wire n_29;
wire n_41;
wire n_55;
wire n_28;
wire n_80;
wire n_97;
wire n_88;
wire n_68;
wire n_104;
wire n_78;
wire n_39;
wire n_63;
wire n_59;
wire n_99;
wire n_35;
wire n_54;
wire n_25;

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

NOR2xp67_ASAP7_75t_L g27 ( 
.A(n_13),
.B(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx5p33_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx5p33_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

NOR2xp67_ASAP7_75t_L g38 ( 
.A(n_20),
.B(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_35),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_R g41 ( 
.A(n_34),
.B(n_11),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_30),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_31),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

CKINVDCx5p33_ASAP7_75t_R g46 ( 
.A(n_35),
.Y(n_46)
);

AOI21x1_ASAP7_75t_L g47 ( 
.A1(n_25),
.A2(n_1),
.B(n_2),
.Y(n_47)
);

CKINVDCx5p33_ASAP7_75t_R g48 ( 
.A(n_28),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_29),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_29),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_36),
.A2(n_24),
.B1(n_22),
.B2(n_33),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_45),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_44),
.Y(n_59)
);

OAI21xp33_ASAP7_75t_SL g60 ( 
.A1(n_50),
.A2(n_40),
.B(n_38),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_40),
.B(n_45),
.C(n_38),
.Y(n_61)
);

AO21x1_ASAP7_75t_L g62 ( 
.A1(n_54),
.A2(n_28),
.B(n_47),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

BUFx8_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

BUFx8_ASAP7_75t_SL g65 ( 
.A(n_58),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_52),
.Y(n_66)
);

NOR2xp67_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_57),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_62),
.A2(n_55),
.B1(n_57),
.B2(n_53),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_69),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

AO21x2_ASAP7_75t_L g75 ( 
.A1(n_70),
.A2(n_73),
.B(n_61),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_69),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_68),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_71),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_77),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_77),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_78),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_82),
.B(n_68),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_68),
.Y(n_89)
);

AOI221xp5_ASAP7_75t_L g90 ( 
.A1(n_83),
.A2(n_24),
.B1(n_22),
.B2(n_33),
.C(n_42),
.Y(n_90)
);

NAND3xp33_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_27),
.C(n_53),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_88),
.A2(n_75),
.B(n_51),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_89),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_90),
.A2(n_47),
.B(n_85),
.Y(n_94)
);

NOR2x1p5_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_84),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_85),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_87),
.Y(n_97)
);

AOI211xp5_ASAP7_75t_L g98 ( 
.A1(n_94),
.A2(n_21),
.B(n_41),
.C(n_74),
.Y(n_98)
);

AOI221xp5_ASAP7_75t_L g99 ( 
.A1(n_93),
.A2(n_97),
.B1(n_96),
.B2(n_21),
.C(n_43),
.Y(n_99)
);

OAI211xp5_ASAP7_75t_L g100 ( 
.A1(n_95),
.A2(n_74),
.B(n_3),
.C(n_5),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_93),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_75),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_100),
.B(n_75),
.Y(n_103)
);

OAI221xp5_ASAP7_75t_L g104 ( 
.A1(n_99),
.A2(n_98),
.B1(n_74),
.B2(n_6),
.C(n_8),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_R g105 ( 
.A(n_103),
.B(n_74),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_102),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_106),
.Y(n_107)
);

OAI22x1_ASAP7_75t_L g108 ( 
.A1(n_107),
.A2(n_74),
.B1(n_105),
.B2(n_104),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_108),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_109),
.A2(n_74),
.B1(n_64),
.B2(n_8),
.Y(n_110)
);

AOI221xp5_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_1),
.B1(n_3),
.B2(n_9),
.C(n_64),
.Y(n_111)
);


endmodule