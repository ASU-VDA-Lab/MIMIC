module fake_jpeg_2590_n_714 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_714);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_714;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_696;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_699;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_543;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_713;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_701;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_704;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_698;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_694;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_697;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_710;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_709;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_708;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_703;
wire n_439;
wire n_262;
wire n_398;
wire n_240;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_695;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_702;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_707;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_705;
wire n_665;
wire n_706;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_700;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_712;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_711;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_19),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_1),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_8),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_5),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_9),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_15),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_16),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_61),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_62),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_63),
.Y(n_144)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

BUFx4f_ASAP7_75t_SL g160 ( 
.A(n_64),
.Y(n_160)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_65),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_66),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_67),
.Y(n_174)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_68),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_69),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_70),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_71),
.Y(n_140)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_24),
.B(n_9),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_72),
.B(n_37),
.C(n_40),
.Y(n_207)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx2_ASAP7_75t_SL g159 ( 
.A(n_73),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx6_ASAP7_75t_L g213 ( 
.A(n_74),
.Y(n_213)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g220 ( 
.A(n_75),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_41),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_76),
.B(n_79),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_77),
.Y(n_188)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_78),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_28),
.B(n_9),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_28),
.B(n_8),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_80),
.B(n_97),
.Y(n_135)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_81),
.Y(n_154)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_82),
.Y(n_137)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_24),
.Y(n_83)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_83),
.Y(n_143)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_84),
.Y(n_189)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_85),
.Y(n_192)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_86),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_87),
.Y(n_197)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_88),
.Y(n_212)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_89),
.Y(n_158)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_90),
.Y(n_227)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_91),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_92),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_93),
.Y(n_162)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_45),
.Y(n_94)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_94),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_95),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g183 ( 
.A(n_96),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_29),
.B(n_8),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_29),
.B(n_59),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_98),
.B(n_107),
.Y(n_142)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_99),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_34),
.B(n_11),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_100),
.B(n_110),
.Y(n_168)
);

INVx4_ASAP7_75t_SL g101 ( 
.A(n_55),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_101),
.B(n_120),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_102),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_103),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_35),
.Y(n_104)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_104),
.Y(n_202)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_105),
.Y(n_173)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_23),
.Y(n_106)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_106),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_57),
.B(n_11),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_56),
.B(n_11),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_108),
.B(n_111),
.Y(n_155)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_51),
.Y(n_109)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_109),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_34),
.B(n_18),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_57),
.B(n_18),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_35),
.Y(n_112)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_112),
.Y(n_221)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_49),
.Y(n_113)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_113),
.Y(n_222)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_22),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_114),
.Y(n_182)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_25),
.Y(n_115)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_115),
.Y(n_232)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_51),
.Y(n_116)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_116),
.Y(n_179)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_49),
.Y(n_117)
);

INVx6_ASAP7_75t_SL g211 ( 
.A(n_117),
.Y(n_211)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_39),
.Y(n_118)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_118),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_34),
.B(n_18),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_119),
.B(n_55),
.Y(n_170)
);

BUFx24_ASAP7_75t_L g120 ( 
.A(n_25),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_49),
.Y(n_121)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_121),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_56),
.B(n_17),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_122),
.B(n_14),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_49),
.Y(n_123)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_123),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_53),
.Y(n_124)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_124),
.Y(n_194)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_22),
.Y(n_125)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_125),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_53),
.Y(n_126)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_126),
.Y(n_204)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_51),
.Y(n_127)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_127),
.Y(n_208)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_22),
.Y(n_128)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_128),
.Y(n_214)
);

BUFx12f_ASAP7_75t_L g129 ( 
.A(n_53),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_129),
.B(n_133),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_53),
.Y(n_130)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_130),
.Y(n_224)
);

BUFx5_ASAP7_75t_L g131 ( 
.A(n_25),
.Y(n_131)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_131),
.Y(n_230)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_39),
.Y(n_132)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_132),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_21),
.Y(n_133)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_25),
.Y(n_134)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_101),
.A2(n_42),
.B1(n_60),
.B2(n_48),
.Y(n_136)
);

OA22x2_ASAP7_75t_L g314 ( 
.A1(n_136),
.A2(n_152),
.B1(n_185),
.B2(n_187),
.Y(n_314)
);

NAND2x1_ASAP7_75t_L g145 ( 
.A(n_100),
.B(n_31),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_145),
.B(n_170),
.Y(n_270)
);

A2O1A1Ixp33_ASAP7_75t_L g146 ( 
.A1(n_72),
.A2(n_59),
.B(n_60),
.C(n_50),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_146),
.B(n_209),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_110),
.B(n_119),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_147),
.B(n_161),
.Y(n_273)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_104),
.A2(n_112),
.B1(n_121),
.B2(n_130),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_150),
.A2(n_206),
.B1(n_231),
.B2(n_0),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_134),
.A2(n_42),
.B1(n_60),
.B2(n_48),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_123),
.Y(n_161)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_164),
.Y(n_238)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_118),
.Y(n_165)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_165),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_62),
.A2(n_27),
.B1(n_47),
.B2(n_46),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_167),
.A2(n_171),
.B1(n_190),
.B2(n_205),
.Y(n_236)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_84),
.Y(n_169)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_169),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_63),
.A2(n_27),
.B1(n_31),
.B2(n_40),
.Y(n_171)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_91),
.Y(n_176)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_176),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_68),
.A2(n_42),
.B1(n_37),
.B2(n_50),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_71),
.B(n_27),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_186),
.B(n_193),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_61),
.A2(n_42),
.B1(n_21),
.B2(n_40),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_65),
.A2(n_93),
.B1(n_89),
.B2(n_120),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_124),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_65),
.B(n_21),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_196),
.B(n_198),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_89),
.B(n_31),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_199),
.B(n_217),
.Y(n_246)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_113),
.Y(n_203)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_203),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_126),
.A2(n_66),
.B1(n_67),
.B2(n_103),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_85),
.A2(n_37),
.B1(n_50),
.B2(n_48),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_207),
.B(n_0),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_64),
.B(n_47),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_69),
.B(n_47),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_70),
.A2(n_44),
.B1(n_46),
.B2(n_36),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_218),
.A2(n_219),
.B1(n_120),
.B2(n_32),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_93),
.A2(n_44),
.B1(n_46),
.B2(n_52),
.Y(n_219)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_74),
.Y(n_225)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_225),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_77),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_226),
.B(n_16),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_87),
.B(n_44),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_229),
.B(n_20),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_92),
.A2(n_52),
.B1(n_36),
.B2(n_32),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_146),
.B(n_52),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_233),
.B(n_301),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_215),
.A2(n_20),
.B1(n_32),
.B2(n_36),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_234),
.Y(n_330)
);

OAI22xp33_ASAP7_75t_L g235 ( 
.A1(n_136),
.A2(n_95),
.B1(n_96),
.B2(n_102),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_235),
.A2(n_245),
.B1(n_260),
.B2(n_293),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_139),
.Y(n_237)
);

INVx6_ASAP7_75t_L g325 ( 
.A(n_237),
.Y(n_325)
);

AND2x2_ASAP7_75t_SL g239 ( 
.A(n_137),
.B(n_129),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_239),
.Y(n_329)
);

INVx2_ASAP7_75t_SL g241 ( 
.A(n_228),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_241),
.Y(n_374)
);

BUFx8_ASAP7_75t_L g243 ( 
.A(n_211),
.Y(n_243)
);

INVx4_ASAP7_75t_SL g339 ( 
.A(n_243),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_205),
.A2(n_155),
.B1(n_218),
.B2(n_168),
.Y(n_245)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_138),
.Y(n_247)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_247),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_159),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_248),
.Y(n_357)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_138),
.Y(n_249)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_249),
.Y(n_366)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_140),
.Y(n_250)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_250),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_228),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_252),
.B(n_272),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_253),
.A2(n_275),
.B1(n_302),
.B2(n_304),
.Y(n_322)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_210),
.Y(n_254)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_254),
.Y(n_369)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_182),
.Y(n_258)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_258),
.Y(n_371)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_141),
.Y(n_259)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_259),
.Y(n_321)
);

OAI22xp33_ASAP7_75t_L g260 ( 
.A1(n_152),
.A2(n_20),
.B1(n_117),
.B2(n_129),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_261),
.B(n_274),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_135),
.B(n_12),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_262),
.B(n_266),
.Y(n_360)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_181),
.Y(n_263)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_263),
.Y(n_373)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_210),
.Y(n_264)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_264),
.Y(n_328)
);

BUFx4f_ASAP7_75t_SL g265 ( 
.A(n_160),
.Y(n_265)
);

INVx13_ASAP7_75t_L g363 ( 
.A(n_265),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_142),
.B(n_12),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_153),
.Y(n_267)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_267),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_230),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_268),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_140),
.Y(n_269)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_269),
.Y(n_347)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_191),
.Y(n_271)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_271),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_160),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_215),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_159),
.A2(n_117),
.B1(n_33),
.B2(n_54),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_194),
.Y(n_276)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_276),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_277),
.Y(n_323)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_151),
.Y(n_278)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_278),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_166),
.B(n_145),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_279),
.B(n_297),
.Y(n_364)
);

INVx5_ASAP7_75t_L g280 ( 
.A(n_189),
.Y(n_280)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_280),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_143),
.B(n_33),
.C(n_54),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_281),
.B(n_294),
.C(n_172),
.Y(n_349)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_157),
.Y(n_282)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_282),
.Y(n_370)
);

OAI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_185),
.A2(n_54),
.B1(n_33),
.B2(n_16),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_283),
.A2(n_315),
.B1(n_241),
.B2(n_243),
.Y(n_331)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_220),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_284),
.B(n_288),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_285),
.B(n_286),
.Y(n_336)
);

INVx2_ASAP7_75t_SL g287 ( 
.A(n_220),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g318 ( 
.A(n_287),
.B(n_303),
.Y(n_318)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_173),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_192),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_289),
.B(n_290),
.Y(n_337)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_204),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g291 ( 
.A1(n_150),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_SL g353 ( 
.A1(n_291),
.A2(n_300),
.B1(n_216),
.B2(n_163),
.Y(n_353)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_222),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_292),
.B(n_295),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_224),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_195),
.B(n_1),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_178),
.Y(n_295)
);

INVx6_ASAP7_75t_L g296 ( 
.A(n_139),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_296),
.B(n_298),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_179),
.B(n_15),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_208),
.B(n_15),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_L g300 ( 
.A1(n_223),
.A2(n_14),
.B1(n_13),
.B2(n_12),
.Y(n_300)
);

INVx6_ASAP7_75t_L g301 ( 
.A(n_144),
.Y(n_301)
);

INVx5_ASAP7_75t_L g302 ( 
.A(n_189),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_214),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_177),
.A2(n_12),
.B1(n_2),
.B2(n_3),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_201),
.Y(n_305)
);

OR2x2_ASAP7_75t_L g338 ( 
.A(n_305),
.B(n_310),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_223),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_306),
.A2(n_221),
.B1(n_172),
.B2(n_188),
.Y(n_342)
);

AO22x2_ASAP7_75t_L g307 ( 
.A1(n_202),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_307)
);

NOR2x1_ASAP7_75t_L g378 ( 
.A(n_307),
.B(n_317),
.Y(n_378)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_158),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_308),
.A2(n_309),
.B1(n_312),
.B2(n_313),
.Y(n_324)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_202),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_180),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_192),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_311),
.B(n_156),
.Y(n_333)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_200),
.Y(n_312)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_158),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g315 ( 
.A(n_160),
.Y(n_315)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_222),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g341 ( 
.A1(n_316),
.A2(n_148),
.B1(n_162),
.B2(n_183),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_212),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_317)
);

INVxp67_ASAP7_75t_SL g413 ( 
.A(n_331),
.Y(n_413)
);

INVx1_ASAP7_75t_SL g406 ( 
.A(n_333),
.Y(n_406)
);

MAJx2_ASAP7_75t_L g334 ( 
.A(n_270),
.B(n_232),
.C(n_227),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_334),
.B(n_365),
.C(n_313),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_341),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_342),
.A2(n_350),
.B1(n_351),
.B2(n_301),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_286),
.A2(n_190),
.B1(n_219),
.B2(n_213),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_343),
.A2(n_352),
.B1(n_380),
.B2(n_293),
.Y(n_393)
);

AOI22xp33_ASAP7_75t_SL g344 ( 
.A1(n_236),
.A2(n_200),
.B1(n_162),
.B2(n_148),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_SL g391 ( 
.A1(n_344),
.A2(n_243),
.B1(n_260),
.B2(n_306),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_257),
.A2(n_154),
.B(n_221),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_345),
.A2(n_379),
.B(n_331),
.Y(n_432)
);

OAI21xp33_ASAP7_75t_L g423 ( 
.A1(n_349),
.A2(n_265),
.B(n_308),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_245),
.A2(n_174),
.B1(n_144),
.B2(n_149),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_235),
.A2(n_149),
.B1(n_174),
.B2(n_188),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_233),
.A2(n_175),
.B1(n_213),
.B2(n_184),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_L g392 ( 
.A1(n_353),
.A2(n_265),
.B1(n_307),
.B2(n_239),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_246),
.B(n_197),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_354),
.B(n_356),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_242),
.B(n_197),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_285),
.B(n_299),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_358),
.B(n_372),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_270),
.B(n_184),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_285),
.B(n_175),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_L g375 ( 
.A1(n_274),
.A2(n_256),
.B1(n_314),
.B2(n_287),
.Y(n_375)
);

OAI22xp33_ASAP7_75t_SL g420 ( 
.A1(n_375),
.A2(n_258),
.B1(n_247),
.B2(n_268),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_294),
.B(n_163),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_376),
.B(n_377),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_294),
.B(n_216),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_270),
.A2(n_154),
.B1(n_183),
.B2(n_7),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_314),
.A2(n_183),
.B1(n_5),
.B2(n_6),
.Y(n_380)
);

FAx1_ASAP7_75t_SL g381 ( 
.A(n_273),
.B(n_5),
.CI(n_281),
.CON(n_381),
.SN(n_381)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_381),
.B(n_314),
.Y(n_383)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_371),
.Y(n_382)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_382),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_383),
.B(n_388),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_320),
.B(n_239),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_384),
.B(n_329),
.C(n_334),
.Y(n_444)
);

INVx4_ASAP7_75t_SL g385 ( 
.A(n_318),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g451 ( 
.A(n_385),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_386),
.B(n_400),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_330),
.A2(n_314),
.B(n_317),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_387),
.A2(n_408),
.B(n_432),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_326),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_371),
.Y(n_389)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_389),
.Y(n_449)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_362),
.Y(n_390)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_390),
.Y(n_441)
);

OAI22xp33_ASAP7_75t_SL g452 ( 
.A1(n_391),
.A2(n_392),
.B1(n_415),
.B2(n_379),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_393),
.A2(n_407),
.B1(n_416),
.B2(n_351),
.Y(n_433)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_362),
.Y(n_394)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_394),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_336),
.A2(n_307),
.B1(n_292),
.B2(n_316),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_396),
.A2(n_398),
.B1(n_403),
.B2(n_418),
.Y(n_455)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_370),
.Y(n_397)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_397),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_336),
.A2(n_307),
.B1(n_276),
.B2(n_271),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_321),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_399),
.B(n_402),
.Y(n_460)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_370),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_323),
.B(n_238),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_401),
.B(n_405),
.Y(n_446)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_340),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_336),
.A2(n_290),
.B1(n_263),
.B2(n_295),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g404 ( 
.A(n_318),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_404),
.B(n_409),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_323),
.B(n_240),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_335),
.A2(n_296),
.B1(n_237),
.B2(n_302),
.Y(n_407)
);

AND2x4_ASAP7_75t_L g408 ( 
.A(n_380),
.B(n_264),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_321),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_338),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_410),
.B(n_411),
.Y(n_447)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_325),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_325),
.Y(n_412)
);

INVx6_ASAP7_75t_L g462 ( 
.A(n_412),
.Y(n_462)
);

CKINVDCx14_ASAP7_75t_R g414 ( 
.A(n_332),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_414),
.Y(n_439)
);

AOI22xp33_ASAP7_75t_SL g415 ( 
.A1(n_343),
.A2(n_269),
.B1(n_280),
.B2(n_250),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_335),
.A2(n_309),
.B1(n_305),
.B2(n_244),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_327),
.A2(n_255),
.B1(n_251),
.B2(n_254),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_420),
.A2(n_374),
.B1(n_386),
.B2(n_404),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_422),
.B(n_423),
.Y(n_436)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_373),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_424),
.B(n_425),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_338),
.Y(n_425)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_348),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_426),
.Y(n_461)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_355),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_427),
.B(n_428),
.Y(n_465)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_355),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_356),
.B(n_249),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_429),
.B(n_430),
.Y(n_472)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_361),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_327),
.A2(n_5),
.B1(n_350),
.B2(n_352),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_431),
.A2(n_342),
.B1(n_346),
.B2(n_361),
.Y(n_459)
);

OAI22xp33_ASAP7_75t_SL g480 ( 
.A1(n_433),
.A2(n_456),
.B1(n_398),
.B2(n_406),
.Y(n_480)
);

A2O1A1O1Ixp25_ASAP7_75t_L g435 ( 
.A1(n_422),
.A2(n_378),
.B(n_320),
.C(n_349),
.D(n_354),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_435),
.A2(n_445),
.B(n_467),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_417),
.B(n_320),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_SL g476 ( 
.A(n_440),
.B(n_448),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_393),
.A2(n_322),
.B1(n_378),
.B2(n_329),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_442),
.A2(n_459),
.B1(n_466),
.B2(n_408),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_417),
.B(n_395),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_443),
.B(n_444),
.C(n_454),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_432),
.A2(n_330),
.B(n_345),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_395),
.B(n_358),
.Y(n_448)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_429),
.Y(n_450)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_450),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_452),
.B(n_469),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_SL g453 ( 
.A1(n_383),
.A2(n_378),
.B(n_381),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_453),
.A2(n_471),
.B(n_419),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_384),
.B(n_365),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_419),
.B(n_372),
.C(n_333),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_458),
.B(n_385),
.C(n_418),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_405),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_463),
.B(n_473),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_396),
.A2(n_359),
.B1(n_374),
.B2(n_381),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_L g467 ( 
.A1(n_387),
.A2(n_318),
.B(n_338),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_413),
.A2(n_364),
.B1(n_376),
.B2(n_377),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g471 ( 
.A1(n_410),
.A2(n_337),
.B(n_364),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_401),
.Y(n_473)
);

A2O1A1Ixp33_ASAP7_75t_L g475 ( 
.A1(n_425),
.A2(n_360),
.B(n_346),
.C(n_357),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_475),
.B(n_388),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_SL g477 ( 
.A(n_443),
.B(n_406),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_SL g549 ( 
.A(n_477),
.B(n_482),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_465),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_478),
.B(n_488),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_480),
.A2(n_491),
.B1(n_513),
.B2(n_459),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_SL g521 ( 
.A(n_481),
.B(n_499),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_SL g482 ( 
.A(n_448),
.B(n_402),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_483),
.A2(n_484),
.B1(n_486),
.B2(n_497),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_442),
.A2(n_408),
.B1(n_407),
.B2(n_416),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_464),
.A2(n_408),
.B1(n_466),
.B2(n_455),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_460),
.B(n_385),
.Y(n_487)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_487),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_465),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_489),
.B(n_436),
.Y(n_527)
);

CKINVDCx14_ASAP7_75t_R g552 ( 
.A(n_490),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_433),
.A2(n_431),
.B1(n_408),
.B2(n_403),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g492 ( 
.A1(n_437),
.A2(n_421),
.B(n_390),
.Y(n_492)
);

OAI21xp5_ASAP7_75t_SL g543 ( 
.A1(n_492),
.A2(n_472),
.B(n_471),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_457),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_495),
.B(n_498),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_SL g496 ( 
.A(n_439),
.B(n_360),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_496),
.B(n_503),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_464),
.A2(n_409),
.B1(n_399),
.B2(n_397),
.Y(n_497)
);

OA22x2_ASAP7_75t_L g498 ( 
.A1(n_456),
.A2(n_400),
.B1(n_394),
.B2(n_428),
.Y(n_498)
);

INVxp33_ASAP7_75t_L g500 ( 
.A(n_446),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_500),
.B(n_463),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_SL g501 ( 
.A(n_454),
.B(n_430),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_501),
.B(n_444),
.Y(n_519)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_474),
.Y(n_502)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_502),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_439),
.B(n_473),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_464),
.A2(n_427),
.B1(n_411),
.B2(n_412),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_504),
.A2(n_506),
.B1(n_461),
.B2(n_468),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_436),
.B(n_347),
.C(n_368),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_505),
.B(n_467),
.C(n_468),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_455),
.A2(n_412),
.B1(n_426),
.B2(n_389),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_457),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_507),
.B(n_510),
.Y(n_555)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_474),
.Y(n_508)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_508),
.Y(n_551)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_460),
.Y(n_509)
);

INVx2_ASAP7_75t_SL g517 ( 
.A(n_509),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_447),
.Y(n_510)
);

INVx4_ASAP7_75t_L g511 ( 
.A(n_462),
.Y(n_511)
);

INVx3_ASAP7_75t_L g536 ( 
.A(n_511),
.Y(n_536)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_441),
.Y(n_512)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_512),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_438),
.A2(n_324),
.B1(n_368),
.B2(n_382),
.Y(n_513)
);

XOR2x2_ASAP7_75t_L g514 ( 
.A(n_440),
.B(n_328),
.Y(n_514)
);

NOR2x1_ASAP7_75t_L g531 ( 
.A(n_514),
.B(n_458),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_446),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_515),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_483),
.A2(n_438),
.B1(n_450),
.B2(n_447),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_516),
.A2(n_550),
.B1(n_493),
.B2(n_478),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g584 ( 
.A1(n_518),
.A2(n_530),
.B1(n_532),
.B2(n_533),
.Y(n_584)
);

XOR2xp5_ASAP7_75t_L g560 ( 
.A(n_519),
.B(n_539),
.Y(n_560)
);

XNOR2x1_ASAP7_75t_L g571 ( 
.A(n_521),
.B(n_531),
.Y(n_571)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_503),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_523),
.B(n_524),
.Y(n_574)
);

CKINVDCx16_ASAP7_75t_R g524 ( 
.A(n_487),
.Y(n_524)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_525),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_499),
.A2(n_437),
.B(n_445),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_L g588 ( 
.A1(n_526),
.A2(n_537),
.B(n_543),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_527),
.B(n_528),
.C(n_535),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_491),
.A2(n_451),
.B1(n_475),
.B2(n_470),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_486),
.A2(n_451),
.B1(n_470),
.B2(n_472),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_485),
.B(n_453),
.C(n_435),
.Y(n_535)
);

OAI21xp5_ASAP7_75t_L g537 ( 
.A1(n_510),
.A2(n_453),
.B(n_435),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_485),
.B(n_469),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_494),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_540),
.B(n_546),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_496),
.B(n_494),
.Y(n_542)
);

CKINVDCx14_ASAP7_75t_R g568 ( 
.A(n_542),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_501),
.B(n_441),
.C(n_347),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_545),
.B(n_554),
.C(n_514),
.Y(n_564)
);

CKINVDCx16_ASAP7_75t_R g546 ( 
.A(n_497),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_482),
.B(n_357),
.Y(n_548)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_548),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_SL g550 ( 
.A1(n_484),
.A2(n_461),
.B1(n_462),
.B2(n_449),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_477),
.B(n_476),
.Y(n_553)
);

XOR2xp5_ASAP7_75t_L g561 ( 
.A(n_553),
.B(n_476),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_505),
.B(n_328),
.C(n_366),
.Y(n_554)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_555),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_556),
.B(n_557),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_555),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_520),
.Y(n_558)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_558),
.Y(n_607)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_528),
.B(n_481),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g593 ( 
.A(n_559),
.B(n_564),
.Y(n_593)
);

MAJx2_ASAP7_75t_L g596 ( 
.A(n_561),
.B(n_577),
.C(n_549),
.Y(n_596)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_563),
.Y(n_597)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_527),
.B(n_489),
.C(n_514),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_565),
.B(n_572),
.C(n_575),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_L g566 ( 
.A1(n_529),
.A2(n_507),
.B1(n_495),
.B2(n_479),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_566),
.A2(n_578),
.B1(n_581),
.B2(n_582),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_520),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_567),
.B(n_586),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_SL g570 ( 
.A1(n_516),
.A2(n_479),
.B1(n_513),
.B2(n_509),
.Y(n_570)
);

XOR2xp5_ASAP7_75t_L g598 ( 
.A(n_570),
.B(n_534),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_539),
.B(n_535),
.C(n_554),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_517),
.Y(n_573)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_573),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_519),
.B(n_493),
.C(n_488),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_545),
.B(n_492),
.C(n_479),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_576),
.B(n_580),
.C(n_541),
.Y(n_613)
);

XOR2xp5_ASAP7_75t_L g577 ( 
.A(n_553),
.B(n_498),
.Y(n_577)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_518),
.A2(n_506),
.B1(n_498),
.B2(n_504),
.Y(n_578)
);

FAx1_ASAP7_75t_SL g579 ( 
.A(n_537),
.B(n_498),
.CI(n_512),
.CON(n_579),
.SN(n_579)
);

FAx1_ASAP7_75t_SL g591 ( 
.A(n_579),
.B(n_526),
.CI(n_543),
.CON(n_591),
.SN(n_591)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_521),
.B(n_502),
.C(n_508),
.Y(n_580)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_552),
.A2(n_511),
.B1(n_449),
.B2(n_434),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_550),
.A2(n_434),
.B1(n_424),
.B2(n_462),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_517),
.Y(n_583)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_583),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_522),
.B(n_373),
.Y(n_586)
);

OAI22xp5_ASAP7_75t_L g587 ( 
.A1(n_547),
.A2(n_530),
.B1(n_532),
.B2(n_538),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_587),
.B(n_544),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_522),
.B(n_348),
.Y(n_590)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_590),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_591),
.B(n_577),
.Y(n_622)
);

NAND3xp33_ASAP7_75t_L g594 ( 
.A(n_574),
.B(n_538),
.C(n_544),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_594),
.B(n_605),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_L g628 ( 
.A1(n_595),
.A2(n_589),
.B1(n_584),
.B2(n_585),
.Y(n_628)
);

XOR2xp5_ASAP7_75t_L g619 ( 
.A(n_596),
.B(n_598),
.Y(n_619)
);

XNOR2xp5_ASAP7_75t_SL g599 ( 
.A(n_559),
.B(n_571),
.Y(n_599)
);

XOR2xp5_ASAP7_75t_L g636 ( 
.A(n_599),
.B(n_606),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g600 ( 
.A1(n_588),
.A2(n_534),
.B(n_517),
.Y(n_600)
);

OAI21xp5_ASAP7_75t_SL g626 ( 
.A1(n_600),
.A2(n_616),
.B(n_563),
.Y(n_626)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_569),
.B(n_531),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_SL g620 ( 
.A(n_602),
.B(n_617),
.Y(n_620)
);

XNOR2xp5_ASAP7_75t_L g605 ( 
.A(n_564),
.B(n_549),
.Y(n_605)
);

XNOR2xp5_ASAP7_75t_SL g606 ( 
.A(n_571),
.B(n_551),
.Y(n_606)
);

XNOR2xp5_ASAP7_75t_L g608 ( 
.A(n_575),
.B(n_576),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_608),
.B(n_611),
.Y(n_627)
);

MAJx2_ASAP7_75t_L g611 ( 
.A(n_560),
.B(n_551),
.C(n_541),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_613),
.B(n_614),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_562),
.B(n_536),
.C(n_366),
.Y(n_614)
);

OAI21xp5_ASAP7_75t_SL g615 ( 
.A1(n_588),
.A2(n_536),
.B(n_363),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_615),
.B(n_339),
.Y(n_640)
);

OAI21xp5_ASAP7_75t_L g616 ( 
.A1(n_558),
.A2(n_566),
.B(n_570),
.Y(n_616)
);

BUFx24_ASAP7_75t_SL g617 ( 
.A(n_568),
.Y(n_617)
);

XOR2xp5_ASAP7_75t_L g618 ( 
.A(n_560),
.B(n_369),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g624 ( 
.A(n_618),
.B(n_573),
.C(n_583),
.Y(n_624)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_609),
.Y(n_621)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_621),
.Y(n_649)
);

OAI21xp5_ASAP7_75t_L g643 ( 
.A1(n_622),
.A2(n_626),
.B(n_638),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_624),
.B(n_640),
.Y(n_661)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_610),
.Y(n_625)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_625),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_628),
.B(n_630),
.Y(n_648)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_612),
.Y(n_629)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_629),
.Y(n_653)
);

CKINVDCx20_ASAP7_75t_R g630 ( 
.A(n_601),
.Y(n_630)
);

MAJIxp5_ASAP7_75t_L g631 ( 
.A(n_614),
.B(n_562),
.C(n_572),
.Y(n_631)
);

MAJIxp5_ASAP7_75t_L g644 ( 
.A(n_631),
.B(n_639),
.C(n_642),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_600),
.B(n_578),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_632),
.B(n_633),
.Y(n_652)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_607),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_603),
.B(n_590),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_634),
.B(n_635),
.Y(n_655)
);

OAI22xp5_ASAP7_75t_SL g635 ( 
.A1(n_592),
.A2(n_579),
.B1(n_581),
.B2(n_582),
.Y(n_635)
);

INVxp67_ASAP7_75t_L g638 ( 
.A(n_597),
.Y(n_638)
);

MAJIxp5_ASAP7_75t_L g639 ( 
.A(n_593),
.B(n_580),
.C(n_565),
.Y(n_639)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_592),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g646 ( 
.A1(n_641),
.A2(n_616),
.B1(n_598),
.B2(n_613),
.Y(n_646)
);

MAJIxp5_ASAP7_75t_L g642 ( 
.A(n_593),
.B(n_561),
.C(n_586),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_L g674 ( 
.A1(n_646),
.A2(n_619),
.B1(n_636),
.B2(n_634),
.Y(n_674)
);

OAI22xp5_ASAP7_75t_L g647 ( 
.A1(n_630),
.A2(n_608),
.B1(n_604),
.B2(n_579),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_647),
.B(n_650),
.Y(n_675)
);

MAJIxp5_ASAP7_75t_L g650 ( 
.A(n_631),
.B(n_604),
.C(n_611),
.Y(n_650)
);

OAI21xp5_ASAP7_75t_SL g651 ( 
.A1(n_626),
.A2(n_591),
.B(n_606),
.Y(n_651)
);

INVxp67_ASAP7_75t_L g663 ( 
.A(n_651),
.Y(n_663)
);

AOI21xp5_ASAP7_75t_SL g654 ( 
.A1(n_632),
.A2(n_591),
.B(n_599),
.Y(n_654)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_654),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_SL g656 ( 
.A(n_623),
.B(n_605),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_SL g669 ( 
.A(n_656),
.B(n_658),
.Y(n_669)
);

OAI22xp5_ASAP7_75t_L g657 ( 
.A1(n_629),
.A2(n_618),
.B1(n_596),
.B2(n_339),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_657),
.B(n_636),
.Y(n_668)
);

BUFx24_ASAP7_75t_SL g658 ( 
.A(n_620),
.Y(n_658)
);

MAJIxp5_ASAP7_75t_L g659 ( 
.A(n_637),
.B(n_319),
.C(n_369),
.Y(n_659)
);

NOR2xp67_ASAP7_75t_SL g679 ( 
.A(n_659),
.B(n_660),
.Y(n_679)
);

MAJIxp5_ASAP7_75t_L g660 ( 
.A(n_639),
.B(n_624),
.C(n_642),
.Y(n_660)
);

OAI21xp5_ASAP7_75t_SL g662 ( 
.A1(n_622),
.A2(n_363),
.B(n_339),
.Y(n_662)
);

XNOR2xp5_ASAP7_75t_L g665 ( 
.A(n_662),
.B(n_625),
.Y(n_665)
);

MAJIxp5_ASAP7_75t_L g664 ( 
.A(n_644),
.B(n_638),
.C(n_641),
.Y(n_664)
);

NOR2xp67_ASAP7_75t_SL g690 ( 
.A(n_664),
.B(n_666),
.Y(n_690)
);

INVx1_ASAP7_75t_SL g682 ( 
.A(n_665),
.Y(n_682)
);

MAJIxp5_ASAP7_75t_L g666 ( 
.A(n_644),
.B(n_627),
.C(n_632),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_650),
.B(n_628),
.Y(n_667)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_667),
.Y(n_689)
);

INVxp67_ASAP7_75t_L g686 ( 
.A(n_668),
.Y(n_686)
);

INVx6_ASAP7_75t_L g670 ( 
.A(n_660),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_670),
.B(n_677),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_661),
.B(n_621),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_671),
.B(n_672),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_648),
.B(n_635),
.Y(n_672)
);

XOR2xp5_ASAP7_75t_L g673 ( 
.A(n_643),
.B(n_654),
.Y(n_673)
);

XOR2xp5_ASAP7_75t_L g681 ( 
.A(n_673),
.B(n_652),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_674),
.B(n_676),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_648),
.B(n_633),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_SL g677 ( 
.A(n_653),
.B(n_619),
.Y(n_677)
);

MAJIxp5_ASAP7_75t_L g680 ( 
.A(n_675),
.B(n_643),
.C(n_655),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_680),
.B(n_684),
.Y(n_693)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_681),
.Y(n_701)
);

XOR2xp5_ASAP7_75t_L g684 ( 
.A(n_666),
.B(n_655),
.Y(n_684)
);

AOI21x1_ASAP7_75t_L g685 ( 
.A1(n_663),
.A2(n_653),
.B(n_651),
.Y(n_685)
);

AOI21xp5_ASAP7_75t_L g696 ( 
.A1(n_685),
.A2(n_691),
.B(n_665),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_670),
.B(n_659),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_688),
.B(n_667),
.Y(n_697)
);

AOI21xp33_ASAP7_75t_L g691 ( 
.A1(n_678),
.A2(n_652),
.B(n_645),
.Y(n_691)
);

AOI21xp33_ASAP7_75t_L g694 ( 
.A1(n_689),
.A2(n_663),
.B(n_673),
.Y(n_694)
);

OAI21xp5_ASAP7_75t_L g706 ( 
.A1(n_694),
.A2(n_696),
.B(n_699),
.Y(n_706)
);

MAJIxp5_ASAP7_75t_L g695 ( 
.A(n_684),
.B(n_664),
.C(n_679),
.Y(n_695)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_695),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_697),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_686),
.B(n_669),
.Y(n_698)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_698),
.Y(n_705)
);

AOI21x1_ASAP7_75t_L g699 ( 
.A1(n_687),
.A2(n_674),
.B(n_662),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_686),
.B(n_649),
.Y(n_700)
);

OAI21xp5_ASAP7_75t_SL g704 ( 
.A1(n_700),
.A2(n_683),
.B(n_692),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_704),
.B(n_681),
.Y(n_708)
);

OAI22xp5_ASAP7_75t_L g707 ( 
.A1(n_702),
.A2(n_701),
.B1(n_695),
.B2(n_693),
.Y(n_707)
);

OAI21x1_ASAP7_75t_SL g711 ( 
.A1(n_707),
.A2(n_708),
.B(n_709),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_705),
.B(n_703),
.Y(n_709)
);

OAI31xp33_ASAP7_75t_SL g710 ( 
.A1(n_708),
.A2(n_706),
.A3(n_694),
.B(n_690),
.Y(n_710)
);

OAI21xp5_ASAP7_75t_L g712 ( 
.A1(n_710),
.A2(n_682),
.B(n_645),
.Y(n_712)
);

A2O1A1Ixp33_ASAP7_75t_L g713 ( 
.A1(n_712),
.A2(n_711),
.B(n_682),
.C(n_367),
.Y(n_713)
);

XNOR2xp5_ASAP7_75t_L g714 ( 
.A(n_713),
.B(n_367),
.Y(n_714)
);


endmodule