module fake_jpeg_997_n_57 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_57);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_57;

wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx8_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx6_ASAP7_75t_SL g22 ( 
.A(n_17),
.Y(n_22)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_17),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_24),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_0),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_17),
.Y(n_27)
);

INVxp67_ASAP7_75t_SL g31 ( 
.A(n_27),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_18),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_28),
.B(n_21),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_26),
.B(n_21),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_33),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_28),
.A2(n_19),
.B1(n_23),
.B2(n_18),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_32),
.A2(n_19),
.B1(n_20),
.B2(n_16),
.Y(n_38)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_31),
.A2(n_22),
.B(n_29),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_35),
.A2(n_0),
.B(n_1),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_16),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_2),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_37),
.B(n_33),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_43),
.C(n_44),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_35),
.A2(n_32),
.B(n_34),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_42),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_44),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_47),
.B(n_3),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_36),
.C(n_38),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_49),
.C(n_8),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_9),
.C(n_14),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_50),
.B(n_4),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_52),
.C(n_11),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_46),
.C(n_10),
.Y(n_52)
);

BUFx24_ASAP7_75t_SL g55 ( 
.A(n_53),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_54),
.C(n_15),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_6),
.Y(n_57)
);


endmodule