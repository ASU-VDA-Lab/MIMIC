module fake_jpeg_7347_n_279 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_279);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_279;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx11_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx24_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_38),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_33),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_40),
.Y(n_54)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_42),
.Y(n_65)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_45),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_18),
.B(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_43),
.A2(n_30),
.B1(n_32),
.B2(n_26),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_59),
.B1(n_24),
.B2(n_22),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_43),
.A2(n_30),
.B1(n_27),
.B2(n_34),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_51),
.A2(n_16),
.B1(n_35),
.B2(n_22),
.Y(n_72)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_61),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_55),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_32),
.B1(n_26),
.B2(n_36),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_57),
.A2(n_16),
.B1(n_35),
.B2(n_37),
.Y(n_82)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_33),
.B1(n_18),
.B2(n_24),
.Y(n_59)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_25),
.B1(n_34),
.B2(n_17),
.Y(n_60)
);

OA22x2_ASAP7_75t_L g80 ( 
.A1(n_60),
.A2(n_37),
.B1(n_27),
.B2(n_36),
.Y(n_80)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_63),
.B(n_41),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_68),
.B(n_75),
.Y(n_109)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_69),
.B(n_70),
.Y(n_111)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_54),
.A2(n_46),
.B(n_39),
.C(n_19),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_71),
.A2(n_13),
.B(n_14),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_72),
.A2(n_80),
.B1(n_96),
.B2(n_98),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_73),
.A2(n_82),
.B1(n_90),
.B2(n_95),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_62),
.B(n_39),
.Y(n_75)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_45),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_77),
.B(n_79),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_55),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_67),
.B(n_39),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_84),
.B(n_85),
.Y(n_138)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_31),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_87),
.B(n_89),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_49),
.B(n_31),
.Y(n_88)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_55),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_51),
.A2(n_29),
.B1(n_23),
.B2(n_21),
.Y(n_90)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_92),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_54),
.B(n_29),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_93),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_50),
.A2(n_23),
.B1(n_21),
.B2(n_20),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_59),
.A2(n_29),
.B1(n_23),
.B2(n_21),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_64),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_60),
.A2(n_25),
.B1(n_1),
.B2(n_0),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_50),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_100),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_60),
.B(n_65),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_60),
.B(n_25),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_101),
.B(n_102),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_50),
.Y(n_102)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_60),
.B(n_25),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g129 ( 
.A(n_104),
.B(n_9),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_66),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_6),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_52),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_107),
.A2(n_63),
.B1(n_61),
.B2(n_58),
.Y(n_112)
);

INVx13_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_108),
.B(n_120),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_112),
.A2(n_113),
.B1(n_124),
.B2(n_136),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_100),
.A2(n_53),
.B1(n_56),
.B2(n_5),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_101),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_116),
.A2(n_125),
.B1(n_128),
.B2(n_130),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_118),
.B(n_134),
.Y(n_144)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_104),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_98),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_128)
);

XOR2x1_ASAP7_75t_L g165 ( 
.A(n_129),
.B(n_132),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_68),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_130)
);

NOR2x1_ASAP7_75t_L g132 ( 
.A(n_71),
.B(n_80),
.Y(n_132)
);

AND2x6_ASAP7_75t_L g134 ( 
.A(n_80),
.B(n_15),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_80),
.A2(n_87),
.B1(n_86),
.B2(n_96),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_137),
.A2(n_13),
.B(n_106),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_131),
.A2(n_91),
.B1(n_92),
.B2(n_99),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_140),
.A2(n_152),
.B1(n_115),
.B2(n_117),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_135),
.B(n_72),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_141),
.B(n_149),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_145),
.A2(n_130),
.B(n_133),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_119),
.B(n_74),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_146),
.B(n_147),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_119),
.B(n_91),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_121),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_153),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_102),
.Y(n_149)
);

AO22x1_ASAP7_75t_L g150 ( 
.A1(n_132),
.A2(n_78),
.B1(n_81),
.B2(n_83),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_155),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_103),
.Y(n_151)
);

NOR2x1_ASAP7_75t_SL g178 ( 
.A(n_151),
.B(n_118),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_110),
.A2(n_122),
.B1(n_126),
.B2(n_139),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_89),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_111),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_159),
.Y(n_172)
);

OAI32xp33_ASAP7_75t_L g158 ( 
.A1(n_113),
.A2(n_105),
.A3(n_81),
.B1(n_78),
.B2(n_85),
.Y(n_158)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_158),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_122),
.B(n_79),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_70),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_160),
.B(n_161),
.C(n_116),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_110),
.B(n_69),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_97),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_162),
.B(n_163),
.Y(n_186)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_114),
.Y(n_163)
);

OAI22x1_ASAP7_75t_SL g164 ( 
.A1(n_134),
.A2(n_129),
.B1(n_112),
.B2(n_137),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_164),
.A2(n_128),
.B1(n_127),
.B2(n_133),
.Y(n_168)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_117),
.Y(n_166)
);

INVx2_ASAP7_75t_SL g190 ( 
.A(n_166),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_129),
.B(n_109),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_114),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_168),
.A2(n_181),
.B1(n_192),
.B2(n_154),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_155),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_174),
.Y(n_196)
);

OAI21xp33_ASAP7_75t_SL g193 ( 
.A1(n_173),
.A2(n_145),
.B(n_158),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_149),
.Y(n_174)
);

NOR2x1_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_118),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_175),
.B(n_189),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_177),
.B(n_191),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_178),
.A2(n_150),
.B(n_142),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_179),
.A2(n_178),
.B(n_175),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_144),
.A2(n_115),
.B1(n_123),
.B2(n_125),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_143),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_183),
.B(n_188),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_184),
.B(n_187),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_163),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_185),
.Y(n_197)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_151),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_108),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_151),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_120),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_164),
.A2(n_141),
.B1(n_161),
.B2(n_148),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_193),
.A2(n_207),
.B1(n_213),
.B2(n_187),
.Y(n_215)
);

NOR3xp33_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_165),
.C(n_167),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_205),
.Y(n_222)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_199),
.B(n_202),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_186),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_200),
.B(n_210),
.Y(n_229)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_184),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_172),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_203),
.B(n_208),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_192),
.B(n_154),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_206),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_182),
.A2(n_150),
.B1(n_166),
.B2(n_157),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_170),
.Y(n_208)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_170),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_211),
.B(n_176),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_169),
.B(n_157),
.Y(n_212)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_212),
.Y(n_216)
);

OAI21xp33_ASAP7_75t_SL g213 ( 
.A1(n_189),
.A2(n_180),
.B(n_179),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_215),
.B(n_201),
.Y(n_236)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_212),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_218),
.B(n_221),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_191),
.C(n_177),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_220),
.C(n_227),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_195),
.B(n_174),
.C(n_180),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_198),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_225),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_209),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_204),
.A2(n_182),
.B1(n_168),
.B2(n_173),
.Y(n_226)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_226),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_183),
.C(n_176),
.Y(n_227)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_228),
.Y(n_242)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_207),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_230),
.B(n_202),
.Y(n_237)
);

INVxp33_ASAP7_75t_L g231 ( 
.A(n_214),
.Y(n_231)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_231),
.Y(n_246)
);

AOI21xp33_ASAP7_75t_SL g233 ( 
.A1(n_223),
.A2(n_210),
.B(n_201),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_233),
.A2(n_237),
.B(n_241),
.Y(n_253)
);

AOI221xp5_ASAP7_75t_L g234 ( 
.A1(n_222),
.A2(n_206),
.B1(n_205),
.B2(n_211),
.C(n_208),
.Y(n_234)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_234),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_240),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_221),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_239),
.B(n_185),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_220),
.B(n_199),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_214),
.Y(n_241)
);

A2O1A1O1Ixp25_ASAP7_75t_L g243 ( 
.A1(n_223),
.A2(n_203),
.B(n_190),
.C(n_197),
.D(n_185),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_245),
.Y(n_248)
);

BUFx12_ASAP7_75t_L g245 ( 
.A(n_216),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_238),
.A2(n_230),
.B1(n_218),
.B2(n_216),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_249),
.A2(n_242),
.B1(n_215),
.B2(n_231),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_219),
.C(n_217),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_254),
.C(n_228),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_227),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_255),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_217),
.C(n_229),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_254),
.B(n_190),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_256),
.B(n_257),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_253),
.B(n_235),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_190),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_258),
.A2(n_259),
.B(n_246),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_236),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_260),
.B(n_250),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_261),
.B(n_251),
.C(n_248),
.Y(n_266)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_264),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_265),
.B(n_266),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_262),
.A2(n_247),
.B(n_245),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_267),
.B(n_243),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_263),
.B(n_261),
.Y(n_268)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_268),
.Y(n_274)
);

OR2x2_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_245),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_270),
.B(n_260),
.Y(n_272)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_272),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_273),
.A2(n_271),
.B(n_226),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_274),
.Y(n_277)
);

AOI21x1_ASAP7_75t_L g278 ( 
.A1(n_277),
.A2(n_239),
.B(n_275),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_197),
.Y(n_279)
);


endmodule