module real_aes_7315_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_755;
wire n_153;
wire n_532;
wire n_316;
wire n_284;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g445 ( .A(n_0), .Y(n_445) );
INVx1_ASAP7_75t_L g501 ( .A(n_1), .Y(n_501) );
INVx1_ASAP7_75t_L g188 ( .A(n_2), .Y(n_188) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_3), .A2(n_37), .B1(n_160), .B2(n_510), .Y(n_509) );
AOI21xp33_ASAP7_75t_L g199 ( .A1(n_4), .A2(n_117), .B(n_200), .Y(n_199) );
AOI22xp5_ASAP7_75t_SL g458 ( .A1(n_5), .A2(n_443), .B1(n_459), .B2(n_747), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_6), .B(n_147), .Y(n_493) );
AND2x6_ASAP7_75t_L g122 ( .A(n_7), .B(n_123), .Y(n_122) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_8), .A2(n_168), .B(n_169), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_9), .B(n_38), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_10), .B(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g205 ( .A(n_11), .Y(n_205) );
INVx1_ASAP7_75t_L g143 ( .A(n_12), .Y(n_143) );
INVx1_ASAP7_75t_L g497 ( .A(n_13), .Y(n_497) );
INVx1_ASAP7_75t_L g176 ( .A(n_14), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_15), .B(n_191), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_16), .B(n_139), .Y(n_560) );
AOI22xp5_ASAP7_75t_L g742 ( .A1(n_17), .A2(n_41), .B1(n_743), .B2(n_744), .Y(n_742) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_17), .Y(n_744) );
AO32x2_ASAP7_75t_L g507 ( .A1(n_18), .A2(n_138), .A3(n_147), .B1(n_479), .B2(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_19), .B(n_160), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_20), .B(n_133), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_21), .B(n_139), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_22), .A2(n_50), .B1(n_160), .B2(n_510), .Y(n_511) );
NAND2xp5_ASAP7_75t_SL g116 ( .A(n_23), .B(n_117), .Y(n_116) );
AOI22xp33_ASAP7_75t_SL g546 ( .A1(n_24), .A2(n_77), .B1(n_160), .B2(n_191), .Y(n_546) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_25), .B(n_160), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_26), .B(n_198), .Y(n_226) );
A2O1A1Ixp33_ASAP7_75t_L g172 ( .A1(n_27), .A2(n_173), .B(n_175), .C(n_177), .Y(n_172) );
BUFx6f_ASAP7_75t_L g121 ( .A(n_28), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_29), .B(n_151), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_30), .B(n_158), .Y(n_189) );
INVx1_ASAP7_75t_L g215 ( .A(n_31), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_32), .B(n_151), .Y(n_523) );
INVx2_ASAP7_75t_L g120 ( .A(n_33), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_34), .B(n_160), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_35), .B(n_151), .Y(n_533) );
A2O1A1Ixp33_ASAP7_75t_L g124 ( .A1(n_36), .A2(n_122), .B(n_125), .C(n_128), .Y(n_124) );
INVx1_ASAP7_75t_L g213 ( .A(n_39), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_40), .B(n_158), .Y(n_249) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_41), .Y(n_743) );
AOI22xp5_ASAP7_75t_L g738 ( .A1(n_42), .A2(n_739), .B1(n_740), .B2(n_746), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_42), .Y(n_746) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_43), .B(n_160), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_44), .A2(n_88), .B1(n_136), .B2(n_510), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_45), .B(n_160), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_46), .B(n_160), .Y(n_498) );
CKINVDCx16_ASAP7_75t_R g216 ( .A(n_47), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_48), .B(n_477), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_49), .B(n_117), .Y(n_161) );
AOI22xp33_ASAP7_75t_SL g558 ( .A1(n_51), .A2(n_60), .B1(n_160), .B2(n_191), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g211 ( .A1(n_52), .A2(n_125), .B1(n_191), .B2(n_212), .Y(n_211) );
CKINVDCx20_ASAP7_75t_R g145 ( .A(n_53), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_54), .B(n_160), .Y(n_478) );
CKINVDCx16_ASAP7_75t_R g184 ( .A(n_55), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_56), .B(n_160), .Y(n_527) );
A2O1A1Ixp33_ASAP7_75t_L g202 ( .A1(n_57), .A2(n_203), .B(n_204), .C(n_206), .Y(n_202) );
CKINVDCx20_ASAP7_75t_R g253 ( .A(n_58), .Y(n_253) );
INVx1_ASAP7_75t_L g201 ( .A(n_59), .Y(n_201) );
INVx1_ASAP7_75t_L g123 ( .A(n_61), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_62), .B(n_160), .Y(n_502) );
INVx1_ASAP7_75t_L g142 ( .A(n_63), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g453 ( .A(n_64), .Y(n_453) );
AOI222xp33_ASAP7_75t_L g103 ( .A1(n_65), .A2(n_104), .B1(n_450), .B2(n_457), .C1(n_750), .C2(n_755), .Y(n_103) );
OAI22xp5_ASAP7_75t_SL g437 ( .A1(n_65), .A2(n_74), .B1(n_438), .B2(n_439), .Y(n_437) );
CKINVDCx16_ASAP7_75t_R g438 ( .A(n_65), .Y(n_438) );
AO32x2_ASAP7_75t_L g543 ( .A1(n_65), .A2(n_147), .A3(n_150), .B1(n_479), .B2(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g475 ( .A(n_66), .Y(n_475) );
INVx1_ASAP7_75t_L g518 ( .A(n_67), .Y(n_518) );
A2O1A1Ixp33_ASAP7_75t_SL g223 ( .A1(n_68), .A2(n_133), .B(n_206), .C(n_224), .Y(n_223) );
INVxp67_ASAP7_75t_L g225 ( .A(n_69), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g519 ( .A(n_70), .B(n_191), .Y(n_519) );
INVx1_ASAP7_75t_L g456 ( .A(n_71), .Y(n_456) );
CKINVDCx20_ASAP7_75t_R g218 ( .A(n_72), .Y(n_218) );
INVx1_ASAP7_75t_L g246 ( .A(n_73), .Y(n_246) );
CKINVDCx16_ASAP7_75t_R g439 ( .A(n_74), .Y(n_439) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_75), .Y(n_448) );
OAI22xp5_ASAP7_75t_SL g434 ( .A1(n_76), .A2(n_90), .B1(n_435), .B2(n_436), .Y(n_434) );
CKINVDCx20_ASAP7_75t_R g435 ( .A(n_76), .Y(n_435) );
A2O1A1Ixp33_ASAP7_75t_L g247 ( .A1(n_78), .A2(n_122), .B(n_125), .C(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_79), .B(n_510), .Y(n_532) );
OAI22xp5_ASAP7_75t_SL g740 ( .A1(n_80), .A2(n_741), .B1(n_742), .B2(n_745), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_80), .Y(n_745) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_81), .B(n_191), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g129 ( .A(n_82), .B(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g140 ( .A(n_83), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_84), .B(n_133), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_85), .B(n_191), .Y(n_488) );
A2O1A1Ixp33_ASAP7_75t_L g186 ( .A1(n_86), .A2(n_122), .B(n_125), .C(n_187), .Y(n_186) );
OR2x2_ASAP7_75t_L g442 ( .A(n_87), .B(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g462 ( .A(n_87), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_89), .A2(n_102), .B1(n_191), .B2(n_192), .Y(n_557) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_90), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_91), .B(n_151), .Y(n_207) );
CKINVDCx20_ASAP7_75t_R g194 ( .A(n_92), .Y(n_194) );
A2O1A1Ixp33_ASAP7_75t_L g153 ( .A1(n_93), .A2(n_122), .B(n_125), .C(n_154), .Y(n_153) );
CKINVDCx20_ASAP7_75t_R g163 ( .A(n_94), .Y(n_163) );
INVx1_ASAP7_75t_L g222 ( .A(n_95), .Y(n_222) );
CKINVDCx16_ASAP7_75t_R g170 ( .A(n_96), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g155 ( .A(n_97), .B(n_130), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_98), .B(n_191), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_99), .B(n_147), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_100), .A2(n_117), .B(n_221), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_101), .B(n_456), .Y(n_455) );
INVxp67_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
AOI21xp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_440), .B(n_447), .Y(n_105) );
XOR2xp5_ASAP7_75t_L g106 ( .A(n_107), .B(n_437), .Y(n_106) );
OAI22xp5_ASAP7_75t_SL g107 ( .A1(n_108), .A2(n_109), .B1(n_433), .B2(n_434), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
OAI22xp5_ASAP7_75t_L g460 ( .A1(n_109), .A2(n_461), .B1(n_462), .B2(n_463), .Y(n_460) );
AND2x2_ASAP7_75t_SL g109 ( .A(n_110), .B(n_402), .Y(n_109) );
NOR3xp33_ASAP7_75t_L g110 ( .A(n_111), .B(n_295), .C(n_368), .Y(n_110) );
OAI211xp5_ASAP7_75t_SL g111 ( .A1(n_112), .A2(n_180), .B(n_227), .C(n_279), .Y(n_111) );
INVxp67_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AND2x2_ASAP7_75t_L g113 ( .A(n_114), .B(n_148), .Y(n_113) );
AND2x2_ASAP7_75t_L g243 ( .A(n_114), .B(n_244), .Y(n_243) );
INVx3_ASAP7_75t_L g262 ( .A(n_114), .Y(n_262) );
INVx2_ASAP7_75t_L g277 ( .A(n_114), .Y(n_277) );
INVx1_ASAP7_75t_L g307 ( .A(n_114), .Y(n_307) );
AND2x2_ASAP7_75t_L g357 ( .A(n_114), .B(n_278), .Y(n_357) );
AOI32xp33_ASAP7_75t_L g384 ( .A1(n_114), .A2(n_312), .A3(n_385), .B1(n_387), .B2(n_388), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_114), .B(n_233), .Y(n_390) );
AND2x2_ASAP7_75t_L g417 ( .A(n_114), .B(n_260), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_114), .B(n_426), .Y(n_425) );
OR2x6_ASAP7_75t_L g114 ( .A(n_115), .B(n_144), .Y(n_114) );
AOI21xp5_ASAP7_75t_SL g115 ( .A1(n_116), .A2(n_124), .B(n_137), .Y(n_115) );
BUFx2_ASAP7_75t_L g168 ( .A(n_117), .Y(n_168) );
AND2x4_ASAP7_75t_L g117 ( .A(n_118), .B(n_122), .Y(n_117) );
NAND2x1p5_ASAP7_75t_L g185 ( .A(n_118), .B(n_122), .Y(n_185) );
AND2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_121), .Y(n_118) );
INVx1_ASAP7_75t_L g477 ( .A(n_119), .Y(n_477) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g126 ( .A(n_120), .Y(n_126) );
INVx1_ASAP7_75t_L g192 ( .A(n_120), .Y(n_192) );
INVx1_ASAP7_75t_L g127 ( .A(n_121), .Y(n_127) );
INVx3_ASAP7_75t_L g131 ( .A(n_121), .Y(n_131) );
INVx1_ASAP7_75t_L g133 ( .A(n_121), .Y(n_133) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_121), .Y(n_158) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_121), .Y(n_174) );
INVx4_ASAP7_75t_SL g178 ( .A(n_122), .Y(n_178) );
BUFx3_ASAP7_75t_L g479 ( .A(n_122), .Y(n_479) );
OAI21xp5_ASAP7_75t_L g485 ( .A1(n_122), .A2(n_486), .B(n_489), .Y(n_485) );
OAI21xp5_ASAP7_75t_L g495 ( .A1(n_122), .A2(n_496), .B(n_500), .Y(n_495) );
OAI21xp5_ASAP7_75t_L g516 ( .A1(n_122), .A2(n_517), .B(n_520), .Y(n_516) );
OAI21xp5_ASAP7_75t_L g525 ( .A1(n_122), .A2(n_526), .B(n_530), .Y(n_525) );
INVx5_ASAP7_75t_L g171 ( .A(n_125), .Y(n_171) );
AND2x6_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
BUFx3_ASAP7_75t_L g136 ( .A(n_126), .Y(n_136) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_126), .Y(n_160) );
INVx1_ASAP7_75t_L g510 ( .A(n_126), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_132), .B(n_134), .Y(n_128) );
O2A1O1Ixp33_ASAP7_75t_L g187 ( .A1(n_130), .A2(n_188), .B(n_189), .C(n_190), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_130), .A2(n_472), .B(n_473), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g486 ( .A1(n_130), .A2(n_487), .B(n_488), .Y(n_486) );
INVx2_ASAP7_75t_L g492 ( .A(n_130), .Y(n_492) );
O2A1O1Ixp5_ASAP7_75t_SL g517 ( .A1(n_130), .A2(n_206), .B(n_518), .C(n_519), .Y(n_517) );
INVx5_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_131), .B(n_205), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_131), .B(n_225), .Y(n_224) );
OAI22xp5_ASAP7_75t_SL g544 ( .A1(n_131), .A2(n_158), .B1(n_545), .B2(n_546), .Y(n_544) );
INVx1_ASAP7_75t_L g529 ( .A(n_133), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_134), .A2(n_249), .B(n_250), .Y(n_248) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g177 ( .A(n_136), .Y(n_177) );
INVx1_ASAP7_75t_L g251 ( .A(n_137), .Y(n_251) );
OA21x2_ASAP7_75t_L g469 ( .A1(n_137), .A2(n_470), .B(n_480), .Y(n_469) );
OA21x2_ASAP7_75t_L g494 ( .A1(n_137), .A2(n_495), .B(n_503), .Y(n_494) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AO21x2_ASAP7_75t_L g182 ( .A1(n_138), .A2(n_183), .B(n_193), .Y(n_182) );
AO21x2_ASAP7_75t_L g209 ( .A1(n_138), .A2(n_210), .B(n_217), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_138), .B(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_139), .Y(n_147) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
AND2x2_ASAP7_75t_SL g151 ( .A(n_140), .B(n_141), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
NOR2xp33_ASAP7_75t_SL g144 ( .A(n_145), .B(n_146), .Y(n_144) );
INVx3_ASAP7_75t_L g198 ( .A(n_146), .Y(n_198) );
AO21x1_ASAP7_75t_L g555 ( .A1(n_146), .A2(n_556), .B(n_559), .Y(n_555) );
NAND3xp33_ASAP7_75t_L g580 ( .A(n_146), .B(n_479), .C(n_556), .Y(n_580) );
INVx4_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
OA21x2_ASAP7_75t_L g219 ( .A1(n_147), .A2(n_220), .B(n_226), .Y(n_219) );
OA21x2_ASAP7_75t_L g484 ( .A1(n_147), .A2(n_485), .B(n_493), .Y(n_484) );
AND2x2_ASAP7_75t_L g306 ( .A(n_148), .B(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g328 ( .A(n_148), .Y(n_328) );
AND2x2_ASAP7_75t_L g413 ( .A(n_148), .B(n_243), .Y(n_413) );
AND2x2_ASAP7_75t_L g416 ( .A(n_148), .B(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g148 ( .A(n_149), .B(n_165), .Y(n_148) );
INVx2_ASAP7_75t_L g235 ( .A(n_149), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_149), .B(n_260), .Y(n_266) );
AND2x2_ASAP7_75t_L g276 ( .A(n_149), .B(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g312 ( .A(n_149), .Y(n_312) );
AO21x2_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_152), .B(n_162), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g164 ( .A(n_151), .Y(n_164) );
OA21x2_ASAP7_75t_L g166 ( .A1(n_151), .A2(n_167), .B(n_179), .Y(n_166) );
OA21x2_ASAP7_75t_L g515 ( .A1(n_151), .A2(n_516), .B(n_523), .Y(n_515) );
OA21x2_ASAP7_75t_L g524 ( .A1(n_151), .A2(n_525), .B(n_533), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_153), .B(n_161), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_156), .B(n_159), .Y(n_154) );
INVx4_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g203 ( .A(n_158), .Y(n_203) );
OAI22xp5_ASAP7_75t_L g508 ( .A1(n_158), .A2(n_492), .B1(n_509), .B2(n_511), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g556 ( .A1(n_158), .A2(n_492), .B1(n_557), .B2(n_558), .Y(n_556) );
HB1xp67_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx3_ASAP7_75t_L g206 ( .A(n_160), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_163), .B(n_164), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_164), .B(n_194), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_164), .B(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g254 ( .A(n_165), .B(n_235), .Y(n_254) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx2_ASAP7_75t_L g236 ( .A(n_166), .Y(n_236) );
AND2x2_ASAP7_75t_L g278 ( .A(n_166), .B(n_260), .Y(n_278) );
AND2x2_ASAP7_75t_L g347 ( .A(n_166), .B(n_244), .Y(n_347) );
O2A1O1Ixp33_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_171), .B(n_172), .C(n_178), .Y(n_169) );
O2A1O1Ixp33_ASAP7_75t_L g200 ( .A1(n_171), .A2(n_178), .B(n_201), .C(n_202), .Y(n_200) );
O2A1O1Ixp33_ASAP7_75t_L g221 ( .A1(n_171), .A2(n_178), .B(n_222), .C(n_223), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_173), .B(n_176), .Y(n_175) );
INVx1_ASAP7_75t_L g499 ( .A(n_173), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_173), .A2(n_521), .B(n_522), .Y(n_520) );
INVx4_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
OAI22xp5_ASAP7_75t_SL g212 ( .A1(n_174), .A2(n_213), .B1(n_214), .B2(n_215), .Y(n_212) );
INVx2_ASAP7_75t_L g214 ( .A(n_174), .Y(n_214) );
OAI22xp33_ASAP7_75t_L g210 ( .A1(n_178), .A2(n_185), .B1(n_211), .B2(n_216), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_181), .B(n_195), .Y(n_180) );
OR2x2_ASAP7_75t_L g241 ( .A(n_181), .B(n_209), .Y(n_241) );
INVx1_ASAP7_75t_L g320 ( .A(n_181), .Y(n_320) );
AND2x2_ASAP7_75t_L g334 ( .A(n_181), .B(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_181), .B(n_208), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_181), .B(n_332), .Y(n_386) );
AND2x2_ASAP7_75t_L g394 ( .A(n_181), .B(n_395), .Y(n_394) );
INVx3_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVx3_ASAP7_75t_L g231 ( .A(n_182), .Y(n_231) );
AND2x2_ASAP7_75t_L g301 ( .A(n_182), .B(n_209), .Y(n_301) );
OAI21xp5_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_185), .B(n_186), .Y(n_183) );
OAI21xp5_ASAP7_75t_L g245 ( .A1(n_185), .A2(n_246), .B(n_247), .Y(n_245) );
O2A1O1Ixp33_ASAP7_75t_L g496 ( .A1(n_190), .A2(n_497), .B(n_498), .C(n_499), .Y(n_496) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx3_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_195), .B(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g428 ( .A(n_195), .Y(n_428) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_208), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_196), .B(n_272), .Y(n_294) );
OR2x2_ASAP7_75t_L g323 ( .A(n_196), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g355 ( .A(n_196), .B(n_335), .Y(n_355) );
INVx1_ASAP7_75t_SL g375 ( .A(n_196), .Y(n_375) );
AND2x2_ASAP7_75t_L g379 ( .A(n_196), .B(n_240), .Y(n_379) );
INVx2_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
AND2x2_ASAP7_75t_SL g232 ( .A(n_197), .B(n_208), .Y(n_232) );
AND2x2_ASAP7_75t_L g239 ( .A(n_197), .B(n_219), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_197), .B(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g282 ( .A(n_197), .B(n_264), .Y(n_282) );
INVx1_ASAP7_75t_SL g289 ( .A(n_197), .Y(n_289) );
BUFx2_ASAP7_75t_L g300 ( .A(n_197), .Y(n_300) );
AND2x2_ASAP7_75t_L g316 ( .A(n_197), .B(n_231), .Y(n_316) );
AND2x2_ASAP7_75t_L g331 ( .A(n_197), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g395 ( .A(n_197), .B(n_209), .Y(n_395) );
OA21x2_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_199), .B(n_207), .Y(n_197) );
O2A1O1Ixp5_ASAP7_75t_L g474 ( .A1(n_203), .A2(n_475), .B(n_476), .C(n_478), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_203), .A2(n_531), .B(n_532), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_208), .B(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g319 ( .A(n_208), .B(n_320), .Y(n_319) );
AOI221xp5_ASAP7_75t_L g336 ( .A1(n_208), .A2(n_337), .B1(n_340), .B2(n_343), .C(n_348), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_208), .B(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g208 ( .A(n_209), .B(n_219), .Y(n_208) );
INVx3_ASAP7_75t_L g264 ( .A(n_209), .Y(n_264) );
BUFx2_ASAP7_75t_L g274 ( .A(n_219), .Y(n_274) );
AND2x2_ASAP7_75t_L g288 ( .A(n_219), .B(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g305 ( .A(n_219), .Y(n_305) );
OR2x2_ASAP7_75t_L g324 ( .A(n_219), .B(n_264), .Y(n_324) );
INVx3_ASAP7_75t_L g332 ( .A(n_219), .Y(n_332) );
AND2x2_ASAP7_75t_L g335 ( .A(n_219), .B(n_264), .Y(n_335) );
AOI221xp5_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_233), .B1(n_237), .B2(n_242), .C(n_255), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_230), .B(n_232), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_230), .B(n_304), .Y(n_429) );
OR2x2_ASAP7_75t_L g432 ( .A(n_230), .B(n_263), .Y(n_432) );
INVx1_ASAP7_75t_SL g230 ( .A(n_231), .Y(n_230) );
OAI221xp5_ASAP7_75t_SL g255 ( .A1(n_231), .A2(n_256), .B1(n_263), .B2(n_265), .C(n_268), .Y(n_255) );
AND2x2_ASAP7_75t_L g272 ( .A(n_231), .B(n_264), .Y(n_272) );
AND2x2_ASAP7_75t_L g280 ( .A(n_231), .B(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_231), .B(n_288), .Y(n_287) );
NAND2x1_ASAP7_75t_L g330 ( .A(n_231), .B(n_331), .Y(n_330) );
OR2x2_ASAP7_75t_L g382 ( .A(n_231), .B(n_324), .Y(n_382) );
AOI22xp5_ASAP7_75t_L g370 ( .A1(n_233), .A2(n_342), .B1(n_371), .B2(n_373), .Y(n_370) );
INVx2_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AOI322xp5_ASAP7_75t_L g279 ( .A1(n_234), .A2(n_243), .A3(n_280), .B1(n_283), .B2(n_286), .C1(n_290), .C2(n_293), .Y(n_279) );
OR2x2_ASAP7_75t_L g291 ( .A(n_234), .B(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_236), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_235), .B(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g270 ( .A(n_235), .B(n_244), .Y(n_270) );
INVx1_ASAP7_75t_L g285 ( .A(n_235), .Y(n_285) );
AND2x2_ASAP7_75t_L g351 ( .A(n_235), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g261 ( .A(n_236), .B(n_262), .Y(n_261) );
INVx2_ASAP7_75t_L g352 ( .A(n_236), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_236), .B(n_260), .Y(n_426) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_239), .B(n_240), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_240), .B(n_375), .Y(n_374) );
INVx3_ASAP7_75t_SL g240 ( .A(n_241), .Y(n_240) );
OR2x2_ASAP7_75t_L g326 ( .A(n_241), .B(n_273), .Y(n_326) );
OR2x2_ASAP7_75t_L g423 ( .A(n_241), .B(n_274), .Y(n_423) );
INVx1_ASAP7_75t_L g404 ( .A(n_242), .Y(n_404) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_254), .Y(n_242) );
INVx4_ASAP7_75t_L g292 ( .A(n_243), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_243), .B(n_311), .Y(n_317) );
INVx2_ASAP7_75t_L g260 ( .A(n_244), .Y(n_260) );
AO21x2_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_251), .B(n_252), .Y(n_244) );
INVx1_ASAP7_75t_L g342 ( .A(n_254), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_254), .B(n_314), .Y(n_383) );
AOI21xp33_ASAP7_75t_L g329 ( .A1(n_256), .A2(n_330), .B(n_333), .Y(n_329) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_261), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g314 ( .A(n_260), .Y(n_314) );
INVx1_ASAP7_75t_L g341 ( .A(n_260), .Y(n_341) );
INVx1_ASAP7_75t_L g267 ( .A(n_261), .Y(n_267) );
AND2x2_ASAP7_75t_L g269 ( .A(n_261), .B(n_270), .Y(n_269) );
AND2x2_ASAP7_75t_L g365 ( .A(n_262), .B(n_351), .Y(n_365) );
AND2x2_ASAP7_75t_L g387 ( .A(n_262), .B(n_347), .Y(n_387) );
BUFx2_ASAP7_75t_L g339 ( .A(n_264), .Y(n_339) );
OR2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
AOI32xp33_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_271), .A3(n_272), .B1(n_273), .B2(n_275), .Y(n_268) );
INVx1_ASAP7_75t_L g349 ( .A(n_269), .Y(n_349) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_269), .A2(n_397), .B1(n_398), .B2(n_400), .Y(n_396) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g302 ( .A(n_272), .B(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_272), .B(n_331), .Y(n_372) );
AND2x2_ASAP7_75t_L g419 ( .A(n_272), .B(n_304), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_273), .B(n_320), .Y(n_367) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g420 ( .A(n_275), .Y(n_420) );
AND2x2_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
INVx1_ASAP7_75t_L g345 ( .A(n_276), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_278), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g392 ( .A(n_278), .B(n_312), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_278), .B(n_307), .Y(n_399) );
INVx1_ASAP7_75t_SL g381 ( .A(n_280), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_281), .B(n_332), .Y(n_359) );
NOR4xp25_ASAP7_75t_L g405 ( .A(n_281), .B(n_304), .C(n_406), .D(n_409), .Y(n_405) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_282), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVxp67_ASAP7_75t_L g362 ( .A(n_285), .Y(n_362) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
OAI21xp33_ASAP7_75t_L g412 ( .A1(n_288), .A2(n_379), .B(n_413), .Y(n_412) );
AND2x4_ASAP7_75t_L g304 ( .A(n_289), .B(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g353 ( .A(n_292), .Y(n_353) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND4xp25_ASAP7_75t_SL g295 ( .A(n_296), .B(n_321), .C(n_336), .D(n_356), .Y(n_295) );
O2A1O1Ixp33_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_302), .B(n_306), .C(n_308), .Y(n_296) );
INVx1_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_301), .Y(n_298) );
INVx1_ASAP7_75t_SL g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g388 ( .A(n_301), .B(n_331), .Y(n_388) );
AND2x2_ASAP7_75t_L g397 ( .A(n_301), .B(n_375), .Y(n_397) );
INVx3_ASAP7_75t_SL g303 ( .A(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_304), .B(n_339), .Y(n_401) );
AND2x2_ASAP7_75t_L g313 ( .A(n_307), .B(n_314), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_315), .B1(n_317), .B2(n_318), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_311), .B(n_313), .Y(n_310) );
AND2x2_ASAP7_75t_L g411 ( .A(n_311), .B(n_357), .Y(n_411) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_313), .B(n_362), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_314), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
O2A1O1Ixp33_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_325), .B(n_327), .C(n_329), .Y(n_321) );
AOI221xp5_ASAP7_75t_L g356 ( .A1(n_322), .A2(n_357), .B1(n_358), .B2(n_360), .C(n_363), .Y(n_356) );
INVx1_ASAP7_75t_SL g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
OAI221xp5_ASAP7_75t_L g414 ( .A1(n_330), .A2(n_415), .B1(n_418), .B2(n_420), .C(n_421), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_331), .B(n_339), .Y(n_338) );
INVx1_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_339), .B(n_408), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
INVx1_ASAP7_75t_L g369 ( .A(n_341), .Y(n_369) );
INVx1_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
OAI22xp5_ASAP7_75t_L g363 ( .A1(n_344), .A2(n_364), .B1(n_366), .B2(n_367), .Y(n_363) );
OR2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AOI21xp33_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_350), .B(n_354), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_351), .B(n_353), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_353), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OAI221xp5_ASAP7_75t_L g427 ( .A1(n_364), .A2(n_390), .B1(n_428), .B2(n_429), .C(n_430), .Y(n_427) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g409 ( .A(n_366), .Y(n_409) );
OAI211xp5_ASAP7_75t_SL g368 ( .A1(n_369), .A2(n_370), .B(n_376), .C(n_396), .Y(n_368) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AOI211xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_379), .B(n_380), .C(n_389), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
A2O1A1Ixp33_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_382), .B(n_383), .C(n_384), .Y(n_380) );
INVx1_ASAP7_75t_L g408 ( .A(n_386), .Y(n_408) );
OAI21xp5_ASAP7_75t_SL g430 ( .A1(n_387), .A2(n_413), .B(n_431), .Y(n_430) );
AOI21xp33_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_391), .B(n_393), .Y(n_389) );
INVx1_ASAP7_75t_SL g391 ( .A(n_392), .Y(n_391) );
INVxp67_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
OAI21xp5_ASAP7_75t_SL g422 ( .A1(n_399), .A2(n_423), .B(n_424), .Y(n_422) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
NOR3xp33_ASAP7_75t_L g402 ( .A(n_403), .B(n_414), .C(n_427), .Y(n_402) );
OAI211xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_405), .B(n_410), .C(n_412), .Y(n_403) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
CKINVDCx14_ASAP7_75t_R g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
OA21x2_ASAP7_75t_L g756 ( .A1(n_441), .A2(n_453), .B(n_454), .Y(n_756) );
BUFx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
HB1xp67_ASAP7_75t_L g449 ( .A(n_442), .Y(n_449) );
INVx1_ASAP7_75t_SL g754 ( .A(n_442), .Y(n_754) );
NOR2x2_ASAP7_75t_L g749 ( .A(n_443), .B(n_462), .Y(n_749) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_446), .Y(n_444) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_448), .B(n_449), .Y(n_447) );
AND2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_454), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NOR2xp33_ASAP7_75t_SL g752 ( .A(n_453), .B(n_455), .Y(n_752) );
INVx1_ASAP7_75t_SL g454 ( .A(n_455), .Y(n_454) );
INVxp67_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
XNOR2xp5_ASAP7_75t_L g459 ( .A(n_460), .B(n_738), .Y(n_459) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
OR3x1_ASAP7_75t_L g464 ( .A(n_465), .B(n_666), .C(n_715), .Y(n_464) );
NAND5xp2_ASAP7_75t_L g465 ( .A(n_466), .B(n_581), .C(n_609), .D(n_639), .E(n_653), .Y(n_465) );
AOI221xp5_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_504), .B1(n_534), .B2(n_539), .C(n_548), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_468), .B(n_481), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_468), .B(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g561 ( .A(n_469), .Y(n_561) );
AND2x2_ASAP7_75t_L g569 ( .A(n_469), .B(n_484), .Y(n_569) );
AND2x2_ASAP7_75t_L g592 ( .A(n_469), .B(n_483), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_469), .B(n_494), .Y(n_607) );
OR2x2_ASAP7_75t_L g616 ( .A(n_469), .B(n_555), .Y(n_616) );
HB1xp67_ASAP7_75t_L g619 ( .A(n_469), .Y(n_619) );
AND2x2_ASAP7_75t_L g727 ( .A(n_469), .B(n_555), .Y(n_727) );
OAI21xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_474), .B(n_479), .Y(n_470) );
O2A1O1Ixp33_ASAP7_75t_L g500 ( .A1(n_476), .A2(n_492), .B(n_501), .C(n_502), .Y(n_500) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_481), .B(n_619), .Y(n_675) );
INVx2_ASAP7_75t_SL g481 ( .A(n_482), .Y(n_481) );
OAI311xp33_ASAP7_75t_L g617 ( .A1(n_482), .A2(n_618), .A3(n_619), .B1(n_620), .C1(n_635), .Y(n_617) );
AND2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_494), .Y(n_482) );
AND2x2_ASAP7_75t_L g578 ( .A(n_483), .B(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g585 ( .A(n_483), .Y(n_585) );
AND2x2_ASAP7_75t_L g706 ( .A(n_483), .B(n_538), .Y(n_706) );
INVx3_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_484), .B(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g562 ( .A(n_484), .B(n_494), .Y(n_562) );
AND2x2_ASAP7_75t_L g614 ( .A(n_484), .B(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g628 ( .A(n_484), .B(n_561), .Y(n_628) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_491), .B(n_492), .Y(n_489) );
INVx2_ASAP7_75t_L g538 ( .A(n_494), .Y(n_538) );
AND2x2_ASAP7_75t_L g577 ( .A(n_494), .B(n_561), .Y(n_577) );
AND2x2_ASAP7_75t_L g504 ( .A(n_505), .B(n_512), .Y(n_504) );
OR2x2_ASAP7_75t_L g672 ( .A(n_505), .B(n_673), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_505), .B(n_678), .Y(n_689) );
INVx2_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g684 ( .A(n_506), .B(n_685), .Y(n_684) );
BUFx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g547 ( .A(n_507), .Y(n_547) );
AND2x2_ASAP7_75t_L g613 ( .A(n_507), .B(n_543), .Y(n_613) );
AND2x2_ASAP7_75t_L g624 ( .A(n_507), .B(n_524), .Y(n_624) );
AND2x2_ASAP7_75t_L g633 ( .A(n_507), .B(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_512), .B(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_512), .B(n_574), .Y(n_618) );
INVx2_ASAP7_75t_SL g512 ( .A(n_513), .Y(n_512) );
OR2x2_ASAP7_75t_L g605 ( .A(n_513), .B(n_564), .Y(n_605) );
OR2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_524), .Y(n_513) );
INVx2_ASAP7_75t_L g541 ( .A(n_514), .Y(n_541) );
AND2x2_ASAP7_75t_L g632 ( .A(n_514), .B(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g551 ( .A(n_515), .Y(n_551) );
OR2x2_ASAP7_75t_L g649 ( .A(n_515), .B(n_650), .Y(n_649) );
HB1xp67_ASAP7_75t_L g712 ( .A(n_515), .Y(n_712) );
AND2x2_ASAP7_75t_L g552 ( .A(n_524), .B(n_547), .Y(n_552) );
INVx1_ASAP7_75t_L g572 ( .A(n_524), .Y(n_572) );
AND2x2_ASAP7_75t_L g593 ( .A(n_524), .B(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g634 ( .A(n_524), .Y(n_634) );
INVx1_ASAP7_75t_L g650 ( .A(n_524), .Y(n_650) );
HB1xp67_ASAP7_75t_L g725 ( .A(n_524), .Y(n_725) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_528), .B(n_529), .Y(n_526) );
INVxp67_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_536), .B(n_638), .Y(n_679) );
OAI22xp5_ASAP7_75t_L g681 ( .A1(n_536), .A2(n_623), .B1(n_672), .B2(n_682), .Y(n_681) );
INVx1_ASAP7_75t_SL g536 ( .A(n_537), .Y(n_536) );
OAI211xp5_ASAP7_75t_SL g715 ( .A1(n_537), .A2(n_716), .B(n_718), .C(n_736), .Y(n_715) );
INVx2_ASAP7_75t_L g568 ( .A(n_538), .Y(n_568) );
AND2x2_ASAP7_75t_L g626 ( .A(n_538), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g637 ( .A(n_538), .B(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_539), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_542), .Y(n_539) );
AND2x2_ASAP7_75t_L g610 ( .A(n_540), .B(n_574), .Y(n_610) );
BUFx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g642 ( .A(n_541), .B(n_633), .Y(n_642) );
AND2x2_ASAP7_75t_L g661 ( .A(n_541), .B(n_575), .Y(n_661) );
AND2x4_ASAP7_75t_L g597 ( .A(n_542), .B(n_571), .Y(n_597) );
AND2x2_ASAP7_75t_L g735 ( .A(n_542), .B(n_711), .Y(n_735) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_547), .Y(n_542) );
BUFx6f_ASAP7_75t_L g564 ( .A(n_543), .Y(n_564) );
INVx1_ASAP7_75t_L g575 ( .A(n_543), .Y(n_575) );
INVx1_ASAP7_75t_L g674 ( .A(n_543), .Y(n_674) );
OR2x2_ASAP7_75t_L g565 ( .A(n_547), .B(n_551), .Y(n_565) );
AND2x2_ASAP7_75t_L g574 ( .A(n_547), .B(n_575), .Y(n_574) );
NOR2xp67_ASAP7_75t_L g594 ( .A(n_547), .B(n_595), .Y(n_594) );
OAI221xp5_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_553), .B1(n_563), .B2(n_566), .C(n_570), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
A2O1A1Ixp33_ASAP7_75t_L g570 ( .A1(n_550), .A2(n_571), .B(n_573), .C(n_576), .Y(n_570) );
AND2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
INVx1_ASAP7_75t_L g595 ( .A(n_551), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_551), .B(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_SL g678 ( .A(n_551), .B(n_572), .Y(n_678) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_551), .Y(n_685) );
AND2x2_ASAP7_75t_L g603 ( .A(n_552), .B(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g640 ( .A(n_552), .B(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_554), .B(n_562), .Y(n_553) );
INVx2_ASAP7_75t_L g631 ( .A(n_554), .Y(n_631) );
AOI222xp33_ASAP7_75t_L g680 ( .A1(n_554), .A2(n_564), .B1(n_681), .B2(n_683), .C1(n_684), .C2(n_686), .Y(n_680) );
AND2x2_ASAP7_75t_L g737 ( .A(n_554), .B(n_706), .Y(n_737) );
AND2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_561), .Y(n_554) );
INVx1_ASAP7_75t_L g627 ( .A(n_555), .Y(n_627) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x4_ASAP7_75t_L g579 ( .A(n_560), .B(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g665 ( .A(n_562), .B(n_599), .Y(n_665) );
AOI21xp33_ASAP7_75t_L g676 ( .A1(n_563), .A2(n_677), .B(n_679), .Y(n_676) );
OR2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
INVx2_ASAP7_75t_L g604 ( .A(n_564), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_564), .B(n_571), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_564), .B(n_717), .Y(n_716) );
INVx1_ASAP7_75t_SL g566 ( .A(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
INVx3_ASAP7_75t_L g630 ( .A(n_568), .Y(n_630) );
OR2x2_ASAP7_75t_L g682 ( .A(n_568), .B(n_604), .Y(n_682) );
AND2x2_ASAP7_75t_L g598 ( .A(n_569), .B(n_599), .Y(n_598) );
AND2x2_ASAP7_75t_L g636 ( .A(n_569), .B(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_569), .B(n_630), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_569), .B(n_626), .Y(n_652) );
AND2x2_ASAP7_75t_L g656 ( .A(n_569), .B(n_638), .Y(n_656) );
INVxp67_ASAP7_75t_L g588 ( .A(n_571), .Y(n_588) );
BUFx3_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
OAI22xp5_ASAP7_75t_L g645 ( .A1(n_573), .A2(n_646), .B1(n_651), .B2(n_652), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_573), .B(n_678), .Y(n_708) );
INVx1_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g694 ( .A(n_574), .B(n_685), .Y(n_694) );
AND2x2_ASAP7_75t_L g723 ( .A(n_574), .B(n_724), .Y(n_723) );
AND2x2_ASAP7_75t_L g728 ( .A(n_574), .B(n_678), .Y(n_728) );
INVx1_ASAP7_75t_L g641 ( .A(n_575), .Y(n_641) );
BUFx2_ASAP7_75t_L g647 ( .A(n_575), .Y(n_647) );
INVx1_ASAP7_75t_L g732 ( .A(n_576), .Y(n_732) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
NAND2x1p5_ASAP7_75t_L g583 ( .A(n_577), .B(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g608 ( .A(n_578), .Y(n_608) );
NOR2x1_ASAP7_75t_L g584 ( .A(n_579), .B(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g591 ( .A(n_579), .B(n_592), .Y(n_591) );
INVx2_ASAP7_75t_L g600 ( .A(n_579), .Y(n_600) );
INVx3_ASAP7_75t_L g638 ( .A(n_579), .Y(n_638) );
OR2x2_ASAP7_75t_L g704 ( .A(n_579), .B(n_705), .Y(n_704) );
AOI211xp5_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_586), .B(n_589), .C(n_601), .Y(n_581) );
AOI221xp5_ASAP7_75t_L g718 ( .A1(n_582), .A2(n_719), .B1(n_726), .B2(n_728), .C(n_729), .Y(n_718) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g589 ( .A(n_590), .B(n_596), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_592), .B(n_630), .Y(n_644) );
AND2x2_ASAP7_75t_L g686 ( .A(n_592), .B(n_626), .Y(n_686) );
INVx1_ASAP7_75t_SL g699 ( .A(n_593), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_593), .B(n_647), .Y(n_702) );
INVx1_ASAP7_75t_L g720 ( .A(n_594), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
AOI221xp5_ASAP7_75t_L g687 ( .A1(n_598), .A2(n_688), .B1(n_690), .B2(n_694), .C(n_695), .Y(n_687) );
AND2x2_ASAP7_75t_L g714 ( .A(n_599), .B(n_706), .Y(n_714) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g698 ( .A(n_600), .Y(n_698) );
AOI21xp33_ASAP7_75t_SL g601 ( .A1(n_602), .A2(n_605), .B(n_606), .Y(n_601) );
INVx1_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
OR2x2_ASAP7_75t_L g669 ( .A(n_604), .B(n_670), .Y(n_669) );
INVx2_ASAP7_75t_L g655 ( .A(n_605), .Y(n_655) );
INVx1_ASAP7_75t_L g683 ( .A(n_606), .Y(n_683) );
OR2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
O2A1O1Ixp33_ASAP7_75t_L g609 ( .A1(n_610), .A2(n_611), .B(n_614), .C(n_617), .Y(n_609) );
OAI31xp33_ASAP7_75t_L g736 ( .A1(n_610), .A2(n_648), .A3(n_735), .B(n_737), .Y(n_736) );
INVxp67_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g710 ( .A(n_613), .B(n_711), .Y(n_710) );
INVx1_ASAP7_75t_SL g731 ( .A(n_613), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_615), .B(n_630), .Y(n_658) );
INVx1_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
OR2x2_ASAP7_75t_L g733 ( .A(n_616), .B(n_630), .Y(n_733) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_625), .B1(n_629), .B2(n_632), .Y(n_620) );
NAND2xp33_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_624), .B(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g660 ( .A(n_624), .B(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g663 ( .A(n_624), .B(n_647), .Y(n_663) );
AND2x2_ASAP7_75t_L g717 ( .A(n_624), .B(n_712), .Y(n_717) );
AND2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_628), .Y(n_625) );
INVx1_ASAP7_75t_L g692 ( .A(n_628), .Y(n_692) );
NOR2xp67_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
OAI32xp33_ASAP7_75t_L g695 ( .A1(n_630), .A2(n_664), .A3(n_696), .B1(n_698), .B2(n_699), .Y(n_695) );
INVx1_ASAP7_75t_L g670 ( .A(n_633), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_633), .B(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g693 ( .A(n_637), .Y(n_693) );
O2A1O1Ixp33_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_642), .B(n_643), .C(n_645), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_641), .B(n_678), .Y(n_677) );
AOI221xp5_ASAP7_75t_L g653 ( .A1(n_642), .A2(n_654), .B1(n_655), .B2(n_656), .C(n_657), .Y(n_653) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g654 ( .A(n_652), .Y(n_654) );
OAI22xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_659), .B1(n_662), .B2(n_664), .Y(n_657) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NAND4xp25_ASAP7_75t_SL g719 ( .A(n_662), .B(n_720), .C(n_721), .D(n_722), .Y(n_719) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
NAND4xp25_ASAP7_75t_SL g666 ( .A(n_667), .B(n_680), .C(n_687), .D(n_700), .Y(n_666) );
O2A1O1Ixp33_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_671), .B(n_675), .C(n_676), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_SL g697 ( .A(n_673), .Y(n_697) );
INVx2_ASAP7_75t_L g721 ( .A(n_678), .Y(n_721) );
OR2x2_ASAP7_75t_L g730 ( .A(n_685), .B(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
OR2x2_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
AOI21xp5_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_703), .B(n_707), .Y(n_700) );
INVxp67_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
AND2x2_ASAP7_75t_L g726 ( .A(n_706), .B(n_727), .Y(n_726) );
AOI21xp33_ASAP7_75t_SL g707 ( .A1(n_708), .A2(n_709), .B(n_713), .Y(n_707) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
CKINVDCx16_ASAP7_75t_R g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
OAI22xp5_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_732), .B1(n_733), .B2(n_734), .Y(n_729) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_SL g747 ( .A(n_748), .Y(n_747) );
INVx3_ASAP7_75t_SL g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
NAND2xp33_ASAP7_75t_L g751 ( .A(n_752), .B(n_753), .Y(n_751) );
INVx1_ASAP7_75t_SL g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_SL g755 ( .A(n_756), .Y(n_755) );
endmodule