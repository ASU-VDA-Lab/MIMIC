module fake_jpeg_5062_n_225 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_225);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_225;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_32),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_41),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_32),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_39),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_40),
.B(n_42),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_32),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_25),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

AND2x2_ASAP7_75t_SL g46 ( 
.A(n_34),
.B(n_32),
.Y(n_46)
);

OR2x2_ASAP7_75t_SL g69 ( 
.A(n_46),
.B(n_68),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_31),
.B1(n_30),
.B2(n_24),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_49),
.A2(n_22),
.B1(n_17),
.B2(n_27),
.Y(n_71)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx2_ASAP7_75t_SL g79 ( 
.A(n_50),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_55),
.Y(n_73)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_58),
.Y(n_78)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_62),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_17),
.Y(n_61)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_61),
.Y(n_75)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_40),
.A2(n_19),
.B(n_24),
.C(n_30),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_63),
.A2(n_29),
.B(n_25),
.C(n_18),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_39),
.A2(n_31),
.B1(n_27),
.B2(n_33),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_65),
.A2(n_23),
.B(n_18),
.Y(n_87)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_20),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_33),
.Y(n_68)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_74),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_71),
.A2(n_77),
.B1(n_87),
.B2(n_13),
.Y(n_109)
);

NAND2x1_ASAP7_75t_SL g72 ( 
.A(n_46),
.B(n_32),
.Y(n_72)
);

OAI21xp33_ASAP7_75t_L g94 ( 
.A1(n_72),
.A2(n_85),
.B(n_62),
.Y(n_94)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_29),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_66),
.Y(n_108)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_47),
.A2(n_21),
.B(n_22),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_82),
.A2(n_52),
.B(n_14),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_68),
.B(n_21),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_83),
.B(n_88),
.Y(n_99)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_91),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_68),
.B(n_0),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_18),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_3),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_0),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_67),
.A2(n_20),
.B1(n_16),
.B2(n_2),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_89),
.A2(n_48),
.B1(n_50),
.B2(n_58),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_0),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_90),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_51),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_98),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_93),
.A2(n_103),
.B1(n_109),
.B2(n_111),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_94),
.Y(n_118)
);

OAI21xp33_ASAP7_75t_L g97 ( 
.A1(n_72),
.A2(n_1),
.B(n_2),
.Y(n_97)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_101),
.A2(n_85),
.B(n_83),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g102 ( 
.A(n_72),
.Y(n_102)
);

INVx4_ASAP7_75t_SL g121 ( 
.A(n_102),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_77),
.A2(n_48),
.B1(n_57),
.B2(n_53),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_110),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_69),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_106),
.B(n_82),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_88),
.A2(n_20),
.B(n_5),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_71),
.Y(n_130)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_4),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_69),
.A2(n_57),
.B1(n_53),
.B2(n_66),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_73),
.B(n_4),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_113),
.Y(n_133)
);

OAI32xp33_ASAP7_75t_L g113 ( 
.A1(n_76),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_87),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_120),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_76),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_119),
.A2(n_111),
.B(n_103),
.Y(n_140)
);

INVx13_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_125),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_124),
.A2(n_99),
.B(n_101),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g125 ( 
.A(n_113),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_126),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_73),
.C(n_80),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_89),
.C(n_81),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_129),
.A2(n_110),
.B(n_105),
.Y(n_137)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_75),
.Y(n_131)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_95),
.B(n_75),
.Y(n_132)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_132),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_142),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_137),
.A2(n_119),
.B(n_134),
.Y(n_168)
);

NOR4xp25_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_102),
.C(n_108),
.D(n_112),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_140),
.Y(n_157)
);

NOR2x1_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_107),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_141),
.A2(n_119),
.B1(n_135),
.B2(n_133),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_128),
.A2(n_93),
.B1(n_70),
.B2(n_74),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_80),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_145),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_100),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_146),
.B(n_154),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_122),
.B(n_78),
.Y(n_147)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_147),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_148),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_150),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_128),
.Y(n_153)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_153),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_91),
.C(n_78),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_118),
.A2(n_13),
.B1(n_15),
.B2(n_7),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_155),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_153),
.A2(n_134),
.B1(n_135),
.B2(n_133),
.Y(n_158)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_158),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_165),
.Y(n_175)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_166),
.B(n_167),
.Y(n_179)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_147),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_168),
.A2(n_173),
.B(n_141),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_120),
.Y(n_170)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_170),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_120),
.Y(n_172)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_172),
.Y(n_176)
);

OA21x2_ASAP7_75t_L g173 ( 
.A1(n_144),
.A2(n_125),
.B(n_130),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_180),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_145),
.Y(n_178)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_178),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_143),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_171),
.A2(n_149),
.B1(n_154),
.B2(n_151),
.Y(n_181)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_181),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_160),
.B(n_151),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_182),
.B(n_186),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_169),
.Y(n_183)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_183),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_159),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_185),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_137),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_140),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_173),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_183),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_189),
.A2(n_190),
.B(n_195),
.Y(n_204)
);

XOR2x2_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_157),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_187),
.B(n_168),
.C(n_163),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_174),
.C(n_178),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_196),
.Y(n_199)
);

AO21x1_ASAP7_75t_L g195 ( 
.A1(n_174),
.A2(n_171),
.B(n_173),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_198),
.B(n_176),
.Y(n_200)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_200),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_193),
.B(n_185),
.C(n_176),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_202),
.Y(n_209)
);

AOI31xp67_ASAP7_75t_SL g202 ( 
.A1(n_190),
.A2(n_155),
.A3(n_161),
.B(n_158),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_205),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_180),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_188),
.A2(n_161),
.B1(n_175),
.B2(n_150),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_206),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_204),
.A2(n_169),
.B1(n_192),
.B2(n_164),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_207),
.A2(n_211),
.B(n_210),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_203),
.A2(n_164),
.B1(n_115),
.B2(n_148),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_212),
.A2(n_179),
.B(n_136),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_189),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_213),
.B(n_126),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_205),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_214),
.B(n_216),
.Y(n_219)
);

FAx1_ASAP7_75t_SL g220 ( 
.A(n_215),
.B(n_209),
.CI(n_129),
.CON(n_220),
.SN(n_220)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_217),
.A2(n_218),
.B(n_211),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_146),
.Y(n_218)
);

MAJx2_ASAP7_75t_L g223 ( 
.A(n_220),
.B(n_221),
.C(n_116),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_142),
.C(n_195),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_222),
.B(n_223),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_90),
.Y(n_225)
);


endmodule