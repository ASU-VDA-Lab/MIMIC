module fake_netlist_6_1798_n_13163 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_127, n_125, n_77, n_106, n_92, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_135, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_13163);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_135;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_13163;

wire n_5643;
wire n_12335;
wire n_12949;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_801;
wire n_4452;
wire n_6566;
wire n_2576;
wire n_5172;
wire n_13045;
wire n_11173;
wire n_4649;
wire n_1674;
wire n_5315;
wire n_741;
wire n_10487;
wire n_6872;
wire n_1351;
wire n_5254;
wire n_11926;
wire n_6441;
wire n_8668;
wire n_1212;
wire n_208;
wire n_6806;
wire n_5362;
wire n_4251;
wire n_2157;
wire n_13146;
wire n_10587;
wire n_5019;
wire n_2332;
wire n_8713;
wire n_7111;
wire n_6141;
wire n_10960;
wire n_3849;
wire n_11111;
wire n_7933;
wire n_7967;
wire n_578;
wire n_5138;
wire n_10931;
wire n_4388;
wire n_4395;
wire n_6960;
wire n_1061;
wire n_3089;
wire n_8169;
wire n_12265;
wire n_9002;
wire n_9130;
wire n_783;
wire n_7180;
wire n_5653;
wire n_11574;
wire n_4978;
wire n_8604;
wire n_5409;
wire n_5301;
wire n_7263;
wire n_13125;
wire n_188;
wire n_1854;
wire n_3088;
wire n_8168;
wire n_3257;
wire n_1342;
wire n_4829;
wire n_5393;
wire n_1387;
wire n_3222;
wire n_7190;
wire n_7504;
wire n_677;
wire n_6126;
wire n_6725;
wire n_4699;
wire n_1151;
wire n_4686;
wire n_12322;
wire n_8899;
wire n_2317;
wire n_5524;
wire n_10236;
wire n_442;
wire n_5345;
wire n_11205;
wire n_11678;
wire n_11776;
wire n_8023;
wire n_11802;
wire n_12251;
wire n_10053;
wire n_1975;
wire n_11650;
wire n_1930;
wire n_3706;
wire n_5818;
wire n_8005;
wire n_8130;
wire n_2179;
wire n_8534;
wire n_5963;
wire n_12179;
wire n_5055;
wire n_1547;
wire n_12570;
wire n_9896;
wire n_11856;
wire n_11905;
wire n_3376;
wire n_4868;
wire n_10020;
wire n_893;
wire n_3801;
wire n_7116;
wire n_5267;
wire n_10202;
wire n_4249;
wire n_11536;
wire n_5950;
wire n_1192;
wire n_3564;
wire n_9104;
wire n_1844;
wire n_6999;
wire n_11046;
wire n_11079;
wire n_1555;
wire n_5548;
wire n_10283;
wire n_5057;
wire n_11065;
wire n_8339;
wire n_8272;
wire n_7161;
wire n_3030;
wire n_830;
wire n_7868;
wire n_5838;
wire n_5725;
wire n_6324;
wire n_447;
wire n_2838;
wire n_5229;
wire n_5325;
wire n_11051;
wire n_3427;
wire n_852;
wire n_11214;
wire n_5101;
wire n_2628;
wire n_3071;
wire n_7000;
wire n_8561;
wire n_11954;
wire n_7398;
wire n_2926;
wire n_1078;
wire n_544;
wire n_10392;
wire n_12882;
wire n_5900;
wire n_4273;
wire n_5545;
wire n_12617;
wire n_8411;
wire n_2321;
wire n_8499;
wire n_2019;
wire n_8236;
wire n_5102;
wire n_13137;
wire n_3345;
wire n_2074;
wire n_6882;
wire n_2919;
wire n_4501;
wire n_9626;
wire n_10775;
wire n_11163;
wire n_2129;
wire n_9526;
wire n_6325;
wire n_4724;
wire n_9840;
wire n_945;
wire n_5598;
wire n_7983;
wire n_10348;
wire n_10863;
wire n_12495;
wire n_9581;
wire n_10719;
wire n_4997;
wire n_2399;
wire n_11419;
wire n_9018;
wire n_4843;
wire n_12095;
wire n_1232;
wire n_8070;
wire n_7389;
wire n_4696;
wire n_6660;
wire n_9055;
wire n_4347;
wire n_11740;
wire n_5259;
wire n_6913;
wire n_8444;
wire n_10015;
wire n_10986;
wire n_7802;
wire n_6948;
wire n_5819;
wire n_2480;
wire n_7008;
wire n_3877;
wire n_12392;
wire n_3929;
wire n_8366;
wire n_9362;
wire n_1455;
wire n_8102;
wire n_11979;
wire n_3048;
wire n_7516;
wire n_7401;
wire n_7596;
wire n_6280;
wire n_6629;
wire n_12767;
wire n_5279;
wire n_2786;
wire n_5894;
wire n_10759;
wire n_8022;
wire n_5930;
wire n_9036;
wire n_9551;
wire n_10262;
wire n_8175;
wire n_8977;
wire n_9658;
wire n_5239;
wire n_567;
wire n_1781;
wire n_1971;
wire n_8953;
wire n_5354;
wire n_8426;
wire n_10239;
wire n_5332;
wire n_9962;
wire n_2004;
wire n_1106;
wire n_4814;
wire n_953;
wire n_3979;
wire n_5908;
wire n_10373;
wire n_3077;
wire n_2873;
wire n_11104;
wire n_3452;
wire n_8913;
wire n_9525;
wire n_3107;
wire n_10816;
wire n_9725;
wire n_155;
wire n_4956;
wire n_11537;
wire n_12707;
wire n_454;
wire n_7686;
wire n_1421;
wire n_3664;
wire n_6914;
wire n_1936;
wire n_5337;
wire n_10335;
wire n_11301;
wire n_5129;
wire n_12424;
wire n_5420;
wire n_1660;
wire n_5070;
wire n_10381;
wire n_6243;
wire n_3047;
wire n_4414;
wire n_6585;
wire n_713;
wire n_11703;
wire n_11699;
wire n_1400;
wire n_2625;
wire n_4646;
wire n_6374;
wire n_2843;
wire n_7651;
wire n_11543;
wire n_10947;
wire n_6628;
wire n_8125;
wire n_3760;
wire n_6015;
wire n_11261;
wire n_10226;
wire n_1560;
wire n_4262;
wire n_734;
wire n_1088;
wire n_6526;
wire n_1894;
wire n_7956;
wire n_7369;
wire n_6570;
wire n_8556;
wire n_7196;
wire n_3347;
wire n_10767;
wire n_5136;
wire n_907;
wire n_8040;
wire n_11821;
wire n_5638;
wire n_13121;
wire n_9100;
wire n_4110;
wire n_6784;
wire n_1658;
wire n_12107;
wire n_10755;
wire n_4950;
wire n_10868;
wire n_9067;
wire n_10161;
wire n_9842;
wire n_4729;
wire n_4268;
wire n_11447;
wire n_6323;
wire n_9614;
wire n_10682;
wire n_6110;
wire n_1967;
wire n_11684;
wire n_3999;
wire n_12652;
wire n_3928;
wire n_6371;
wire n_8079;
wire n_10699;
wire n_2613;
wire n_3535;
wire n_4751;
wire n_8595;
wire n_7846;
wire n_2708;
wire n_1648;
wire n_9400;
wire n_5151;
wire n_1911;
wire n_8142;
wire n_11627;
wire n_2011;
wire n_5684;
wire n_8598;
wire n_13139;
wire n_10022;
wire n_5729;
wire n_7256;
wire n_281;
wire n_6404;
wire n_12209;
wire n_7331;
wire n_7856;
wire n_7774;
wire n_564;
wire n_5680;
wire n_6674;
wire n_9680;
wire n_6148;
wire n_6951;
wire n_11659;
wire n_7625;
wire n_279;
wire n_686;
wire n_4102;
wire n_1641;
wire n_3871;
wire n_9106;
wire n_12775;
wire n_2735;
wire n_4662;
wire n_8869;
wire n_7863;
wire n_4671;
wire n_6989;
wire n_3959;
wire n_2268;
wire n_8381;
wire n_1367;
wire n_5504;
wire n_1336;
wire n_5522;
wire n_5828;
wire n_7342;
wire n_4314;
wire n_9520;
wire n_2080;
wire n_8958;
wire n_12833;
wire n_323;
wire n_5099;
wire n_12090;
wire n_6896;
wire n_7770;
wire n_10606;
wire n_8421;
wire n_11164;
wire n_7623;
wire n_6968;
wire n_7217;
wire n_1381;
wire n_331;
wire n_1699;
wire n_2093;
wire n_12371;
wire n_4296;
wire n_10114;
wire n_12203;
wire n_10357;
wire n_7147;
wire n_2770;
wire n_8115;
wire n_608;
wire n_2101;
wire n_4507;
wire n_8389;
wire n_9398;
wire n_5902;
wire n_11497;
wire n_512;
wire n_3484;
wire n_12359;
wire n_4677;
wire n_792;
wire n_12915;
wire n_5063;
wire n_6196;
wire n_9037;
wire n_1328;
wire n_2917;
wire n_13149;
wire n_2616;
wire n_5275;
wire n_5306;
wire n_12548;
wire n_12742;
wire n_3923;
wire n_9042;
wire n_11768;
wire n_3900;
wire n_8412;
wire n_9267;
wire n_3488;
wire n_939;
wire n_2811;
wire n_3732;
wire n_6485;
wire n_8987;
wire n_11805;
wire n_10177;
wire n_6107;
wire n_9652;
wire n_2832;
wire n_4226;
wire n_5493;
wire n_1762;
wire n_8849;
wire n_11944;
wire n_9059;
wire n_1910;
wire n_1075;
wire n_3980;
wire n_2998;
wire n_5346;
wire n_4366;
wire n_3446;
wire n_5252;
wire n_5309;
wire n_7796;
wire n_237;
wire n_6282;
wire n_6863;
wire n_6994;
wire n_12770;
wire n_1895;
wire n_10012;
wire n_4294;
wire n_12985;
wire n_4698;
wire n_4445;
wire n_13013;
wire n_4810;
wire n_7564;
wire n_11635;
wire n_3859;
wire n_2692;
wire n_175;
wire n_9446;
wire n_11129;
wire n_12951;
wire n_10204;
wire n_6768;
wire n_9453;
wire n_6383;
wire n_7234;
wire n_3914;
wire n_4456;
wire n_8119;
wire n_10296;
wire n_3397;
wire n_8641;
wire n_11637;
wire n_12988;
wire n_3575;
wire n_8151;
wire n_8118;
wire n_12393;
wire n_9718;
wire n_9128;
wire n_2469;
wire n_10281;
wire n_9038;
wire n_9872;
wire n_10310;
wire n_11139;
wire n_8748;
wire n_3927;
wire n_8436;
wire n_5452;
wire n_12685;
wire n_6794;
wire n_3888;
wire n_6151;
wire n_8718;
wire n_7110;
wire n_764;
wire n_5476;
wire n_2764;
wire n_12831;
wire n_9935;
wire n_2895;
wire n_6431;
wire n_8659;
wire n_6990;
wire n_733;
wire n_2922;
wire n_8223;
wire n_3882;
wire n_4856;
wire n_10097;
wire n_3492;
wire n_4369;
wire n_2068;
wire n_9135;
wire n_7849;
wire n_8915;
wire n_12667;
wire n_4331;
wire n_7297;
wire n_9866;
wire n_10018;
wire n_4972;
wire n_1290;
wire n_4993;
wire n_7298;
wire n_5536;
wire n_9129;
wire n_9858;
wire n_10141;
wire n_2072;
wire n_12427;
wire n_1354;
wire n_7533;
wire n_586;
wire n_423;
wire n_7221;
wire n_4375;
wire n_1701;
wire n_10656;
wire n_6575;
wire n_6055;
wire n_8727;
wire n_8224;
wire n_2678;
wire n_11295;
wire n_3935;
wire n_5130;
wire n_4291;
wire n_11662;
wire n_5532;
wire n_5897;
wire n_1726;
wire n_8246;
wire n_4613;
wire n_8952;
wire n_13014;
wire n_2434;
wire n_9070;
wire n_2878;
wire n_11708;
wire n_3012;
wire n_3875;
wire n_10266;
wire n_5609;
wire n_1167;
wire n_2428;
wire n_4717;
wire n_10827;
wire n_10897;
wire n_4877;
wire n_3247;
wire n_871;
wire n_5922;
wire n_210;
wire n_10449;
wire n_7569;
wire n_2641;
wire n_7734;
wire n_7062;
wire n_7823;
wire n_7861;
wire n_9477;
wire n_5658;
wire n_4731;
wire n_8955;
wire n_12172;
wire n_12147;
wire n_12923;
wire n_3052;
wire n_178;
wire n_7039;
wire n_355;
wire n_8577;
wire n_12384;
wire n_11349;
wire n_8594;
wire n_5046;
wire n_8428;
wire n_9829;
wire n_2749;
wire n_11260;
wire n_3298;
wire n_8848;
wire n_12825;
wire n_2254;
wire n_5058;
wire n_10685;
wire n_1926;
wire n_11351;
wire n_3273;
wire n_4467;
wire n_12083;
wire n_7077;
wire n_12014;
wire n_1747;
wire n_195;
wire n_5667;
wire n_780;
wire n_8259;
wire n_12540;
wire n_10607;
wire n_2624;
wire n_5865;
wire n_12249;
wire n_8349;
wire n_6836;
wire n_2350;
wire n_5042;
wire n_5305;
wire n_11998;
wire n_4681;
wire n_8164;
wire n_4072;
wire n_10628;
wire n_4752;
wire n_4220;
wire n_835;
wire n_928;
wire n_5281;
wire n_11775;
wire n_8776;
wire n_7905;
wire n_9143;
wire n_8287;
wire n_2092;
wire n_10256;
wire n_7753;
wire n_10368;
wire n_1654;
wire n_6771;
wire n_10769;
wire n_7950;
wire n_9947;
wire n_1750;
wire n_1462;
wire n_9088;
wire n_8607;
wire n_2514;
wire n_10138;
wire n_12117;
wire n_604;
wire n_11706;
wire n_6248;
wire n_11800;
wire n_10183;
wire n_10375;
wire n_6952;
wire n_10452;
wire n_5314;
wire n_1588;
wire n_6795;
wire n_11464;
wire n_7806;
wire n_3942;
wire n_3997;
wire n_12960;
wire n_13033;
wire n_11642;
wire n_2468;
wire n_4381;
wire n_11143;
wire n_7595;
wire n_5144;
wire n_7648;
wire n_515;
wire n_2096;
wire n_3968;
wire n_10383;
wire n_4466;
wire n_4418;
wire n_11074;
wire n_6831;
wire n_8066;
wire n_3434;
wire n_4510;
wire n_6776;
wire n_12131;
wire n_12851;
wire n_5795;
wire n_11934;
wire n_12349;
wire n_4473;
wire n_6043;
wire n_5552;
wire n_7452;
wire n_5226;
wire n_9269;
wire n_10320;
wire n_6715;
wire n_514;
wire n_6714;
wire n_687;
wire n_11308;
wire n_890;
wire n_7677;
wire n_10903;
wire n_5457;
wire n_8416;
wire n_10396;
wire n_2812;
wire n_190;
wire n_4518;
wire n_10724;
wire n_8404;
wire n_8997;
wire n_6584;
wire n_11084;
wire n_9988;
wire n_1709;
wire n_7009;
wire n_8453;
wire n_10693;
wire n_12740;
wire n_2393;
wire n_2657;
wire n_9113;
wire n_7149;
wire n_5291;
wire n_2921;
wire n_2136;
wire n_10363;
wire n_2409;
wire n_2252;
wire n_3237;
wire n_949;
wire n_8949;
wire n_10831;
wire n_3500;
wire n_3834;
wire n_9131;
wire n_11553;
wire n_10517;
wire n_12578;
wire n_12795;
wire n_4589;
wire n_2075;
wire n_10323;
wire n_12194;
wire n_2972;
wire n_10842;
wire n_3542;
wire n_7519;
wire n_7400;
wire n_10876;
wire n_2763;
wire n_11511;
wire n_2762;
wire n_9137;
wire n_11180;
wire n_9724;
wire n_11146;
wire n_9281;
wire n_3192;
wire n_8995;
wire n_10883;
wire n_760;
wire n_10101;
wire n_1546;
wire n_9393;
wire n_4394;
wire n_6581;
wire n_12709;
wire n_2279;
wire n_161;
wire n_6010;
wire n_1296;
wire n_3352;
wire n_8711;
wire n_3073;
wire n_7013;
wire n_12771;
wire n_5343;
wire n_12125;
wire n_12505;
wire n_2150;
wire n_1294;
wire n_3696;
wire n_1420;
wire n_4082;
wire n_7290;
wire n_12278;
wire n_595;
wire n_1779;
wire n_524;
wire n_10820;
wire n_4921;
wire n_9687;
wire n_1858;
wire n_4329;
wire n_5135;
wire n_7303;
wire n_3021;
wire n_6616;
wire n_8306;
wire n_10123;
wire n_10781;
wire n_7488;
wire n_2558;
wire n_7315;
wire n_9886;
wire n_10651;
wire n_9426;
wire n_8887;
wire n_1164;
wire n_4697;
wire n_4288;
wire n_4289;
wire n_11866;
wire n_3763;
wire n_6185;
wire n_2712;
wire n_11450;
wire n_12522;
wire n_5529;
wire n_3733;
wire n_7889;
wire n_10943;
wire n_12344;
wire n_6042;
wire n_9102;
wire n_1487;
wire n_11526;
wire n_9578;
wire n_3614;
wire n_874;
wire n_382;
wire n_5183;
wire n_13109;
wire n_8500;
wire n_7438;
wire n_2145;
wire n_7337;
wire n_7268;
wire n_11851;
wire n_898;
wire n_4964;
wire n_9489;
wire n_12804;
wire n_5957;
wire n_6965;
wire n_12116;
wire n_10728;
wire n_4228;
wire n_3423;
wire n_6357;
wire n_925;
wire n_1932;
wire n_1101;
wire n_9144;
wire n_10094;
wire n_6800;
wire n_10084;
wire n_4636;
wire n_10468;
wire n_7461;
wire n_8285;
wire n_4322;
wire n_10655;
wire n_3644;
wire n_9797;
wire n_6955;
wire n_8483;
wire n_1249;
wire n_4946;
wire n_2706;
wire n_4767;
wire n_4287;
wire n_2693;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_9521;
wire n_8332;
wire n_9478;
wire n_1451;
wire n_9932;
wire n_13040;
wire n_320;
wire n_639;
wire n_963;
wire n_2767;
wire n_11370;
wire n_6509;
wire n_7278;
wire n_4576;
wire n_11253;
wire n_7454;
wire n_11379;
wire n_10670;
wire n_5929;
wire n_12861;
wire n_9020;
wire n_4615;
wire n_5787;
wire n_11981;
wire n_1139;
wire n_3179;
wire n_1018;
wire n_3400;
wire n_9895;
wire n_1521;
wire n_8741;
wire n_12918;
wire n_1366;
wire n_4000;
wire n_9351;
wire n_11585;
wire n_5445;
wire n_2897;
wire n_13140;
wire n_4389;
wire n_3970;
wire n_5342;
wire n_5501;
wire n_6839;
wire n_7232;
wire n_4345;
wire n_7377;
wire n_996;
wire n_532;
wire n_173;
wire n_6646;
wire n_8648;
wire n_12388;
wire n_1376;
wire n_12102;
wire n_9189;
wire n_413;
wire n_4664;
wire n_2170;
wire n_4156;
wire n_948;
wire n_7098;
wire n_7069;
wire n_12560;
wire n_7904;
wire n_11691;
wire n_6033;
wire n_977;
wire n_11541;
wire n_536;
wire n_3158;
wire n_1788;
wire n_8851;
wire n_8921;
wire n_4873;
wire n_9410;
wire n_9801;
wire n_2643;
wire n_5748;
wire n_3782;
wire n_9356;
wire n_12865;
wire n_8773;
wire n_6097;
wire n_6369;
wire n_10712;
wire n_1835;
wire n_8394;
wire n_3470;
wire n_11155;
wire n_5076;
wire n_581;
wire n_5870;
wire n_4713;
wire n_9175;
wire n_7093;
wire n_4098;
wire n_6508;
wire n_5026;
wire n_4476;
wire n_7168;
wire n_432;
wire n_3700;
wire n_12013;
wire n_11835;
wire n_4995;
wire n_7542;
wire n_7970;
wire n_7091;
wire n_3166;
wire n_10959;
wire n_3104;
wire n_6809;
wire n_11233;
wire n_3435;
wire n_842;
wire n_5636;
wire n_2239;
wire n_7840;
wire n_10972;
wire n_4310;
wire n_6359;
wire n_7782;
wire n_1432;
wire n_12231;
wire n_5212;
wire n_10024;
wire n_10945;
wire n_989;
wire n_8800;
wire n_10845;
wire n_7080;
wire n_2689;
wire n_1473;
wire n_6636;
wire n_5286;
wire n_2191;
wire n_8229;
wire n_1246;
wire n_4528;
wire n_8410;
wire n_5811;
wire n_899;
wire n_10711;
wire n_7739;
wire n_7624;
wire n_1035;
wire n_4914;
wire n_6766;
wire n_4939;
wire n_7629;
wire n_499;
wire n_1426;
wire n_3418;
wire n_705;
wire n_9735;
wire n_9186;
wire n_10818;
wire n_1004;
wire n_1529;
wire n_5530;
wire n_2473;
wire n_5397;
wire n_10624;
wire n_4634;
wire n_12552;
wire n_2069;
wire n_11069;
wire n_2362;
wire n_4096;
wire n_2539;
wire n_2698;
wire n_4123;
wire n_5595;
wire n_9941;
wire n_7003;
wire n_11951;
wire n_12222;
wire n_11900;
wire n_3119;
wire n_5427;
wire n_10788;
wire n_3735;
wire n_2297;
wire n_11369;
wire n_4379;
wire n_10563;
wire n_486;
wire n_8810;
wire n_5388;
wire n_4718;
wire n_9802;
wire n_1448;
wire n_5901;
wire n_6538;
wire n_5962;
wire n_3631;
wire n_5599;
wire n_8107;
wire n_648;
wire n_11108;
wire n_7010;
wire n_9728;
wire n_12883;
wire n_11004;
wire n_12992;
wire n_2445;
wire n_5324;
wire n_2057;
wire n_6519;
wire n_2103;
wire n_8983;
wire n_10422;
wire n_11686;
wire n_3770;
wire n_9818;
wire n_2772;
wire n_7219;
wire n_6530;
wire n_9662;
wire n_12896;
wire n_4440;
wire n_8774;
wire n_4402;
wire n_10566;
wire n_927;
wire n_10178;
wire n_5052;
wire n_7299;
wire n_12367;
wire n_4541;
wire n_12104;
wire n_5009;
wire n_4872;
wire n_929;
wire n_6402;
wire n_12469;
wire n_9936;
wire n_12563;
wire n_4551;
wire n_2857;
wire n_6195;
wire n_13132;
wire n_7326;
wire n_7243;
wire n_9530;
wire n_10115;
wire n_6609;
wire n_5326;
wire n_7471;
wire n_10455;
wire n_11778;
wire n_1183;
wire n_7067;
wire n_12793;
wire n_4627;
wire n_4079;
wire n_2494;
wire n_5300;
wire n_9909;
wire n_11393;
wire n_8620;
wire n_8691;
wire n_12406;
wire n_3342;
wire n_6748;
wire n_7741;
wire n_998;
wire n_5035;
wire n_9466;
wire n_717;
wire n_7790;
wire n_11719;
wire n_6149;
wire n_10052;
wire n_10109;
wire n_1383;
wire n_7484;
wire n_3390;
wire n_3656;
wire n_7002;
wire n_1424;
wire n_10448;
wire n_6414;
wire n_11196;
wire n_1000;
wire n_11963;
wire n_12428;
wire n_8424;
wire n_9571;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_7528;
wire n_8026;
wire n_9470;
wire n_3810;
wire n_552;
wire n_4798;
wire n_9638;
wire n_2532;
wire n_1388;
wire n_3006;
wire n_216;
wire n_10265;
wire n_8174;
wire n_12655;
wire n_7941;
wire n_912;
wire n_11175;
wire n_5010;
wire n_11483;
wire n_2296;
wire n_3633;
wire n_5352;
wire n_11995;
wire n_5089;
wire n_2849;
wire n_11371;
wire n_1201;
wire n_1398;
wire n_884;
wire n_10040;
wire n_5394;
wire n_4592;
wire n_9405;
wire n_1395;
wire n_6264;
wire n_2199;
wire n_2661;
wire n_8861;
wire n_731;
wire n_5359;
wire n_8644;
wire n_1955;
wire n_8907;
wire n_931;
wire n_474;
wire n_312;
wire n_1791;
wire n_12304;
wire n_11080;
wire n_10984;
wire n_958;
wire n_5137;
wire n_6902;
wire n_3331;
wire n_5104;
wire n_10100;
wire n_1897;
wire n_2064;
wire n_7117;
wire n_13138;
wire n_9894;
wire n_5741;
wire n_8324;
wire n_2773;
wire n_6205;
wire n_9441;
wire n_6380;
wire n_10906;
wire n_7478;
wire n_7913;
wire n_12001;
wire n_5405;
wire n_7136;
wire n_6754;
wire n_7883;
wire n_5288;
wire n_7456;
wire n_589;
wire n_3606;
wire n_1310;
wire n_12692;
wire n_819;
wire n_1334;
wire n_3591;
wire n_7939;
wire n_2788;
wire n_964;
wire n_8503;
wire n_9612;
wire n_4756;
wire n_8196;
wire n_10380;
wire n_10790;
wire n_6449;
wire n_2797;
wire n_6723;
wire n_7458;
wire n_9108;
wire n_9787;
wire n_10846;
wire n_7436;
wire n_6440;
wire n_4746;
wire n_6461;
wire n_3892;
wire n_4970;
wire n_4069;
wire n_211;
wire n_2748;
wire n_8446;
wire n_5194;
wire n_9376;
wire n_9786;
wire n_1834;
wire n_9033;
wire n_2331;
wire n_12933;
wire n_2292;
wire n_7435;
wire n_12908;
wire n_3441;
wire n_9537;
wire n_11297;
wire n_3534;
wire n_6997;
wire n_10509;
wire n_5952;
wire n_3964;
wire n_12996;
wire n_2416;
wire n_311;
wire n_5947;
wire n_8923;
wire n_12643;
wire n_1877;
wire n_3944;
wire n_6736;
wire n_6124;
wire n_7685;
wire n_7363;
wire n_8192;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_5985;
wire n_8197;
wire n_556;
wire n_2209;
wire n_3605;
wire n_6622;
wire n_11946;
wire n_9443;
wire n_1602;
wire n_11521;
wire n_9996;
wire n_11742;
wire n_4633;
wire n_6891;
wire n_7800;
wire n_10031;
wire n_3306;
wire n_12827;
wire n_12678;
wire n_276;
wire n_9115;
wire n_3026;
wire n_12235;
wire n_221;
wire n_4584;
wire n_3090;
wire n_5232;
wire n_11833;
wire n_3724;
wire n_7663;
wire n_4276;
wire n_11897;
wire n_12204;
wire n_10898;
wire n_5116;
wire n_2990;
wire n_3847;
wire n_1773;
wire n_5001;
wire n_2552;
wire n_1053;
wire n_5176;
wire n_7443;
wire n_7747;
wire n_9779;
wire n_9938;
wire n_11285;
wire n_8082;
wire n_12098;
wire n_4428;
wire n_8730;
wire n_1533;
wire n_3323;
wire n_7917;
wire n_7261;
wire n_266;
wire n_9023;
wire n_12579;
wire n_6528;
wire n_2274;
wire n_9203;
wire n_9977;
wire n_7532;
wire n_8051;
wire n_9613;
wire n_11818;
wire n_5761;
wire n_518;
wire n_9242;
wire n_6773;
wire n_4618;
wire n_12611;
wire n_7375;
wire n_4679;
wire n_1745;
wire n_914;
wire n_3479;
wire n_11262;
wire n_4496;
wire n_7968;
wire n_6382;
wire n_7455;
wire n_317;
wire n_12713;
wire n_12880;
wire n_13144;
wire n_4805;
wire n_1679;
wire n_8651;
wire n_3454;
wire n_2160;
wire n_9141;
wire n_5760;
wire n_6885;
wire n_9201;
wire n_10732;
wire n_2146;
wire n_6531;
wire n_10952;
wire n_2131;
wire n_488;
wire n_10851;
wire n_11027;
wire n_11852;
wire n_10660;
wire n_7430;
wire n_5472;
wire n_3547;
wire n_10221;
wire n_9559;
wire n_9299;
wire n_8377;
wire n_11803;
wire n_9937;
wire n_5679;
wire n_11162;
wire n_7912;
wire n_9913;
wire n_2575;
wire n_5100;
wire n_9286;
wire n_8015;
wire n_5973;
wire n_7921;
wire n_10044;
wire n_7728;
wire n_4410;
wire n_1933;
wire n_8281;
wire n_10819;
wire n_1179;
wire n_324;
wire n_3816;
wire n_4807;
wire n_8842;
wire n_4411;
wire n_9184;
wire n_3214;
wire n_1243;
wire n_9704;
wire n_301;
wire n_2928;
wire n_5166;
wire n_9046;
wire n_6339;
wire n_1917;
wire n_8024;
wire n_1580;
wire n_7730;
wire n_12562;
wire n_8814;
wire n_8530;
wire n_11428;
wire n_2822;
wire n_11592;
wire n_4180;
wire n_9193;
wire n_1281;
wire n_8467;
wire n_11677;
wire n_7281;
wire n_3109;
wire n_9717;
wire n_3354;
wire n_2572;
wire n_7711;
wire n_1520;
wire n_3126;
wire n_11090;
wire n_8984;
wire n_3663;
wire n_2863;
wire n_1419;
wire n_3299;
wire n_5688;
wire n_6417;
wire n_9290;
wire n_351;
wire n_5740;
wire n_259;
wire n_1731;
wire n_5820;
wire n_5648;
wire n_2135;
wire n_5745;
wire n_4707;
wire n_1645;
wire n_1832;
wire n_4676;
wire n_9403;
wire n_10996;
wire n_9875;
wire n_5180;
wire n_8956;
wire n_6763;
wire n_858;
wire n_2049;
wire n_5182;
wire n_7858;
wire n_11561;
wire n_8676;
wire n_956;
wire n_5534;
wire n_8003;
wire n_663;
wire n_4880;
wire n_8785;
wire n_9853;
wire n_3566;
wire n_7448;
wire n_6542;
wire n_2781;
wire n_4126;
wire n_410;
wire n_2829;
wire n_1696;
wire n_3845;
wire n_6556;
wire n_1594;
wire n_8692;
wire n_664;
wire n_1869;
wire n_7230;
wire n_6889;
wire n_9183;
wire n_3804;
wire n_7989;
wire n_4207;
wire n_9778;
wire n_5196;
wire n_6199;
wire n_2016;
wire n_9823;
wire n_5171;
wire n_12937;
wire n_10698;
wire n_10852;
wire n_4470;
wire n_6726;
wire n_12374;
wire n_9529;
wire n_580;
wire n_4813;
wire n_5542;
wire n_1030;
wire n_3901;
wire n_1937;
wire n_7011;
wire n_465;
wire n_8998;
wire n_1790;
wire n_10538;
wire n_5261;
wire n_12848;
wire n_11425;
wire n_12158;
wire n_10870;
wire n_4014;
wire n_4704;
wire n_11066;
wire n_341;
wire n_1744;
wire n_828;
wire n_10315;
wire n_2142;
wire n_4252;
wire n_607;
wire n_9123;
wire n_4028;
wire n_6576;
wire n_6471;
wire n_2448;
wire n_8906;
wire n_5949;
wire n_11455;
wire n_4048;
wire n_4596;
wire n_12368;
wire n_4444;
wire n_5255;
wire n_3756;
wire n_8482;
wire n_6478;
wire n_7952;
wire n_11867;
wire n_3406;
wire n_820;
wire n_951;
wire n_6100;
wire n_12796;
wire n_6516;
wire n_952;
wire n_3919;
wire n_8462;
wire n_6977;
wire n_9380;
wire n_10062;
wire n_7660;
wire n_6915;
wire n_12529;
wire n_2263;
wire n_12103;
wire n_7834;
wire n_11716;
wire n_5185;
wire n_6911;
wire n_8409;
wire n_6599;
wire n_974;
wire n_8979;
wire n_6522;
wire n_4952;
wire n_2656;
wire n_5023;
wire n_2375;
wire n_5906;
wire n_1934;
wire n_8429;
wire n_8930;
wire n_10514;
wire n_628;
wire n_5660;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_7890;
wire n_12785;
wire n_3973;
wire n_2756;
wire n_11950;
wire n_7245;
wire n_5334;
wire n_6024;
wire n_9347;
wire n_807;
wire n_4761;
wire n_6675;
wire n_6270;
wire n_12461;
wire n_1275;
wire n_2884;
wire n_6808;
wire n_485;
wire n_1510;
wire n_7620;
wire n_11415;
wire n_11886;
wire n_7265;
wire n_7986;
wire n_5783;
wire n_7006;
wire n_6931;
wire n_6207;
wire n_3120;
wire n_5821;
wire n_6245;
wire n_6079;
wire n_7948;
wire n_3797;
wire n_238;
wire n_9082;
wire n_10925;
wire n_2024;
wire n_1595;
wire n_4770;
wire n_202;
wire n_9879;
wire n_1749;
wire n_11158;
wire n_3474;
wire n_9861;
wire n_11390;
wire n_6963;
wire n_8685;
wire n_2549;
wire n_4690;
wire n_11669;
wire n_1669;
wire n_1024;
wire n_3864;
wire n_8264;
wire n_5556;
wire n_4932;
wire n_8250;
wire n_8492;
wire n_7381;
wire n_12078;
wire n_10601;
wire n_5456;
wire n_9158;
wire n_248;
wire n_2302;
wire n_8135;
wire n_10618;
wire n_1667;
wire n_9594;
wire n_7837;
wire n_9832;
wire n_7717;
wire n_9518;
wire n_8445;
wire n_1037;
wire n_6427;
wire n_6580;
wire n_5143;
wire n_9898;
wire n_3592;
wire n_11739;
wire n_468;
wire n_5500;
wire n_10497;
wire n_4230;
wire n_6412;
wire n_9445;
wire n_2637;
wire n_1639;
wire n_7627;
wire n_183;
wire n_9803;
wire n_3967;
wire n_7601;
wire n_6437;
wire n_8298;
wire n_3195;
wire n_466;
wire n_2526;
wire n_6346;
wire n_4274;
wire n_5215;
wire n_7860;
wire n_8408;
wire n_12639;
wire n_3277;
wire n_2548;
wire n_5386;
wire n_991;
wire n_10661;
wire n_7335;
wire n_4189;
wire n_9815;
wire n_8895;
wire n_9495;
wire n_3817;
wire n_10028;
wire n_7811;
wire n_340;
wire n_13158;
wire n_1108;
wire n_11676;
wire n_11044;
wire n_11771;
wire n_12266;
wire n_3659;
wire n_2559;
wire n_2595;
wire n_2177;
wire n_12175;
wire n_5003;
wire n_10512;
wire n_11384;
wire n_4827;
wire n_1601;
wire n_12287;
wire n_1960;
wire n_2694;
wire n_11679;
wire n_8450;
wire n_3648;
wire n_8273;
wire n_1686;
wire n_9867;
wire n_6059;
wire n_7499;
wire n_12353;
wire n_3042;
wire n_6065;
wire n_9688;
wire n_9761;
wire n_7292;
wire n_12398;
wire n_5094;
wire n_4610;
wire n_10967;
wire n_9087;
wire n_4472;
wire n_5433;
wire n_7870;
wire n_9043;
wire n_6075;
wire n_12991;
wire n_3228;
wire n_3657;
wire n_7397;
wire n_3081;
wire n_10789;
wire n_11134;
wire n_12705;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_6117;
wire n_7977;
wire n_8886;
wire n_12847;
wire n_10434;
wire n_7211;
wire n_12869;
wire n_13047;
wire n_10933;
wire n_11828;
wire n_8312;
wire n_5618;
wire n_6781;
wire n_6861;
wire n_12326;
wire n_1586;
wire n_7847;
wire n_8506;
wire n_2264;
wire n_3464;
wire n_6494;
wire n_380;
wire n_6133;
wire n_3723;
wire n_11548;
wire n_13041;
wire n_1190;
wire n_13154;
wire n_8963;
wire n_12404;
wire n_7822;
wire n_397;
wire n_4380;
wire n_6453;
wire n_5978;
wire n_11606;
wire n_11889;
wire n_9307;
wire n_4990;
wire n_5247;
wire n_4996;
wire n_6127;
wire n_10762;
wire n_11342;
wire n_4398;
wire n_2498;
wire n_11452;
wire n_11362;
wire n_8078;
wire n_7785;
wire n_6217;
wire n_4515;
wire n_1891;
wire n_5031;
wire n_1213;
wire n_6006;
wire n_2235;
wire n_10797;
wire n_11266;
wire n_4193;
wire n_7289;
wire n_3570;
wire n_12309;
wire n_7926;
wire n_5082;
wire n_6598;
wire n_7399;
wire n_1673;
wire n_5338;
wire n_3828;
wire n_12479;
wire n_172;
wire n_7354;
wire n_8352;
wire n_12502;
wire n_2392;
wire n_3424;
wire n_4131;
wire n_10360;
wire n_239;
wire n_7960;
wire n_9450;
wire n_2298;
wire n_2326;
wire n_1539;
wire n_490;
wire n_3594;
wire n_5689;
wire n_7482;
wire n_1043;
wire n_12912;
wire n_10312;
wire n_4090;
wire n_12211;
wire n_6115;
wire n_4165;
wire n_12454;
wire n_8143;
wire n_2305;
wire n_2120;
wire n_4626;
wire n_9223;
wire n_10480;
wire n_6048;
wire n_4144;
wire n_6416;
wire n_2964;
wire n_10131;
wire n_352;
wire n_12537;
wire n_6838;
wire n_10068;
wire n_6867;
wire n_9693;
wire n_11988;
wire n_12600;
wire n_12921;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_5931;
wire n_2371;
wire n_6139;
wire n_1361;
wire n_11957;
wire n_10633;
wire n_12133;
wire n_662;
wire n_6256;
wire n_7965;
wire n_3262;
wire n_6613;
wire n_11438;
wire n_11244;
wire n_4008;
wire n_12919;
wire n_3356;
wire n_5221;
wire n_10273;
wire n_5641;
wire n_1642;
wire n_12215;
wire n_11416;
wire n_10209;
wire n_3210;
wire n_6361;
wire n_937;
wire n_9880;
wire n_4689;
wire n_8183;
wire n_1682;
wire n_11348;
wire n_4547;
wire n_11245;
wire n_9685;
wire n_6085;
wire n_7474;
wire n_11169;
wire n_11685;
wire n_5731;
wire n_12422;
wire n_12467;
wire n_11607;
wire n_8650;
wire n_6329;
wire n_6678;
wire n_11546;
wire n_3329;
wire n_8662;
wire n_330;
wire n_10503;
wire n_9694;
wire n_3826;
wire n_4905;
wire n_7158;
wire n_1406;
wire n_4601;
wire n_9905;
wire n_962;
wire n_9948;
wire n_10465;
wire n_12429;
wire n_10590;
wire n_3647;
wire n_3681;
wire n_1883;
wire n_4300;
wire n_1288;
wire n_8526;
wire n_1186;
wire n_4623;
wire n_7325;
wire n_10887;
wire n_9456;
wire n_5007;
wire n_7044;
wire n_3320;
wire n_9710;
wire n_6370;
wire n_8623;
wire n_11113;
wire n_9923;
wire n_2518;
wire n_5883;
wire n_7166;
wire n_6554;
wire n_12146;
wire n_7356;
wire n_5754;
wire n_6759;
wire n_10786;
wire n_3988;
wire n_6560;
wire n_11319;
wire n_1720;
wire n_3476;
wire n_7028;
wire n_4842;
wire n_204;
wire n_482;
wire n_7838;
wire n_9890;
wire n_5629;
wire n_3439;
wire n_4135;
wire n_11492;
wire n_7873;
wire n_2688;
wire n_394;
wire n_1845;
wire n_1489;
wire n_6535;
wire n_12731;
wire n_12399;
wire n_942;
wire n_12342;
wire n_7518;
wire n_2798;
wire n_7414;
wire n_9817;
wire n_9744;
wire n_6147;
wire n_2852;
wire n_9199;
wire n_10063;
wire n_12640;
wire n_1524;
wire n_9548;
wire n_8973;
wire n_11160;
wire n_6448;
wire n_7791;
wire n_1964;
wire n_12378;
wire n_8419;
wire n_9782;
wire n_1920;
wire n_2753;
wire n_12533;
wire n_1496;
wire n_3292;
wire n_2007;
wire n_2039;
wire n_9862;
wire n_5434;
wire n_5934;
wire n_7431;
wire n_1225;
wire n_12616;
wire n_11385;
wire n_1544;
wire n_1485;
wire n_12319;
wire n_10805;
wire n_11355;
wire n_11674;
wire n_1846;
wire n_12535;
wire n_3437;
wire n_12178;
wire n_4111;
wire n_12653;
wire n_6643;
wire n_533;
wire n_12327;
wire n_7146;
wire n_9471;
wire n_3712;
wire n_4608;
wire n_879;
wire n_2310;
wire n_11346;
wire n_2506;
wire n_10091;
wire n_11638;
wire n_6157;
wire n_4859;
wire n_9363;
wire n_12047;
wire n_2626;
wire n_12930;
wire n_12587;
wire n_5880;
wire n_1567;
wire n_4037;
wire n_8351;
wire n_8430;
wire n_10747;
wire n_12058;
wire n_9069;
wire n_13110;
wire n_3562;
wire n_5852;
wire n_2973;
wire n_9422;
wire n_8603;
wire n_5218;
wire n_8249;
wire n_7052;
wire n_11343;
wire n_12348;
wire n_3665;
wire n_273;
wire n_10496;
wire n_3007;
wire n_12257;
wire n_3528;
wire n_12575;
wire n_5960;
wire n_11451;
wire n_4571;
wire n_10843;
wire n_3698;
wire n_7888;
wire n_11823;
wire n_5358;
wire n_6397;
wire n_3355;
wire n_2454;
wire n_8234;
wire n_2114;
wire n_3174;
wire n_5321;
wire n_9960;
wire n_1066;
wire n_10997;
wire n_1948;
wire n_157;
wire n_4215;
wire n_9010;
wire n_10998;
wire n_9003;
wire n_2154;
wire n_9280;
wire n_6073;
wire n_7502;
wire n_1484;
wire n_12418;
wire n_6331;
wire n_5290;
wire n_4185;
wire n_3752;
wire n_7312;
wire n_7919;
wire n_2283;
wire n_5145;
wire n_4219;
wire n_1229;
wire n_11269;
wire n_10800;
wire n_7085;
wire n_1373;
wire n_11491;
wire n_12065;
wire n_3958;
wire n_9341;
wire n_6939;
wire n_7848;
wire n_11408;
wire n_3985;
wire n_2427;
wire n_11772;
wire n_4196;
wire n_1447;
wire n_4774;
wire n_2056;
wire n_5210;
wire n_6689;
wire n_10993;
wire n_7632;
wire n_4242;
wire n_5109;
wire n_3389;
wire n_12519;
wire n_9172;
wire n_12769;
wire n_4232;
wire n_4190;
wire n_4902;
wire n_3000;
wire n_6405;
wire n_7580;
wire n_5149;
wire n_8980;
wire n_12641;
wire n_13007;
wire n_5571;
wire n_2680;
wire n_11311;
wire n_10112;
wire n_1047;
wire n_10765;
wire n_3375;
wire n_3899;
wire n_6698;
wire n_11792;
wire n_1385;
wire n_7304;
wire n_3713;
wire n_1931;
wire n_9734;
wire n_502;
wire n_2668;
wire n_7288;
wire n_8558;
wire n_10489;
wire n_1257;
wire n_7707;
wire n_3197;
wire n_7223;
wire n_12421;
wire n_7833;
wire n_12113;
wire n_4987;
wire n_2128;
wire n_5512;
wire n_7274;
wire n_9297;
wire n_10159;
wire n_10495;
wire n_9004;
wire n_4736;
wire n_2398;
wire n_1725;
wire n_3743;
wire n_6206;
wire n_9068;
wire n_8136;
wire n_834;
wire n_5033;
wire n_9808;
wire n_4035;
wire n_2695;
wire n_3818;
wire n_6610;
wire n_7445;
wire n_3124;
wire n_10612;
wire n_11086;
wire n_1741;
wire n_7466;
wire n_1002;
wire n_10260;
wire n_6529;
wire n_11293;
wire n_1949;
wire n_3759;
wire n_545;
wire n_2671;
wire n_4516;
wire n_12285;
wire n_6750;
wire n_6363;
wire n_2715;
wire n_1804;
wire n_11710;
wire n_8619;
wire n_251;
wire n_2508;
wire n_11568;
wire n_3511;
wire n_2054;
wire n_6290;
wire n_10253;
wire n_7429;
wire n_11766;
wire n_6025;
wire n_11038;
wire n_1337;
wire n_9150;
wire n_10134;
wire n_11603;
wire n_1477;
wire n_7277;
wire n_6455;
wire n_12683;
wire n_11271;
wire n_12455;
wire n_13099;
wire n_2614;
wire n_12015;
wire n_8146;
wire n_4492;
wire n_2833;
wire n_2758;
wire n_8813;
wire n_5607;
wire n_11562;
wire n_3694;
wire n_7695;
wire n_2937;
wire n_10194;
wire n_7179;
wire n_10356;
wire n_7122;
wire n_10173;
wire n_12157;
wire n_7869;
wire n_7165;
wire n_4789;
wire n_5999;
wire n_8910;
wire n_12311;
wire n_4376;
wire n_6203;
wire n_1001;
wire n_6408;
wire n_2241;
wire n_6555;
wire n_9448;
wire n_7683;
wire n_10739;
wire n_13064;
wire n_6150;
wire n_7630;
wire n_10077;
wire n_4708;
wire n_8470;
wire n_4657;
wire n_9587;
wire n_12031;
wire n_1690;
wire n_5341;
wire n_1191;
wire n_8643;
wire n_1076;
wire n_4512;
wire n_9278;
wire n_10671;
wire n_1378;
wire n_855;
wire n_10889;
wire n_10010;
wire n_10193;
wire n_1377;
wire n_11718;
wire n_8565;
wire n_10821;
wire n_11170;
wire n_695;
wire n_11758;
wire n_12126;
wire n_8550;
wire n_4081;
wire n_1542;
wire n_9396;
wire n_4542;
wire n_6892;
wire n_11094;
wire n_4462;
wire n_7061;
wire n_11680;
wire n_12480;
wire n_10599;
wire n_9667;
wire n_6401;
wire n_7322;
wire n_1716;
wire n_278;
wire n_9053;
wire n_11658;
wire n_11893;
wire n_6685;
wire n_11639;
wire n_12226;
wire n_4931;
wire n_9739;
wire n_10573;
wire n_4536;
wire n_9480;
wire n_5562;
wire n_3303;
wire n_978;
wire n_4324;
wire n_7051;
wire n_10850;
wire n_384;
wire n_8477;
wire n_9185;
wire n_1976;
wire n_7880;
wire n_9793;
wire n_11692;
wire n_4382;
wire n_12195;
wire n_2905;
wire n_13115;
wire n_1291;
wire n_11759;
wire n_8230;
wire n_12549;
wire n_6679;
wire n_8092;
wire n_749;
wire n_1824;
wire n_3954;
wire n_5911;
wire n_11601;
wire n_11971;
wire n_2122;
wire n_11456;
wire n_12314;
wire n_10546;
wire n_5622;
wire n_2140;
wire n_3503;
wire n_9919;
wire n_3160;
wire n_12135;
wire n_1065;
wire n_6574;
wire n_11116;
wire n_12604;
wire n_6571;
wire n_5577;
wire n_9541;
wire n_11286;
wire n_1255;
wire n_568;
wire n_8876;
wire n_5124;
wire n_143;
wire n_9151;
wire n_3951;
wire n_8829;
wire n_823;
wire n_7824;
wire n_9359;
wire n_1074;
wire n_698;
wire n_3569;
wire n_739;
wire n_7094;
wire n_3874;
wire n_2528;
wire n_5123;
wire n_7097;
wire n_4639;
wire n_5413;
wire n_8140;
wire n_8971;
wire n_8060;
wire n_1338;
wire n_1097;
wire n_10558;
wire n_3027;
wire n_781;
wire n_4083;
wire n_7036;
wire n_9579;
wire n_9475;
wire n_11124;
wire n_6392;
wire n_1810;
wire n_182;
wire n_5915;
wire n_8527;
wire n_573;
wire n_12899;
wire n_9049;
wire n_7351;
wire n_1583;
wire n_4480;
wire n_1730;
wire n_9352;
wire n_2295;
wire n_2746;
wire n_389;
wire n_814;
wire n_7608;
wire n_5779;
wire n_1643;
wire n_2020;
wire n_6260;
wire n_6832;
wire n_7394;
wire n_11045;
wire n_7909;
wire n_7413;
wire n_4171;
wire n_6303;
wire n_3652;
wire n_8935;
wire n_222;
wire n_11340;
wire n_10734;
wire n_6286;
wire n_7675;
wire n_8267;
wire n_4023;
wire n_11903;
wire n_7027;
wire n_1105;
wire n_7992;
wire n_6912;
wire n_11560;
wire n_721;
wire n_10330;
wire n_1461;
wire n_742;
wire n_8276;
wire n_691;
wire n_3617;
wire n_10395;
wire n_7175;
wire n_2076;
wire n_6019;
wire n_10174;
wire n_11435;
wire n_3567;
wire n_11465;
wire n_377;
wire n_1598;
wire n_7524;
wire n_4344;
wire n_2935;
wire n_8027;
wire n_4705;
wire n_4046;
wire n_11564;
wire n_3807;
wire n_8925;
wire n_6214;
wire n_12946;
wire n_9978;
wire n_11914;
wire n_11265;
wire n_9370;
wire n_11125;
wire n_918;
wire n_9670;
wire n_13136;
wire n_1114;
wire n_763;
wire n_4027;
wire n_12916;
wire n_3154;
wire n_9334;
wire n_7783;
wire n_6692;
wire n_1227;
wire n_2485;
wire n_3898;
wire n_10276;
wire n_12331;
wire n_3520;
wire n_191;
wire n_8978;
wire n_10594;
wire n_8093;
wire n_12531;
wire n_8245;
wire n_6036;
wire n_8471;
wire n_4391;
wire n_12521;
wire n_11302;
wire n_946;
wire n_12910;
wire n_9956;
wire n_1303;
wire n_9800;
wire n_8454;
wire n_6552;
wire n_4095;
wire n_8327;
wire n_11382;
wire n_13096;
wire n_9413;
wire n_12727;
wire n_10991;
wire n_2881;
wire n_10098;
wire n_1116;
wire n_11745;
wire n_1570;
wire n_1702;
wire n_8891;
wire n_1219;
wire n_3551;
wire n_4947;
wire n_3064;
wire n_11690;
wire n_9487;
wire n_1780;
wire n_3897;
wire n_11707;
wire n_1689;
wire n_5591;
wire n_11373;
wire n_3372;
wire n_7697;
wire n_1944;
wire n_6403;
wire n_7306;
wire n_1347;
wire n_7947;
wire n_795;
wire n_10118;
wire n_1221;
wire n_7470;
wire n_7547;
wire n_6013;
wire n_7733;
wire n_1245;
wire n_7693;
wire n_9557;
wire n_3215;
wire n_6491;
wire n_448;
wire n_3853;
wire n_4740;
wire n_4631;
wire n_11412;
wire n_6348;
wire n_6744;
wire n_1561;
wire n_13039;
wire n_13130;
wire n_8582;
wire n_10441;
wire n_1112;
wire n_5518;
wire n_6982;
wire n_10002;
wire n_2081;
wire n_2168;
wire n_5068;
wire n_6293;
wire n_6661;
wire n_234;
wire n_9124;
wire n_5847;
wire n_7345;
wire n_6049;
wire n_1460;
wire n_911;
wire n_8847;
wire n_9762;
wire n_11242;
wire n_8957;
wire n_7385;
wire n_10923;
wire n_5159;
wire n_2862;
wire n_472;
wire n_2615;
wire n_4068;
wire n_6558;
wire n_4625;
wire n_11149;
wire n_10841;
wire n_2474;
wire n_3703;
wire n_12635;
wire n_12227;
wire n_12258;
wire n_2444;
wire n_2437;
wire n_12313;
wire n_3962;
wire n_2743;
wire n_4766;
wire n_8488;
wire n_9271;
wire n_4863;
wire n_2267;
wire n_9543;
wire n_3035;
wire n_668;
wire n_4166;
wire n_11396;
wire n_8356;
wire n_1821;
wire n_6136;
wire n_9660;
wire n_11443;
wire n_9483;
wire n_1058;
wire n_3378;
wire n_6855;
wire n_3745;
wire n_3362;
wire n_10665;
wire n_4744;
wire n_12906;
wire n_8888;
wire n_11810;
wire n_4188;
wire n_5357;
wire n_2934;
wire n_3667;
wire n_6091;
wire n_3523;
wire n_2222;
wire n_712;
wire n_13093;
wire n_13062;
wire n_9328;
wire n_7857;
wire n_3176;
wire n_7481;
wire n_12583;
wire n_6551;
wire n_7691;
wire n_7907;
wire n_5541;
wire n_5568;
wire n_10576;
wire n_6312;
wire n_8747;
wire n_2505;
wire n_9539;
wire n_334;
wire n_4817;
wire n_11532;
wire n_6668;
wire n_9415;
wire n_4115;
wire n_2999;
wire n_2014;
wire n_9385;
wire n_1239;
wire n_3697;
wire n_1584;
wire n_9147;
wire n_470;
wire n_11209;
wire n_7653;
wire n_3680;
wire n_5381;
wire n_8354;
wire n_2408;
wire n_9785;
wire n_5723;
wire n_6859;
wire n_5918;
wire n_3468;
wire n_6959;
wire n_8353;
wire n_8922;
wire n_6388;
wire n_5045;
wire n_10237;
wire n_11053;
wire n_11790;
wire n_9027;
wire n_1972;
wire n_12159;
wire n_9434;
wire n_12750;
wire n_4383;
wire n_10902;
wire n_6995;
wire n_4491;
wire n_12889;
wire n_5696;
wire n_8348;
wire n_7032;
wire n_455;
wire n_8211;
wire n_12050;
wire n_12922;
wire n_363;
wire n_12250;
wire n_4486;
wire n_9515;
wire n_10420;
wire n_6971;
wire n_1816;
wire n_11304;
wire n_9642;
wire n_393;
wire n_503;
wire n_9233;
wire n_6131;
wire n_9681;
wire n_5848;
wire n_3024;
wire n_7475;
wire n_10485;
wire n_12105;
wire n_4612;
wire n_12385;
wire n_6435;
wire n_10536;
wire n_5673;
wire n_5443;
wire n_2531;
wire n_6351;
wire n_9079;
wire n_9382;
wire n_10282;
wire n_5163;
wire n_6212;
wire n_7668;
wire n_9775;
wire n_307;
wire n_10444;
wire n_4529;
wire n_500;
wire n_3361;
wire n_11377;
wire n_714;
wire n_3478;
wire n_8653;
wire n_8018;
wire n_3936;
wire n_1349;
wire n_291;
wire n_8920;
wire n_10913;
wire n_7937;
wire n_9176;
wire n_6829;
wire n_2723;
wire n_10950;
wire n_5485;
wire n_7819;
wire n_10631;
wire n_5823;
wire n_7305;
wire n_2800;
wire n_3496;
wire n_13160;
wire n_11071;
wire n_5473;
wire n_10072;
wire n_6682;
wire n_6334;
wire n_6823;
wire n_10708;
wire n_10703;
wire n_9089;
wire n_9666;
wire n_4390;
wire n_12248;
wire n_8678;
wire n_3096;
wire n_10565;
wire n_10011;
wire n_2651;
wire n_8884;
wire n_8803;
wire n_2095;
wire n_3239;
wire n_8942;
wire n_7993;
wire n_7181;
wire n_9865;
wire n_3161;
wire n_2799;
wire n_5537;
wire n_10978;
wire n_8222;
wire n_6822;
wire n_4062;
wire n_3902;
wire n_3295;
wire n_11715;
wire n_4396;
wire n_8553;
wire n_7071;
wire n_1998;
wire n_9706;
wire n_1574;
wire n_3101;
wire n_240;
wire n_10642;
wire n_756;
wire n_1981;
wire n_4233;
wire n_1606;
wire n_12181;
wire n_10187;
wire n_3374;
wire n_10387;
wire n_11014;
wire n_2640;
wire n_253;
wire n_1552;
wire n_3288;
wire n_583;
wire n_2918;
wire n_8751;
wire n_4307;
wire n_3992;
wire n_11864;
wire n_3876;
wire n_11007;
wire n_11224;
wire n_249;
wire n_11006;
wire n_9564;
wire n_3125;
wire n_7391;
wire n_8790;
wire n_9230;
wire n_6617;
wire n_4293;
wire n_10219;
wire n_941;
wire n_3552;
wire n_1031;
wire n_7511;
wire n_6533;
wire n_11924;
wire n_10768;
wire n_10316;
wire n_9795;
wire n_849;
wire n_4684;
wire n_3116;
wire n_9591;
wire n_6429;
wire n_6407;
wire n_4091;
wire n_1753;
wire n_6389;
wire n_5027;
wire n_3095;
wire n_6137;
wire n_10364;
wire n_2471;
wire n_10479;
wire n_11422;
wire n_8338;
wire n_6983;
wire n_10494;
wire n_8398;
wire n_4412;
wire n_2807;
wire n_8178;
wire n_6801;
wire n_1921;
wire n_12489;
wire n_8491;
wire n_3618;
wire n_4580;
wire n_1055;
wire n_2217;
wire n_2197;
wire n_4758;
wire n_5630;
wire n_4781;
wire n_10065;
wire n_12046;
wire n_10212;
wire n_9283;
wire n_8700;
wire n_4148;
wire n_2461;
wire n_271;
wire n_12030;
wire n_12738;
wire n_206;
wire n_4057;
wire n_633;
wire n_1170;
wire n_5379;
wire n_13025;
wire n_5335;
wire n_11599;
wire n_12565;
wire n_308;
wire n_10268;
wire n_3444;
wire n_1040;
wire n_3059;
wire n_6113;
wire n_9468;
wire n_10070;
wire n_12601;
wire n_9425;
wire n_12917;
wire n_2634;
wire n_1761;
wire n_11172;
wire n_10089;
wire n_5424;
wire n_12415;
wire n_8750;
wire n_1890;
wire n_3017;
wire n_1805;
wire n_2477;
wire n_5505;
wire n_5868;
wire n_10305;
wire n_8560;
wire n_10559;
wire n_2308;
wire n_2333;
wire n_8439;
wire n_3001;
wire n_9641;
wire n_1089;
wire n_12755;
wire n_10004;
wire n_12807;
wire n_12059;
wire n_12488;
wire n_3795;
wire n_7321;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_5289;
wire n_8200;
wire n_11110;
wire n_7154;
wire n_5018;
wire n_6129;
wire n_6518;
wire n_8304;
wire n_3896;
wire n_3815;
wire n_11418;
wire n_6655;
wire n_8674;
wire n_12981;
wire n_5274;
wire n_9138;
wire n_3274;
wire n_5401;
wire n_12977;
wire n_7584;
wire n_9958;
wire n_4457;
wire n_7537;
wire n_10516;
wire n_4093;
wire n_1616;
wire n_8675;
wire n_6254;
wire n_1862;
wire n_5989;
wire n_10892;
wire n_339;
wire n_434;
wire n_10493;
wire n_288;
wire n_12567;
wire n_9367;
wire n_7320;
wire n_4928;
wire n_5769;
wire n_10405;
wire n_4794;
wire n_722;
wire n_5613;
wire n_8212;
wire n_5612;
wire n_2223;
wire n_4197;
wire n_7964;
wire n_4482;
wire n_629;
wire n_1621;
wire n_9016;
wire n_2547;
wire n_2415;
wire n_13101;
wire n_11887;
wire n_6278;
wire n_6786;
wire n_7022;
wire n_10026;
wire n_11545;
wire n_9729;
wire n_5073;
wire n_12691;
wire n_827;
wire n_8846;
wire n_8315;
wire n_12471;
wire n_11033;
wire n_12451;
wire n_4834;
wire n_11040;
wire n_12665;
wire n_11754;
wire n_11850;
wire n_9194;
wire n_8760;
wire n_9756;
wire n_12592;
wire n_4762;
wire n_192;
wire n_5581;
wire n_9029;
wire n_9411;
wire n_11672;
wire n_3113;
wire n_6837;
wire n_10353;
wire n_992;
wire n_3813;
wire n_3660;
wire n_10847;
wire n_12651;
wire n_3766;
wire n_1613;
wire n_10451;
wire n_11043;
wire n_1458;
wire n_5303;
wire n_12507;
wire n_7486;
wire n_12240;
wire n_6756;
wire n_9414;
wire n_1027;
wire n_3266;
wire n_12003;
wire n_3574;
wire n_9615;
wire n_7023;
wire n_7496;
wire n_1189;
wire n_11277;
wire n_223;
wire n_4154;
wire n_12165;
wire n_4907;
wire n_5077;
wire n_5034;
wire n_726;
wire n_10866;
wire n_7410;
wire n_9940;
wire n_10779;
wire n_8563;
wire n_6200;
wire n_4504;
wire n_365;
wire n_3844;
wire n_8777;
wire n_1237;
wire n_2534;
wire n_4975;
wire n_11061;
wire n_11763;
wire n_8465;
wire n_6670;
wire n_3741;
wire n_10653;
wire n_11534;
wire n_11587;
wire n_8535;
wire n_5375;
wire n_12280;
wire n_6373;
wire n_9221;
wire n_12492;
wire n_2451;
wire n_12972;
wire n_5370;
wire n_2243;
wire n_4898;
wire n_4815;
wire n_5784;
wire n_5601;
wire n_9811;
wire n_3443;
wire n_7899;
wire n_8631;
wire n_509;
wire n_4819;
wire n_1209;
wire n_7906;
wire n_5248;
wire n_9951;
wire n_1708;
wire n_7131;
wire n_805;
wire n_396;
wire n_6411;
wire n_350;
wire n_2051;
wire n_9424;
wire n_9586;
wire n_10285;
wire n_4370;
wire n_8909;
wire n_11032;
wire n_2359;
wire n_5112;
wire n_480;
wire n_142;
wire n_1402;
wire n_1691;
wire n_3332;
wire n_4134;
wire n_10507;
wire n_10520;
wire n_7302;
wire n_11968;
wire n_11843;
wire n_1238;
wire n_2570;
wire n_4092;
wire n_10045;
wire n_11174;
wire n_4645;
wire n_7797;
wire n_3668;
wire n_11335;
wire n_11629;
wire n_6381;
wire n_7030;
wire n_6656;
wire n_9730;
wire n_7687;
wire n_2491;
wire n_1264;
wire n_9554;
wire n_10294;
wire n_4755;
wire n_4359;
wire n_4960;
wire n_10106;
wire n_4087;
wire n_1700;
wire n_5635;
wire n_7582;
wire n_9934;
wire n_4933;
wire n_10541;
wire n_5091;
wire n_3487;
wire n_4591;
wire n_6546;
wire n_5528;
wire n_287;
wire n_4302;
wire n_9234;
wire n_10674;
wire n_5111;
wire n_8959;
wire n_11698;
wire n_6534;
wire n_3340;
wire n_10614;
wire n_230;
wire n_5227;
wire n_7809;
wire n_11785;
wire n_461;
wire n_873;
wire n_10417;
wire n_3946;
wire n_12841;
wire n_6265;
wire n_12855;
wire n_2989;
wire n_5778;
wire n_8425;
wire n_11257;
wire n_8087;
wire n_9910;
wire n_3395;
wire n_7060;
wire n_7607;
wire n_10217;
wire n_8938;
wire n_4474;
wire n_5665;
wire n_2509;
wire n_11801;
wire n_2513;
wire n_12073;
wire n_6898;
wire n_6596;
wire n_3757;
wire n_5363;
wire n_4178;
wire n_10743;
wire n_5165;
wire n_1704;
wire n_2247;
wire n_250;
wire n_1711;
wire n_4884;
wire n_10853;
wire n_1579;
wire n_7867;
wire n_9651;
wire n_3275;
wire n_10249;
wire n_8361;
wire n_836;
wire n_6135;
wire n_7761;
wire n_10705;
wire n_8007;
wire n_9246;
wire n_10338;
wire n_522;
wire n_10270;
wire n_3678;
wire n_6814;
wire n_10557;
wire n_3440;
wire n_11115;
wire n_8669;
wire n_12978;
wire n_8001;
wire n_2094;
wire n_7525;
wire n_1511;
wire n_2356;
wire n_7257;
wire n_12363;
wire n_9372;
wire n_7553;
wire n_1422;
wire n_7529;
wire n_1772;
wire n_4692;
wire n_6791;
wire n_616;
wire n_8496;
wire n_3165;
wire n_11915;
wire n_1119;
wire n_6824;
wire n_5788;
wire n_11016;
wire n_9326;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_11788;
wire n_1620;
wire n_2739;
wire n_12544;
wire n_1735;
wire n_3890;
wire n_1541;
wire n_1300;
wire n_641;
wire n_13036;
wire n_3750;
wire n_1313;
wire n_3607;
wire n_7650;
wire n_12476;
wire n_3316;
wire n_8568;
wire n_516;
wire n_6903;
wire n_2418;
wire n_2864;
wire n_13009;
wire n_13043;
wire n_8852;
wire n_4311;
wire n_12023;
wire n_1180;
wire n_8637;
wire n_2703;
wire n_6168;
wire n_6881;
wire n_3371;
wire n_4722;
wire n_4606;
wire n_10339;
wire n_9908;
wire n_10908;
wire n_9486;
wire n_6450;
wire n_9544;
wire n_13002;
wire n_3261;
wire n_666;
wire n_12620;
wire n_12632;
wire n_9831;
wire n_7520;
wire n_4187;
wire n_6309;
wire n_940;
wire n_7903;
wire n_9697;
wire n_2058;
wire n_11303;
wire n_405;
wire n_213;
wire n_2660;
wire n_11877;
wire n_6733;
wire n_8864;
wire n_7384;
wire n_8456;
wire n_5317;
wire n_1094;
wire n_5430;
wire n_5942;
wire n_8610;
wire n_7894;
wire n_4962;
wire n_4563;
wire n_9902;
wire n_7137;
wire n_494;
wire n_5056;
wire n_8362;
wire n_4820;
wire n_2394;
wire n_5540;
wire n_11750;
wire n_9900;
wire n_6300;
wire n_8256;
wire n_3532;
wire n_9920;
wire n_7055;
wire n_7202;
wire n_5716;
wire n_8520;
wire n_9310;
wire n_10132;
wire n_3948;
wire n_9039;
wire n_12598;
wire n_11854;
wire n_12416;
wire n_8573;
wire n_12055;
wire n_12091;
wire n_2124;
wire n_8704;
wire n_4619;
wire n_381;
wire n_7639;
wire n_8265;
wire n_5762;
wire n_6132;
wire n_4327;
wire n_1961;
wire n_5211;
wire n_5336;
wire n_11609;
wire n_3765;
wire n_5447;
wire n_4125;
wire n_7743;
wire n_9294;
wire n_5036;
wire n_12811;
wire n_4221;
wire n_3297;
wire n_12186;
wire n_11747;
wire n_6179;
wire n_6395;
wire n_10327;
wire n_12494;
wire n_13032;
wire n_976;
wire n_7605;
wire n_7054;
wire n_3067;
wire n_11556;
wire n_2155;
wire n_11001;
wire n_9512;
wire n_10437;
wire n_11529;
wire n_2686;
wire n_5327;
wire n_10021;
wire n_9146;
wire n_2364;
wire n_9125;
wire n_4392;
wire n_9170;
wire n_9139;
wire n_11858;
wire n_2996;
wire n_7433;
wire n_9616;
wire n_8131;
wire n_3803;
wire n_2085;
wire n_8941;
wire n_917;
wire n_5014;
wire n_5747;
wire n_3639;
wire n_9073;
wire n_10075;
wire n_12733;
wire n_10423;
wire n_12897;
wire n_12623;
wire n_11444;
wire n_5192;
wire n_4334;
wire n_659;
wire n_3351;
wire n_6171;
wire n_8775;
wire n_808;
wire n_12272;
wire n_9302;
wire n_5519;
wire n_11798;
wire n_9062;
wire n_11895;
wire n_4047;
wire n_6269;
wire n_5753;
wire n_3413;
wire n_7092;
wire n_6980;
wire n_11213;
wire n_12245;
wire n_1193;
wire n_9171;
wire n_10886;
wire n_5233;
wire n_3412;
wire n_8279;
wire n_12213;
wire n_9358;
wire n_6654;
wire n_12191;
wire n_9580;
wire n_8019;
wire n_9972;
wire n_3791;
wire n_13003;
wire n_6083;
wire n_13091;
wire n_12909;
wire n_3164;
wire n_4575;
wire n_6434;
wire n_6387;
wire n_551;
wire n_699;
wire n_4320;
wire n_9565;
wire n_9157;
wire n_8257;
wire n_13072;
wire n_10192;
wire n_7832;
wire n_3884;
wire n_9465;
wire n_9540;
wire n_9324;
wire n_5808;
wire n_451;
wire n_8390;
wire n_11137;
wire n_8898;
wire n_7726;
wire n_8807;
wire n_5436;
wire n_5139;
wire n_757;
wire n_594;
wire n_5231;
wire n_2190;
wire n_6120;
wire n_8613;
wire n_6068;
wire n_6933;
wire n_8521;
wire n_3438;
wire n_166;
wire n_4141;
wire n_10436;
wire n_8464;
wire n_6547;
wire n_8799;
wire n_12794;
wire n_5193;
wire n_6423;
wire n_9442;
wire n_2850;
wire n_572;
wire n_6342;
wire n_6641;
wire n_1481;
wire n_6984;
wire n_1441;
wire n_3373;
wire n_5789;
wire n_10763;
wire n_2104;
wire n_7441;
wire n_9957;
wire n_513;
wire n_10124;
wire n_12483;
wire n_12759;
wire n_11793;
wire n_7106;
wire n_7213;
wire n_12112;
wire n_13060;
wire n_3883;
wire n_10245;
wire n_5961;
wire n_10905;
wire n_261;
wire n_11235;
wire n_9449;
wire n_5866;
wire n_9050;
wire n_3728;
wire n_6507;
wire n_2925;
wire n_4499;
wire n_6399;
wire n_9313;
wire n_6687;
wire n_5822;
wire n_9173;
wire n_433;
wire n_5195;
wire n_6690;
wire n_6121;
wire n_7412;
wire n_9959;
wire n_12144;
wire n_3949;
wire n_5726;
wire n_9563;
wire n_11015;
wire n_2792;
wire n_9160;
wire n_219;
wire n_5364;
wire n_9974;
wire n_12129;
wire n_11166;
wire n_3315;
wire n_7031;
wire n_9285;
wire n_263;
wire n_5533;
wire n_7763;
wire n_3798;
wire n_788;
wire n_9631;
wire n_1543;
wire n_8033;
wire n_1599;
wire n_329;
wire n_4257;
wire n_4458;
wire n_6194;
wire n_2674;
wire n_5103;
wire n_4641;
wire n_8393;
wire n_7133;
wire n_12032;
wire n_4720;
wire n_10784;
wire n_12202;
wire n_4893;
wire n_3857;
wire n_1876;
wire n_4107;
wire n_8463;
wire n_8153;
wire n_243;
wire n_12815;
wire n_1873;
wire n_3630;
wire n_6524;
wire n_3518;
wire n_10944;
wire n_10211;
wire n_12835;
wire n_10129;
wire n_10431;
wire n_1866;
wire n_9945;
wire n_8661;
wire n_12431;
wire n_2130;
wire n_7424;
wire n_1413;
wire n_1330;
wire n_3714;
wire n_7523;
wire n_2228;
wire n_8654;
wire n_5039;
wire n_11855;
wire n_2455;
wire n_2876;
wire n_4772;
wire n_6790;
wire n_8746;
wire n_11241;
wire n_5953;
wire n_12870;
wire n_11183;
wire n_10019;
wire n_3099;
wire n_11156;
wire n_8531;
wire n_11508;
wire n_10611;
wire n_12093;
wire n_7141;
wire n_5198;
wire n_11581;
wire n_10715;
wire n_4468;
wire n_5718;
wire n_4161;
wire n_6505;
wire n_1663;
wire n_6459;
wire n_12333;
wire n_12636;
wire n_8379;
wire n_8609;
wire n_4172;
wire n_3403;
wire n_11227;
wire n_7626;
wire n_13100;
wire n_2714;
wire n_2245;
wire n_4961;
wire n_7310;
wire n_4454;
wire n_1107;
wire n_12334;
wire n_2457;
wire n_3294;
wire n_6686;
wire n_4119;
wire n_6001;
wire n_7311;
wire n_9209;
wire n_3686;
wire n_7669;
wire n_11218;
wire n_4502;
wire n_12119;
wire n_11787;
wire n_12618;
wire n_5958;
wire n_8793;
wire n_12355;
wire n_8103;
wire n_318;
wire n_9767;
wire n_2971;
wire n_1713;
wire n_9838;
wire n_10195;
wire n_715;
wire n_4277;
wire n_4526;
wire n_9300;
wire n_1265;
wire n_11500;
wire n_3490;
wire n_4849;
wire n_12943;
wire n_530;
wire n_277;
wire n_4319;
wire n_7327;
wire n_3369;
wire n_12938;
wire n_13057;
wire n_8873;
wire n_8367;
wire n_11891;
wire n_618;
wire n_7367;
wire n_199;
wire n_5792;
wire n_11021;
wire n_3581;
wire n_12401;
wire n_8543;
wire n_3069;
wire n_6183;
wire n_6023;
wire n_13055;
wire n_7323;
wire n_11544;
wire n_7189;
wire n_7301;
wire n_12173;
wire n_13067;
wire n_10730;
wire n_6258;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_6905;
wire n_10243;
wire n_612;
wire n_9700;
wire n_10564;
wire n_8682;
wire n_3725;
wire n_8089;
wire n_9218;
wire n_6704;
wire n_3933;
wire n_8533;
wire n_9118;
wire n_11122;
wire n_6657;
wire n_7655;
wire n_5554;
wire n_1175;
wire n_7244;
wire n_10745;
wire n_7368;
wire n_2311;
wire n_429;
wire n_1012;
wire n_3691;
wire n_10596;
wire n_5553;
wire n_4485;
wire n_8011;
wire n_4066;
wire n_903;
wire n_7633;
wire n_4146;
wire n_5711;
wire n_12140;
wire n_9437;
wire n_1802;
wire n_1504;
wire n_10263;
wire n_4340;
wire n_5790;
wire n_286;
wire n_11509;
wire n_8640;
wire n_254;
wire n_8063;
wire n_3961;
wire n_11960;
wire n_4855;
wire n_12599;
wire n_1801;
wire n_2347;
wire n_3917;
wire n_6186;
wire n_7878;
wire n_6803;
wire n_9514;
wire n_12411;
wire n_816;
wire n_6210;
wire n_8437;
wire n_6500;
wire n_8427;
wire n_8032;
wire n_10280;
wire n_1188;
wire n_12465;
wire n_7427;
wire n_10605;
wire n_2206;
wire n_4004;
wire n_11029;
wire n_2967;
wire n_13118;
wire n_5404;
wire n_9933;
wire n_11449;
wire n_2916;
wire n_11190;
wire n_5739;
wire n_10951;
wire n_12152;
wire n_4292;
wire n_9892;
wire n_8570;
wire n_6163;
wire n_11794;
wire n_7628;
wire n_9462;
wire n_9074;
wire n_5972;
wire n_10519;
wire n_2467;
wire n_5549;
wire n_9408;
wire n_267;
wire n_3145;
wire n_6785;
wire n_6553;
wire n_1124;
wire n_1624;
wire n_10163;
wire n_10454;
wire n_3983;
wire n_4940;
wire n_5444;
wire n_3538;
wire n_12568;
wire n_3280;
wire n_8039;
wire n_12501;
wire n_5757;
wire n_12970;
wire n_1515;
wire n_8916;
wire n_8902;
wire n_961;
wire n_7557;
wire n_10087;
wire n_4356;
wire n_3510;
wire n_2824;
wire n_593;
wire n_8843;
wire n_9891;
wire n_10146;
wire n_7128;
wire n_9946;
wire n_12959;
wire n_637;
wire n_2377;
wire n_701;
wire n_6849;
wire n_9885;
wire n_7594;
wire n_950;
wire n_12330;
wire n_8129;
wire n_8162;
wire n_7457;
wire n_10643;
wire n_8744;
wire n_3009;
wire n_10504;
wire n_5824;
wire n_3719;
wire n_2525;
wire n_7788;
wire n_4361;
wire n_10872;
wire n_5488;
wire n_6760;
wire n_10701;
wire n_3827;
wire n_891;
wire n_5154;
wire n_2067;
wire n_10658;
wire n_11590;
wire n_11238;
wire n_7752;
wire n_3889;
wire n_2687;
wire n_12591;
wire n_12466;
wire n_1630;
wire n_2887;
wire n_9509;
wire n_4245;
wire n_4136;
wire n_8286;
wire n_3526;
wire n_2194;
wire n_12798;
wire n_2619;
wire n_5329;
wire n_9925;
wire n_4367;
wire n_9757;
wire n_5637;
wire n_9015;
wire n_10874;
wire n_6825;
wire n_1987;
wire n_10008;
wire n_7586;
wire n_6452;
wire n_11831;
wire n_507;
wire n_9628;
wire n_968;
wire n_7767;
wire n_8294;
wire n_2271;
wire n_1008;
wire n_9419;
wire n_12279;
wire n_12243;
wire n_6611;
wire n_8562;
wire n_2583;
wire n_4560;
wire n_12614;
wire n_11378;
wire n_2606;
wire n_4899;
wire n_10250;
wire n_5728;
wire n_5471;
wire n_1033;
wire n_462;
wire n_1052;
wire n_2794;
wire n_10032;
wire n_10592;
wire n_11433;
wire n_5164;
wire n_9277;
wire n_9257;
wire n_2391;
wire n_304;
wire n_2431;
wire n_7207;
wire n_8218;
wire n_9806;
wire n_5843;
wire n_8170;
wire n_9159;
wire n_11558;
wire n_7744;
wire n_2078;
wire n_7021;
wire n_2932;
wire n_1767;
wire n_3431;
wire n_10595;
wire n_7748;
wire n_8537;
wire n_3450;
wire n_6827;
wire n_10126;
wire n_12041;
wire n_449;
wire n_4663;
wire n_11713;
wire n_2893;
wire n_11073;
wire n_1208;
wire n_5484;
wire n_6355;
wire n_2954;
wire n_12566;
wire n_12931;
wire n_2728;
wire n_1072;
wire n_815;
wire n_6227;
wire n_7215;
wire n_7485;
wire n_13074;
wire n_3421;
wire n_9066;
wire n_3183;
wire n_2493;
wire n_4802;
wire n_2705;
wire n_5523;
wire n_10302;
wire n_11974;
wire n_1067;
wire n_12881;
wire n_3405;
wire n_8016;
wire n_8671;
wire n_5423;
wire n_12546;
wire n_255;
wire n_10645;
wire n_13058;
wire n_284;
wire n_1952;
wire n_5074;
wire n_10604;
wire n_11096;
wire n_12036;
wire n_12876;
wire n_4044;
wire n_6564;
wire n_3436;
wire n_11161;
wire n_9671;
wire n_8709;
wire n_8782;
wire n_1026;
wire n_1880;
wire n_3442;
wire n_3366;
wire n_2631;
wire n_12911;
wire n_289;
wire n_12491;
wire n_6468;
wire n_3937;
wire n_10080;
wire n_11216;
wire n_12228;
wire n_10570;
wire n_1293;
wire n_9857;
wire n_3159;
wire n_4701;
wire n_10966;
wire n_12781;
wire n_10057;
wire n_794;
wire n_12929;
wire n_10882;
wire n_727;
wire n_894;
wire n_685;
wire n_9338;
wire n_13071;
wire n_353;
wire n_6857;
wire n_3240;
wire n_8144;
wire n_12261;
wire n_3576;
wire n_10435;
wire n_1863;
wire n_9542;
wire n_12536;
wire n_3385;
wire n_10795;
wire n_10921;
wire n_7171;
wire n_4851;
wire n_6442;
wire n_12061;
wire n_12106;
wire n_3293;
wire n_872;
wire n_3922;
wire n_11085;
wire n_8049;
wire n_5204;
wire n_7762;
wire n_5333;
wire n_9467;
wire n_7068;
wire n_7925;
wire n_7186;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_10609;
wire n_11157;
wire n_4991;
wire n_5594;
wire n_2554;
wire n_12291;
wire n_9097;
wire n_5422;
wire n_6871;
wire n_12124;
wire n_11755;
wire n_1513;
wire n_9783;
wire n_9510;
wire n_9389;
wire n_1913;
wire n_12074;
wire n_4934;
wire n_9404;
wire n_837;
wire n_8357;
wire n_6904;
wire n_10912;
wire n_5087;
wire n_9916;
wire n_12645;
wire n_5526;
wire n_5292;
wire n_2517;
wire n_2713;
wire n_9314;
wire n_11918;
wire n_7017;
wire n_11748;
wire n_12433;
wire n_12745;
wire n_7777;
wire n_9752;
wire n_12138;
wire n_5000;
wire n_2765;
wire n_5403;
wire n_12887;
wire n_2590;
wire n_5551;
wire n_7652;
wire n_3150;
wire n_10220;
wire n_10341;
wire n_11347;
wire n_8701;
wire n_2060;
wire n_4479;
wire n_2608;
wire n_10550;
wire n_6499;
wire n_7830;
wire n_4011;
wire n_5131;
wire n_12217;
wire n_12365;
wire n_1959;
wire n_3133;
wire n_7138;
wire n_12097;
wire n_5257;
wire n_8097;
wire n_9679;
wire n_765;
wire n_1492;
wire n_8084;
wire n_9306;
wire n_8645;
wire n_1340;
wire n_4753;
wire n_4688;
wire n_8712;
wire n_10232;
wire n_4058;
wire n_10461;
wire n_631;
wire n_8289;
wire n_11178;
wire n_2262;
wire n_3611;
wire n_3082;
wire n_4848;
wire n_7966;
wire n_8591;
wire n_5059;
wire n_156;
wire n_8837;
wire n_5887;
wire n_8811;
wire n_843;
wire n_8824;
wire n_11673;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_11432;
wire n_7191;
wire n_3799;
wire n_7712;
wire n_2574;
wire n_4475;
wire n_10412;
wire n_5242;
wire n_10326;
wire n_12650;
wire n_5219;
wire n_8417;
wire n_2675;
wire n_6276;
wire n_9721;
wire n_11344;
wire n_5631;
wire n_3537;
wire n_10499;
wire n_8340;
wire n_4443;
wire n_3887;
wire n_6008;
wire n_1022;
wire n_12487;
wire n_12658;
wire n_614;
wire n_9197;
wire n_7997;
wire n_6420;
wire n_5854;
wire n_11387;
wire n_11333;
wire n_2667;
wire n_5460;
wire n_4587;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_1571;
wire n_2948;
wire n_1577;
wire n_8455;
wire n_7208;
wire n_12288;
wire n_12859;
wire n_2119;
wire n_7283;
wire n_947;
wire n_9210;
wire n_12185;
wire n_1117;
wire n_7961;
wire n_12130;
wire n_9770;
wire n_13120;
wire n_1992;
wire n_5686;
wire n_5899;
wire n_6893;
wire n_7406;
wire n_8681;
wire n_11417;
wire n_8905;
wire n_13008;
wire n_3223;
wire n_10617;
wire n_12271;
wire n_12704;
wire n_3140;
wire n_7807;
wire n_3185;
wire n_4749;
wire n_9592;
wire n_2605;
wire n_5155;
wire n_7680;
wire n_9180;
wire n_10922;
wire n_10544;
wire n_12958;
wire n_926;
wire n_13030;
wire n_3654;
wire n_1849;
wire n_2848;
wire n_919;
wire n_8172;
wire n_9917;
wire n_10718;
wire n_12056;
wire n_1698;
wire n_8106;
wire n_9502;
wire n_4100;
wire n_6447;
wire n_4264;
wire n_12238;
wire n_11952;
wire n_5981;
wire n_3788;
wire n_9625;
wire n_4891;
wire n_5937;
wire n_777;
wire n_6422;
wire n_1299;
wire n_6751;
wire n_5339;
wire n_12976;
wire n_3837;
wire n_2718;
wire n_1436;
wire n_1384;
wire n_11087;
wire n_11477;
wire n_3325;
wire n_2238;
wire n_9873;
wire n_6040;
wire n_11888;
wire n_8375;
wire n_4085;
wire n_4464;
wire n_8612;
wire n_13042;
wire n_4624;
wire n_4818;
wire n_6851;
wire n_6460;
wire n_8345;
wire n_10095;
wire n_4659;
wire n_10309;
wire n_3600;
wire n_8459;
wire n_11773;
wire n_12608;
wire n_6741;
wire n_5217;
wire n_5465;
wire n_11099;
wire n_5015;
wire n_8974;
wire n_4339;
wire n_8268;
wire n_1178;
wire n_2338;
wire n_3324;
wire n_6160;
wire n_9871;
wire n_6650;
wire n_8221;
wire n_10050;
wire n_11682;
wire n_7066;
wire n_9164;
wire n_8255;
wire n_7183;
wire n_796;
wire n_1195;
wire n_7789;
wire n_10306;
wire n_184;
wire n_10878;
wire n_8461;
wire n_7606;
wire n_6192;
wire n_1811;
wire n_6368;
wire n_10056;
wire n_7140;
wire n_7193;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_6039;
wire n_2144;
wire n_1284;
wire n_1604;
wire n_4487;
wire n_11919;
wire n_6583;
wire n_4866;
wire n_4889;
wire n_1142;
wire n_10450;
wire n_623;
wire n_1048;
wire n_5721;
wire n_11414;
wire n_11472;
wire n_3638;
wire n_9114;
wire n_11978;
wire n_4816;
wire n_12520;
wire n_8515;
wire n_10529;
wire n_2110;
wire n_5719;
wire n_1502;
wire n_5773;
wire n_1659;
wire n_5482;
wire n_3393;
wire n_8812;
wire n_13020;
wire n_6012;
wire n_12254;
wire n_3451;
wire n_9392;
wire n_13148;
wire n_1418;
wire n_10429;
wire n_1250;
wire n_292;
wire n_4937;
wire n_11459;
wire n_10904;
wire n_11317;
wire n_5277;
wire n_8792;
wire n_12436;
wire n_3615;
wire n_7344;
wire n_9888;
wire n_11470;
wire n_11538;
wire n_3072;
wire n_3087;
wire n_10037;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_12808;
wire n_4222;
wire n_6707;
wire n_9698;
wire n_4874;
wire n_4401;
wire n_889;
wire n_12744;
wire n_2710;
wire n_6064;
wire n_11136;
wire n_9903;
wire n_3142;
wire n_4015;
wire n_1966;
wire n_5793;
wire n_477;
wire n_9644;
wire n_11353;
wire n_6787;
wire n_11102;
wire n_11620;
wire n_8523;
wire n_1110;
wire n_10179;
wire n_2213;
wire n_9228;
wire n_11539;
wire n_4976;
wire n_7710;
wire n_12143;
wire n_2389;
wire n_9499;
wire n_4709;
wire n_11899;
wire n_7892;
wire n_2132;
wire n_2892;
wire n_6647;
wire n_4120;
wire n_6275;
wire n_9522;
wire n_1564;
wire n_5578;
wire n_11215;
wire n_4658;
wire n_231;
wire n_2860;
wire n_2330;
wire n_5296;
wire n_11076;
wire n_1457;
wire n_9366;
wire n_505;
wire n_11890;
wire n_3718;
wire n_7915;
wire n_5893;
wire n_7750;
wire n_1787;
wire n_9077;
wire n_6769;
wire n_11597;
wire n_537;
wire n_1993;
wire n_9148;
wire n_2281;
wire n_11054;
wire n_11806;
wire n_8406;
wire n_6277;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_10754;
wire n_1919;
wire n_5742;
wire n_5207;
wire n_11050;
wire n_3705;
wire n_3211;
wire n_12443;
wire n_6463;
wire n_3909;
wire n_5676;
wire n_11683;
wire n_8554;
wire n_546;
wire n_10920;
wire n_9275;
wire n_386;
wire n_10223;
wire n_1220;
wire n_6051;
wire n_1893;
wire n_8896;
wire n_2301;
wire n_4665;
wire n_3582;
wire n_11484;
wire n_11126;
wire n_4223;
wire n_7206;
wire n_7538;
wire n_2387;
wire n_5674;
wire n_12934;
wire n_3270;
wire n_5539;
wire n_6895;
wire n_2846;
wire n_5282;
wire n_970;
wire n_10295;
wire n_2488;
wire n_1980;
wire n_5464;
wire n_9409;
wire n_6799;
wire n_2237;
wire n_1060;
wire n_10336;
wire n_1951;
wire n_10228;
wire n_444;
wire n_12555;
wire n_4362;
wire n_1252;
wire n_3311;
wire n_3913;
wire n_1223;
wire n_7716;
wire n_6487;
wire n_11646;
wire n_511;
wire n_5121;
wire n_8758;
wire n_9768;
wire n_6026;
wire n_6070;
wire n_1286;
wire n_8818;
wire n_2115;
wire n_4430;
wire n_3302;
wire n_8617;
wire n_4348;
wire n_12980;
wire n_9881;
wire n_12530;
wire n_5013;
wire n_1597;
wire n_6807;
wire n_8954;
wire n_9463;
wire n_7251;
wire n_4489;
wire n_4839;
wire n_7254;
wire n_12212;
wire n_10466;
wire n_2596;
wire n_12973;
wire n_3163;
wire n_7540;
wire n_775;
wire n_11953;
wire n_4404;
wire n_13123;
wire n_1153;
wire n_5589;
wire n_439;
wire n_13077;
wire n_6563;
wire n_12234;
wire n_10776;
wire n_12624;
wire n_1531;
wire n_7882;
wire n_2828;
wire n_453;
wire n_8552;
wire n_10425;
wire n_7554;
wire n_2384;
wire n_8069;
wire n_7558;
wire n_4261;
wire n_4204;
wire n_8373;
wire n_10848;
wire n_759;
wire n_2724;
wire n_426;
wire n_6481;
wire n_2585;
wire n_5628;
wire n_4825;
wire n_2352;
wire n_7765;
wire n_11482;
wire n_1625;
wire n_3986;
wire n_5006;
wire n_4513;
wire n_7816;
wire n_12151;
wire n_4006;
wire n_2226;
wire n_11089;
wire n_2801;
wire n_9997;
wire n_6341;
wire n_10164;
wire n_6384;
wire n_1901;
wire n_3869;
wire n_7421;
wire n_2556;
wire n_10166;
wire n_7489;
wire n_4747;
wire n_7541;
wire n_6906;
wire n_1647;
wire n_5251;
wire n_3753;
wire n_2306;
wire n_12033;
wire n_1614;
wire n_1892;
wire n_11839;
wire n_3742;
wire n_9844;
wire n_3683;
wire n_8318;
wire n_4801;
wire n_12826;
wire n_401;
wire n_3260;
wire n_10366;
wire n_2550;
wire n_8341;
wire n_9970;
wire n_11193;
wire n_11365;
wire n_3175;
wire n_9595;
wire n_7188;
wire n_3736;
wire n_5475;
wire n_11217;
wire n_7334;
wire n_6923;
wire n_5807;
wire n_4448;
wire n_1096;
wire n_9287;
wire n_7991;
wire n_13051;
wire n_6233;
wire n_2227;
wire n_10877;
wire n_6377;
wire n_11524;
wire n_9265;
wire n_12402;
wire n_5216;
wire n_3284;
wire n_12214;
wire n_10225;
wire n_4869;
wire n_8239;
wire n_427;
wire n_8926;
wire n_6257;
wire n_2159;
wire n_4386;
wire n_688;
wire n_2315;
wire n_1077;
wire n_4132;
wire n_10361;
wire n_11228;
wire n_2995;
wire n_5273;
wire n_7898;
wire n_10766;
wire n_1437;
wire n_4438;
wire n_4844;
wire n_8383;
wire n_10086;
wire n_4836;
wire n_5439;
wire n_7143;
wire n_9789;
wire n_10424;
wire n_12621;
wire n_4955;
wire n_8965;
wire n_11290;
wire n_4149;
wire n_5936;
wire n_12518;
wire n_9608;
wire n_4355;
wire n_7646;
wire n_501;
wire n_2276;
wire n_3234;
wire n_9052;
wire n_856;
wire n_2803;
wire n_8817;
wire n_379;
wire n_8190;
wire n_1668;
wire n_2777;
wire n_11488;
wire n_12162;
wire n_3202;
wire n_2830;
wire n_3220;
wire n_6587;
wire n_1129;
wire n_7781;
wire n_6987;
wire n_602;
wire n_7360;
wire n_11037;
wire n_2181;
wire n_11702;
wire n_6069;
wire n_171;
wire n_2911;
wire n_7497;
wire n_169;
wire n_4655;
wire n_11372;
wire n_1429;
wire n_5706;
wire n_2826;
wire n_7665;
wire n_9354;
wire n_3429;
wire n_10501;
wire n_10817;
wire n_11829;
wire n_2379;
wire n_11517;
wire n_326;
wire n_7793;
wire n_587;
wire n_8355;
wire n_3554;
wire n_1593;
wire n_6991;
wire n_10556;
wire n_1202;
wire n_12741;
wire n_7671;
wire n_7101;
wire n_9436;
wire n_1635;
wire n_7530;
wire n_8489;
wire n_13150;
wire n_5431;
wire n_7248;
wire n_4067;
wire n_4357;
wire n_10350;
wire n_11551;
wire n_12541;
wire n_7204;
wire n_12730;
wire n_9860;
wire n_8649;
wire n_12510;
wire n_12852;
wire n_6887;
wire n_11756;
wire n_10567;
wire n_7578;
wire n_3462;
wire n_7654;
wire n_2851;
wire n_13152;
wire n_8303;
wire n_6153;
wire n_4374;
wire n_5132;
wire n_6637;
wire n_9022;
wire n_8369;
wire n_9238;
wire n_358;
wire n_160;
wire n_8059;
wire n_10230;
wire n_6633;
wire n_12675;
wire n_2420;
wire n_5627;
wire n_9103;
wire n_11031;
wire n_5774;
wire n_11665;
wire n_6579;
wire n_3722;
wire n_186;
wire n_4846;
wire n_4400;
wire n_5798;
wire n_2984;
wire n_11138;
wire n_575;
wire n_11731;
wire n_5187;
wire n_5875;
wire n_9839;
wire n_12821;
wire n_4024;
wire n_8831;
wire n_1508;
wire n_5621;
wire n_5608;
wire n_7900;
wire n_732;
wire n_6569;
wire n_2983;
wire n_6335;
wire n_7120;
wire n_8728;
wire n_2240;
wire n_392;
wire n_10807;
wire n_12478;
wire n_12233;
wire n_2538;
wire n_724;
wire n_3250;
wire n_6789;
wire n_8386;
wire n_12100;
wire n_8853;
wire n_1042;
wire n_4582;
wire n_1728;
wire n_6252;
wire n_557;
wire n_1871;
wire n_4860;
wire n_6211;
wire n_845;
wire n_10511;
wire n_140;
wire n_5844;
wire n_8862;
wire n_3414;
wire n_10580;
wire n_1549;
wire n_4870;
wire n_6164;
wire n_768;
wire n_7576;
wire n_6173;
wire n_8081;
wire n_9675;
wire n_7786;
wire n_11023;
wire n_3651;
wire n_7313;
wire n_10058;
wire n_2102;
wire n_2563;
wire n_10873;
wire n_4989;
wire n_7676;
wire n_11454;
wire n_7757;
wire n_7609;
wire n_3449;
wire n_1683;
wire n_2598;
wire n_1916;
wire n_8900;
wire n_597;
wire n_12523;
wire n_280;
wire n_6934;
wire n_6630;
wire n_10484;
wire n_1187;
wire n_9017;
wire n_4304;
wire n_4558;
wire n_1403;
wire n_6737;
wire n_11744;
wire n_4488;
wire n_3767;
wire n_8396;
wire n_6612;
wire n_8478;
wire n_6606;
wire n_2544;
wire n_6695;
wire n_3550;
wire n_12395;
wire n_8865;
wire n_10288;
wire n_10337;
wire n_4211;
wire n_7779;
wire n_8999;
wire n_6189;
wire n_10388;
wire n_1206;
wire n_11626;
wire n_12148;
wire n_4016;
wire n_11072;
wire n_5867;
wire n_621;
wire n_750;
wire n_5508;
wire n_4656;
wire n_6479;
wire n_10791;
wire n_10506;
wire n_12907;
wire n_3839;
wire n_8497;
wire n_2823;
wire n_10770;
wire n_8820;
wire n_6410;
wire n_9318;
wire n_6158;
wire n_11917;
wire n_5597;
wire n_9028;
wire n_4915;
wire n_4328;
wire n_9492;
wire n_6413;
wire n_6090;
wire n_8020;
wire n_1057;
wire n_9374;
wire n_7419;
wire n_6506;
wire n_2785;
wire n_235;
wire n_5515;
wire n_1997;
wire n_5662;
wire n_2636;
wire n_3131;
wire n_12132;
wire n_710;
wire n_1818;
wire n_3730;
wire n_6935;
wire n_9727;
wire n_10413;
wire n_1298;
wire n_10593;
wire n_13019;
wire n_5862;
wire n_12703;
wire n_13079;
wire n_4397;
wire n_3399;
wire n_2088;
wire n_12182;
wire n_1611;
wire n_12670;
wire n_5050;
wire n_10636;
wire n_12043;
wire n_2740;
wire n_746;
wire n_4808;
wire n_7667;
wire n_5697;
wire n_3416;
wire n_10203;
wire n_3498;
wire n_10980;
wire n_9174;
wire n_5767;
wire n_2401;
wire n_8992;
wire n_1589;
wire n_12708;
wire n_4712;
wire n_8880;
wire n_10369;
wire n_8690;
wire n_2309;
wire n_2900;
wire n_6234;
wire n_2957;
wire n_1740;
wire n_2737;
wire n_6821;
wire n_3994;
wire n_5462;
wire n_9983;
wire n_1497;
wire n_9375;
wire n_10082;
wire n_6688;
wire n_5980;
wire n_8580;
wire n_7818;
wire n_9993;
wire n_8770;
wire n_11721;
wire n_3672;
wire n_7182;
wire n_5318;
wire n_7365;
wire n_6608;
wire n_10467;
wire n_3533;
wire n_9109;
wire n_1622;
wire n_9849;
wire n_6105;
wire n_4725;
wire n_6022;
wire n_11207;
wire n_9856;
wire n_10964;
wire n_4406;
wire n_1694;
wire n_1535;
wire n_3382;
wire n_3132;
wire n_5498;
wire n_2571;
wire n_12493;
wire n_3138;
wire n_13135;
wire n_8075;
wire n_6798;
wire n_10838;
wire n_10530;
wire n_5053;
wire n_7896;
wire n_7841;
wire n_9458;
wire n_12482;
wire n_9237;
wire n_11668;
wire n_7885;
wire n_6860;
wire n_6557;
wire n_8466;
wire n_6753;
wire n_12137;
wire n_2171;
wire n_6527;
wire n_7341;
wire n_11328;
wire n_2988;
wire n_9349;
wire n_12306;
wire n_4908;
wire n_3136;
wire n_1350;
wire n_11200;
wire n_12088;
wire n_11091;
wire n_8094;
wire n_4109;
wire n_4192;
wire n_10940;
wire n_6639;
wire n_4824;
wire n_2037;
wire n_2808;
wire n_4567;
wire n_12096;
wire n_6430;
wire n_12508;
wire n_5150;
wire n_782;
wire n_809;
wire n_8832;
wire n_10987;
wire n_3819;
wire n_4778;
wire n_5477;
wire n_12684;
wire n_1797;
wire n_5175;
wire n_8839;
wire n_7996;
wire n_986;
wire n_2050;
wire n_4595;
wire n_2164;
wire n_4174;
wire n_12891;
wire n_402;
wire n_1870;
wire n_11098;
wire n_11615;
wire n_10533;
wire n_1171;
wire n_11059;
wire n_460;
wire n_5987;
wire n_5179;
wire n_7957;
wire n_1827;
wire n_11965;
wire n_4904;
wire n_10938;
wire n_2187;
wire n_10176;
wire n_7517;
wire n_1152;
wire n_6627;
wire n_8080;
wire n_450;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_5988;
wire n_5585;
wire n_12324;
wire n_12345;
wire n_6058;
wire n_711;
wire n_7745;
wire n_12941;
wire n_3105;
wire n_2872;
wire n_6666;
wire n_3692;
wire n_10927;
wire n_12200;
wire n_4616;
wire n_8321;
wire n_8772;
wire n_8735;
wire n_9954;
wire n_4982;
wire n_370;
wire n_1695;
wire n_11722;
wire n_2046;
wire n_2272;
wire n_8592;
wire n_8786;
wire n_11204;
wire n_8684;
wire n_6190;
wire n_2760;
wire n_1979;
wire n_4643;
wire n_6249;
wire n_2738;
wire n_972;
wire n_12694;
wire n_12701;
wire n_8083;
wire n_12310;
wire n_5348;
wire n_11060;
wire n_10578;
wire n_6594;
wire n_1332;
wire n_9805;
wire n_5480;
wire n_10155;
wire n_4323;
wire n_624;
wire n_8157;
wire n_2346;
wire n_4831;
wire n_7095;
wire n_936;
wire n_3045;
wire n_3821;
wire n_11461;
wire n_10714;
wire n_11701;
wire n_6969;
wire n_885;
wire n_7459;
wire n_6161;
wire n_6615;
wire n_2342;
wire n_2167;
wire n_2970;
wire n_8206;
wire n_3676;
wire n_4896;
wire n_7294;
wire n_2882;
wire n_3675;
wire n_4916;
wire n_4017;
wire n_4260;
wire n_3666;
wire n_9110;
wire n_11811;
wire n_10569;
wire n_2541;
wire n_8622;
wire n_2940;
wire n_5904;
wire n_4739;
wire n_7184;
wire n_9617;
wire n_6607;
wire n_599;
wire n_9335;
wire n_6062;
wire n_7908;
wire n_12550;
wire n_1974;
wire n_4122;
wire n_9452;
wire n_7974;
wire n_7551;
wire n_11427;
wire n_11980;
wire n_10051;
wire n_934;
wire n_4209;
wire n_11255;
wire n_10414;
wire n_8104;
wire n_8344;
wire n_2768;
wire n_3858;
wire n_1341;
wire n_5284;
wire n_11720;
wire n_4298;
wire n_12673;
wire n_2314;
wire n_8120;
wire n_3502;
wire n_8513;
wire n_10120;
wire n_9474;
wire n_5461;
wire n_3003;
wire n_9075;
wire n_12961;
wire n_6482;
wire n_9427;
wire n_11496;
wire n_4128;
wire n_10746;
wire n_12225;
wire n_9188;
wire n_6294;
wire n_543;
wire n_5147;
wire n_9611;
wire n_4271;
wire n_4644;
wire n_9021;
wire n_1355;
wire n_8779;
wire n_9810;
wire n_2258;
wire n_8621;
wire n_5503;
wire n_325;
wire n_5845;
wire n_9250;
wire n_5945;
wire n_804;
wire n_9550;
wire n_11212;
wire n_12884;
wire n_13145;
wire n_10697;
wire n_11714;
wire n_11263;
wire n_10641;
wire n_2390;
wire n_6246;
wire n_8868;
wire n_959;
wire n_2562;
wire n_8134;
wire n_4716;
wire n_4312;
wire n_12207;
wire n_1343;
wire n_1522;
wire n_9975;
wire n_2734;
wire n_7250;
wire n_1782;
wire n_5600;
wire n_5755;
wire n_8762;
wire n_12011;
wire n_8043;
wire n_8694;
wire n_707;
wire n_1900;
wire n_5048;
wire n_6053;
wire n_11994;
wire n_7252;
wire n_3246;
wire n_1548;
wire n_3381;
wire n_1155;
wire n_9207;
wire n_2195;
wire n_3208;
wire n_4944;
wire n_11860;
wire n_11990;
wire n_12837;
wire n_10103;
wire n_5245;
wire n_4343;
wire n_6843;
wire n_10926;
wire n_4715;
wire n_6123;
wire n_8897;
wire n_11000;
wire n_10626;
wire n_6901;
wire n_4935;
wire n_4694;
wire n_11503;
wire n_8191;
wire n_10325;
wire n_6841;
wire n_4672;
wire n_10153;
wire n_8101;
wire n_5054;
wire n_10298;
wire n_2962;
wire n_8171;
wire n_8376;
wire n_5448;
wire n_6922;
wire n_9006;
wire n_2939;
wire n_7698;
wire n_5749;
wire n_1672;
wire n_6774;
wire n_12854;
wire n_6271;
wire n_6489;
wire n_8600;
wire n_1925;
wire n_4407;
wire n_7402;
wire n_8431;
wire n_8710;
wire n_737;
wire n_12806;
wire n_4045;
wire n_3517;
wire n_2945;
wire n_3893;
wire n_3061;
wire n_4598;
wire n_3932;
wire n_3469;
wire n_8599;
wire n_2960;
wire n_8549;
wire n_10172;
wire n_5993;
wire n_8054;
wire n_11273;
wire n_10400;
wire n_6716;
wire n_9637;
wire n_11636;
wire n_138;
wire n_3258;
wire n_9418;
wire n_8616;
wire n_4524;
wire n_3143;
wire n_6020;
wire n_12472;
wire n_9177;
wire n_9060;
wire n_13105;
wire n_11947;
wire n_9096;
wire n_9081;
wire n_11697;
wire n_333;
wire n_13076;
wire n_4084;
wire n_3149;
wire n_6844;
wire n_9236;
wire n_11762;
wire n_11969;
wire n_12950;
wire n_8628;
wire n_7914;
wire n_3365;
wire n_6521;
wire n_7891;
wire n_3379;
wire n_13028;
wire n_8857;
wire n_8517;
wire n_459;
wire n_4850;
wire n_8547;
wire n_10156;
wire n_4424;
wire n_9040;
wire n_7113;
wire n_9607;
wire n_3008;
wire n_1751;
wire n_6162;
wire n_10433;
wire n_2840;
wire n_6779;
wire n_8010;
wire n_285;
wire n_3939;
wire n_4776;
wire n_6432;
wire n_9116;
wire n_1375;
wire n_10774;
wire n_3972;
wire n_12332;
wire n_4153;
wire n_10901;
wire n_11034;
wire n_11983;
wire n_10549;
wire n_10839;
wire n_12115;
wire n_11813;
wire n_3506;
wire n_1650;
wire n_1962;
wire n_3855;
wire n_7216;
wire n_12762;
wire n_11499;
wire n_1928;
wire n_10825;
wire n_3091;
wire n_4317;
wire n_8275;
wire n_4723;
wire n_6198;
wire n_4269;
wire n_5418;
wire n_6543;
wire n_9830;
wire n_6762;
wire n_6178;
wire n_9621;
wire n_4088;
wire n_3398;
wire n_5685;
wire n_10761;
wire n_2761;
wire n_2793;
wire n_3776;
wire n_3711;
wire n_4235;
wire n_5459;
wire n_9035;
wire n_11579;
wire n_1019;
wire n_10398;
wire n_8291;
wire n_4170;
wire n_4143;
wire n_729;
wire n_876;
wire n_774;
wire n_11535;
wire n_3642;
wire n_12558;
wire n_2845;
wire n_4650;
wire n_11984;
wire n_11948;
wire n_7706;
wire n_438;
wire n_4719;
wire n_5173;
wire n_7477;
wire n_1860;
wire n_5016;
wire n_1904;
wire n_12975;
wire n_2874;
wire n_1200;
wire n_2588;
wire n_11402;
wire n_479;
wire n_6458;
wire n_1353;
wire n_1777;
wire n_4967;
wire n_7642;
wire n_9678;
wire n_11401;
wire n_8247;
wire n_6577;
wire n_12506;
wire n_6740;
wire n_3308;
wire n_12718;
wire n_1113;
wire n_1600;
wire n_12956;
wire n_2253;
wire n_11510;
wire n_6315;
wire n_2366;
wire n_10581;
wire n_12638;
wire n_4912;
wire n_4799;
wire n_2261;
wire n_9284;
wire n_12736;
wire n_4423;
wire n_5086;
wire n_5283;
wire n_9111;
wire n_2210;
wire n_7156;
wire n_4735;
wire n_9163;
wire n_3602;
wire n_187;
wire n_3300;
wire n_2978;
wire n_12086;
wire n_2516;
wire n_1050;
wire n_1411;
wire n_5170;
wire n_7604;
wire n_6910;
wire n_6262;
wire n_2827;
wire n_1177;
wire n_7703;
wire n_3515;
wire n_1150;
wire n_9606;
wire n_6319;
wire n_566;
wire n_1023;
wire n_2951;
wire n_10470;
wire n_1118;
wire n_11589;
wire n_194;
wire n_2949;
wire n_10297;
wire n_11246;
wire n_12553;
wire n_1807;
wire n_12350;
wire n_12542;
wire n_5028;
wire n_5839;
wire n_1814;
wire n_1631;
wire n_1879;
wire n_6536;
wire n_12747;
wire n_256;
wire n_440;
wire n_6175;
wire n_3806;
wire n_7040;
wire n_10625;
wire n_8827;
wire n_8280;
wire n_12561;
wire n_12390;
wire n_5514;
wire n_2931;
wire n_209;
wire n_367;
wire n_8388;
wire n_12849;
wire n_2569;
wire n_10235;
wire n_11312;
wire n_3866;
wire n_6978;
wire n_9589;
wire n_5351;
wire n_5909;
wire n_9344;
wire n_671;
wire n_12805;
wire n_10865;
wire n_9549;
wire n_6093;
wire n_11649;
wire n_4543;
wire n_10445;
wire n_740;
wire n_7378;
wire n_703;
wire n_10738;
wire n_12866;
wire n_4157;
wire n_9798;
wire n_6845;
wire n_8988;
wire n_9190;
wire n_6947;
wire n_11612;
wire n_4229;
wire n_9482;
wire n_5293;
wire n_12447;
wire n_12296;
wire n_8203;
wire n_6099;
wire n_12900;
wire n_3865;
wire n_4073;
wire n_1324;
wire n_8569;
wire n_3629;
wire n_1435;
wire n_5400;
wire n_3920;
wire n_969;
wire n_4892;
wire n_3255;
wire n_6140;
wire n_8877;
wire n_9412;
wire n_1401;
wire n_7498;
wire n_10679;
wire n_1516;
wire n_11323;
wire n_10799;
wire n_3846;
wire n_6321;
wire n_12914;
wire n_11916;
wire n_180;
wire n_3512;
wire n_6819;
wire n_5201;
wire n_2029;
wire n_7501;
wire n_9506;
wire n_10136;
wire n_10421;
wire n_5890;
wire n_6415;
wire n_10976;
wire n_6465;
wire n_9447;
wire n_4439;
wire n_1394;
wire n_10585;
wire n_12764;
wire n_1326;
wire n_4783;
wire n_11356;
wire n_1379;
wire n_214;
wire n_12948;
wire n_7931;
wire n_8688;
wire n_10828;
wire n_9092;
wire n_10034;
wire n_935;
wire n_9451;
wire n_4910;
wire n_11148;
wire n_12409;
wire n_11625;
wire n_12300;
wire n_1130;
wire n_6899;
wire n_3083;
wire n_7549;
wire n_10692;
wire n_7373;
wire n_7895;
wire n_11281;
wire n_13056;
wire n_676;
wire n_832;
wire n_11280;
wire n_12337;
wire n_6592;
wire n_3049;
wire n_8686;
wire n_12239;
wire n_8871;
wire n_9712;
wire n_6626;
wire n_8585;
wire n_8951;
wire n_5389;
wire n_5142;
wire n_11114;
wire n_9011;
wire n_8418;
wire n_3830;
wire n_7740;
wire n_8403;
wire n_3679;
wire n_5891;
wire n_13050;
wire n_7613;
wire n_3541;
wire n_11493;
wire n_6101;
wire n_9220;
wire n_3117;
wire n_5935;
wire n_7556;
wire n_10528;
wire n_10860;
wire n_12763;
wire n_4930;
wire n_372;
wire n_8588;
wire n_314;
wire n_378;
wire n_11339;
wire n_5623;
wire n_12273;
wire n_8564;
wire n_11943;
wire n_6944;
wire n_9121;
wire n_10471;
wire n_338;
wire n_1283;
wire n_2385;
wire n_4112;
wire n_12712;
wire n_506;
wire n_11220;
wire n_360;
wire n_2149;
wire n_9012;
wire n_2396;
wire n_4557;
wire n_13012;
wire n_4917;
wire n_8698;
wire n_895;
wire n_8924;
wire n_12584;
wire n_2450;
wire n_3739;
wire n_4432;
wire n_2284;
wire n_10376;
wire n_12752;
wire n_4352;
wire n_7515;
wire n_6928;
wire n_4416;
wire n_10880;
wire n_4593;
wire n_7238;
wire n_344;
wire n_9994;
wire n_2769;
wire n_4465;
wire n_3622;
wire n_8780;
wire n_7309;
wire n_5114;
wire n_7958;
wire n_4980;
wire n_8047;
wire n_11596;
wire n_1392;
wire n_8559;
wire n_5693;
wire n_4495;
wire n_6273;
wire n_11885;
wire n_5117;
wire n_1924;
wire n_5663;
wire n_525;
wire n_2463;
wire n_3363;
wire n_7572;
wire n_8214;
wire n_10224;
wire n_11955;
wire n_12777;
wire n_1677;
wire n_5990;
wire n_611;
wire n_7043;
wire n_10777;
wire n_3721;
wire n_11462;
wire n_3062;
wire n_11732;
wire n_2679;
wire n_5024;
wire n_9391;
wire n_7760;
wire n_4559;
wire n_8514;
wire n_9134;
wire n_9753;
wire n_12819;
wire n_8722;
wire n_11654;
wire n_12268;
wire n_10214;
wire n_8589;
wire n_8241;
wire n_838;
wire n_12077;
wire n_3969;
wire n_12982;
wire n_3336;
wire n_7573;
wire n_4160;
wire n_8442;
wire n_4231;
wire n_6281;
wire n_11619;
wire n_10649;
wire n_7364;
wire n_2952;
wire n_5647;
wire n_1017;
wire n_13133;
wire n_4256;
wire n_2779;
wire n_4938;
wire n_5396;
wire n_9572;
wire n_8608;
wire n_5203;
wire n_12874;
wire n_12534;
wire n_6846;
wire n_10469;
wire n_445;
wire n_11194;
wire n_9229;
wire n_11480;
wire n_6311;
wire n_930;
wire n_7590;
wire n_9342;
wire n_12237;
wire n_2620;
wire n_5162;
wire n_6134;
wire n_9329;
wire n_1945;
wire n_5426;
wire n_10175;
wire n_1656;
wire n_5803;
wire n_11481;
wire n_2112;
wire n_1464;
wire n_2430;
wire n_653;
wire n_9868;
wire n_11375;
wire n_1414;
wire n_5285;
wire n_11267;
wire n_9602;
wire n_7048;
wire n_6886;
wire n_2721;
wire n_944;
wire n_4335;
wire n_9311;
wire n_12275;
wire n_2034;
wire n_576;
wire n_6593;
wire n_8630;
wire n_270;
wire n_2683;
wire n_12376;
wire n_563;
wire n_9884;
wire n_5365;
wire n_13114;
wire n_9876;
wire n_8583;
wire n_2744;
wire n_1011;
wire n_4521;
wire n_1566;
wire n_8405;
wire n_8145;
wire n_10447;
wire n_9260;
wire n_7176;
wire n_8928;
wire n_7682;
wire n_9353;
wire n_11350;
wire n_13054;
wire n_626;
wire n_990;
wire n_11925;
wire n_6231;
wire n_8948;
wire n_10406;
wire n_8672;
wire n_3204;
wire n_1104;
wire n_5715;
wire n_12509;
wire n_4920;
wire n_8295;
wire n_6932;
wire n_6746;
wire n_11985;
wire n_498;
wire n_8447;
wire n_7901;
wire n_870;
wire n_5395;
wire n_1253;
wire n_10522;
wire n_366;
wire n_6443;
wire n_5709;
wire n_7658;
wire n_11782;
wire n_1693;
wire n_6446;
wire n_10278;
wire n_10055;
wire n_10979;
wire n_7980;
wire n_3256;
wire n_348;
wire n_3802;
wire n_6996;
wire n_8828;
wire n_9430;
wire n_7218;
wire n_376;
wire n_11407;
wire n_2118;
wire n_2111;
wire n_390;
wire n_9750;
wire n_9749;
wire n_2915;
wire n_12710;
wire n_1148;
wire n_6749;
wire n_2188;
wire n_9263;
wire n_11082;
wire n_8440;
wire n_1989;
wire n_7005;
wire n_10408;
wire n_2802;
wire n_8572;
wire n_10798;
wire n_10965;
wire n_7732;
wire n_6337;
wire n_3643;
wire n_6181;
wire n_7447;
wire n_2425;
wire n_9776;
wire n_11911;
wire n_6777;
wire n_4265;
wire n_11987;
wire n_11442;
wire n_8227;
wire n_12936;
wire n_12721;
wire n_2950;
wire n_5634;
wire n_5672;
wire n_719;
wire n_8475;
wire n_3060;
wire n_11730;
wire n_10482;
wire n_3098;
wire n_6924;
wire n_8029;
wire n_9804;
wire n_4105;
wire n_1851;
wire n_1090;
wire n_4861;
wire n_9304;
wire n_5799;
wire n_8859;
wire n_8380;
wire n_4064;
wire n_7405;
wire n_12039;
wire n_4926;
wire n_1518;
wire n_11388;
wire n_1362;
wire n_11651;
wire n_3123;
wire n_8314;
wire n_3380;
wire n_9386;
wire n_10154;
wire n_5617;
wire n_1829;
wire n_7922;
wire n_13089;
wire n_10377;
wire n_5580;
wire n_5266;
wire n_1450;
wire n_4828;
wire n_1638;
wire n_9926;
wire n_10033;
wire n_3038;
wire n_570;
wire n_11121;
wire n_11270;
wire n_1789;
wire n_12329;
wire n_6310;
wire n_11689;
wire n_620;
wire n_10003;
wire n_519;
wire n_8311;
wire n_2523;
wire n_10858;
wire n_10321;
wire n_5450;
wire n_2413;
wire n_3769;
wire n_12253;
wire n_1482;
wire n_11147;
wire n_12928;
wire n_5310;
wire n_9661;
wire n_9843;
wire n_9877;
wire n_8764;
wire n_3863;
wire n_3669;
wire n_6953;
wire n_3130;
wire n_4316;
wire n_5722;
wire n_4640;
wire n_5122;
wire n_13001;
wire n_5390;
wire n_9901;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_2805;
wire n_5593;
wire n_12990;
wire n_6683;
wire n_4769;
wire n_10683;
wire n_5764;
wire n_9834;
wire n_8934;
wire n_13059;
wire n_2282;
wire n_6365;
wire n_4628;
wire n_6920;
wire n_9921;
wire n_2047;
wire n_12318;
wire n_8407;
wire n_6229;
wire n_5385;
wire n_8567;
wire n_11817;
wire n_1609;
wire n_8729;
wire n_11288;
wire n_12772;
wire n_10359;
wire n_3344;
wire n_5237;
wire n_2334;
wire n_5133;
wire n_409;
wire n_11042;
wire n_1763;
wire n_5322;
wire n_6907;
wire n_10726;
wire n_3989;
wire n_7144;
wire n_2490;
wire n_7089;
wire n_7286;
wire n_11479;
wire n_11737;
wire n_4460;
wire n_4108;
wire n_8048;
wire n_635;
wire n_12028;
wire n_3786;
wire n_3841;
wire n_7072;
wire n_13016;
wire n_11272;
wire n_13095;
wire n_4254;
wire n_8253;
wire n_6177;
wire n_1996;
wire n_6332;
wire n_2867;
wire n_1442;
wire n_2726;
wire n_4303;
wire n_5853;
wire n_12048;
wire n_8283;
wire n_5982;
wire n_1158;
wire n_10930;
wire n_2248;
wire n_11600;
wire n_8749;
wire n_8088;
wire n_7403;
wire n_10722;
wire n_5011;
wire n_10666;
wire n_7338;
wire n_5917;
wire n_7129;
wire n_2662;
wire n_4909;
wire n_3147;
wire n_12057;
wire n_6696;
wire n_753;
wire n_3925;
wire n_9882;
wire n_9527;
wire n_3180;
wire n_8566;
wire n_7343;
wire n_2795;
wire n_12766;
wire n_3472;
wire n_8516;
wire n_8302;
wire n_10637;
wire n_8317;
wire n_5376;
wire n_12229;
wire n_5106;
wire n_269;
wire n_6116;
wire n_9205;
wire n_359;
wire n_9511;
wire n_8167;
wire n_7859;
wire n_7492;
wire n_7872;
wire n_6730;
wire n_7972;
wire n_11254;
wire n_1479;
wire n_4768;
wire n_11617;
wire n_1675;
wire n_9071;
wire n_7916;
wire n_3717;
wire n_9368;
wire n_10415;
wire n_7694;
wire n_5561;
wire n_7480;
wire n_13069;
wire n_11711;
wire n_5410;
wire n_571;
wire n_2215;
wire n_12362;
wire n_404;
wire n_8944;
wire n_6167;
wire n_158;
wire n_1884;
wire n_11931;
wire n_8008;
wire n_10023;
wire n_10999;
wire n_6170;
wire n_665;
wire n_8109;
wire n_9459;
wire n_2055;
wire n_5156;
wire n_12780;
wire n_2553;
wire n_6307;
wire n_149;
wire n_10410;
wire n_632;
wire n_6094;
wire n_9098;
wire n_2038;
wire n_7987;
wire n_7483;
wire n_4447;
wire n_9133;
wire n_12664;
wire n_7434;
wire n_4826;
wire n_3445;
wire n_9009;
wire n_6155;
wire n_7269;
wire n_9777;
wire n_373;
wire n_9504;
wire n_8975;
wire n_6267;
wire n_9063;
wire n_7787;
wire n_1833;
wire n_3903;
wire n_12360;
wire n_5998;
wire n_1494;
wire n_2325;
wire n_9268;
wire n_1850;
wire n_5304;
wire n_3854;
wire n_3235;
wire n_6568;
wire n_8673;
wire n_7507;
wire n_7159;
wire n_11305;
wire n_5378;
wire n_6028;
wire n_9101;
wire n_1417;
wire n_10456;
wire n_6261;
wire n_3673;
wire n_4281;
wire n_5916;
wire n_681;
wire n_11907;
wire n_4648;
wire n_10096;
wire n_3094;
wire n_10025;
wire n_412;
wire n_10627;
wire n_10475;
wire n_10189;
wire n_8697;
wire n_6299;
wire n_6813;
wire n_965;
wire n_8825;
wire n_1428;
wire n_12969;
wire n_1576;
wire n_1856;
wire n_11753;
wire n_2077;
wire n_7425;
wire n_12260;
wire n_12016;
wire n_6669;
wire n_8581;
wire n_8266;
wire n_5691;
wire n_1059;
wire n_12457;
wire n_4951;
wire n_8981;
wire n_422;
wire n_8420;
wire n_4957;
wire n_8297;
wire n_11150;
wire n_3079;
wire n_165;
wire n_4360;
wire n_8771;
wire n_10881;
wire n_540;
wire n_4039;
wire n_457;
wire n_3070;
wire n_3800;
wire n_4566;
wire n_3263;
wire n_12939;
wire n_6316;
wire n_6292;
wire n_4853;
wire n_9726;
wire n_1748;
wire n_10404;
wire n_8639;
wire n_8058;
wire n_8138;
wire n_9308;
wire n_3504;
wire n_6638;
wire n_12779;
wire n_11838;
wire n_10508;
wire n_531;
wire n_7719;
wire n_4272;
wire n_10811;
wire n_8333;
wire n_2930;
wire n_5615;
wire n_1025;
wire n_6220;
wire n_7562;
wire n_3111;
wire n_12816;
wire n_336;
wire n_6985;
wire n_7619;
wire n_12783;
wire n_7170;
wire n_9211;
wire n_12019;
wire n_1885;
wire n_8176;
wire n_8124;
wire n_8823;
wire n_7366;
wire n_9395;
wire n_5269;
wire n_10891;
wire n_11457;
wire n_12751;
wire n_9026;
wire n_3054;
wire n_10803;
wire n_1538;
wire n_8147;
wire n_1240;
wire n_5468;
wire n_6188;
wire n_4730;
wire n_5399;
wire n_8127;
wire n_9402;
wire n_1234;
wire n_5262;
wire n_10700;
wire n_3254;
wire n_3684;
wire n_7938;
wire n_4670;
wire n_10968;
wire n_4882;
wire n_11695;
wire n_4620;
wire n_3152;
wire n_8458;
wire n_4738;
wire n_3579;
wire n_5421;
wire n_7935;
wire n_6772;
wire n_8113;
wire n_3335;
wire n_9716;
wire n_4177;
wire n_3783;
wire n_700;
wire n_1307;
wire n_3178;
wire n_11453;
wire n_4127;
wire n_5206;
wire n_6077;
wire n_1003;
wire n_5713;
wire n_11512;
wire n_5256;
wire n_168;
wire n_6318;
wire n_2353;
wire n_11970;
wire n_4099;
wire n_7918;
wire n_4517;
wire n_4168;
wire n_5188;
wire n_6916;
wire n_1738;
wire n_4490;
wire n_1575;
wire n_6651;
wire n_12308;
wire n_10290;
wire n_1923;
wire n_10783;
wire n_2260;
wire n_10147;
wire n_11862;
wire n_12163;
wire n_10725;
wire n_3952;
wire n_11523;
wire n_7845;
wire n_12688;
wire n_5550;
wire n_12944;
wire n_3911;
wire n_8290;
wire n_7536;
wire n_7472;
wire n_9433;
wire n_9737;
wire n_9298;
wire n_11660;
wire n_1688;
wire n_4285;
wire n_3465;
wire n_10812;
wire n_1743;
wire n_12297;
wire n_6366;
wire n_6230;
wire n_2997;
wire n_6604;
wire n_1991;
wire n_2386;
wire n_5161;
wire n_5373;
wire n_1724;
wire n_10001;
wire n_3708;
wire n_11107;
wire n_4078;
wire n_9301;
wire n_12145;
wire n_3046;
wire n_11088;
wire n_2956;
wire n_5573;
wire n_1553;
wire n_5939;
wire n_5509;
wire n_5382;
wire n_6391;
wire n_8160;
wire n_10284;
wire n_12757;
wire n_12054;
wire n_5659;
wire n_8099;
wire n_11595;
wire n_8840;
wire n_3619;
wire n_11405;
wire n_1415;
wire n_5881;
wire n_8522;
wire n_12971;
wire n_1370;
wire n_7942;
wire n_1786;
wire n_8578;
wire n_6473;
wire n_7222;
wire n_13103;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_10046;
wire n_12328;
wire n_2291;
wire n_415;
wire n_11318;
wire n_9083;
wire n_1371;
wire n_7725;
wire n_383;
wire n_2886;
wire n_2974;
wire n_4213;
wire n_10977;
wire n_200;
wire n_11299;
wire n_2184;
wire n_10397;
wire n_2982;
wire n_6483;
wire n_1803;
wire n_10615;
wire n_10994;
wire n_11542;
wire n_4065;
wire n_5863;
wire n_229;
wire n_7647;
wire n_10385;
wire n_10936;
wire n_8626;
wire n_2645;
wire n_12442;
wire n_3904;
wire n_8611;
wire n_8036;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_8819;
wire n_11485;
wire n_12426;
wire n_2630;
wire n_1444;
wire n_9835;
wire n_1603;
wire n_7300;
wire n_12839;
wire n_6697;
wire n_9054;
wire n_7875;
wire n_13153;
wire n_6975;
wire n_2470;
wire n_4446;
wire n_1263;
wire n_10532;
wire n_4417;
wire n_5466;
wire n_7643;
wire n_13073;
wire n_11048;
wire n_4733;
wire n_6728;
wire n_6729;
wire n_4764;
wire n_1261;
wire n_3879;
wire n_11240;
wire n_2286;
wire n_4743;
wire n_10207;
wire n_2018;
wire n_3080;
wire n_1903;
wire n_1143;
wire n_10401;
wire n_11634;
wire n_12580;
wire n_5955;
wire n_7242;
wire n_10013;
wire n_10771;
wire n_658;
wire n_1874;
wire n_11487;
wire n_2865;
wire n_2825;
wire n_8441;
wire n_11441;
wire n_2013;
wire n_6076;
wire n_8933;
wire n_2044;
wire n_3023;
wire n_3232;
wire n_693;
wire n_1056;
wire n_7778;
wire n_758;
wire n_12844;
wire n_5851;
wire n_7073;
wire n_2256;
wire n_9755;
wire n_11287;
wire n_943;
wire n_4060;
wire n_5110;
wire n_9774;
wire n_8397;
wire n_4879;
wire n_10139;
wire n_6390;
wire n_5796;
wire n_10104;
wire n_772;
wire n_8726;
wire n_12986;
wire n_11381;
wire n_2806;
wire n_6665;
wire n_8797;
wire n_10723;
wire n_7224;
wire n_12441;
wire n_770;
wire n_9117;
wire n_9720;
wire n_3028;
wire n_7746;
wire n_3662;
wire n_9381;
wire n_2981;
wire n_10169;
wire n_6958;
wire n_3076;
wire n_12049;
wire n_12690;
wire n_886;
wire n_7563;
wire n_343;
wire n_12475;
wire n_3624;
wire n_1345;
wire n_1820;
wire n_4556;
wire n_12516;
wire n_11765;
wire n_6549;
wire n_539;
wire n_8414;
wire n_6297;
wire n_6523;
wire n_6653;
wire n_8434;
wire n_12302;
wire n_10477;
wire n_6096;
wire n_4117;
wire n_7853;
wire n_12526;
wire n_4687;
wire n_2836;
wire n_7531;
wire n_12377;
wire n_638;
wire n_1404;
wire n_8890;
wire n_5492;
wire n_5995;
wire n_9965;
wire n_8615;
wire n_11062;
wire n_2378;
wire n_7721;
wire n_887;
wire n_7192;
wire n_5905;
wire n_11933;
wire n_11206;
wire n_9887;
wire n_9149;
wire n_2655;
wire n_4600;
wire n_11593;
wire n_7035;
wire n_6193;
wire n_6501;
wire n_1467;
wire n_8316;
wire n_4250;
wire n_9990;
wire n_5829;
wire n_3906;
wire n_10005;
wire n_224;
wire n_11786;
wire n_12737;
wire n_8057;
wire n_12905;
wire n_11426;
wire n_4954;
wire n_5191;
wire n_1231;
wire n_2599;
wire n_8505;
wire n_9273;
wire n_3963;
wire n_3368;
wire n_7884;
wire n_9345;
wire n_11258;
wire n_11550;
wire n_2370;
wire n_2612;
wire n_8970;
wire n_7527;
wire n_7417;
wire n_13061;
wire n_9682;
wire n_2591;
wire n_4881;
wire n_1815;
wire n_12513;
wire n_2214;
wire n_4253;
wire n_10640;
wire n_407;
wire n_913;
wire n_6582;
wire n_5734;
wire n_2593;
wire n_4255;
wire n_867;
wire n_4071;
wire n_10729;
wire n_12545;
wire n_7388;
wire n_3568;
wire n_1230;
wire n_3850;
wire n_11657;
wire n_9924;
wire n_8717;
wire n_5770;
wire n_1333;
wire n_2496;
wire n_5705;
wire n_3313;
wire n_4605;
wire n_9064;
wire n_3189;
wire n_7635;
wire n_5525;
wire n_13102;
wire n_163;
wire n_1644;
wire n_11268;
wire n_12753;
wire n_2725;
wire n_2277;
wire n_4691;
wire n_7090;
wire n_9254;
wire n_1558;
wire n_12894;
wire n_1732;
wire n_2300;
wire n_3943;
wire n_8571;
wire n_11641;
wire n_11501;
wire n_4305;
wire n_7227;
wire n_10492;
wire n_7415;
wire n_11211;
wire n_824;
wire n_6745;
wire n_6972;
wire n_12514;
wire n_10048;
wire n_4297;
wire n_8030;
wire n_9247;
wire n_6052;
wire n_8378;
wire n_8687;
wire n_2907;
wire n_577;
wire n_5374;
wire n_10526;
wire n_5575;
wire n_8725;
wire n_12010;
wire n_1843;
wire n_619;
wire n_5675;
wire n_9738;
wire n_9570;
wire n_12026;
wire n_4227;
wire n_521;
wire n_2778;
wire n_12356;
wire n_11857;
wire n_395;
wire n_1909;
wire n_6240;
wire n_11077;
wire n_8243;
wire n_6347;
wire n_8633;
wire n_5020;
wire n_9846;
wire n_7689;
wire n_9593;
wire n_6511;
wire n_606;
wire n_5297;
wire n_7121;
wire n_1123;
wire n_1309;
wire n_9469;
wire n_10764;
wire n_9677;
wire n_2961;
wire n_916;
wire n_3934;
wire n_4033;
wire n_4415;
wire n_6515;
wire n_7099;
wire n_483;
wire n_6804;
wire n_1970;
wire n_8449;
wire n_6358;
wire n_630;
wire n_2059;
wire n_2669;
wire n_4094;
wire n_6603;
wire n_4765;
wire n_2546;
wire n_3193;
wire n_2522;
wire n_476;
wire n_4364;
wire n_7534;
wire n_9406;
wire n_11313;
wire n_1957;
wire n_8201;
wire n_8967;
wire n_4354;
wire n_6986;
wire n_4732;
wire n_3912;
wire n_10438;
wire n_9322;
wire n_3118;
wire n_8801;
wire n_5959;
wire n_11201;
wire n_3720;
wire n_10531;
wire n_1907;
wire n_2529;
wire n_8031;
wire n_8918;
wire n_264;
wire n_12878;
wire n_9348;
wire n_12188;
wire n_860;
wire n_8219;
wire n_1530;
wire n_8696;
wire n_4745;
wire n_938;
wire n_1302;
wire n_6396;
wire n_8932;
wire n_5642;
wire n_9232;
wire n_10575;
wire n_12630;
wire n_4581;
wire n_6890;
wire n_549;
wire n_11028;
wire n_12171;
wire n_4377;
wire n_12299;
wire n_12022;
wire n_9249;
wire n_12935;
wire n_7827;
wire n_2143;
wire n_8180;
wire n_905;
wire n_10741;
wire n_6109;
wire n_10760;
wire n_4792;
wire n_12425;
wire n_9444;
wire n_7731;
wire n_1680;
wire n_3842;
wire n_10772;
wire n_322;
wire n_993;
wire n_11527;
wire n_689;
wire n_2031;
wire n_7114;
wire n_4878;
wire n_1605;
wire n_3514;
wire n_11327;
wire n_10915;
wire n_4979;
wire n_1988;
wire n_9535;
wire n_558;
wire n_6770;
wire n_2654;
wire n_7943;
wire n_3036;
wire n_11743;
wire n_8892;
wire n_12199;
wire n_5302;
wire n_12000;
wire n_966;
wire n_4511;
wire n_2908;
wire n_9707;
wire n_12490;
wire n_3357;
wire n_692;
wire n_5639;
wire n_5781;
wire n_1233;
wire n_3895;
wire n_487;
wire n_8943;
wire n_8486;
wire n_241;
wire n_10279;
wire n_4520;
wire n_5299;
wire n_12829;
wire n_3455;
wire n_4118;
wire n_4503;
wire n_2176;
wire n_10680;
wire n_2459;
wire n_10127;
wire n_1111;
wire n_3599;
wire n_5543;
wire n_1251;
wire n_5361;
wire n_11610;
wire n_7081;
wire n_2711;
wire n_11814;
wire n_7132;
wire n_12255;
wire n_12739;
wire n_13015;
wire n_4199;
wire n_5885;
wire n_6663;
wire n_1912;
wire n_9723;
wire n_5356;
wire n_12609;
wire n_7319;
wire n_4441;
wire n_1982;
wire n_3872;
wire n_3772;
wire n_5458;
wire n_7644;
wire n_1312;
wire n_11176;
wire n_11473;
wire n_9883;
wire n_11135;
wire n_8155;
wire n_11360;
wire n_5668;
wire n_11275;
wire n_11868;
wire n_5038;
wire n_268;
wire n_1760;
wire n_5330;
wire n_4585;
wire n_7199;
wire n_2664;
wire n_1664;
wire n_1722;
wire n_10039;
wire n_11726;
wire n_10854;
wire n_11358;
wire n_5463;
wire n_3022;
wire n_8098;
wire n_12574;
wire n_12700;
wire n_247;
wire n_12904;
wire n_9191;
wire n_8833;
wire n_5489;
wire n_1165;
wire n_5892;
wire n_7828;
wire n_10142;
wire n_4773;
wire n_7940;
wire n_9918;
wire n_7910;
wire n_5654;
wire n_6782;
wire n_2008;
wire n_6009;
wire n_2192;
wire n_3281;
wire n_2345;
wire n_9034;
wire n_328;
wire n_1386;
wire n_6503;
wire n_6376;
wire n_4427;
wire n_7084;
wire n_5923;
wire n_9390;
wire n_5113;
wire n_12017;
wire n_12888;
wire n_10069;
wire n_5479;
wire n_3549;
wire n_5714;
wire n_8541;
wire n_2804;
wire n_2453;
wire n_8074;
wire n_8485;
wire n_8860;
wire n_2676;
wire n_5510;
wire n_3940;
wire n_6621;
wire n_11958;
wire n_7001;
wire n_9650;
wire n_4822;
wire n_1214;
wire n_13070;
wire n_690;
wire n_850;
wire n_8271;
wire n_5692;
wire n_8473;
wire n_4800;
wire n_9266;
wire n_1157;
wire n_3453;
wire n_12728;
wire n_5555;
wire n_3410;
wire n_10027;
wire n_12784;
wire n_1752;
wire n_1813;
wire n_3768;
wire n_4958;
wire n_2810;
wire n_4043;
wire n_2319;
wire n_5441;
wire n_6783;
wire n_9664;
wire n_825;
wire n_12458;
wire n_12259;
wire n_6066;
wire n_12877;
wire n_8699;
wire n_3785;
wire n_6897;
wire n_2963;
wire n_10616;
wire n_8587;
wire n_9619;
wire n_11171;
wire n_5366;
wire n_2602;
wire n_6925;
wire n_6878;
wire n_3873;
wire n_8225;
wire n_9078;
wire n_9536;
wire n_2980;
wire n_696;
wire n_4886;
wire n_9931;
wire n_1082;
wire n_1317;
wire n_3227;
wire n_2733;
wire n_3289;
wire n_6296;
wire n_9187;
wire n_7708;
wire n_4055;
wire n_12610;
wire n_2178;
wire n_11671;
wire n_10328;
wire n_5968;
wire n_11251;
wire n_12293;
wire n_11063;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_10753;
wire n_6497;
wire n_8319;
wire n_9989;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_7108;
wire n_12853;
wire n_6470;
wire n_12942;
wire n_11598;
wire n_1796;
wire n_8368;
wire n_9259;
wire n_8322;
wire n_7333;
wire n_11879;
wire n_2082;
wire n_3519;
wire n_6187;
wire n_7876;
wire n_12397;
wire n_8546;
wire n_10963;
wire n_8300;
wire n_7371;
wire n_9378;
wire n_8152;
wire n_678;
wire n_10826;
wire n_7463;
wire n_12206;
wire n_8525;
wire n_6573;
wire n_9656;
wire n_7634;
wire n_5078;
wire n_3707;
wire n_283;
wire n_8148;
wire n_11400;
wire n_8150;
wire n_3578;
wire n_909;
wire n_11440;
wire n_12596;
wire n_6693;
wire n_10483;
wire n_12160;
wire n_4737;
wire n_590;
wire n_11563;
wire n_4925;
wire n_9620;
wire n_4116;
wire n_5415;
wire n_8986;
wire n_362;
wire n_7285;
wire n_11337;
wire n_12444;
wire n_12005;
wire n_5419;
wire n_11243;
wire n_1990;
wire n_3805;
wire n_8929;
wire n_9360;
wire n_12697;
wire n_7260;
wire n_2943;
wire n_5205;
wire n_12778;
wire n_12485;
wire n_6409;
wire n_11939;
wire n_1634;
wire n_3252;
wire n_627;
wire n_3253;
wire n_7954;
wire n_9824;
wire n_1465;
wire n_11119;
wire n_342;
wire n_2622;
wire n_7951;
wire n_2658;
wire n_7552;
wire n_8096;
wire n_2665;
wire n_11468;
wire n_12166;
wire n_2133;
wire n_1712;
wire n_6130;
wire n_4603;
wire n_8233;
wire n_7273;
wire n_9683;
wire n_1523;
wire n_10646;
wire n_7231;
wire n_1627;
wire n_5080;
wire n_5976;
wire n_11704;
wire n_3128;
wire n_1527;
wire n_495;
wire n_5732;
wire n_5372;
wire n_11878;
wire n_2691;
wire n_840;
wire n_2913;
wire n_4471;
wire n_7772;
wire n_7449;
wire n_2230;
wire n_8763;
wire n_12800;
wire n_1969;
wire n_2690;
wire n_5208;
wire n_8679;
wire n_1565;
wire n_7239;
wire n_1493;
wire n_9848;
wire n_11962;
wire n_5690;
wire n_9227;
wire n_8187;
wire n_10751;
wire n_7050;
wire n_10240;
wire n_10691;
wire n_8996;
wire n_9399;
wire n_2573;
wire n_2646;
wire n_2535;
wire n_9561;
wire n_6623;
wire n_10378;
wire n_12070;
wire n_9714;
wire n_1364;
wire n_9740;
wire n_3078;
wire n_9773;
wire n_2436;
wire n_10313;
wire n_615;
wire n_3838;
wire n_12947;
wire n_5371;
wire n_4651;
wire n_9745;
wire n_3941;
wire n_3793;
wire n_10216;
wire n_11928;
wire n_8139;
wire n_9764;
wire n_4854;
wire n_5071;
wire n_3789;
wire n_605;
wire n_1514;
wire n_7597;
wire n_10150;
wire n_12354;
wire n_5801;
wire n_12666;
wire n_6047;
wire n_12581;
wire n_8292;
wire n_12631;
wire n_3037;
wire n_1646;
wire n_10133;
wire n_3729;
wire n_8601;
wire n_10773;
wire n_4994;
wire n_6652;
wire n_9377;
wire n_2537;
wire n_11932;
wire n_10971;
wire n_8830;
wire n_5347;
wire n_4483;
wire n_6970;
wire n_6921;
wire n_5168;
wire n_4661;
wire n_1308;
wire n_13027;
wire n_12867;
wire n_4988;
wire n_7674;
wire n_9826;
wire n_3171;
wire n_12607;
wire n_7568;
wire n_6354;
wire n_7272;
wire n_3608;
wire n_12075;
wire n_4540;
wire n_11942;
wire n_6344;
wire n_2097;
wire n_12305;
wire n_12123;
wire n_3459;
wire n_9772;
wire n_12170;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_3358;
wire n_6021;
wire n_7949;
wire n_7724;
wire n_3499;
wire n_9630;
wire n_6624;
wire n_6956;
wire n_4284;
wire n_12966;
wire n_6305;
wire n_9255;
wire n_1005;
wire n_1947;
wire n_10231;
wire n_8310;
wire n_6209;
wire n_12547;
wire n_9758;
wire n_3426;
wire n_11922;
wire n_4971;
wire n_8936;
wire n_5656;
wire n_7126;
wire n_1469;
wire n_5125;
wire n_5857;
wire n_12358;
wire n_7329;
wire n_8646;
wire n_7408;
wire n_9691;
wire n_12997;
wire n_10259;
wire n_2650;
wire n_7107;
wire n_5652;
wire n_6457;
wire n_8597;
wire n_10488;
wire n_987;
wire n_7690;
wire n_8969;
wire n_7123;
wire n_10752;
wire n_11577;
wire n_5499;
wire n_720;
wire n_8117;
wire n_10067;
wire n_153;
wire n_3229;
wire n_3348;
wire n_1707;
wire n_10399;
wire n_11223;
wire n_10213;
wire n_12498;
wire n_656;
wire n_11475;
wire n_8208;
wire n_6950;
wire n_10038;
wire n_9048;
wire n_5228;
wire n_797;
wire n_11010;
wire n_2933;
wire n_10274;
wire n_9590;
wire n_2717;
wire n_1723;
wire n_11588;
wire n_1878;
wire n_189;
wire n_738;
wire n_2012;
wire n_6694;
wire n_3497;
wire n_6880;
wire n_5066;
wire n_9168;
wire n_7418;
wire n_2842;
wire n_3580;
wire n_11221;
wire n_12387;
wire n_2335;
wire n_9497;
wire n_8536;
wire n_9435;
wire n_7229;
wire n_8350;
wire n_529;
wire n_2307;
wire n_3704;
wire n_11448;
wire n_684;
wire n_9219;
wire n_5507;
wire n_1809;
wire n_5569;
wire n_8028;
wire n_4280;
wire n_8328;
wire n_8914;
wire n_1181;
wire n_12576;
wire n_7258;
wire n_5190;
wire n_8391;
wire n_10579;
wire n_10832;
wire n_3173;
wire n_3677;
wire n_8336;
wire n_6856;
wire n_3996;
wire n_1049;
wire n_6466;
wire n_7864;
wire n_6727;
wire n_4097;
wire n_1666;
wire n_10584;
wire n_803;
wire n_4218;
wire n_5392;
wire n_1717;
wire n_1817;
wire n_12862;
wire n_2449;
wire n_11445;
wire n_13151;
wire n_3880;
wire n_3685;
wire n_8216;
wire n_11552;
wire n_2868;
wire n_10332;
wire n_7709;
wire n_11874;
wire n_2231;
wire n_3609;
wire n_9982;
wire n_10171;
wire n_1228;
wire n_5455;
wire n_417;
wire n_5442;
wire n_6386;
wire n_12803;
wire n_5948;
wire n_7804;
wire n_4459;
wire n_4545;
wire n_12656;
wire n_9852;
wire n_272;
wire n_6820;
wire n_2896;
wire n_11623;
wire n_8313;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_5511;
wire n_2898;
wire n_7656;
wire n_6208;
wire n_5295;
wire n_6739;
wire n_2368;
wire n_8041;
wire n_10676;
wire n_8202;
wire n_8263;
wire n_458;
wire n_4175;
wire n_10299;
wire n_10540;
wire n_5490;
wire n_11936;
wire n_6438;
wire n_12845;
wire n_10374;
wire n_11645;
wire n_3200;
wire n_4771;
wire n_10200;
wire n_7332;
wire n_12734;
wire n_3259;
wire n_2524;
wire n_10382;
wire n_3167;
wire n_2460;
wire n_5836;
wire n_7185;
wire n_6291;
wire n_11489;
wire n_3867;
wire n_10269;
wire n_3593;
wire n_4455;
wire n_8374;
wire n_12262;
wire n_1073;
wire n_9169;
wire n_252;
wire n_4514;
wire n_5834;
wire n_3191;
wire n_10229;
wire n_5584;
wire n_7512;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_4806;
wire n_7386;
wire n_9939;
wire n_7766;
wire n_11018;
wire n_8738;
wire n_10981;
wire n_9126;
wire n_6469;
wire n_6700;
wire n_12797;
wire n_2682;
wire n_3032;
wire n_6223;
wire n_11376;
wire n_6758;
wire n_9438;
wire n_11398;
wire n_5160;
wire n_7808;
wire n_6544;
wire n_8798;
wire n_9481;
wire n_9600;
wire n_2877;
wire n_9122;
wire n_11274;
wire n_8085;
wire n_5098;
wire n_1021;
wire n_8123;
wire n_10344;
wire n_7955;
wire n_811;
wire n_683;
wire n_1207;
wire n_5707;
wire n_12012;
wire n_5140;
wire n_4992;
wire n_12512;
wire n_5197;
wire n_7287;
wire n_9927;
wire n_5497;
wire n_10076;
wire n_11515;
wire n_8721;
wire n_880;
wire n_12820;
wire n_6464;
wire n_9912;
wire n_6356;
wire n_3505;
wire n_3577;
wire n_3540;
wire n_11554;
wire n_7637;
wire n_2432;
wire n_10148;
wire n_150;
wire n_1478;
wire n_10318;
wire n_4796;
wire n_3598;
wire n_4442;
wire n_2581;
wire n_1363;
wire n_3777;
wire n_4203;
wire n_3641;
wire n_7127;
wire n_767;
wire n_1837;
wire n_2218;
wire n_4533;
wire n_831;
wire n_9635;
wire n_5481;
wire n_12890;
wire n_3590;
wire n_8666;
wire n_2435;
wire n_5344;
wire n_954;
wire n_9264;
wire n_4419;
wire n_8326;
wire n_8670;
wire n_5308;
wire n_1410;
wire n_5184;
wire n_5794;
wire n_7638;
wire n_11972;
wire n_12284;
wire n_1382;
wire n_5408;
wire n_7801;
wire n_1736;
wire n_9155;
wire n_4053;
wire n_10234;
wire n_8460;
wire n_1483;
wire n_3848;
wire n_10416;
wire n_1372;
wire n_3327;
wire n_1719;
wire n_8836;
wire n_7959;
wire n_319;
wire n_7019;
wire n_8181;
wire n_2701;
wire n_2511;
wire n_11325;
wire n_8254;
wire n_4167;
wire n_8071;
wire n_1427;
wire n_2745;
wire n_7735;
wire n_8004;
wire n_1080;
wire n_6667;
wire n_7409;
wire n_5271;
wire n_10735;
wire n_10583;
wire n_10731;
wire n_9878;
wire n_562;
wire n_5964;
wire n_6004;
wire n_10806;
wire n_2323;
wire n_9825;
wire n_2784;
wire n_5494;
wire n_7444;
wire n_11628;
wire n_162;
wire n_5234;
wire n_4431;
wire n_7546;
wire n_2421;
wire n_1136;
wire n_6272;
wire n_4387;
wire n_2618;
wire n_6588;
wire n_3265;
wire n_11549;
wire n_2464;
wire n_1125;
wire n_4042;
wire n_3755;
wire n_5128;
wire n_12286;
wire n_9001;
wire n_2224;
wire n_10393;
wire n_11498;
wire n_13081;
wire n_2329;
wire n_1092;
wire n_10513;
wire n_12252;
wire n_441;
wire n_5467;
wire n_10439;
wire n_7296;
wire n_8013;
wire n_4299;
wire n_12627;
wire n_4890;
wire n_146;
wire n_1784;
wire n_7575;
wire n_3571;
wire n_9045;
wire n_7083;
wire n_193;
wire n_1775;
wire n_12281;
wire n_11237;
wire n_2410;
wire n_7720;
wire n_6222;
wire n_11643;
wire n_1093;
wire n_9373;
wire n_1783;
wire n_6268;
wire n_2929;
wire n_4176;
wire n_5827;
wire n_5199;
wire n_12347;
wire n_6456;
wire n_11103;
wire n_11809;
wire n_296;
wire n_11181;
wire n_9967;
wire n_7521;
wire n_651;
wire n_3407;
wire n_5992;
wire n_217;
wire n_12968;
wire n_5313;
wire n_10663;
wire n_1185;
wire n_3856;
wire n_4236;
wire n_9971;
wire n_7187;
wire n_3425;
wire n_215;
wire n_10894;
wire n_3894;
wire n_9524;
wire n_12277;
wire n_3127;
wire n_1831;
wire n_12698;
wire n_2621;
wire n_3623;
wire n_5312;
wire n_6467;
wire n_9243;
wire n_9182;
wire n_9282;
wire n_5079;
wire n_9365;
wire n_6540;
wire n_6625;
wire n_10909;
wire n_1453;
wire n_6336;
wire n_10083;
wire n_6796;
wire n_2502;
wire n_3646;
wire n_10347;
wire n_9224;
wire n_5513;
wire n_5614;
wire n_497;
wire n_12417;
wire n_11871;
wire n_6541;
wire n_12410;
wire n_4830;
wire n_4706;
wire n_1315;
wire n_5225;
wire n_4570;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_10208;
wire n_7722;
wire n_3188;
wire n_1459;
wire n_2462;
wire n_3243;
wire n_1135;
wire n_2889;
wire n_8487;
wire n_4034;
wire n_4056;
wire n_9240;
wire n_10804;
wire n_8293;
wire n_6486;
wire n_4622;
wire n_3960;
wire n_1470;
wire n_8141;
wire n_12294;
wire n_7603;
wire n_10667;
wire n_4887;
wire n_8438;
wire n_10548;
wire n_11020;
wire n_12957;
wire n_2732;
wire n_4693;
wire n_13141;
wire n_4206;
wire n_11616;
wire n_8791;
wire n_11920;
wire n_2249;
wire n_10793;
wire n_8288;
wire n_1091;
wire n_2000;
wire n_3862;
wire n_4267;
wire n_5835;
wire n_10481;
wire n_6732;
wire n_7979;
wire n_6876;
wire n_2270;
wire n_1425;
wire n_12786;
wire n_5049;
wire n_12711;
wire n_11675;
wire n_983;
wire n_12219;
wire n_10678;
wire n_6757;
wire n_9573;
wire n_5846;
wire n_906;
wire n_1390;
wire n_2289;
wire n_8657;
wire n_1733;
wire n_8006;
wire n_8296;
wire n_10440;
wire n_7636;
wire n_9799;
wire n_10391;
wire n_9695;
wire n_2955;
wire n_11083;
wire n_5592;
wire n_6954;
wire n_2158;
wire n_6938;
wire n_4609;
wire n_7866;
wire n_1855;
wire n_11306;
wire n_3051;
wire n_9784;
wire n_11198;
wire n_3367;
wire n_7205;
wire n_385;
wire n_1687;
wire n_8757;
wire n_1439;
wire n_2328;
wire n_7990;
wire n_7020;
wire n_2859;
wire n_10036;
wire n_2202;
wire n_13035;
wire n_13021;
wire n_1331;
wire n_736;
wire n_613;
wire n_5278;
wire n_11728;
wire n_12893;
wire n_8596;
wire n_3314;
wire n_3525;
wire n_2100;
wire n_5157;
wire n_11840;
wire n_3016;
wire n_2993;
wire n_4754;
wire n_4647;
wire n_9556;
wire n_1134;
wire n_3688;
wire n_11292;
wire n_8590;
wire n_8720;
wire n_10261;
wire n_13157;
wire n_4003;
wire n_5708;
wire n_554;
wire n_1995;
wire n_3751;
wire n_5223;
wire n_6298;
wire n_12205;
wire n_11989;
wire n_4894;
wire n_5474;
wire n_12289;
wire n_4113;
wire n_10813;
wire n_1889;
wire n_10757;
wire n_4760;
wire n_5649;
wire n_11326;
wire n_13046;
wire n_6421;
wire n_435;
wire n_1905;
wire n_11870;
wire n_9827;
wire n_7407;
wire n_3466;
wire n_10907;
wire n_762;
wire n_5704;
wire n_11431;
wire n_4983;
wire n_1778;
wire n_7148;
wire n_6328;
wire n_5956;
wire n_11283;
wire n_5287;
wire n_6236;
wire n_9417;
wire n_11834;
wire n_1079;
wire n_2139;
wire n_12020;
wire n_419;
wire n_5083;
wire n_7214;
wire n_4509;
wire n_6007;
wire n_3907;
wire n_1103;
wire n_2875;
wire n_6144;
wire n_11506;
wire n_10135;
wire n_13161;
wire n_3338;
wire n_144;
wire n_4217;
wire n_6197;
wire n_6658;
wire n_4906;
wire n_2219;
wire n_6835;
wire n_1203;
wire n_8834;
wire n_3636;
wire n_11624;
wire n_2327;
wire n_8826;
wire n_11352;
wire n_999;
wire n_5516;
wire n_1254;
wire n_2841;
wire n_6247;
wire n_7075;
wire n_4897;
wire n_10822;
wire n_11234;
wire n_10919;
wire n_7104;
wire n_9152;
wire n_7124;
wire n_12099;
wire n_12858;
wire n_3539;
wire n_3291;
wire n_7467;
wire n_4399;
wire n_2304;
wire n_8364;
wire n_7799;
wire n_2487;
wire n_5698;
wire n_11092;
wire n_3276;
wire n_2597;
wire n_9534;
wire n_3194;
wire n_5084;
wire n_5771;
wire n_7544;
wire n_13053;
wire n_9792;
wire n_7513;
wire n_10720;
wire n_9336;
wire n_10535;
wire n_3572;
wire n_11836;
wire n_349;
wire n_6602;
wire n_10924;
wire n_3886;
wire n_6708;
wire n_11186;
wire n_8854;
wire n_8917;
wire n_9647;
wire n_6645;
wire n_9742;
wire n_11236;
wire n_10727;
wire n_10885;
wire n_6484;
wire n_4710;
wire n_4420;
wire n_443;
wire n_892;
wire n_3637;
wire n_6242;
wire n_12527;
wire n_4574;
wire n_12379;
wire n_1468;
wire n_2855;
wire n_1859;
wire n_9312;
wire n_2156;
wire n_9019;
wire n_1718;
wire n_8985;
wire n_7692;
wire n_12067;
wire n_9214;
wire n_12932;
wire n_5174;
wire n_4234;
wire n_12477;
wire n_7469;
wire n_5538;
wire n_4101;
wire n_3548;
wire n_7776;
wire n_5017;
wire n_10418;
wire n_1768;
wire n_10895;
wire n_3974;
wire n_198;
wire n_1847;
wire n_3634;
wire n_10875;
wire n_11736;
wire n_11977;
wire n_7560;
wire n_9864;
wire n_8548;
wire n_10672;
wire n_7645;
wire n_11846;
wire n_1397;
wire n_3236;
wire n_11696;
wire n_12400;
wire n_901;
wire n_3141;
wire n_2755;
wire n_923;
wire n_5096;
wire n_11734;
wire n_1841;
wire n_4660;
wire n_9533;
wire n_9494;
wire n_12114;
wire n_5241;
wire n_11770;
wire n_10308;
wire n_11608;
wire n_1623;
wire n_11507;
wire n_9145;
wire n_1015;
wire n_7082;
wire n_12092;
wire n_3112;
wire n_12295;
wire n_10623;
wire n_9754;
wire n_4797;
wire n_3108;
wire n_6285;
wire n_9315;
wire n_11320;
wire n_4270;
wire n_11837;
wire n_5428;
wire n_4151;
wire n_7451;
wire n_4945;
wire n_8260;
wire n_3417;
wire n_9000;
wire n_5677;
wire n_9454;
wire n_4124;
wire n_6734;
wire n_7476;
wire n_10864;
wire n_10586;
wire n_5570;
wire n_11938;
wire n_6418;
wire n_8742;
wire n_12626;
wire n_785;
wire n_8307;
wire n_5153;
wire n_11967;
wire n_9383;
wire n_9253;
wire n_609;
wire n_10571;
wire n_4611;
wire n_8874;
wire n_5927;
wire n_7392;
wire n_11996;
wire n_9566;
wire n_11338;
wire n_7495;
wire n_5435;
wire n_2337;
wire n_12174;
wire n_9765;
wire n_1356;
wire n_3213;
wire n_9807;
wire n_4333;
wire n_3820;
wire n_5200;
wire n_8706;
wire n_9057;
wire n_6400;
wire n_2607;
wire n_7666;
wire n_7945;
wire n_8894;
wire n_2890;
wire n_1168;
wire n_5115;
wire n_6941;
wire n_12053;
wire n_1943;
wire n_5566;
wire n_11250;
wire n_7829;
wire n_12619;
wire n_3249;
wire n_1320;
wire n_7543;
wire n_8680;
wire n_11289;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_7877;
wire n_7963;
wire n_9672;
wire n_2499;
wire n_12582;
wire n_4152;
wire n_5487;
wire n_8855;
wire n_6398;
wire n_10394;
wire n_8885;
wire n_8329;
wire n_302;
wire n_5486;
wire n_9503;
wire n_12423;
wire n_137;
wire n_11391;
wire n_1596;
wire n_5092;
wire n_5244;
wire n_1734;
wire n_3172;
wire n_8270;
wire n_4832;
wire n_12714;
wire n_2902;
wire n_5889;
wire n_11738;
wire n_3217;
wire n_7284;
wire n_12153;
wire n_1983;
wire n_7264;
wire n_5391;
wire n_11522;
wire n_1938;
wire n_9763;
wire n_7737;
wire n_6537;
wire n_8614;
wire n_2472;
wire n_7328;
wire n_10702;
wire n_11070;
wire n_10958;
wire n_9479;
wire n_3394;
wire n_9162;
wire n_9568;
wire n_1715;
wire n_3536;
wire n_12405;
wire n_8816;
wire n_1443;
wire n_1272;
wire n_2894;
wire n_3957;
wire n_3710;
wire n_9119;
wire n_4195;
wire n_10319;
wire n_5849;
wire n_9654;
wire n_9181;
wire n_11648;
wire n_4554;
wire n_10322;
wire n_7135;
wire n_6578;
wire n_6224;
wire n_3040;
wire n_9859;
wire n_8802;
wire n_3279;
wire n_8555;
wire n_5240;
wire n_10695;
wire n_8636;
wire n_7024;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_6092;
wire n_10879;
wire n_5951;
wire n_6241;
wire n_6589;
wire n_1692;
wire n_1084;
wire n_6614;
wire n_8508;
wire n_5912;
wire n_8667;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_10639;
wire n_3501;
wire n_3475;
wire n_374;
wire n_1705;
wire n_8121;
wire n_3905;
wire n_8207;
wire n_9645;
wire n_9276;
wire n_8035;
wire n_12554;
wire n_8323;
wire n_11653;
wire n_12722;
wire n_6735;
wire n_7754;
wire n_4680;
wire n_3013;
wire n_10491;
wire n_921;
wire n_12037;
wire n_579;
wire n_2789;
wire n_5152;
wire n_5265;
wire n_12792;
wire n_2257;
wire n_11717;
wire n_9943;
wire n_4927;
wire n_5574;
wire n_12391;
wire n_9821;
wire n_11112;
wire n_4258;
wire n_1828;
wire n_2699;
wire n_7152;
wire n_11723;
wire n_2200;
wire n_9575;
wire n_650;
wire n_6165;
wire n_8320;
wire n_9796;
wire n_10409;
wire n_1940;
wire n_4548;
wire n_11822;
wire n_4862;
wire n_10521;
wire n_9610;
wire n_1405;
wire n_2376;
wire n_11830;
wire n_12438;
wire n_5469;
wire n_8766;
wire n_456;
wire n_12364;
wire n_3878;
wire n_12420;
wire n_12838;
wire n_9165;
wire n_6567;
wire n_2670;
wire n_313;
wire n_2700;
wire n_12323;
wire n_5910;
wire n_5895;
wire n_1041;
wire n_5804;
wire n_9508;
wire n_12539;
wire n_12776;
wire n_10527;
wire n_565;
wire n_3134;
wire n_5965;
wire n_9596;
wire n_1569;
wire n_3115;
wire n_1062;
wire n_7240;
wire n_7570;
wire n_896;
wire n_4553;
wire n_3278;
wire n_7033;
wire n_2084;
wire n_4875;
wire n_10476;
wire n_9966;
wire n_13156;
wire n_7817;
wire n_5682;
wire n_10710;
wire n_5387;
wire n_654;
wire n_5557;
wire n_411;
wire n_11394;
wire n_2458;
wire n_8850;
wire n_1222;
wire n_11906;
wire n_3050;
wire n_9928;
wire n_11820;
wire n_2673;
wire n_2456;
wire n_8002;
wire n_9741;
wire n_2527;
wire n_2635;
wire n_1637;
wire n_3307;
wire n_11486;
wire n_1407;
wire n_1795;
wire n_2871;
wire n_12677;
wire n_420;
wire n_4321;
wire n_10180;
wire n_4183;
wire n_8370;
wire n_7237;
wire n_164;
wire n_5681;
wire n_10650;
wire n_12120;
wire n_9090;
wire n_12021;
wire n_10157;
wire n_6877;
wire n_7423;
wire n_12873;
wire n_12008;
wire n_10402;
wire n_12515;
wire n_6949;
wire n_7566;
wire n_6119;
wire n_11940;
wire n_1271;
wire n_4145;
wire n_1545;
wire n_4821;
wire n_4901;
wire n_3121;
wire n_9217;
wire n_9261;
wire n_9166;
wire n_12901;
wire n_1640;
wire n_4040;
wire n_10518;
wire n_8301;
wire n_2406;
wire n_12895;
wire n_7617;
wire n_12223;
wire n_12045;
wire n_806;
wire n_9771;
wire n_584;
wire n_2141;
wire n_5316;
wire n_7718;
wire n_244;
wire n_6940;
wire n_9893;
wire n_12276;
wire n_548;
wire n_7396;
wire n_282;
wire n_10942;
wire n_12726;
wire n_12668;
wire n_5703;
wire n_7835;
wire n_11430;
wire n_833;
wire n_13010;
wire n_523;
wire n_6320;
wire n_8126;
wire n_345;
wire n_11239;
wire n_7998;
wire n_10362;
wire n_9239;
wire n_3930;
wire n_4943;
wire n_799;
wire n_10953;
wire n_12432;
wire n_3044;
wire n_4757;
wire n_7561;
wire n_6810;
wire n_7842;
wire n_2196;
wire n_2629;
wire n_12352;
wire n_2809;
wire n_787;
wire n_2172;
wire n_6202;
wire n_9969;
wire n_10099;
wire n_11437;
wire n_4682;
wire n_9961;
wire n_12898;
wire n_12879;
wire n_5564;
wire n_11869;
wire n_12559;
wire n_5620;
wire n_7163;
wire n_4530;
wire n_1528;
wire n_1146;
wire n_10343;
wire n_2021;
wire n_10836;
wire n_4942;
wire n_9899;
wire n_9258;
wire n_159;
wire n_1086;
wire n_13004;
wire n_10181;
wire n_10286;
wire n_5406;
wire n_2125;
wire n_8072;
wire n_10371;
wire n_2561;
wire n_8277;
wire n_7236;
wire n_652;
wire n_4604;
wire n_13117;
wire n_10257;
wire n_1906;
wire n_3305;
wire n_2992;
wire n_7130;
wire n_5724;
wire n_1241;
wire n_7201;
wire n_11219;
wire n_3157;
wire n_4841;
wire n_10047;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_2422;
wire n_1914;
wire n_1318;
wire n_5806;
wire n_10949;
wire n_3457;
wire n_4338;
wire n_10486;
wire n_11282;
wire n_11226;
wire n_306;
wire n_3762;
wire n_8724;
wire n_5738;
wire n_3005;
wire n_11413;
wire n_3151;
wire n_3411;
wire n_4840;
wire n_1029;
wire n_4519;
wire n_3779;
wire n_2388;
wire n_5355;
wire n_3984;
wire n_5320;
wire n_7491;
wire n_5353;
wire n_9995;
wire n_1706;
wire n_5710;
wire n_5186;
wire n_9076;
wire n_11232;
wire n_1498;
wire n_12351;
wire n_12693;
wire n_2417;
wire n_9105;
wire n_6792;
wire n_1210;
wire n_12080;
wire n_5093;
wire n_1556;
wire n_4052;
wire n_9316;
wire n_5979;
wire n_9636;
wire n_9668;
wire n_3558;
wire n_10372;
wire n_7559;
wire n_1984;
wire n_2236;
wire n_5438;
wire n_6044;
wire n_8867;
wire n_9491;
wire n_4326;
wire n_12702;
wire n_1269;
wire n_2083;
wire n_2834;
wire n_5517;
wire n_3207;
wire n_11276;
wire n_5605;
wire n_12439;
wire n_2441;
wire n_3401;
wire n_10744;
wire n_12648;
wire n_3242;
wire n_11008;
wire n_9870;
wire n_9833;
wire n_3613;
wire n_6125;
wire n_7314;
wire n_655;
wire n_9095;
wire n_4726;
wire n_7678;
wire n_1045;
wire n_5907;
wire n_11334;
wire n_786;
wire n_1559;
wire n_6045;
wire n_13075;
wire n_13129;
wire n_1872;
wire n_9914;
wire n_8132;
wire n_6731;
wire n_9178;
wire n_7526;
wire n_5040;
wire n_6063;
wire n_10736;
wire n_10917;
wire n_1325;
wire n_6504;
wire n_3761;
wire n_11575;
wire n_4315;
wire n_2923;
wire n_2888;
wire n_7004;
wire n_7821;
wire n_1727;
wire n_12407;
wire n_8308;
wire n_6154;
wire n_11284;
wire n_6943;
wire n_4301;
wire n_10597;
wire n_11827;
wire n_151;
wire n_13049;
wire n_3744;
wire n_8165;
wire n_12038;
wire n_4788;
wire n_8400;
wire n_10458;
wire n_2041;
wire n_8210;
wire n_11656;
wire n_12644;
wire n_1360;
wire n_5977;
wire n_10446;
wire n_13134;
wire n_11826;
wire n_7879;
wire n_10271;
wire n_3814;
wire n_3781;
wire n_1908;
wire n_10888;
wire n_2484;
wire n_10116;
wire n_2126;
wire n_7696;
wire n_11570;
wire n_6003;
wire n_12952;
wire n_6684;
wire n_3843;
wire n_1098;
wire n_5746;
wire n_6600;
wire n_11764;
wire n_13063;
wire n_2045;
wire n_817;
wire n_5451;
wire n_9323;
wire n_3687;
wire n_2216;
wire n_5402;
wire n_6673;
wire n_10696;
wire n_7355;
wire n_6961;
wire n_3543;
wire n_9331;
wire n_3621;
wire n_6031;
wire n_9922;
wire n_10170;
wire n_12024;
wire n_8331;
wire n_11909;
wire n_13084;
wire n_8217;
wire n_10603;
wire n_12004;
wire n_2903;
wire n_6962;
wire n_3216;
wire n_332;
wire n_12830;
wire n_12637;
wire n_3808;
wire n_8858;
wire n_7887;
wire n_7246;
wire n_398;
wire n_4365;
wire n_6060;
wire n_1882;
wire n_7929;
wire n_10255;
wire n_10572;
wire n_3726;
wire n_12009;
wire n_1007;
wire n_1929;
wire n_2369;
wire n_1592;
wire n_2719;
wire n_7270;
wire n_591;
wire n_11490;
wire n_3758;
wire n_8689;
wire n_10648;
wire n_5417;
wire n_6967;
wire n_2587;
wire n_10113;
wire n_7550;
wire n_3199;
wire n_12414;
wire n_680;
wire n_9760;
wire n_10690;
wire n_3339;
wire n_6853;
wire n_10188;
wire n_6742;
wire n_4923;
wire n_2400;
wire n_5864;
wire n_10686;
wire n_9841;
wire n_6691;
wire n_8743;
wire n_7087;
wire n_12681;
wire n_8753;
wire n_1953;
wire n_6191;
wire n_4741;
wire n_10689;
wire n_6172;
wire n_3343;
wire n_12634;
wire n_10974;
wire n_13022;
wire n_11067;
wire n_2752;
wire n_8627;
wire n_9513;
wire n_9863;
wire n_12680;
wire n_11613;
wire n_4885;
wire n_10233;
wire n_12034;
wire n_751;
wire n_10500;
wire n_10555;
wire n_5432;
wire n_1399;
wire n_10314;
wire n_4550;
wire n_6988;
wire n_4652;
wire n_11929;
wire n_10810;
wire n_11075;
wire n_7851;
wire n_6894;
wire n_12176;
wire n_9791;
wire n_10311;
wire n_9179;
wire n_2358;
wire n_5453;
wire n_3658;
wire n_9140;
wire n_8752;
wire n_6834;
wire n_4900;
wire n_2163;
wire n_2186;
wire n_2815;
wire n_3034;
wire n_11177;
wire n_4408;
wire n_4577;
wire n_4748;
wire n_643;
wire n_5842;
wire n_6817;
wire n_10937;
wire n_13126;
wire n_6927;
wire n_12134;
wire n_400;
wire n_12449;
wire n_337;
wire n_5814;
wire n_2814;
wire n_7798;
wire n_5253;
wire n_5209;
wire n_10857;
wire n_11310;
wire n_12094;
wire n_6215;
wire n_789;
wire n_3231;
wire n_11165;
wire n_4212;
wire n_9736;
wire n_2979;
wire n_5699;
wire n_181;
wire n_5531;
wire n_5765;
wire n_12823;
wire n_2953;
wire n_12517;
wire n_6517;
wire n_327;
wire n_6284;
wire n_4295;
wire n_5943;
wire n_10167;
wire n_7862;
wire n_12193;
wire n_9225;
wire n_12524;
wire n_2946;
wire n_11923;
wire n_12071;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_10630;
wire n_8105;
wire n_6088;
wire n_9031;
wire n_5777;
wire n_4225;
wire n_6883;
wire n_10061;
wire n_8808;
wire n_12963;
wire n_10428;
wire n_13087;
wire n_300;
wire n_11865;
wire n_12366;
wire n_8528;
wire n_747;
wire n_8204;
wire n_13024;
wire n_11733;
wire n_11068;
wire n_11035;
wire n_2565;
wire n_5495;
wire n_10694;
wire n_1389;
wire n_12339;
wire n_10602;
wire n_535;
wire n_7100;
wire n_12729;
wire n_3583;
wire n_12198;
wire n_3860;
wire n_11041;
wire n_9420;
wire n_3851;
wire n_5655;
wire n_6393;
wire n_9708;
wire n_5064;
wire n_7825;
wire n_10079;
wire n_12242;
wire n_7119;
wire n_5610;
wire n_8154;
wire n_7212;
wire n_6966;
wire n_8889;
wire n_3015;
wire n_2175;
wire n_601;
wire n_2182;
wire n_9790;
wire n_10502;
wire n_11973;
wire n_11131;
wire n_4009;
wire n_1848;
wire n_5002;
wire n_5759;
wire n_10778;
wire n_6722;
wire n_1506;
wire n_3473;
wire n_1652;
wire n_6035;
wire n_957;
wire n_1994;
wire n_7874;
wire n_8490;
wire n_7622;
wire n_10329;
wire n_9014;
wire n_9979;
wire n_8509;
wire n_8767;
wire n_11123;
wire n_8512;
wire n_9505;
wire n_8634;
wire n_9531;
wire n_2566;
wire n_6364;
wire n_387;
wire n_744;
wire n_971;
wire n_8635;
wire n_2702;
wire n_3241;
wire n_7420;
wire n_7102;
wire n_2906;
wire n_4342;
wire n_12605;
wire n_10855;
wire n_7995;
wire n_6114;
wire n_4568;
wire n_1205;
wire n_11003;
wire n_6061;
wire n_10662;
wire n_5559;
wire n_1258;
wire n_2438;
wire n_6253;
wire n_7831;
wire n_2914;
wire n_12828;
wire n_12723;
wire n_10258;
wire n_5786;
wire n_8532;
wire n_12661;
wire n_10227;
wire n_10588;
wire n_8624;
wire n_8991;
wire n_11022;
wire n_10574;
wire n_8065;
wire n_10247;
wire n_3100;
wire n_2180;
wire n_11140;
wire n_2858;
wire n_5377;
wire n_3573;
wire n_6201;
wire n_1016;
wire n_8796;
wire n_12218;
wire n_4106;
wire n_5737;
wire n_1501;
wire n_3604;
wire n_12343;
wire n_10733;
wire n_4373;
wire n_8518;
wire n_10472;
wire n_8919;
wire n_12597;
wire n_12316;
wire n_197;
wire n_4711;
wire n_11478;
wire n_12834;
wire n_3068;
wire n_10066;
wire n_13017;
wire n_12236;
wire n_12902;
wire n_2685;
wire n_6419;
wire n_1083;
wire n_7784;
wire n_9272;
wire n_8372;
wire n_5768;
wire n_3553;
wire n_10088;
wire n_13038;
wire n_2465;
wire n_2275;
wire n_7225;
wire n_8077;
wire n_2568;
wire n_12892;
wire n_2022;
wire n_3811;
wire n_11294;
wire n_910;
wire n_3494;
wire n_1721;
wire n_9812;
wire n_6900;
wire n_6244;
wire n_1737;
wire n_9337;
wire n_3486;
wire n_4086;
wire n_752;
wire n_908;
wire n_6755;
wire n_9432;
wire n_6565;
wire n_10289;
wire n_9949;
wire n_7361;
wire n_1028;
wire n_6942;
wire n_7705;
wire n_11819;
wire n_2106;
wire n_2265;
wire n_7228;
wire n_5350;
wire n_13037;
wire n_5470;
wire n_2032;
wire n_4812;
wire n_7932;
wire n_4409;
wire n_9576;
wire n_11573;
wire n_10145;
wire n_7509;
wire n_5872;
wire n_6862;
wire n_7058;
wire n_11005;
wire n_5858;
wire n_4629;
wire n_6255;
wire n_4638;
wire n_708;
wire n_1973;
wire n_6840;
wire n_13005;
wire n_3181;
wire n_6338;
wire n_8262;
wire n_8423;
wire n_5700;
wire n_1500;
wire n_6037;
wire n_7981;
wire n_9577;
wire n_9874;
wire n_3699;
wire n_12588;
wire n_854;
wire n_4913;
wire n_12589;
wire n_2312;
wire n_5874;
wire n_6266;
wire n_6488;
wire n_904;
wire n_8337;
wire n_709;
wire n_1266;
wire n_2242;
wire n_9231;
wire n_11844;
wire n_7164;
wire n_3328;
wire n_6635;
wire n_7973;
wire n_6815;
wire n_185;
wire n_11364;
wire n_3868;
wire n_9569;
wire n_1276;
wire n_12790;
wire n_4266;
wire n_8632;
wire n_2466;
wire n_2530;
wire n_7018;
wire n_5873;
wire n_12247;
wire n_7975;
wire n_12699;
wire n_9719;
wire n_10009;
wire n_8358;
wire n_1085;
wire n_9552;
wire n_12927;
wire n_11100;
wire n_2042;
wire n_9279;
wire n_11902;
wire n_771;
wire n_6317;
wire n_475;
wire n_924;
wire n_8199;
wire n_298;
wire n_1582;
wire n_492;
wire n_5588;
wire n_11993;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_1149;
wire n_3170;
wire n_10443;
wire n_8656;
wire n_7167;
wire n_265;
wire n_10756;
wire n_12813;
wire n_6480;
wire n_3645;
wire n_10918;
wire n_13122;
wire n_5075;
wire n_11797;
wire n_3682;
wire n_3304;
wire n_2592;
wire n_4968;
wire n_3771;
wire n_12765;
wire n_7865;
wire n_2666;
wire n_1585;
wire n_12663;
wire n_10384;
wire n_1799;
wire n_9289;
wire n_2564;
wire n_5085;
wire n_11315;
wire n_5736;
wire n_4259;
wire n_2433;
wire n_829;
wire n_6561;
wire n_7978;
wire n_7820;
wire n_2035;
wire n_12706;
wire n_11127;
wire n_10293;
wire n_8881;
wire n_7844;
wire n_7134;
wire n_9633;
wire n_11153;
wire n_12312;
wire n_3422;
wire n_10074;
wire n_4572;
wire n_859;
wire n_3086;
wire n_2033;
wire n_406;
wire n_4104;
wire n_4845;
wire n_9547;
wire n_13097;
wire n_6875;
wire n_10934;
wire n_1770;
wire n_10197;
wire n_878;
wire n_8346;
wire n_5120;
wire n_3285;
wire n_4208;
wire n_8761;
wire n_13112;
wire n_9085;
wire n_9632;
wire n_10042;
wire n_8226;
wire n_11949;
wire n_8402;
wire n_10478;
wire n_7079;
wire n_9690;
wire n_9084;
wire n_981;
wire n_5928;
wire n_12256;
wire n_4089;
wire n_5478;
wire n_6016;
wire n_1144;
wire n_2071;
wire n_11746;
wire n_11812;
wire n_3219;
wire n_9371;
wire n_3702;
wire n_9711;
wire n_8754;
wire n_9431;
wire n_9847;
wire n_2233;
wire n_4779;
wire n_7267;
wire n_481;
wire n_10367;
wire n_3233;
wire n_4599;
wire n_12315;
wire n_997;
wire n_11505;
wire n_4437;
wire n_5222;
wire n_9889;
wire n_10867;
wire n_7850;
wire n_7316;
wire n_12375;
wire n_12556;
wire n_3310;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_12998;
wire n_7812;
wire n_1198;
wire n_7103;
wire n_13143;
wire n_9080;
wire n_4061;
wire n_8133;
wire n_10168;
wire n_7460;
wire n_6176;
wire n_2174;
wire n_436;
wire n_9519;
wire n_11363;
wire n_3881;
wire n_6367;
wire n_12156;
wire n_13128;
wire n_4508;
wire n_4727;
wire n_4594;
wire n_11530;
wire n_12671;
wire n_2426;
wire n_10621;
wire n_2478;
wire n_7056;
wire n_9731;
wire n_8193;
wire n_6572;
wire n_8714;
wire n_12445;
wire n_1133;
wire n_4429;
wire n_9604;
wire n_7962;
wire n_12856;
wire n_4642;
wire n_4051;
wire n_1051;
wire n_10085;
wire n_7813;
wire n_7755;
wire n_7514;
wire n_7649;
wire n_11151;
wire n_8182;
wire n_4865;
wire n_12525;
wire n_8387;
wire n_6080;
wire n_1039;
wire n_6078;
wire n_10613;
wire n_10716;
wire n_12076;
wire n_2043;
wire n_1480;
wire n_6056;
wire n_6717;
wire n_5832;
wire n_10664;
wire n_7473;
wire n_7200;
wire n_11359;
wire n_3206;
wire n_1305;
wire n_2578;
wire n_2363;
wire n_7688;
wire n_4562;
wire n_553;
wire n_3383;
wire n_8707;
wire n_12357;
wire n_4903;
wire n_3709;
wire n_10561;
wire n_11434;
wire n_3738;
wire n_9208;
wire n_11791;
wire n_7611;
wire n_6873;
wire n_4186;
wire n_8494;
wire n_5812;
wire n_2540;
wire n_973;
wire n_5743;
wire n_12468;
wire n_9429;
wire n_8544;
wire n_11848;
wire n_3610;
wire n_11152;
wire n_4998;
wire n_10749;
wire n_3330;
wire n_11632;
wire n_7795;
wire n_12180;
wire n_2065;
wire n_2879;
wire n_8788;
wire n_967;
wire n_4522;
wire n_10122;
wire n_10935;
wire n_7038;
wire n_10992;
wire n_2001;
wire n_7723;
wire n_4341;
wire n_11621;
wire n_679;
wire n_1629;
wire n_10160;
wire n_10560;
wire n_9327;
wire n_7404;
wire n_12857;
wire n_5368;
wire n_4263;
wire n_225;
wire n_1260;
wire n_1819;
wire n_309;
wire n_8177;
wire n_3555;
wire n_9854;
wire n_7059;
wire n_11667;
wire n_12025;
wire n_7450;
wire n_8962;
wire n_915;
wire n_9538;
wire n_5971;
wire n_6327;
wire n_7362;
wire n_812;
wire n_12208;
wire n_6145;
wire n_1131;
wire n_11964;
wire n_3155;
wire n_6539;
wire n_6926;
wire n_1006;
wire n_3110;
wire n_7271;
wire n_1632;
wire n_7826;
wire n_9713;
wire n_11298;
wire n_5933;
wire n_257;
wire n_1888;
wire n_8993;
wire n_6204;
wire n_1311;
wire n_7076;
wire n_4780;
wire n_10300;
wire n_670;
wire n_9588;
wire n_11403;
wire n_2697;
wire n_11741;
wire n_12383;
wire n_11912;
wire n_3908;
wire n_4973;
wire n_6842;
wire n_3467;
wire n_12773;
wire n_6866;
wire n_1887;
wire n_9044;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_4803;
wire n_2512;
wire n_3950;
wire n_9423;
wire n_12381;
wire n_9387;
wire n_6030;
wire n_1242;
wire n_2086;
wire n_2927;
wire n_4750;
wire n_12962;
wire n_6451;
wire n_9813;
wire n_3039;
wire n_9127;
wire n_1226;
wire n_6514;
wire n_3740;
wire n_9794;
wire n_5996;
wire n_11666;
wire n_12459;
wire n_2166;
wire n_2899;
wire n_3186;
wire n_640;
wire n_1322;
wire n_7105;
wire n_10140;
wire n_12612;
wire n_9244;
wire n_9869;
wire n_11142;
wire n_1958;
wire n_315;
wire n_7049;
wire n_5903;
wire n_5986;
wire n_1197;
wire n_3065;
wire n_2632;
wire n_6710;
wire n_4984;
wire n_8278;
wire n_12885;
wire n_11644;
wire n_2579;
wire n_6345;
wire n_2105;
wire n_9715;
wire n_1423;
wire n_8618;
wire n_3387;
wire n_12108;
wire n_9094;
wire n_13108;
wire n_364;
wire n_5782;
wire n_7535;
wire n_3420;
wire n_5041;
wire n_1915;
wire n_4275;
wire n_10862;
wire n_11531;
wire n_4283;
wire n_4959;
wire n_900;
wire n_8248;
wire n_9056;
wire n_11357;
wire n_8911;
wire n_4426;
wire n_9407;
wire n_2912;
wire n_11476;
wire n_2659;
wire n_4425;
wire n_3409;
wire n_9985;
wire n_4449;
wire n_2116;
wire n_12089;
wire n_12496;
wire n_2320;
wire n_11824;
wire n_12814;
wire n_7057;
wire n_1013;
wire n_1259;
wire n_11959;
wire n_11367;
wire n_2183;
wire n_3002;
wire n_6957;
wire n_9361;
wire n_649;
wire n_1612;
wire n_11921;
wire n_4809;
wire n_8495;
wire n_12676;
wire n_8783;
wire n_12987;
wire n_11566;
wire n_1199;
wire n_3392;
wire n_8529;
wire n_8733;
wire n_12603;
wire n_8990;
wire n_6050;
wire n_625;
wire n_7976;
wire n_6444;
wire n_10254;
wire n_226;
wire n_7944;
wire n_13080;
wire n_11208;
wire n_7262;
wire n_212;
wire n_3773;
wire n_8647;
wire n_11374;
wire n_12967;
wire n_12452;
wire n_2003;
wire n_8574;
wire n_1038;
wire n_1581;
wire n_7016;
wire n_10782;
wire n_12292;
wire n_12232;
wire n_3301;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_11859;
wire n_12818;
wire n_10386;
wire n_12128;
wire n_6379;
wire n_798;
wire n_2324;
wire n_11420;
wire n_12754;
wire n_12500;
wire n_5563;
wire n_245;
wire n_1348;
wire n_11026;
wire n_8044;
wire n_2977;
wire n_1739;
wire n_5840;
wire n_6719;
wire n_7178;
wire n_9439;
wire n_1380;
wire n_9553;
wire n_11633;
wire n_11467;
wire n_2847;
wire n_7506;
wire n_2557;
wire n_12672;
wire n_8551;
wire n_12063;
wire n_11630;
wire n_8330;
wire n_12760;
wire n_1009;
wire n_2405;
wire n_4050;
wire n_1160;
wire n_883;
wire n_2647;
wire n_6232;
wire n_9132;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_5717;
wire n_6017;
wire n_9696;
wire n_10861;
wire n_2521;
wire n_9120;
wire n_8879;
wire n_1099;
wire n_11203;
wire n_471;
wire n_11159;
wire n_424;
wire n_8052;
wire n_12168;
wire n_4578;
wire n_2211;
wire n_6362;
wire n_4777;
wire n_11956;
wire n_11975;
wire n_12121;
wire n_5720;
wire n_9332;
wire n_369;
wire n_8903;
wire n_11030;
wire n_2672;
wire n_4702;
wire n_12590;
wire n_2299;
wire n_4179;
wire n_4895;
wire n_5871;
wire n_12924;
wire n_7142;
wire n_141;
wire n_1285;
wire n_12577;
wire n_10182;
wire n_12732;
wire n_1985;
wire n_6326;
wire n_12649;
wire n_5898;
wire n_7125;
wire n_6858;
wire n_9252;
wire n_9464;
wire n_1172;
wire n_6649;
wire n_6283;
wire n_4026;
wire n_10073;
wire n_4531;
wire n_3282;
wire n_11655;
wire n_1590;
wire n_3626;
wire n_1532;
wire n_2313;
wire n_5072;
wire n_11017;
wire n_7241;
wire n_7247;
wire n_12843;
wire n_12069;
wire n_10419;
wire n_7172;
wire n_3106;
wire n_1140;
wire n_1670;
wire n_10333;
wire n_2344;
wire n_12430;
wire n_10317;
wire n_2365;
wire n_4666;
wire n_7893;
wire n_6213;
wire n_3031;
wire n_4029;
wire n_375;
wire n_7235;
wire n_8540;
wire n_2447;
wire n_11248;
wire n_12613;
wire n_6239;
wire n_12270;
wire n_9915;
wire n_4617;
wire n_2340;
wire n_9325;
wire n_9196;
wire n_4010;
wire n_5896;
wire n_1649;
wire n_4555;
wire n_5882;
wire n_5940;
wire n_6089;
wire n_5650;
wire n_7588;
wire n_9384;
wire n_4969;
wire n_6057;
wire n_6216;
wire n_10017;
wire n_7340;
wire n_12557;
wire n_6974;
wire n_11141;
wire n_5105;
wire n_12695;
wire n_10893;
wire n_1572;
wire n_4308;
wire n_11093;
wire n_5021;
wire n_9251;
wire n_3463;
wire n_11576;
wire n_8939;
wire n_428;
wire n_9973;
wire n_5263;
wire n_11117;
wire n_2510;
wire n_1954;
wire n_6713;
wire n_12139;
wire n_8064;
wire n_9030;
wire n_7657;
wire n_822;
wire n_8468;
wire n_2791;
wire n_4325;
wire n_3251;
wire n_4602;
wire n_5044;
wire n_9665;
wire n_10201;
wire n_5134;
wire n_7096;
wire n_2212;
wire n_3063;
wire n_1163;
wire n_2729;
wire n_12210;
wire n_2582;
wire n_1798;
wire n_1550;
wire n_8778;
wire n_11197;
wire n_491;
wire n_3998;
wire n_7442;
wire n_1591;
wire n_3632;
wire n_10093;
wire n_3122;
wire n_5567;
wire n_8343;
wire n_1344;
wire n_6174;
wire n_12006;
wire n_2730;
wire n_2495;
wire n_7999;
wire n_10128;
wire n_10675;
wire n_6087;
wire n_371;
wire n_7593;
wire n_12246;
wire n_5249;
wire n_2090;
wire n_2603;
wire n_8068;
wire n_9955;
wire n_538;
wire n_3829;
wire n_10539;
wire n_4164;
wire n_2173;
wire n_5625;
wire n_9007;
wire n_10143;
wire n_7764;
wire n_11777;
wire n_1471;
wire n_4919;
wire n_3737;
wire n_10107;
wire n_5969;
wire n_3655;
wire n_10196;
wire n_10121;
wire n_8198;
wire n_493;
wire n_3825;
wire n_3225;
wire n_2880;
wire n_13085;
wire n_2108;
wire n_7780;
wire n_6828;
wire n_5158;
wire n_7255;
wire n_8693;
wire n_12189;
wire n_1211;
wire n_11469;
wire n_6454;
wire n_5022;
wire n_12625;
wire n_9270;
wire n_8452;
wire n_7041;
wire n_7307;
wire n_11518;
wire n_12177;
wire n_10742;
wire n_5670;
wire n_10829;
wire n_8557;
wire n_1280;
wire n_6918;
wire n_6041;
wire n_9099;
wire n_12389;
wire n_9309;
wire n_3296;
wire n_7350;
wire n_10620;
wire n_10303;
wire n_10814;
wire n_5276;
wire n_9627;
wire n_11252;
wire n_8012;
wire n_1445;
wire n_7672;
wire n_11494;
wire n_2551;
wire n_6664;
wire n_1526;
wire n_5047;
wire n_196;
wire n_7318;
wire n_2985;
wire n_1978;
wire n_6472;
wire n_10218;
wire n_574;
wire n_8114;
wire n_13131;
wire n_3792;
wire n_4202;
wire n_12995;
wire n_1446;
wire n_3938;
wire n_4791;
wire n_11154;
wire n_3507;
wire n_11700;
wire n_5879;
wire n_8062;
wire n_4403;
wire n_11883;
wire n_5238;
wire n_11256;
wire n_11832;
wire n_6166;
wire n_5855;
wire n_3269;
wire n_12370;
wire n_3531;
wire n_9136;
wire n_6375;
wire n_12860;
wire n_473;
wire n_10975;
wire n_11901;
wire n_6352;
wire n_12974;
wire n_1054;
wire n_9460;
wire n_559;
wire n_8542;
wire n_12136;
wire n_10859;
wire n_13078;
wire n_7063;
wire n_1956;
wire n_11652;
wire n_7047;
wire n_4139;
wire n_6632;
wire n_4549;
wire n_11056;
wire n_8576;
wire n_6238;
wire n_1986;
wire n_10542;
wire n_8038;
wire n_2397;
wire n_3931;
wire n_4349;
wire n_10681;
wire n_6081;
wire n_9732;
wire n_10459;
wire n_11572;
wire n_5141;
wire n_2113;
wire n_1918;
wire n_11894;
wire n_3603;
wire n_10222;
wire n_6724;
wire n_13113;
wire n_10524;
wire n_5429;
wire n_6545;
wire n_813;
wire n_11583;
wire n_8716;
wire n_11336;
wire n_6705;
wire n_3822;
wire n_9766;
wire n_12758;
wire n_8629;
wire n_4163;
wire n_818;
wire n_9517;
wire n_10463;
wire n_5535;
wire n_645;
wire n_7074;
wire n_3910;
wire n_3812;
wire n_9204;
wire n_8734;
wire n_9476;
wire n_9689;
wire n_11849;
wire n_12142;
wire n_2633;
wire n_10659;
wire n_6591;
wire n_2207;
wire n_7585;
wire n_12564;
wire n_4948;
wire n_5268;
wire n_9780;
wire n_6946;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_6002;
wire n_2198;
wire n_3319;
wire n_541;
wire n_10403;
wire n_12983;
wire n_2073;
wire n_2273;
wire n_7037;
wire n_6289;
wire n_3748;
wire n_3272;
wire n_11784;
wire n_6424;
wire n_4941;
wire n_5506;
wire n_5298;
wire n_11399;
wire n_9025;
wire n_8524;
wire n_3396;
wire n_11210;
wire n_7599;
wire n_7928;
wire n_8768;
wire n_4393;
wire n_10884;
wire n_12886;
wire n_1162;
wire n_6532;
wire n_821;
wire n_4372;
wire n_1068;
wire n_7293;
wire n_13000;
wire n_982;
wire n_12035;
wire n_13006;
wire n_5640;
wire n_11191;
wire n_12791;
wire n_7600;
wire n_10547;
wire n_408;
wire n_932;
wire n_2831;
wire n_4318;
wire n_6778;
wire n_4158;
wire n_3317;
wire n_3978;
wire n_6721;
wire n_5560;
wire n_6644;
wire n_2123;
wire n_1697;
wire n_6512;
wire n_979;
wire n_4074;
wire n_3716;
wire n_4795;
wire n_5544;
wire n_12810;
wire n_6108;
wire n_8258;
wire n_10370;
wire n_4918;
wire n_3824;
wire n_9597;
wire n_5067;
wire n_11322;
wire n_5744;
wire n_4013;
wire n_11892;
wire n_12122;
wire n_6703;
wire n_5384;
wire n_4544;
wire n_3248;
wire n_354;
wire n_5841;
wire n_12241;
wire n_12396;
wire n_7614;
wire n_9343;
wire n_2941;
wire n_1278;
wire n_547;
wire n_7839;
wire n_5108;
wire n_8299;
wire n_12473;
wire n_7347;
wire n_4032;
wire n_1064;
wire n_6086;
wire n_9837;
wire n_1396;
wire n_11421;
wire n_11057;
wire n_634;
wire n_2355;
wire n_4147;
wire n_10896;
wire n_10969;
wire n_136;
wire n_4477;
wire n_11966;
wire n_12748;
wire n_3168;
wire n_7383;
wire n_2751;
wire n_6805;
wire n_4337;
wire n_8863;
wire n_4130;
wire n_10562;
wire n_5941;
wire n_2009;
wire n_7759;
wire n_12184;
wire n_10210;
wire n_1793;
wire n_3601;
wire n_5611;
wire n_6340;
wire n_10054;
wire n_3092;
wire n_1289;
wire n_6219;
wire n_3055;
wire n_6706;
wire n_7479;
wire n_3966;
wire n_10355;
wire n_11853;
wire n_12571;
wire n_9692;
wire n_2866;
wire n_7395;
wire n_10598;
wire n_13034;
wire n_8947;
wire n_4742;
wire n_1014;
wire n_3734;
wire n_9609;
wire n_10717;
wire n_11118;
wire n_10029;
wire n_1703;
wire n_7078;
wire n_2580;
wire n_8188;
wire n_6761;
wire n_882;
wire n_8972;
wire n_10007;
wire n_3649;
wire n_11751;
wire n_2821;
wire n_11423;
wire n_1875;
wire n_11725;
wire n_1865;
wire n_5701;
wire n_3746;
wire n_6067;
wire n_10801;
wire n_9206;
wire n_12674;
wire n_8510;
wire n_11410;
wire n_3384;
wire n_12230;
wire n_9567;
wire n_1950;
wire n_6811;
wire n_9061;
wire n_1563;
wire n_11495;
wire n_3419;
wire n_9942;
wire n_11712;
wire n_9703;
wire n_1297;
wire n_1662;
wire n_4478;
wire n_7372;
wire n_1359;
wire n_2818;
wire n_5367;
wire n_3794;
wire n_12220;
wire n_674;
wire n_3921;
wire n_6868;
wire n_8664;
wire n_922;
wire n_10704;
wire n_1335;
wire n_11520;
wire n_11622;
wire n_1927;
wire n_4838;
wire n_5970;
wire n_12169;
wire n_12283;
wire n_12336;
wire n_7174;
wire n_9421;
wire n_5202;
wire n_10740;
wire n_10457;
wire n_12543;
wire n_702;
wire n_4965;
wire n_347;
wire n_8021;
wire n_3346;
wire n_9705;
wire n_7803;
wire n_1896;
wire n_11012;
wire n_2965;
wire n_6111;
wire n_3058;
wire n_12595;
wire n_9624;
wire n_3861;
wire n_9701;
wire n_675;
wire n_11502;
wire n_11429;
wire n_1540;
wire n_1977;
wire n_10389;
wire n_11631;
wire n_3891;
wire n_2193;
wire n_6659;
wire n_4523;
wire n_1655;
wire n_9709;
wire n_242;
wire n_6011;
wire n_9416;
wire n_1886;
wire n_9295;
wire n_4371;
wire n_6225;
wire n_11842;
wire n_12463;
wire n_10990;
wire n_2994;
wire n_11640;
wire n_5502;
wire n_12263;
wire n_3428;
wire n_3153;
wire n_4552;
wire n_6218;
wire n_3689;
wire n_8982;
wire n_877;
wire n_9929;
wire n_12920;
wire n_10264;
wire n_5850;
wire n_4673;
wire n_2519;
wire n_9953;
wire n_7086;
wire n_728;
wire n_3415;
wire n_1063;
wire n_6648;
wire n_4607;
wire n_12528;
wire n_10955;
wire n_11389;
wire n_7927;
wire n_6182;
wire n_9013;
wire n_7226;
wire n_12717;
wire n_4041;
wire n_2947;
wire n_6520;
wire n_12660;
wire n_3918;
wire n_9634;
wire n_9532;
wire n_11011;
wire n_5876;
wire n_9998;
wire n_11795;
wire n_5521;
wire n_1965;
wire n_4837;
wire n_2476;
wire n_9850;
wire n_6601;
wire n_10916;
wire n_598;
wire n_12141;
wire n_8584;
wire n_11547;
wire n_11557;
wire n_9346;
wire n_7920;
wire n_437;
wire n_12774;
wire n_7810;
wire n_8501;
wire n_4169;
wire n_11904;
wire n_8480;
wire n_697;
wire n_10301;
wire n_3271;
wire n_295;
wire n_5088;
wire n_4248;
wire n_8034;
wire n_388;
wire n_13018;
wire n_484;
wire n_7025;
wire n_9364;
wire n_8228;
wire n_2976;
wire n_2152;
wire n_2652;
wire n_8076;
wire n_6826;
wire n_1825;
wire n_1757;
wire n_170;
wire n_1792;
wire n_5856;
wire n_11395;
wire n_8484;
wire n_9472;
wire n_9836;
wire n_1412;
wire n_2497;
wire n_10929;
wire n_9107;
wire n_3809;
wire n_11279;
wire n_11724;
wire n_13044;
wire n_11789;
wire n_3139;
wire n_11525;
wire n_8100;
wire n_4070;
wire n_11999;
wire n_13086;
wire n_10837;
wire n_3545;
wire n_3885;
wire n_1369;
wire n_881;
wire n_10554;
wire n_8014;
wire n_3993;
wire n_8994;
wire n_8091;
wire n_8413;
wire n_4685;
wire n_12746;
wire n_4031;
wire n_5837;
wire n_148;
wire n_4675;
wire n_10149;
wire n_10970;
wire n_7768;
wire n_2663;
wire n_8638;
wire n_5825;
wire n_4018;
wire n_5491;
wire n_2987;
wire n_694;
wire n_2938;
wire n_3780;
wire n_5496;
wire n_5802;
wire n_7982;
wire n_12190;
wire n_12787;
wire n_8804;
wire n_297;
wire n_3337;
wire n_11383;
wire n_12799;
wire n_4002;
wire n_11847;
wire n_11976;
wire n_3209;
wire n_5178;
wire n_1044;
wire n_9317;
wire n_12657;
wire n_2165;
wire n_9769;
wire n_5547;
wire n_1391;
wire n_8158;
wire n_12511;
wire n_2750;
wire n_11167;
wire n_2775;
wire n_6879;
wire n_12532;
wire n_1295;
wire n_8469;
wire n_7567;
wire n_10238;
wire n_8765;
wire n_3477;
wire n_8433;
wire n_10102;
wire n_2349;
wire n_8931;
wire n_5596;
wire n_6074;
wire n_2684;
wire n_5983;
wire n_8213;
wire n_3146;
wire n_1495;
wire n_1438;
wire n_3953;
wire n_4588;
wire n_1100;
wire n_10534;
wire n_11825;
wire n_585;
wire n_4653;
wire n_4435;
wire n_10932;
wire n_10619;
wire n_7684;
wire n_11049;
wire n_5604;
wire n_1756;
wire n_8451;
wire n_1128;
wire n_5411;
wire n_673;
wire n_8334;
wire n_12743;
wire n_4019;
wire n_1071;
wire n_8731;
wire n_10589;
wire n_11611;
wire n_11681;
wire n_8385;
wire n_10890;
wire n_9156;
wire n_11202;
wire n_1968;
wire n_4728;
wire n_4999;
wire n_4385;
wire n_6642;
wire n_6847;
wire n_10707;
wire n_4922;
wire n_10552;
wire n_10248;
wire n_865;
wire n_3616;
wire n_5815;
wire n_7370;
wire n_9748;
wire n_6595;
wire n_4191;
wire n_7771;
wire n_9350;
wire n_12408;
wire n_11780;
wire n_5695;
wire n_6027;
wire n_2870;
wire n_8539;
wire n_10205;
wire n_2151;
wire n_7026;
wire n_7701;
wire n_7053;
wire n_1839;
wire n_2341;
wire n_9226;
wire n_1765;
wire n_3727;
wire n_5235;
wire n_10110;
wire n_2707;
wire n_6306;
wire n_11230;
wire n_6720;
wire n_11930;
wire n_10608;
wire n_11688;
wire n_6888;
wire n_826;
wire n_7173;
wire n_4350;
wire n_3747;
wire n_7042;
wire n_12715;
wire n_1714;
wire n_11709;
wire n_12434;
wire n_12628;
wire n_8122;
wire n_718;
wire n_6095;
wire n_8432;
wire n_11663;
wire n_5331;
wire n_4330;
wire n_7592;
wire n_542;
wire n_11331;
wire n_5311;
wire n_305;
wire n_12979;
wire n_9528;
wire n_6590;
wire n_2089;
wire n_10638;
wire n_7583;
wire n_12201;
wire n_3522;
wire n_6559;
wire n_12499;
wire n_2747;
wire n_3924;
wire n_9112;
wire n_12448;
wire n_791;
wire n_4621;
wire n_4216;
wire n_11876;
wire n_5797;
wire n_510;
wire n_9235;
wire n_10610;
wire n_11187;
wire n_4240;
wire n_12761;
wire n_3491;
wire n_5572;
wire n_1488;
wire n_9333;
wire n_704;
wire n_2148;
wire n_7151;
wire n_4162;
wire n_5565;
wire n_8950;
wire n_2339;
wire n_10758;
wire n_2861;
wire n_10190;
wire n_1999;
wire n_2731;
wire n_622;
wire n_5520;
wire n_147;
wire n_3353;
wire n_11804;
wire n_3018;
wire n_3975;
wire n_5800;
wire n_6562;
wire n_5984;
wire n_1838;
wire n_6287;
wire n_2638;
wire n_12809;
wire n_4785;
wire n_8347;
wire n_4683;
wire n_1766;
wire n_1776;
wire n_7353;
wire n_2002;
wire n_9330;
wire n_12538;
wire n_2138;
wire n_7758;
wire n_4021;
wire n_2414;
wire n_12446;
wire n_9490;
wire n_3014;
wire n_1771;
wire n_2316;
wire n_12029;
wire n_4103;
wire n_9355;
wire n_11052;
wire n_5060;
wire n_9523;
wire n_3148;
wire n_4022;
wire n_4986;
wire n_5888;
wire n_5669;
wire n_9024;
wire n_9574;
wire n_11694;
wire n_5772;
wire n_7571;
wire n_9582;
wire n_145;
wire n_2208;
wire n_4775;
wire n_5884;
wire n_10060;
wire n_6671;
wire n_11009;
wire n_6812;
wire n_12361;
wire n_4864;
wire n_9686;
wire n_9288;
wire n_9488;
wire n_5758;
wire n_10748;
wire n_4674;
wire n_13068;
wire n_4481;
wire n_6308;
wire n_7897;
wire n_11446;
wire n_10910;
wire n_1304;
wire n_10162;
wire n_294;
wire n_8242;
wire n_3775;
wire n_4669;
wire n_7118;
wire n_2134;
wire n_1176;
wire n_8284;
wire n_9964;
wire n_11540;
wire n_7792;
wire n_8161;
wire n_9702;
wire n_7510;
wire n_9819;
wire n_6662;
wire n_11291;
wire n_8184;
wire n_425;
wire n_5603;
wire n_9154;
wire n_6525;
wire n_7422;
wire n_13107;
wire n_1431;
wire n_3312;
wire n_3835;
wire n_6738;
wire n_4286;
wire n_12307;
wire n_13119;
wire n_5763;
wire n_2958;
wire n_10014;
wire n_8703;
wire n_7109;
wire n_12642;
wire n_3731;
wire n_1822;
wire n_2936;
wire n_3224;
wire n_12484;
wire n_6128;
wire n_2489;
wire n_6029;
wire n_1087;
wire n_8822;
wire n_10677;
wire n_12187;
wire n_657;
wire n_5751;
wire n_2771;
wire n_3020;
wire n_5264;
wire n_4525;
wire n_12321;
wire n_5924;
wire n_1505;
wire n_9992;
wire n_290;
wire n_11247;
wire n_7253;
wire n_8384;
wire n_5712;
wire n_6445;
wire n_3557;
wire n_2610;
wire n_12669;
wire n_13106;
wire n_3129;
wire n_8476;
wire n_6702;
wire n_11927;
wire n_3620;
wire n_11179;
wire n_478;
wire n_6701;
wire n_7339;
wire n_3832;
wire n_2520;
wire n_8359;
wire n_7380;
wire n_4484;
wire n_3693;
wire n_446;
wire n_8545;
wire n_8736;
wire n_9051;
wire n_4497;
wire n_7749;
wire n_10105;
wire n_1568;
wire n_2372;
wire n_1490;
wire n_10078;
wire n_11514;
wire n_12470;
wire n_12994;
wire n_11321;
wire n_9500;
wire n_8705;
wire n_10215;
wire n_526;
wire n_11779;
wire n_2251;
wire n_7508;
wire n_3674;
wire n_2959;
wire n_2501;
wire n_3203;
wire n_5694;
wire n_9455;
wire n_10251;
wire n_4871;
wire n_8708;
wire n_10834;
wire n_293;
wire n_7574;
wire n_1070;
wire n_2403;
wire n_2837;
wire n_4700;
wire n_4883;
wire n_9980;
wire n_1665;
wire n_4306;
wire n_11882;
wire n_11647;
wire n_154;
wire n_4224;
wire n_12064;
wire n_10706;
wire n_2127;
wire n_12462;
wire n_6005;
wire n_3341;
wire n_8872;
wire n_12696;
wire n_4453;
wire n_9555;
wire n_11133;
wire n_3559;
wire n_5449;
wire n_4005;
wire n_6169;
wire n_8238;
wire n_3546;
wire n_1358;
wire n_3661;
wire n_12735;
wire n_7713;
wire n_4564;
wire n_11222;
wire n_9200;
wire n_5146;
wire n_10709;
wire n_3056;
wire n_745;
wire n_2424;
wire n_12646;
wire n_3201;
wire n_10871;
wire n_3447;
wire n_7352;
wire n_3971;
wire n_5926;
wire n_716;
wire n_1774;
wire n_1475;
wire n_2354;
wire n_3103;
wire n_4573;
wire n_5398;
wire n_5860;
wire n_10304;
wire n_6936;
wire n_2589;
wire n_4535;
wire n_10244;
wire n_7704;
wire n_11571;
wire n_7487;
wire n_9986;
wire n_755;
wire n_8844;
wire n_13147;
wire n_6302;
wire n_527;
wire n_2442;
wire n_7641;
wire n_3627;
wire n_6106;
wire n_3480;
wire n_1368;
wire n_7203;
wire n_12999;
wire n_9397;
wire n_1137;
wire n_7169;
wire n_10407;
wire n_11259;
wire n_7670;
wire n_12682;
wire n_3612;
wire n_9673;
wire n_4695;
wire n_6848;
wire n_2545;
wire n_8642;
wire n_3509;
wire n_10043;
wire n_9855;
wire n_10568;
wire n_11875;
wire n_11941;
wire n_5919;
wire n_4368;
wire n_8159;
wire n_12111;
wire n_8912;
wire n_2966;
wire n_2294;
wire n_1942;
wire n_7439;
wire n_1314;
wire n_600;
wire n_9496;
wire n_3196;
wire n_8110;
wire n_864;
wire n_5319;
wire n_2504;
wire n_10796;
wire n_2623;
wire n_10016;
wire n_9008;
wire n_12903;
wire n_12079;
wire n_399;
wire n_6343;
wire n_12593;
wire n_1440;
wire n_5270;
wire n_2063;
wire n_10030;
wire n_8805;
wire n_1534;
wire n_6850;
wire n_12864;
wire n_5005;
wire n_9653;
wire n_11602;
wire n_10272;
wire n_8989;
wire n_9640;
wire n_6098;
wire n_12413;
wire n_6014;
wire n_7209;
wire n_7112;
wire n_1339;
wire n_2475;
wire n_11307;
wire n_5181;
wire n_6979;
wire n_7815;
wire n_403;
wire n_7934;
wire n_9545;
wire n_723;
wire n_3144;
wire n_8111;
wire n_3244;
wire n_596;
wire n_9629;
wire n_9603;
wire n_11578;
wire n_6865;
wire n_10432;
wire n_1141;
wire n_1268;
wire n_12719;
wire n_7276;
wire n_10342;
wire n_8056;
wire n_3287;
wire n_3322;
wire n_1755;
wire n_5043;
wire n_8739;
wire n_9674;
wire n_6747;
wire n_2357;
wire n_2025;
wire n_5583;
wire n_4654;
wire n_6433;
wire n_10462;
wire n_12725;
wire n_3640;
wire n_642;
wire n_1159;
wire n_995;
wire n_3481;
wire n_6640;
wire n_11769;
wire n_8856;
wire n_2250;
wire n_3033;
wire n_303;
wire n_6142;
wire n_9930;
wire n_11908;
wire n_12925;
wire n_5775;
wire n_6462;
wire n_7769;
wire n_2374;
wire n_416;
wire n_1681;
wire n_6034;
wire n_520;
wire n_9781;
wire n_418;
wire n_10291;
wire n_13159;
wire n_4597;
wire n_9659;
wire n_3364;
wire n_3226;
wire n_2780;
wire n_4020;
wire n_7233;
wire n_8732;
wire n_11913;
wire n_7602;
wire n_9296;
wire n_7034;
wire n_9897;
wire n_5220;
wire n_9241;
wire n_11341;
wire n_1618;
wire n_7390;
wire n_10787;
wire n_4867;
wire n_10669;
wire n_6870;
wire n_6221;
wire n_8231;
wire n_8185;
wire n_11466;
wire n_6279;
wire n_5061;
wire n_6775;
wire n_1653;
wire n_9291;
wire n_7881;
wire n_12290;
wire n_4063;
wire n_9906;
wire n_9369;
wire n_11982;
wire n_4237;
wire n_2601;
wire n_5029;
wire n_5127;
wire n_12317;
wire n_6071;
wire n_2920;
wire n_773;
wire n_11873;
wire n_7598;
wire n_9583;
wire n_12440;
wire n_920;
wire n_1374;
wire n_10185;
wire n_11182;
wire n_8908;
wire n_2648;
wire n_3212;
wire n_10092;
wire n_8220;
wire n_6833;
wire n_12150;
wire n_6793;
wire n_1169;
wire n_6767;
wire n_11815;
wire n_6295;
wire n_1617;
wire n_12782;
wire n_3370;
wire n_3386;
wire n_335;
wire n_4721;
wire n_11231;
wire n_463;
wire n_3093;
wire n_8090;
wire n_8053;
wire n_10184;
wire n_10111;
wire n_11991;
wire n_848;
wire n_12875;
wire n_274;
wire n_6385;
wire n_11354;
wire n_11807;
wire n_9262;
wire n_7426;
wire n_4247;
wire n_8137;
wire n_7045;
wire n_12027;
wire n_9851;
wire n_11799;
wire n_3169;
wire n_8740;
wire n_8009;
wire n_7852;
wire n_3205;
wire n_1881;
wire n_1267;
wire n_9987;
wire n_1806;
wire n_10983;
wire n_7984;
wire n_11727;
wire n_6788;
wire n_2023;
wire n_7014;
wire n_12192;
wire n_12633;
wire n_2204;
wire n_2720;
wire n_496;
wire n_10430;
wire n_8305;
wire n_4614;
wire n_177;
wire n_3360;
wire n_2087;
wire n_10277;
wire n_1636;
wire n_3956;
wire n_8163;
wire n_4001;
wire n_7220;
wire n_1323;
wire n_6709;
wire n_2627;
wire n_4422;
wire n_960;
wire n_10948;
wire n_11749;
wire n_6712;
wire n_6550;
wire n_10525;
wire n_9507;
wire n_11528;
wire n_7416;
wire n_11300;
wire n_6143;
wire n_778;
wire n_3004;
wire n_8841;
wire n_3870;
wire n_5177;
wire n_9657;
wire n_12551;
wire n_12196;
wire n_5483;
wire n_3625;
wire n_1764;
wire n_6743;
wire n_12497;
wire n_4632;
wire n_10354;
wire n_1610;
wire n_12412;
wire n_3084;
wire n_11880;
wire n_5785;
wire n_2343;
wire n_793;
wire n_7465;
wire n_5967;
wire n_4546;
wire n_10049;
wire n_12724;
wire n_4583;
wire n_4963;
wire n_3749;
wire n_6672;
wire n_9457;
wire n_2942;
wire n_4966;
wire n_9485;
wire n_5780;
wire n_4714;
wire n_7679;
wire n_5037;
wire n_2515;
wire n_7936;
wire n_8966;
wire n_316;
wire n_6084;
wire n_11249;
wire n_1551;
wire n_4847;
wire n_10287;
wire n_4054;
wire n_8538;
wire n_11039;
wire n_7738;
wire n_2555;
wire n_12101;
wire n_10119;
wire n_11145;
wire n_3586;
wire n_12606;
wire n_11986;
wire n_3653;
wire n_8395;
wire n_10900;
wire n_5966;
wire n_2201;
wire n_725;
wire n_10349;
wire n_6634;
wire n_3349;
wire n_4668;
wire n_5213;
wire n_8961;
wire n_10849;
wire n_7462;
wire n_4635;
wire n_368;
wire n_994;
wire n_5735;
wire n_12118;
wire n_7490;
wire n_11380;
wire n_2278;
wire n_7545;
wire n_1020;
wire n_10792;
wire n_11513;
wire n_8625;
wire n_1273;
wire n_7464;
wire n_7160;
wire n_8937;
wire n_4214;
wire n_9809;
wire n_6919;
wire n_10750;
wire n_3448;
wire n_7805;
wire n_10995;
wire n_617;
wire n_13092;
wire n_7115;
wire n_7295;
wire n_2924;
wire n_12087;
wire n_9192;
wire n_1036;
wire n_3595;
wire n_7348;
wire n_1138;
wire n_5752;
wire n_1661;
wire n_11618;
wire n_12594;
wire n_5360;
wire n_10673;
wire n_12460;
wire n_6681;
wire n_6104;
wire n_8179;
wire n_10537;
wire n_421;
wire n_11861;
wire n_3991;
wire n_6548;
wire n_3516;
wire n_3926;
wire n_6082;
wire n_6993;
wire n_1095;
wire n_8511;
wire n_6973;
wire n_12081;
wire n_1270;
wire n_10426;
wire n_4405;
wire n_610;
wire n_4413;
wire n_9558;
wire n_11594;
wire n_1852;
wire n_7453;
wire n_9167;
wire n_12082;
wire n_8715;
wire n_9655;
wire n_10241;
wire n_12474;
wire n_4036;
wire n_10684;
wire n_4759;
wire n_2153;
wire n_7162;
wire n_3670;
wire n_2381;
wire n_11436;
wire n_12346;
wire n_2052;
wire n_179;
wire n_4667;
wire n_5081;
wire n_517;
wire n_11729;
wire n_4182;
wire n_667;
wire n_3230;
wire n_8371;
wire n_8702;
wire n_8116;
wire n_1279;
wire n_1115;
wire n_7946;
wire n_8195;
wire n_1499;
wire n_8806;
wire n_11458;
wire n_12989;
wire n_12244;
wire n_504;
wire n_1409;
wire n_5877;
wire n_9991;
wire n_11670;
wire n_11366;
wire n_11872;
wire n_7681;
wire n_8845;
wire n_11504;
wire n_6018;
wire n_6619;
wire n_5189;
wire n_1503;
wire n_7702;
wire n_6676;
wire n_2819;
wire n_8149;
wire n_10823;
wire n_3041;
wire n_4637;
wire n_9976;
wire n_2423;
wire n_8042;
wire n_11516;
wire n_603;
wire n_10390;
wire n_12464;
wire n_11106;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_8392;
wire n_9560;
wire n_8095;
wire n_7210;
wire n_5869;
wire n_10830;
wire n_2439;
wire n_11132;
wire n_2404;
wire n_1182;
wire n_6718;
wire n_3635;
wire n_5118;
wire n_7503;
wire n_10824;
wire n_4155;
wire n_6854;
wire n_4238;
wire n_3011;
wire n_2061;
wire n_2757;
wire n_4977;
wire n_167;
wire n_5632;
wire n_8519;
wire n_5582;
wire n_5425;
wire n_5886;
wire n_8269;
wire n_1216;
wire n_2716;
wire n_6032;
wire n_9047;
wire n_12953;
wire n_2452;
wire n_12842;
wire n_3650;
wire n_8968;
wire n_12481;
wire n_9319;
wire n_9215;
wire n_11406;
wire n_5446;
wire n_11316;
wire n_3010;
wire n_7855;
wire n_3043;
wire n_11047;
wire n_8050;
wire n_12450;
wire n_5224;
wire n_12817;
wire n_4590;
wire n_8399;
wire n_2543;
wire n_5090;
wire n_3137;
wire n_9599;
wire n_11767;
wire n_2486;
wire n_3560;
wire n_10985;
wire n_11559;
wire n_9072;
wire n_3177;
wire n_4929;
wire n_9401;
wire n_5678;
wire n_12435;
wire n_9428;
wire n_10340;
wire n_10946;
wire n_11586;
wire n_6981;
wire n_2220;
wire n_7065;
wire n_2577;
wire n_12149;
wire n_9216;
wire n_1262;
wire n_3238;
wire n_218;
wire n_3529;
wire n_12002;
wire n_12836;
wire n_4835;
wire n_11519;
wire n_11109;
wire n_13065;
wire n_11229;
wire n_2232;
wire n_11591;
wire n_11961;
wire n_11195;
wire n_4038;
wire n_6122;
wire n_11225;
wire n_11397;
wire n_2790;
wire n_7911;
wire n_9747;
wire n_6765;
wire n_4565;
wire n_5414;
wire n_4159;
wire n_12840;
wire n_3784;
wire n_7330;
wire n_5437;
wire n_8883;
wire n_220;
wire n_10634;
wire n_8586;
wire n_12846;
wire n_9202;
wire n_4586;
wire n_11058;
wire n_9058;
wire n_1608;
wire n_7336;
wire n_11471;
wire n_2373;
wire n_1472;
wire n_7446;
wire n_3628;
wire n_8401;
wire n_7854;
wire n_10351;
wire n_5454;
wire n_8186;
wire n_10577;
wire n_800;
wire n_4734;
wire n_7493;
wire n_10961;
wire n_12940;
wire n_10460;
wire n_10780;
wire n_7357;
wire n_1491;
wire n_8756;
wire n_11324;
wire n_8737;
wire n_1840;
wire n_10334;
wire n_4434;
wire n_12945;
wire n_5307;
wire n_7923;
wire n_10379;
wire n_2244;
wire n_10151;
wire n_6439;
wire n_11614;
wire n_4290;
wire n_8602;
wire n_2586;
wire n_1684;
wire n_2446;
wire n_1346;
wire n_8240;
wire n_12850;
wire n_7714;
wire n_1352;
wire n_5407;
wire n_10411;
wire n_9484;
wire n_12984;
wire n_10989;
wire n_2017;
wire n_8422;
wire n_3029;
wire n_10939;
wire n_12224;
wire n_3597;
wire n_5913;
wire n_7088;
wire n_1046;
wire n_2560;
wire n_9305;
wire n_9394;
wire n_9999;
wire n_2704;
wire n_1145;
wire n_1121;
wire n_8878;
wire n_11144;
wire n_10090;
wire n_6406;
wire n_11361;
wire n_7440;
wire n_1102;
wire n_1963;
wire n_6945;
wire n_8112;
wire n_258;
wire n_11567;
wire n_3790;
wire n_10962;
wire n_7029;
wire n_2766;
wire n_260;
wire n_11128;
wire n_9622;
wire n_9292;
wire n_10721;
wire n_8593;
wire n_356;
wire n_12197;
wire n_10186;
wire n_3318;
wire n_4833;
wire n_11580;
wire n_11841;
wire n_11025;
wire n_12007;
wire n_5062;
wire n_6618;
wire n_6474;
wire n_13082;
wire n_10191;
wire n_5230;
wire n_5944;
wire n_6226;
wire n_152;
wire n_4888;
wire n_13094;
wire n_7317;
wire n_10856;
wire n_12403;
wire n_776;
wire n_321;
wire n_1823;
wire n_2479;
wire n_3350;
wire n_6000;
wire n_2782;
wire n_12679;
wire n_9584;
wire n_3977;
wire n_227;
wire n_8194;
wire n_9461;
wire n_11168;
wire n_8055;
wire n_8579;
wire n_6816;
wire n_10914;
wire n_10911;
wire n_10928;
wire n_12756;
wire n_8360;
wire n_3588;
wire n_4279;
wire n_5008;
wire n_12018;
wire n_6425;
wire n_1456;
wire n_5004;
wire n_5294;
wire n_6493;
wire n_9845;
wire n_6502;
wire n_6250;
wire n_7374;
wire n_6288;
wire n_5974;
wire n_11937;
wire n_12872;
wire n_7522;
wire n_6492;
wire n_2229;
wire n_10071;
wire n_8755;
wire n_4133;
wire n_4527;
wire n_2288;
wire n_6046;
wire n_11460;
wire n_2099;
wire n_8251;
wire n_5323;
wire n_11565;
wire n_3388;
wire n_4790;
wire n_1946;
wire n_4181;
wire n_3184;
wire n_12372;
wire n_9618;
wire n_6118;
wire n_5810;
wire n_4561;
wire n_4461;
wire n_464;
wire n_3245;
wire n_3075;
wire n_7046;
wire n_11192;
wire n_11808;
wire n_4007;
wire n_10956;
wire n_4949;
wire n_6852;
wire n_2642;
wire n_4239;
wire n_8677;
wire n_13052;
wire n_7468;
wire n_9091;
wire n_11013;
wire n_2383;
wire n_5991;
wire n_4184;
wire n_1676;
wire n_1830;
wire n_2351;
wire n_1319;
wire n_5069;
wire n_12453;
wire n_12572;
wire n_2986;
wire n_5702;
wire n_10035;
wire n_6251;
wire n_9828;
wire n_2536;
wire n_3915;
wire n_139;
wire n_1633;
wire n_9699;
wire n_12340;
wire n_3489;
wire n_8108;
wire n_2835;
wire n_5243;
wire n_1416;
wire n_5914;
wire n_2820;
wire n_2293;
wire n_12955;
wire n_12068;
wire n_10252;
wire n_5250;
wire n_11555;
wire n_3074;
wire n_6869;
wire n_3102;
wire n_10041;
wire n_9321;
wire n_5590;
wire n_10345;
wire n_2026;
wire n_1282;
wire n_10059;
wire n_5260;
wire n_8325;
wire n_9751;
wire n_7621;
wire n_8498;
wire n_7359;
wire n_550;
wire n_3321;
wire n_2567;
wire n_5809;
wire n_2322;
wire n_10543;
wire n_275;
wire n_2727;
wire n_3377;
wire n_7924;
wire n_560;
wire n_4782;
wire n_12394;
wire n_1321;
wire n_7659;
wire n_2533;
wire n_569;
wire n_3530;
wire n_9161;
wire n_9005;
wire n_2869;
wire n_8875;
wire n_4378;
wire n_5349;
wire n_8274;
wire n_9585;
wire n_7153;
wire n_11101;
wire n_1235;
wire n_2759;
wire n_12954;
wire n_7836;
wire n_2361;
wire n_10737;
wire n_1292;
wire n_12662;
wire n_2266;
wire n_4876;
wire n_6146;
wire n_8504;
wire n_346;
wire n_10464;
wire n_10644;
wire n_7280;
wire n_12801;
wire n_5813;
wire n_9293;
wire n_12503;
wire n_10365;
wire n_790;
wire n_5833;
wire n_11781;
wire n_2611;
wire n_2901;
wire n_11055;
wire n_7886;
wire n_4358;
wire n_10982;
wire n_5616;
wire n_5805;
wire n_9648;
wire n_2653;
wire n_12871;
wire n_6884;
wire n_7664;
wire n_7012;
wire n_299;
wire n_1248;
wire n_12965;
wire n_13029;
wire n_10591;
wire n_11845;
wire n_12486;
wire n_902;
wire n_2189;
wire n_2246;
wire n_6631;
wire n_12788;
wire n_12369;
wire n_4469;
wire n_9498;
wire n_7376;
wire n_7577;
wire n_7308;
wire n_5169;
wire n_431;
wire n_5816;
wire n_3156;
wire n_10809;
wire n_8927;
wire n_10899;
wire n_672;
wire n_9639;
wire n_11898;
wire n_10137;
wire n_12084;
wire n_12686;
wire n_6228;
wire n_11997;
wire n_1941;
wire n_3483;
wire n_11884;
wire n_5416;
wire n_8946;
wire n_6711;
wire n_13090;
wire n_12822;
wire n_706;
wire n_1794;
wire n_1236;
wire n_11863;
wire n_4493;
wire n_4924;
wire n_7279;
wire n_7971;
wire n_9646;
wire n_8017;
wire n_743;
wire n_766;
wire n_12264;
wire n_11761;
wire n_430;
wire n_1746;
wire n_8474;
wire n_9984;
wire n_3524;
wire n_8232;
wire n_7275;
wire n_489;
wire n_2885;
wire n_8795;
wire n_7195;
wire n_10600;
wire n_10794;
wire n_6102;
wire n_636;
wire n_9649;
wire n_8904;
wire n_11199;
wire n_6274;
wire n_10833;
wire n_8838;
wire n_11264;
wire n_12109;
wire n_10629;
wire n_9562;
wire n_3097;
wire n_7007;
wire n_660;
wire n_2062;
wire n_7070;
wire n_4539;
wire n_2975;
wire n_8382;
wire n_4421;
wire n_13023;
wire n_7610;
wire n_6072;
wire n_12303;
wire n_2839;
wire n_9501;
wire n_11896;
wire n_2856;
wire n_4793;
wire n_4498;
wire n_10006;
wire n_2070;
wire n_11757;
wire n_7259;
wire n_12320;
wire n_1607;
wire n_12274;
wire n_1454;
wire n_9759;
wire n_6353;
wire n_4953;
wire n_12622;
wire n_11185;
wire n_6992;
wire n_2348;
wire n_2944;
wire n_8128;
wire n_12659;
wire n_6818;
wire n_3831;
wire n_869;
wire n_1154;
wire n_646;
wire n_528;
wire n_391;
wire n_10206;
wire n_1329;
wire n_6322;
wire n_5167;
wire n_5661;
wire n_5932;
wire n_5830;
wire n_3589;
wire n_262;
wire n_11345;
wire n_12380;
wire n_897;
wire n_846;
wire n_2066;
wire n_7539;
wire n_841;
wire n_1476;
wire n_12586;
wire n_3391;
wire n_12629;
wire n_8794;
wire n_11760;
wire n_7616;
wire n_508;
wire n_1800;
wire n_9733;
wire n_12868;
wire n_12282;
wire n_8189;
wire n_6498;
wire n_1463;
wire n_8481;
wire n_10275;
wire n_11081;
wire n_3458;
wire n_7775;
wire n_13011;
wire n_4505;
wire n_11392;
wire n_9981;
wire n_3190;
wire n_1562;
wire n_7930;
wire n_5558;
wire n_1826;
wire n_8787;
wire n_5687;
wire n_7661;
wire n_6378;
wire n_5383;
wire n_5126;
wire n_1759;
wire n_8205;
wire n_5051;
wire n_9907;
wire n_13088;
wire n_5587;
wire n_6976;
wire n_10941;
wire n_11024;
wire n_6304;
wire n_5236;
wire n_12269;
wire n_853;
wire n_7640;
wire n_9816;
wire n_10498;
wire n_875;
wire n_11424;
wire n_12585;
wire n_5012;
wire n_1678;
wire n_11463;
wire n_10292;
wire n_661;
wire n_6864;
wire n_8605;
wire n_11278;
wire n_7969;
wire n_10358;
wire n_3787;
wire n_1256;
wire n_7548;
wire n_3585;
wire n_10635;
wire n_3565;
wire n_9944;
wire n_4450;
wire n_5954;
wire n_6156;
wire n_12832;
wire n_12913;
wire n_5025;
wire n_933;
wire n_6998;
wire n_8067;
wire n_7587;
wire n_7064;
wire n_4173;
wire n_12301;
wire n_3135;
wire n_12338;
wire n_9643;
wire n_7615;
wire n_5651;
wire n_6930;
wire n_4630;
wire n_9605;
wire n_12802;
wire n_12154;
wire n_8000;
wire n_11569;
wire n_10064;
wire n_1217;
wire n_7197;
wire n_5645;
wire n_9676;
wire n_3990;
wire n_11881;
wire n_7393;
wire n_11332;
wire n_6917;
wire n_6937;
wire n_7591;
wire n_310;
wire n_1628;
wire n_9963;
wire n_5766;
wire n_11404;
wire n_2109;
wire n_7727;
wire n_7358;
wire n_988;
wire n_2796;
wire n_7324;
wire n_2507;
wire n_9950;
wire n_5878;
wire n_5671;
wire n_10152;
wire n_11935;
wire n_4534;
wire n_1536;
wire n_6301;
wire n_9788;
wire n_1204;
wire n_1132;
wire n_6929;
wire n_233;
wire n_11309;
wire n_1327;
wire n_8719;
wire n_955;
wire n_8045;
wire n_10785;
wire n_7729;
wire n_246;
wire n_2787;
wire n_2969;
wire n_2395;
wire n_12341;
wire n_12615;
wire n_1554;
wire n_4494;
wire n_6436;
wire n_5412;
wire n_8209;
wire n_10802;
wire n_769;
wire n_2380;
wire n_4786;
wire n_10815;
wire n_7565;
wire n_1120;
wire n_6699;
wire n_12926;
wire n_9213;
wire n_555;
wire n_4579;
wire n_7291;
wire n_7631;
wire n_669;
wire n_8784;
wire n_2290;
wire n_7382;
wire n_4811;
wire n_2048;
wire n_176;
wire n_6874;
wire n_7387;
wire n_6259;
wire n_9212;
wire n_9340;
wire n_2005;
wire n_12167;
wire n_9473;
wire n_4857;
wire n_13026;
wire n_10490;
wire n_7437;
wire n_6677;
wire n_12161;
wire n_3432;
wire n_12085;
wire n_2736;
wire n_2883;
wire n_11735;
wire n_1408;
wire n_7618;
wire n_4282;
wire n_1196;
wire n_10647;
wire n_3493;
wire n_9320;
wire n_10523;
wire n_8769;
wire n_8575;
wire n_6764;
wire n_12298;
wire n_10081;
wire n_863;
wire n_3774;
wire n_5733;
wire n_10324;
wire n_6780;
wire n_11189;
wire n_8815;
wire n_11582;
wire n_12569;
wire n_2910;
wire n_6620;
wire n_6597;
wire n_12044;
wire n_748;
wire n_3268;
wire n_1785;
wire n_9303;
wire n_1147;
wire n_11105;
wire n_1754;
wire n_3057;
wire n_11705;
wire n_3701;
wire n_5148;
wire n_8261;
wire n_2584;
wire n_7673;
wire n_1812;
wire n_6830;
wire n_866;
wire n_12456;
wire n_13104;
wire n_8655;
wire n_7282;
wire n_2287;
wire n_452;
wire n_9968;
wire n_10808;
wire n_11474;
wire n_6586;
wire n_6333;
wire n_10474;
wire n_7139;
wire n_8745;
wire n_12689;
wire n_5791;
wire n_5727;
wire n_10657;
wire n_8086;
wire n_761;
wire n_5946;
wire n_8789;
wire n_5997;
wire n_2492;
wire n_7953;
wire n_3778;
wire n_6428;
wire n_5328;
wire n_7379;
wire n_10687;
wire n_9722;
wire n_12042;
wire n_12155;
wire n_5657;
wire n_174;
wire n_1173;
wire n_8901;
wire n_11078;
wire n_11130;
wire n_8695;
wire n_4974;
wire n_12373;
wire n_5975;
wire n_4911;
wire n_8173;
wire n_11664;
wire n_12072;
wire n_12110;
wire n_4436;
wire n_8363;
wire n_5119;
wire n_10652;
wire n_4569;
wire n_10545;
wire n_9669;
wire n_1174;
wire n_8665;
wire n_13098;
wire n_6510;
wire n_8282;
wire n_3334;
wire n_9388;
wire n_5938;
wire n_6237;
wire n_12040;
wire n_11752;
wire n_12216;
wire n_12654;
wire n_5602;
wire n_647;
wire n_9379;
wire n_11992;
wire n_5097;
wire n_844;
wire n_4985;
wire n_7751;
wire n_2117;
wire n_2234;
wire n_10869;
wire n_3823;
wire n_4384;
wire n_3114;
wire n_2741;
wire n_13142;
wire n_7581;
wire n_888;
wire n_13116;
wire n_11783;
wire n_6360;
wire n_2203;
wire n_2255;
wire n_3584;
wire n_5246;
wire n_10453;
wire n_236;
wire n_12386;
wire n_4858;
wire n_4678;
wire n_9952;
wire n_2649;
wire n_3556;
wire n_9911;
wire n_12183;
wire n_3836;
wire n_5579;
wire n_8835;
wire n_414;
wire n_1922;
wire n_9256;
wire n_10668;
wire n_10346;
wire n_12419;
wire n_5750;
wire n_10688;
wire n_4823;
wire n_5831;
wire n_4309;
wire n_4363;
wire n_7742;
wire n_9274;
wire n_1215;
wire n_12964;
wire n_839;
wire n_10473;
wire n_5107;
wire n_3456;
wire n_5095;
wire n_8493;
wire n_7346;
wire n_10331;
wire n_11439;
wire n_779;
wire n_1537;
wire n_10957;
wire n_2205;
wire n_4243;
wire n_7579;
wire n_12863;
wire n_10352;
wire n_4025;
wire n_11188;
wire n_7428;
wire n_3404;
wire n_1122;
wire n_5666;
wire n_12221;
wire n_4059;
wire n_9195;
wire n_10442;
wire n_1509;
wire n_11687;
wire n_4121;
wire n_3290;
wire n_1109;
wire n_8870;
wire n_7150;
wire n_7155;
wire n_8252;
wire n_11774;
wire n_4313;
wire n_3309;
wire n_4142;
wire n_3671;
wire n_2015;
wire n_6475;
wire n_7015;
wire n_3982;
wire n_7699;
wire n_8507;
wire n_6314;
wire n_8415;
wire n_10632;
wire n_9623;
wire n_6103;
wire n_2609;
wire n_1161;
wire n_5546;
wire n_7249;
wire n_10713;
wire n_3796;
wire n_232;
wire n_6394;
wire n_8781;
wire n_6964;
wire n_3840;
wire n_3461;
wire n_6680;
wire n_3408;
wire n_7985;
wire n_10954;
wire n_4246;
wire n_12267;
wire n_7432;
wire n_8365;
wire n_3513;
wire n_3690;
wire n_1184;
wire n_2483;
wire n_4532;
wire n_228;
wire n_8893;
wire n_1525;
wire n_6372;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_11329;
wire n_5994;
wire n_6495;
wire n_7194;
wire n_9516;
wire n_4244;
wire n_2147;
wire n_592;
wire n_13162;
wire n_2503;
wire n_4049;
wire n_6752;
wire n_1156;
wire n_12768;
wire n_8976;
wire n_6426;
wire n_2600;
wire n_984;
wire n_7505;
wire n_5626;
wire n_3508;
wire n_8025;
wire n_8502;
wire n_10165;
wire n_8244;
wire n_10130;
wire n_7612;
wire n_8156;
wire n_11661;
wire n_7494;
wire n_868;
wire n_4353;
wire n_11120;
wire n_9222;
wire n_735;
wire n_13031;
wire n_8435;
wire n_6350;
wire n_8882;
wire n_4787;
wire n_7736;
wire n_10622;
wire n_5633;
wire n_13155;
wire n_9546;
wire n_469;
wire n_1218;
wire n_5664;
wire n_7589;
wire n_5921;
wire n_6797;
wire n_3596;
wire n_4537;
wire n_4346;
wire n_8759;
wire n_4351;
wire n_6159;
wire n_7814;
wire n_7177;
wire n_357;
wire n_13066;
wire n_8660;
wire n_2429;
wire n_11296;
wire n_8479;
wire n_985;
wire n_12993;
wire n_2440;
wire n_13124;
wire n_6054;
wire n_11095;
wire n_3521;
wire n_11314;
wire n_8723;
wire n_802;
wire n_11019;
wire n_561;
wire n_8606;
wire n_9663;
wire n_980;
wire n_2681;
wire n_6235;
wire n_7843;
wire n_8235;
wire n_13083;
wire n_1651;
wire n_2360;
wire n_3764;
wire n_12647;
wire n_7662;
wire n_4784;
wire n_6152;
wire n_4075;
wire n_9820;
wire n_7773;
wire n_7902;
wire n_5340;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_9743;
wire n_6496;
wire n_3066;
wire n_7756;
wire n_2844;
wire n_12749;
wire n_8342;
wire n_8940;
wire n_2303;
wire n_1619;
wire n_13048;
wire n_11584;
wire n_2285;
wire n_5280;
wire n_8448;
wire n_8472;
wire n_7700;
wire n_4451;
wire n_4332;
wire n_810;
wire n_7555;
wire n_10000;
wire n_1194;
wire n_4538;
wire n_4506;
wire n_10158;
wire n_2742;
wire n_10582;
wire n_12066;
wire n_12812;
wire n_3695;
wire n_10427;
wire n_11816;
wire n_12060;
wire n_3976;
wire n_10199;
wire n_7988;
wire n_8658;
wire n_3563;
wire n_6513;
wire n_10246;
wire n_2367;
wire n_7500;
wire n_11910;
wire n_201;
wire n_3198;
wire n_11693;
wire n_3495;
wire n_1034;
wire n_5925;
wire n_2909;
wire n_9248;
wire n_754;
wire n_6138;
wire n_5369;
wire n_8866;
wire n_10835;
wire n_9822;
wire n_8061;
wire n_975;
wire n_5730;
wire n_11411;
wire n_5576;
wire n_11184;
wire n_11386;
wire n_11945;
wire n_11604;
wire n_3359;
wire n_12164;
wire n_5272;
wire n_11368;
wire n_10125;
wire n_12824;
wire n_13111;
wire n_6330;
wire n_10117;
wire n_9065;
wire n_467;
wire n_3187;
wire n_12716;
wire n_10844;
wire n_3218;
wire n_8457;
wire n_6802;
wire n_10654;
wire n_9086;
wire n_9153;
wire n_10505;
wire n_9339;
wire n_582;
wire n_10198;
wire n_861;
wire n_7157;
wire n_11064;
wire n_6909;
wire n_6908;
wire n_857;
wire n_8237;
wire n_7411;
wire n_9601;
wire n_9093;
wire n_11409;
wire n_2107;
wire n_2040;
wire n_2968;
wire n_4201;
wire n_4336;
wire n_7266;
wire n_2221;
wire n_8046;
wire n_588;
wire n_7871;
wire n_5646;
wire n_12051;
wire n_11097;
wire n_12437;
wire n_5624;
wire n_4852;
wire n_1010;
wire n_4210;
wire n_4981;
wire n_10840;
wire n_12052;
wire n_6477;
wire n_9746;
wire n_6263;
wire n_10515;
wire n_8073;
wire n_1166;
wire n_5440;
wire n_2891;
wire n_6490;
wire n_11533;
wire n_11605;
wire n_2709;
wire n_8652;
wire n_9198;
wire n_8821;
wire n_534;
wire n_7198;
wire n_1578;
wire n_8335;
wire n_1861;
wire n_9904;
wire n_10242;
wire n_9142;
wire n_9440;
wire n_10144;
wire n_3955;
wire n_9684;
wire n_1557;
wire n_2280;
wire n_3945;
wire n_6184;
wire n_730;
wire n_5817;
wire n_5214;
wire n_203;
wire n_10973;
wire n_1898;
wire n_2443;
wire n_4936;
wire n_4205;
wire n_2162;
wire n_1868;
wire n_207;
wire n_2079;
wire n_9493;
wire n_4763;
wire n_3587;
wire n_4278;
wire n_5586;
wire n_11036;
wire n_8663;
wire n_3433;
wire n_11330;
wire n_12720;
wire n_4463;
wire n_7794;
wire n_10267;
wire n_205;
wire n_2185;
wire n_6038;
wire n_10551;
wire n_5861;
wire n_1836;
wire n_3833;
wire n_10553;
wire n_2774;
wire n_13127;
wire n_3162;
wire n_1274;
wire n_8309;
wire n_1486;
wire n_3333;
wire n_4129;
wire n_5258;
wire n_8945;
wire n_11002;
wire n_6605;
wire n_12687;
wire n_5032;
wire n_8964;
wire n_10988;
wire n_1899;
wire n_9032;
wire n_9814;
wire n_6313;
wire n_784;
wire n_4804;
wire n_5619;
wire n_6112;
wire n_3965;
wire n_7145;
wire n_9041;
wire n_5859;
wire n_12325;
wire n_5380;
wire n_4500;
wire n_9245;
wire n_5065;
wire n_862;
wire n_5776;
wire n_8166;
wire n_2098;
wire n_3085;
wire n_4433;
wire n_5606;
wire n_9357;
wire n_5644;
wire n_11796;
wire n_2813;
wire n_1935;
wire n_5826;
wire n_2027;
wire n_10108;
wire n_2091;
wire n_8960;
wire n_12789;
wire n_5920;
wire n_2991;
wire n_10307;
wire n_5030;
wire n_4194;
wire n_7994;
wire n_1449;
wire n_4703;
wire n_8443;
wire n_361;
wire n_7349;
wire n_9598;
wire n_8215;
wire n_7715;
wire n_2419;
wire n_6180;
wire n_8683;
wire n_8809;
wire n_5683;
wire n_6349;
wire n_10510;
wire n_2677;
wire n_12127;
wire n_12382;
wire n_12504;
wire n_3182;
wire n_5756;
wire n_12602;
wire n_3283;
wire n_5527;
wire n_6476;
wire n_8037;
wire n_12062;
wire n_1742;
wire n_4030;
wire n_12573;

INVx1_ASAP7_75t_L g136 ( 
.A(n_94),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_36),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_28),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_7),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_105),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_92),
.Y(n_142)
);

BUFx10_ASAP7_75t_L g143 ( 
.A(n_98),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_69),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_131),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_79),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g147 ( 
.A(n_101),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_6),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_112),
.Y(n_149)
);

BUFx2_ASAP7_75t_SL g150 ( 
.A(n_66),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_114),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_26),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_73),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_55),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_110),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_20),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

INVxp33_ASAP7_75t_L g158 ( 
.A(n_20),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_62),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_23),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_67),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_42),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_2),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_7),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_43),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_49),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_27),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_18),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_58),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_29),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_106),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_118),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_133),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_14),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g175 ( 
.A(n_52),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_119),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_54),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_38),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_1),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_72),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_113),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_70),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_17),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_84),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_132),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_93),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_89),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_44),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_117),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_115),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_13),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_5),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_53),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_1),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_14),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_103),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_65),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_33),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_56),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_86),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_40),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_15),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_34),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_10),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_111),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_134),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_16),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_75),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_91),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_30),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_122),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_39),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_50),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_81),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_97),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_127),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_121),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_4),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_57),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_124),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_48),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_126),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_3),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_90),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_6),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_87),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_8),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_2),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_64),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_17),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_10),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_76),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_24),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_13),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_18),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_37),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_8),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_31),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_104),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_96),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_78),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_125),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_15),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_128),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_116),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_68),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_59),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_41),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_107),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_85),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_47),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_5),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_46),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_25),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_129),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_16),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_51),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_135),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_100),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_83),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_35),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_120),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_77),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_82),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_130),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_109),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_22),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_19),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_102),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_168),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_168),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_140),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_148),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_268),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_244),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_175),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_187),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_175),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_175),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_268),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_163),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_268),
.Y(n_282)
);

NOR2xp67_ASAP7_75t_L g283 ( 
.A(n_164),
.B(n_0),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_268),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_174),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_229),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_183),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_202),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_223),
.Y(n_289)
);

BUFx8_ASAP7_75t_SL g290 ( 
.A(n_227),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_175),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_153),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_234),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_243),
.Y(n_294)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_179),
.Y(n_295)
);

NOR2xp67_ASAP7_75t_L g296 ( 
.A(n_252),
.B(n_0),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_256),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_188),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_244),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_191),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_192),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_195),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_136),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_137),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_204),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_139),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_207),
.Y(n_307)
);

CKINVDCx14_ASAP7_75t_R g308 ( 
.A(n_143),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_218),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_225),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_228),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_157),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_295),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_274),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_292),
.Y(n_315)
);

NOR2xp67_ASAP7_75t_L g316 ( 
.A(n_272),
.B(n_159),
.Y(n_316)
);

INVxp33_ASAP7_75t_SL g317 ( 
.A(n_286),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_280),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_277),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_282),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_290),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_282),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_284),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_308),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_272),
.Y(n_325)
);

NOR2xp67_ASAP7_75t_L g326 ( 
.A(n_273),
.B(n_263),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_284),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_303),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_304),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_273),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_275),
.B(n_188),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_295),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_306),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_312),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_281),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_285),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_287),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_288),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_289),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_293),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_275),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_281),
.Y(n_342)
);

INVxp67_ASAP7_75t_SL g343 ( 
.A(n_299),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_300),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_294),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_297),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g347 ( 
.A(n_270),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_300),
.B(n_153),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_271),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_298),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_298),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_276),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_276),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_301),
.B(n_238),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_301),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_302),
.B(n_254),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_302),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_305),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_278),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_305),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_349),
.Y(n_361)
);

OAI21x1_ASAP7_75t_L g362 ( 
.A1(n_352),
.A2(n_291),
.B(n_278),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_353),
.B(n_279),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_336),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_359),
.B(n_279),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_314),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_325),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_318),
.Y(n_368)
);

AND2x6_ASAP7_75t_L g369 ( 
.A(n_331),
.B(n_239),
.Y(n_369)
);

AND2x4_ASAP7_75t_L g370 ( 
.A(n_343),
.B(n_283),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_322),
.B(n_291),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_337),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_338),
.Y(n_373)
);

AND2x2_ASAP7_75t_SL g374 ( 
.A(n_341),
.B(n_189),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_350),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_317),
.B(n_307),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_322),
.B(n_175),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_339),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_320),
.B(n_175),
.Y(n_379)
);

AND2x4_ASAP7_75t_L g380 ( 
.A(n_347),
.B(n_296),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_323),
.B(n_175),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_340),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_344),
.Y(n_383)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_350),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_345),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_327),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_350),
.B(n_351),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_358),
.Y(n_388)
);

AND2x4_ASAP7_75t_L g389 ( 
.A(n_346),
.B(n_160),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_328),
.Y(n_390)
);

AND2x4_ASAP7_75t_L g391 ( 
.A(n_316),
.B(n_173),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_329),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_333),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_350),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_334),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_313),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_332),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_354),
.Y(n_398)
);

AND2x2_ASAP7_75t_SL g399 ( 
.A(n_356),
.B(n_236),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_326),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_317),
.B(n_239),
.Y(n_401)
);

AND2x4_ASAP7_75t_L g402 ( 
.A(n_330),
.B(n_177),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_360),
.B(n_241),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_335),
.B(n_241),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_319),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_335),
.Y(n_406)
);

BUFx2_ASAP7_75t_L g407 ( 
.A(n_342),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_355),
.Y(n_408)
);

INVx2_ASAP7_75t_SL g409 ( 
.A(n_355),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_342),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_319),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_357),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_357),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_324),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_324),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_348),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_315),
.Y(n_417)
);

INVx2_ASAP7_75t_SL g418 ( 
.A(n_315),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_321),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_321),
.Y(n_420)
);

OA21x2_ASAP7_75t_L g421 ( 
.A1(n_352),
.A2(n_206),
.B(n_205),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_350),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_350),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_349),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_314),
.Y(n_425)
);

OA21x2_ASAP7_75t_L g426 ( 
.A1(n_352),
.A2(n_203),
.B(n_200),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_349),
.Y(n_427)
);

OA21x2_ASAP7_75t_L g428 ( 
.A1(n_352),
.A2(n_193),
.B(n_186),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_343),
.B(n_185),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_341),
.B(n_307),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_349),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_317),
.B(n_309),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_331),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_352),
.B(n_215),
.Y(n_434)
);

AND2x4_ASAP7_75t_L g435 ( 
.A(n_343),
.B(n_217),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_314),
.Y(n_436)
);

BUFx8_ASAP7_75t_L g437 ( 
.A(n_349),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_350),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_350),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_352),
.B(n_220),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_350),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_314),
.Y(n_442)
);

BUFx8_ASAP7_75t_L g443 ( 
.A(n_349),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_349),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_349),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_350),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_314),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_350),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_341),
.B(n_309),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_350),
.Y(n_450)
);

OR2x2_ASAP7_75t_L g451 ( 
.A(n_341),
.B(n_310),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_349),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_354),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_352),
.B(n_222),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_314),
.Y(n_455)
);

BUFx12f_ASAP7_75t_L g456 ( 
.A(n_319),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_352),
.B(n_224),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_349),
.Y(n_458)
);

AND2x4_ASAP7_75t_L g459 ( 
.A(n_343),
.B(n_240),
.Y(n_459)
);

OAI21x1_ASAP7_75t_L g460 ( 
.A1(n_352),
.A2(n_259),
.B(n_265),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_325),
.Y(n_461)
);

NAND3xp33_ASAP7_75t_L g462 ( 
.A(n_331),
.B(n_154),
.C(n_211),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_349),
.Y(n_463)
);

OA21x2_ASAP7_75t_L g464 ( 
.A1(n_352),
.A2(n_161),
.B(n_226),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_331),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_314),
.Y(n_466)
);

CKINVDCx11_ASAP7_75t_R g467 ( 
.A(n_321),
.Y(n_467)
);

OA21x2_ASAP7_75t_L g468 ( 
.A1(n_352),
.A2(n_214),
.B(n_201),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_350),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_314),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_352),
.B(n_150),
.Y(n_471)
);

INVx4_ASAP7_75t_L g472 ( 
.A(n_350),
.Y(n_472)
);

OA21x2_ASAP7_75t_L g473 ( 
.A1(n_352),
.A2(n_149),
.B(n_199),
.Y(n_473)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_349),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_349),
.Y(n_475)
);

AND2x4_ASAP7_75t_L g476 ( 
.A(n_343),
.B(n_165),
.Y(n_476)
);

BUFx2_ASAP7_75t_L g477 ( 
.A(n_342),
.Y(n_477)
);

AOI22x1_ASAP7_75t_SL g478 ( 
.A1(n_321),
.A2(n_227),
.B1(n_165),
.B2(n_249),
.Y(n_478)
);

AND2x4_ASAP7_75t_L g479 ( 
.A(n_343),
.B(n_178),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_352),
.B(n_147),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_343),
.B(n_178),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_349),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_349),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_343),
.B(n_181),
.Y(n_484)
);

AND2x4_ASAP7_75t_L g485 ( 
.A(n_343),
.B(n_181),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_352),
.B(n_184),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_349),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_349),
.Y(n_488)
);

INVx5_ASAP7_75t_L g489 ( 
.A(n_350),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_350),
.Y(n_490)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_331),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_352),
.B(n_232),
.Y(n_492)
);

AO22x2_ASAP7_75t_L g493 ( 
.A1(n_401),
.A2(n_194),
.B1(n_156),
.B2(n_258),
.Y(n_493)
);

AO22x2_ASAP7_75t_L g494 ( 
.A1(n_401),
.A2(n_158),
.B1(n_4),
.B2(n_9),
.Y(n_494)
);

NAND3x1_ASAP7_75t_L g495 ( 
.A(n_376),
.B(n_158),
.C(n_249),
.Y(n_495)
);

OAI22xp33_ASAP7_75t_SL g496 ( 
.A1(n_404),
.A2(n_310),
.B1(n_311),
.B2(n_267),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g497 ( 
.A1(n_399),
.A2(n_245),
.B1(n_311),
.B2(n_176),
.Y(n_497)
);

NAND3x1_ASAP7_75t_L g498 ( 
.A(n_376),
.B(n_245),
.C(n_143),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_386),
.Y(n_499)
);

OAI22xp33_ASAP7_75t_SL g500 ( 
.A1(n_404),
.A2(n_453),
.B1(n_403),
.B2(n_398),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_399),
.A2(n_237),
.B1(n_235),
.B2(n_231),
.Y(n_501)
);

BUFx6f_ASAP7_75t_SL g502 ( 
.A(n_405),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_453),
.B(n_144),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_364),
.Y(n_504)
);

AO22x2_ASAP7_75t_L g505 ( 
.A1(n_478),
.A2(n_3),
.B1(n_9),
.B2(n_11),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_432),
.B(n_230),
.Y(n_506)
);

OAI22xp33_ASAP7_75t_L g507 ( 
.A1(n_433),
.A2(n_145),
.B1(n_144),
.B2(n_266),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_362),
.Y(n_508)
);

AO22x2_ASAP7_75t_L g509 ( 
.A1(n_406),
.A2(n_11),
.B1(n_12),
.B2(n_19),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_403),
.B(n_145),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_433),
.A2(n_172),
.B1(n_262),
.B2(n_261),
.Y(n_511)
);

OR2x2_ASAP7_75t_L g512 ( 
.A(n_396),
.B(n_12),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_458),
.Y(n_513)
);

OAI22xp33_ASAP7_75t_L g514 ( 
.A1(n_465),
.A2(n_171),
.B1(n_260),
.B2(n_257),
.Y(n_514)
);

INVx2_ASAP7_75t_SL g515 ( 
.A(n_370),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_432),
.B(n_143),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_372),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_430),
.B(n_170),
.Y(n_518)
);

OAI22xp33_ASAP7_75t_SL g519 ( 
.A1(n_400),
.A2(n_180),
.B1(n_255),
.B2(n_253),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_465),
.A2(n_491),
.B1(n_370),
.B2(n_380),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_491),
.A2(n_167),
.B1(n_251),
.B2(n_250),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_449),
.B(n_166),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_380),
.B(n_162),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_397),
.A2(n_169),
.B1(n_248),
.B2(n_247),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_476),
.B(n_152),
.Y(n_525)
);

OR2x6_ASAP7_75t_L g526 ( 
.A(n_418),
.B(n_21),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_366),
.Y(n_527)
);

AO22x2_ASAP7_75t_L g528 ( 
.A1(n_408),
.A2(n_21),
.B1(n_22),
.B2(n_155),
.Y(n_528)
);

INVx1_ASAP7_75t_SL g529 ( 
.A(n_451),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_405),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_429),
.A2(n_182),
.B1(n_246),
.B2(n_242),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_476),
.B(n_151),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_373),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g534 ( 
.A(n_405),
.Y(n_534)
);

AO22x2_ASAP7_75t_L g535 ( 
.A1(n_412),
.A2(n_146),
.B1(n_233),
.B2(n_221),
.Y(n_535)
);

OAI22xp33_ASAP7_75t_L g536 ( 
.A1(n_392),
.A2(n_142),
.B1(n_219),
.B2(n_216),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_479),
.B(n_138),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_378),
.Y(n_538)
);

AO22x1_ASAP7_75t_L g539 ( 
.A1(n_369),
.A2(n_402),
.B1(n_392),
.B2(n_389),
.Y(n_539)
);

INVx8_ASAP7_75t_L g540 ( 
.A(n_456),
.Y(n_540)
);

OAI22xp33_ASAP7_75t_L g541 ( 
.A1(n_480),
.A2(n_141),
.B1(n_213),
.B2(n_212),
.Y(n_541)
);

AO22x2_ASAP7_75t_L g542 ( 
.A1(n_413),
.A2(n_264),
.B1(n_210),
.B2(n_209),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_368),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_425),
.Y(n_544)
);

OAI22xp33_ASAP7_75t_SL g545 ( 
.A1(n_382),
.A2(n_208),
.B1(n_198),
.B2(n_197),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_479),
.B(n_196),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_429),
.A2(n_190),
.B1(n_45),
.B2(n_60),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_436),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_481),
.Y(n_549)
);

AO22x2_ASAP7_75t_L g550 ( 
.A1(n_409),
.A2(n_402),
.B1(n_417),
.B2(n_484),
.Y(n_550)
);

OAI22xp33_ASAP7_75t_L g551 ( 
.A1(n_480),
.A2(n_32),
.B1(n_61),
.B2(n_63),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_481),
.B(n_71),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_385),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_484),
.B(n_74),
.Y(n_554)
);

OAI22xp33_ASAP7_75t_L g555 ( 
.A1(n_486),
.A2(n_80),
.B1(n_88),
.B2(n_95),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_L g556 ( 
.A1(n_485),
.A2(n_99),
.B1(n_462),
.B2(n_435),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_485),
.B(n_374),
.Y(n_557)
);

OR2x2_ASAP7_75t_L g558 ( 
.A(n_407),
.B(n_410),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_390),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_374),
.B(n_435),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_459),
.A2(n_391),
.B1(n_462),
.B2(n_393),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_459),
.B(n_391),
.Y(n_562)
);

INVx2_ASAP7_75t_SL g563 ( 
.A(n_474),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_395),
.A2(n_361),
.B1(n_488),
.B2(n_487),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_424),
.A2(n_431),
.B1(n_444),
.B2(n_483),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_389),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_427),
.Y(n_567)
);

OR2x6_ASAP7_75t_L g568 ( 
.A(n_411),
.B(n_477),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_367),
.B(n_461),
.Y(n_569)
);

OAI22xp33_ASAP7_75t_L g570 ( 
.A1(n_486),
.A2(n_492),
.B1(n_482),
.B2(n_475),
.Y(n_570)
);

NAND3x1_ASAP7_75t_L g571 ( 
.A(n_420),
.B(n_445),
.C(n_452),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_442),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_463),
.B(n_388),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_447),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_SL g575 ( 
.A1(n_383),
.A2(n_416),
.B1(n_414),
.B2(n_415),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_455),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_411),
.B(n_492),
.Y(n_577)
);

OR2x2_ASAP7_75t_L g578 ( 
.A(n_416),
.B(n_419),
.Y(n_578)
);

AO22x2_ASAP7_75t_L g579 ( 
.A1(n_466),
.A2(n_470),
.B1(n_471),
.B2(n_387),
.Y(n_579)
);

OAI22xp33_ASAP7_75t_SL g580 ( 
.A1(n_471),
.A2(n_381),
.B1(n_379),
.B2(n_387),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_411),
.B(n_468),
.Y(n_581)
);

NAND3x1_ASAP7_75t_L g582 ( 
.A(n_379),
.B(n_381),
.C(n_467),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_464),
.A2(n_473),
.B1(n_468),
.B2(n_369),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_384),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_464),
.B(n_473),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_434),
.B(n_457),
.Y(n_586)
);

AO22x2_ASAP7_75t_L g587 ( 
.A1(n_434),
.A2(n_440),
.B1(n_454),
.B2(n_457),
.Y(n_587)
);

AO22x2_ASAP7_75t_L g588 ( 
.A1(n_440),
.A2(n_454),
.B1(n_394),
.B2(n_377),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g589 ( 
.A1(n_369),
.A2(n_384),
.B1(n_472),
.B2(n_490),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g590 ( 
.A1(n_369),
.A2(n_472),
.B1(n_490),
.B2(n_439),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_375),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_421),
.B(n_428),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_377),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_421),
.B(n_428),
.Y(n_594)
);

OAI22xp33_ASAP7_75t_L g595 ( 
.A1(n_363),
.A2(n_365),
.B1(n_371),
.B2(n_426),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_371),
.Y(n_596)
);

AND2x2_ASAP7_75t_SL g597 ( 
.A(n_416),
.B(n_426),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_375),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_363),
.Y(n_599)
);

BUFx10_ASAP7_75t_L g600 ( 
.A(n_467),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_375),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_365),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_422),
.A2(n_423),
.B1(n_490),
.B2(n_438),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_422),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_422),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_423),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_423),
.B(n_446),
.Y(n_607)
);

OAI22xp33_ASAP7_75t_R g608 ( 
.A1(n_437),
.A2(n_443),
.B1(n_460),
.B2(n_441),
.Y(n_608)
);

OAI22xp33_ASAP7_75t_SL g609 ( 
.A1(n_489),
.A2(n_437),
.B1(n_443),
.B2(n_439),
.Y(n_609)
);

INVx1_ASAP7_75t_SL g610 ( 
.A(n_438),
.Y(n_610)
);

AO22x2_ASAP7_75t_L g611 ( 
.A1(n_438),
.A2(n_439),
.B1(n_441),
.B2(n_446),
.Y(n_611)
);

NAND2xp33_ASAP7_75t_SL g612 ( 
.A(n_441),
.B(n_446),
.Y(n_612)
);

AOI22xp5_ASAP7_75t_L g613 ( 
.A1(n_448),
.A2(n_450),
.B1(n_469),
.B2(n_489),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_448),
.A2(n_450),
.B1(n_469),
.B2(n_489),
.Y(n_614)
);

NAND3x1_ASAP7_75t_L g615 ( 
.A(n_448),
.B(n_450),
.C(n_469),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g616 ( 
.A1(n_489),
.A2(n_399),
.B1(n_317),
.B2(n_453),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_364),
.Y(n_617)
);

AO22x2_ASAP7_75t_L g618 ( 
.A1(n_401),
.A2(n_453),
.B1(n_398),
.B2(n_404),
.Y(n_618)
);

OAI22xp33_ASAP7_75t_R g619 ( 
.A1(n_376),
.A2(n_432),
.B1(n_354),
.B2(n_356),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_364),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_364),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_L g622 ( 
.A1(n_399),
.A2(n_317),
.B1(n_453),
.B2(n_398),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_SL g623 ( 
.A1(n_399),
.A2(n_292),
.B1(n_227),
.B2(n_348),
.Y(n_623)
);

OAI22xp33_ASAP7_75t_SL g624 ( 
.A1(n_401),
.A2(n_317),
.B1(n_404),
.B2(n_453),
.Y(n_624)
);

OAI22xp33_ASAP7_75t_SL g625 ( 
.A1(n_401),
.A2(n_317),
.B1(n_404),
.B2(n_453),
.Y(n_625)
);

OAI22xp5_ASAP7_75t_SL g626 ( 
.A1(n_399),
.A2(n_292),
.B1(n_227),
.B2(n_348),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_405),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_386),
.Y(n_628)
);

INVx2_ASAP7_75t_SL g629 ( 
.A(n_370),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_399),
.A2(n_317),
.B1(n_453),
.B2(n_398),
.Y(n_630)
);

AOI22xp5_ASAP7_75t_L g631 ( 
.A1(n_399),
.A2(n_317),
.B1(n_453),
.B2(n_398),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_433),
.B(n_465),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_386),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_386),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_399),
.A2(n_317),
.B1(n_453),
.B2(n_398),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_399),
.A2(n_317),
.B1(n_453),
.B2(n_398),
.Y(n_636)
);

INVx2_ASAP7_75t_L g637 ( 
.A(n_386),
.Y(n_637)
);

OAI22xp33_ASAP7_75t_SL g638 ( 
.A1(n_401),
.A2(n_317),
.B1(n_404),
.B2(n_453),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_L g639 ( 
.A1(n_399),
.A2(n_317),
.B1(n_453),
.B2(n_398),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_453),
.B(n_398),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_453),
.B(n_398),
.Y(n_641)
);

AOI22xp5_ASAP7_75t_L g642 ( 
.A1(n_399),
.A2(n_317),
.B1(n_453),
.B2(n_398),
.Y(n_642)
);

OR2x2_ASAP7_75t_L g643 ( 
.A(n_398),
.B(n_401),
.Y(n_643)
);

AO22x2_ASAP7_75t_L g644 ( 
.A1(n_401),
.A2(n_453),
.B1(n_398),
.B2(n_404),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_364),
.Y(n_645)
);

OAI22xp33_ASAP7_75t_SL g646 ( 
.A1(n_401),
.A2(n_317),
.B1(n_404),
.B2(n_453),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_433),
.B(n_465),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_364),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_398),
.B(n_453),
.Y(n_649)
);

OAI22xp33_ASAP7_75t_L g650 ( 
.A1(n_401),
.A2(n_453),
.B1(n_398),
.B2(n_317),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_386),
.Y(n_651)
);

INVx5_ASAP7_75t_L g652 ( 
.A(n_369),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_386),
.Y(n_653)
);

OA22x2_ASAP7_75t_L g654 ( 
.A1(n_401),
.A2(n_453),
.B1(n_398),
.B2(n_332),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_398),
.B(n_453),
.Y(n_655)
);

OR2x6_ASAP7_75t_L g656 ( 
.A(n_418),
.B(n_405),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_453),
.B(n_398),
.Y(n_657)
);

OA22x2_ASAP7_75t_L g658 ( 
.A1(n_401),
.A2(n_453),
.B1(n_398),
.B2(n_332),
.Y(n_658)
);

OAI22xp33_ASAP7_75t_L g659 ( 
.A1(n_401),
.A2(n_453),
.B1(n_398),
.B2(n_317),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_433),
.B(n_465),
.Y(n_660)
);

OAI22xp33_ASAP7_75t_R g661 ( 
.A1(n_376),
.A2(n_432),
.B1(n_286),
.B2(n_156),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_399),
.A2(n_317),
.B1(n_453),
.B2(n_398),
.Y(n_662)
);

OR2x6_ASAP7_75t_L g663 ( 
.A(n_418),
.B(n_405),
.Y(n_663)
);

AOI22xp5_ASAP7_75t_L g664 ( 
.A1(n_399),
.A2(n_317),
.B1(n_453),
.B2(n_398),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_386),
.Y(n_665)
);

INVx3_ASAP7_75t_L g666 ( 
.A(n_458),
.Y(n_666)
);

AO22x2_ASAP7_75t_L g667 ( 
.A1(n_401),
.A2(n_453),
.B1(n_398),
.B2(n_404),
.Y(n_667)
);

INVxp67_ASAP7_75t_SL g668 ( 
.A(n_375),
.Y(n_668)
);

AOI22xp5_ASAP7_75t_L g669 ( 
.A1(n_399),
.A2(n_317),
.B1(n_453),
.B2(n_398),
.Y(n_669)
);

OAI22xp33_ASAP7_75t_L g670 ( 
.A1(n_401),
.A2(n_453),
.B1(n_398),
.B2(n_317),
.Y(n_670)
);

BUFx3_ASAP7_75t_L g671 ( 
.A(n_458),
.Y(n_671)
);

OA22x2_ASAP7_75t_L g672 ( 
.A1(n_401),
.A2(n_453),
.B1(n_398),
.B2(n_332),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_L g673 ( 
.A1(n_399),
.A2(n_317),
.B1(n_453),
.B2(n_398),
.Y(n_673)
);

OAI22xp33_ASAP7_75t_SL g674 ( 
.A1(n_401),
.A2(n_317),
.B1(n_404),
.B2(n_453),
.Y(n_674)
);

OR2x2_ASAP7_75t_L g675 ( 
.A(n_398),
.B(n_401),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_386),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_386),
.Y(n_677)
);

AND2x4_ASAP7_75t_L g678 ( 
.A(n_458),
.B(n_474),
.Y(n_678)
);

OAI22xp33_ASAP7_75t_SL g679 ( 
.A1(n_401),
.A2(n_317),
.B1(n_404),
.B2(n_453),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_386),
.Y(n_680)
);

AO22x2_ASAP7_75t_L g681 ( 
.A1(n_401),
.A2(n_453),
.B1(n_398),
.B2(n_404),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_SL g682 ( 
.A(n_399),
.B(n_367),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_453),
.B(n_398),
.Y(n_683)
);

OAI22xp33_ASAP7_75t_SL g684 ( 
.A1(n_401),
.A2(n_317),
.B1(n_404),
.B2(n_453),
.Y(n_684)
);

OAI22xp33_ASAP7_75t_R g685 ( 
.A1(n_376),
.A2(n_432),
.B1(n_286),
.B2(n_156),
.Y(n_685)
);

AOI22xp5_ASAP7_75t_L g686 ( 
.A1(n_399),
.A2(n_317),
.B1(n_453),
.B2(n_398),
.Y(n_686)
);

AOI22xp5_ASAP7_75t_L g687 ( 
.A1(n_399),
.A2(n_317),
.B1(n_453),
.B2(n_398),
.Y(n_687)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_399),
.A2(n_317),
.B1(n_453),
.B2(n_398),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_364),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_453),
.B(n_398),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_386),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_386),
.Y(n_692)
);

OAI22xp33_ASAP7_75t_L g693 ( 
.A1(n_401),
.A2(n_453),
.B1(n_398),
.B2(n_317),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_398),
.B(n_453),
.Y(n_694)
);

AOI22xp5_ASAP7_75t_L g695 ( 
.A1(n_399),
.A2(n_317),
.B1(n_453),
.B2(n_398),
.Y(n_695)
);

OAI22xp33_ASAP7_75t_SL g696 ( 
.A1(n_401),
.A2(n_317),
.B1(n_404),
.B2(n_453),
.Y(n_696)
);

OAI22xp33_ASAP7_75t_SL g697 ( 
.A1(n_401),
.A2(n_317),
.B1(n_404),
.B2(n_453),
.Y(n_697)
);

OR2x2_ASAP7_75t_L g698 ( 
.A(n_398),
.B(n_401),
.Y(n_698)
);

OA22x2_ASAP7_75t_L g699 ( 
.A1(n_401),
.A2(n_453),
.B1(n_398),
.B2(n_332),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_386),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_386),
.Y(n_701)
);

OAI22xp5_ASAP7_75t_SL g702 ( 
.A1(n_399),
.A2(n_292),
.B1(n_227),
.B2(n_348),
.Y(n_702)
);

AO22x2_ASAP7_75t_L g703 ( 
.A1(n_401),
.A2(n_453),
.B1(n_398),
.B2(n_404),
.Y(n_703)
);

AO22x2_ASAP7_75t_L g704 ( 
.A1(n_401),
.A2(n_453),
.B1(n_398),
.B2(n_404),
.Y(n_704)
);

OAI22xp33_ASAP7_75t_L g705 ( 
.A1(n_401),
.A2(n_453),
.B1(n_398),
.B2(n_317),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_386),
.Y(n_706)
);

AOI22xp5_ASAP7_75t_L g707 ( 
.A1(n_399),
.A2(n_317),
.B1(n_453),
.B2(n_398),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_458),
.Y(n_708)
);

OAI22xp33_ASAP7_75t_L g709 ( 
.A1(n_401),
.A2(n_453),
.B1(n_398),
.B2(n_317),
.Y(n_709)
);

OAI22xp5_ASAP7_75t_SL g710 ( 
.A1(n_399),
.A2(n_292),
.B1(n_227),
.B2(n_348),
.Y(n_710)
);

AOI22xp5_ASAP7_75t_L g711 ( 
.A1(n_399),
.A2(n_317),
.B1(n_453),
.B2(n_398),
.Y(n_711)
);

OAI22xp5_ASAP7_75t_L g712 ( 
.A1(n_398),
.A2(n_453),
.B1(n_401),
.B2(n_433),
.Y(n_712)
);

AOI22xp5_ASAP7_75t_L g713 ( 
.A1(n_399),
.A2(n_317),
.B1(n_453),
.B2(n_398),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_386),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_398),
.B(n_453),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_453),
.B(n_398),
.Y(n_716)
);

OR2x6_ASAP7_75t_L g717 ( 
.A(n_418),
.B(n_405),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_386),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_386),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_399),
.A2(n_317),
.B1(n_453),
.B2(n_398),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_399),
.A2(n_317),
.B1(n_453),
.B2(n_398),
.Y(n_721)
);

OAI22xp33_ASAP7_75t_L g722 ( 
.A1(n_401),
.A2(n_453),
.B1(n_398),
.B2(n_317),
.Y(n_722)
);

OA22x2_ASAP7_75t_L g723 ( 
.A1(n_401),
.A2(n_453),
.B1(n_398),
.B2(n_332),
.Y(n_723)
);

BUFx10_ASAP7_75t_L g724 ( 
.A(n_376),
.Y(n_724)
);

OR2x6_ASAP7_75t_L g725 ( 
.A(n_418),
.B(n_405),
.Y(n_725)
);

AOI22xp5_ASAP7_75t_L g726 ( 
.A1(n_399),
.A2(n_317),
.B1(n_453),
.B2(n_398),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_364),
.Y(n_727)
);

AOI22xp5_ASAP7_75t_L g728 ( 
.A1(n_399),
.A2(n_317),
.B1(n_453),
.B2(n_398),
.Y(n_728)
);

AOI22xp5_ASAP7_75t_L g729 ( 
.A1(n_399),
.A2(n_317),
.B1(n_453),
.B2(n_398),
.Y(n_729)
);

OAI22xp33_ASAP7_75t_L g730 ( 
.A1(n_401),
.A2(n_453),
.B1(n_398),
.B2(n_317),
.Y(n_730)
);

AOI22xp5_ASAP7_75t_L g731 ( 
.A1(n_399),
.A2(n_317),
.B1(n_453),
.B2(n_398),
.Y(n_731)
);

OAI22xp5_ASAP7_75t_SL g732 ( 
.A1(n_399),
.A2(n_292),
.B1(n_227),
.B2(n_348),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_364),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_433),
.B(n_465),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_398),
.B(n_453),
.Y(n_735)
);

AO22x2_ASAP7_75t_L g736 ( 
.A1(n_401),
.A2(n_453),
.B1(n_398),
.B2(n_404),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_364),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_433),
.B(n_465),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_386),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_367),
.Y(n_740)
);

AOI22xp5_ASAP7_75t_L g741 ( 
.A1(n_399),
.A2(n_317),
.B1(n_453),
.B2(n_398),
.Y(n_741)
);

OA22x2_ASAP7_75t_L g742 ( 
.A1(n_401),
.A2(n_453),
.B1(n_398),
.B2(n_332),
.Y(n_742)
);

AO22x2_ASAP7_75t_L g743 ( 
.A1(n_401),
.A2(n_453),
.B1(n_398),
.B2(n_404),
.Y(n_743)
);

AO22x2_ASAP7_75t_L g744 ( 
.A1(n_401),
.A2(n_453),
.B1(n_398),
.B2(n_404),
.Y(n_744)
);

AO22x2_ASAP7_75t_L g745 ( 
.A1(n_401),
.A2(n_453),
.B1(n_398),
.B2(n_404),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_399),
.A2(n_317),
.B1(n_453),
.B2(n_398),
.Y(n_746)
);

OAI22xp33_ASAP7_75t_L g747 ( 
.A1(n_401),
.A2(n_453),
.B1(n_398),
.B2(n_317),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_398),
.B(n_453),
.Y(n_748)
);

OAI22xp33_ASAP7_75t_L g749 ( 
.A1(n_401),
.A2(n_453),
.B1(n_398),
.B2(n_317),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_364),
.Y(n_750)
);

OR2x6_ASAP7_75t_L g751 ( 
.A(n_418),
.B(n_405),
.Y(n_751)
);

AO22x2_ASAP7_75t_L g752 ( 
.A1(n_401),
.A2(n_453),
.B1(n_398),
.B2(n_404),
.Y(n_752)
);

OR2x6_ASAP7_75t_L g753 ( 
.A(n_418),
.B(n_405),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_398),
.B(n_453),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_398),
.B(n_453),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_398),
.B(n_453),
.Y(n_756)
);

OAI22xp33_ASAP7_75t_SL g757 ( 
.A1(n_401),
.A2(n_317),
.B1(n_404),
.B2(n_453),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_399),
.A2(n_317),
.B1(n_453),
.B2(n_398),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_364),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_386),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_386),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_398),
.B(n_453),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_364),
.Y(n_763)
);

OAI22xp33_ASAP7_75t_L g764 ( 
.A1(n_401),
.A2(n_453),
.B1(n_398),
.B2(n_317),
.Y(n_764)
);

AO22x2_ASAP7_75t_L g765 ( 
.A1(n_401),
.A2(n_453),
.B1(n_398),
.B2(n_404),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_386),
.Y(n_766)
);

OAI22xp5_ASAP7_75t_L g767 ( 
.A1(n_398),
.A2(n_453),
.B1(n_401),
.B2(n_433),
.Y(n_767)
);

OAI22xp33_ASAP7_75t_L g768 ( 
.A1(n_401),
.A2(n_453),
.B1(n_398),
.B2(n_317),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_398),
.B(n_453),
.Y(n_769)
);

AOI22xp5_ASAP7_75t_L g770 ( 
.A1(n_399),
.A2(n_317),
.B1(n_453),
.B2(n_398),
.Y(n_770)
);

INVx1_ASAP7_75t_SL g771 ( 
.A(n_430),
.Y(n_771)
);

OAI22xp33_ASAP7_75t_SL g772 ( 
.A1(n_401),
.A2(n_317),
.B1(n_404),
.B2(n_453),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_399),
.A2(n_317),
.B1(n_453),
.B2(n_398),
.Y(n_773)
);

AOI22x1_ASAP7_75t_L g774 ( 
.A1(n_433),
.A2(n_491),
.B1(n_465),
.B2(n_398),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_399),
.A2(n_317),
.B1(n_453),
.B2(n_398),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_386),
.Y(n_776)
);

OAI22xp33_ASAP7_75t_L g777 ( 
.A1(n_401),
.A2(n_453),
.B1(n_398),
.B2(n_317),
.Y(n_777)
);

OAI22xp5_ASAP7_75t_SL g778 ( 
.A1(n_399),
.A2(n_292),
.B1(n_227),
.B2(n_348),
.Y(n_778)
);

OAI22xp33_ASAP7_75t_L g779 ( 
.A1(n_401),
.A2(n_453),
.B1(n_398),
.B2(n_317),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_364),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_364),
.Y(n_781)
);

OAI22xp5_ASAP7_75t_SL g782 ( 
.A1(n_399),
.A2(n_292),
.B1(n_227),
.B2(n_348),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_399),
.A2(n_317),
.B1(n_453),
.B2(n_398),
.Y(n_783)
);

OAI22xp33_ASAP7_75t_L g784 ( 
.A1(n_401),
.A2(n_453),
.B1(n_398),
.B2(n_317),
.Y(n_784)
);

OAI22xp33_ASAP7_75t_L g785 ( 
.A1(n_401),
.A2(n_453),
.B1(n_398),
.B2(n_317),
.Y(n_785)
);

INVx3_ASAP7_75t_L g786 ( 
.A(n_458),
.Y(n_786)
);

AND2x2_ASAP7_75t_SL g787 ( 
.A(n_399),
.B(n_374),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_386),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_386),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_398),
.B(n_453),
.Y(n_790)
);

OAI22xp33_ASAP7_75t_R g791 ( 
.A1(n_376),
.A2(n_432),
.B1(n_354),
.B2(n_356),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_386),
.Y(n_792)
);

OAI22xp5_ASAP7_75t_SL g793 ( 
.A1(n_399),
.A2(n_292),
.B1(n_227),
.B2(n_348),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_386),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_398),
.B(n_453),
.Y(n_795)
);

AOI22xp5_ASAP7_75t_L g796 ( 
.A1(n_399),
.A2(n_317),
.B1(n_453),
.B2(n_398),
.Y(n_796)
);

AOI22xp5_ASAP7_75t_L g797 ( 
.A1(n_399),
.A2(n_317),
.B1(n_453),
.B2(n_398),
.Y(n_797)
);

OA22x2_ASAP7_75t_L g798 ( 
.A1(n_401),
.A2(n_453),
.B1(n_398),
.B2(n_332),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_504),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_517),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_508),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_500),
.B(n_624),
.Y(n_802)
);

AND2x6_ASAP7_75t_L g803 ( 
.A(n_585),
.B(n_592),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_533),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_586),
.B(n_599),
.Y(n_805)
);

BUFx6f_ASAP7_75t_L g806 ( 
.A(n_530),
.Y(n_806)
);

OAI22xp33_ASAP7_75t_L g807 ( 
.A1(n_643),
.A2(n_698),
.B1(n_675),
.B2(n_622),
.Y(n_807)
);

INVx3_ASAP7_75t_L g808 ( 
.A(n_591),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_538),
.Y(n_809)
);

AND2x2_ASAP7_75t_SL g810 ( 
.A(n_787),
.B(n_682),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_553),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_559),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_567),
.Y(n_813)
);

HB1xp67_ASAP7_75t_SL g814 ( 
.A(n_740),
.Y(n_814)
);

INVx5_ASAP7_75t_L g815 ( 
.A(n_652),
.Y(n_815)
);

INVx3_ASAP7_75t_L g816 ( 
.A(n_598),
.Y(n_816)
);

CKINVDCx20_ASAP7_75t_R g817 ( 
.A(n_623),
.Y(n_817)
);

BUFx6f_ASAP7_75t_SL g818 ( 
.A(n_600),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_602),
.B(n_640),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_625),
.B(n_638),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_601),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_617),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_620),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_641),
.B(n_657),
.Y(n_824)
);

NAND2xp33_ASAP7_75t_SL g825 ( 
.A(n_552),
.B(n_554),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_683),
.B(n_690),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_649),
.B(n_655),
.Y(n_827)
);

INVx1_ASAP7_75t_SL g828 ( 
.A(n_694),
.Y(n_828)
);

CKINVDCx6p67_ASAP7_75t_R g829 ( 
.A(n_502),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_584),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_621),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_716),
.B(n_650),
.Y(n_832)
);

INVx3_ASAP7_75t_L g833 ( 
.A(n_604),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_645),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_648),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_659),
.B(n_670),
.Y(n_836)
);

OR2x2_ASAP7_75t_L g837 ( 
.A(n_632),
.B(n_647),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_605),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_689),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_727),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_596),
.B(n_593),
.Y(n_841)
);

BUFx6f_ASAP7_75t_SL g842 ( 
.A(n_568),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_530),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_733),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_737),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_715),
.B(n_735),
.Y(n_846)
);

BUFx10_ASAP7_75t_L g847 ( 
.A(n_573),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_748),
.B(n_754),
.Y(n_848)
);

BUFx6f_ASAP7_75t_L g849 ( 
.A(n_534),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_750),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_755),
.B(n_756),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_762),
.B(n_769),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_759),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_763),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_780),
.Y(n_855)
);

BUFx6f_ASAP7_75t_L g856 ( 
.A(n_534),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_607),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_781),
.Y(n_858)
);

AOI22xp5_ASAP7_75t_L g859 ( 
.A1(n_619),
.A2(n_791),
.B1(n_597),
.B2(n_577),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_693),
.B(n_705),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_790),
.B(n_795),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_611),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_569),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_499),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_709),
.B(n_722),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_570),
.B(n_712),
.Y(n_866)
);

INVx2_ASAP7_75t_SL g867 ( 
.A(n_627),
.Y(n_867)
);

AOI22xp33_ASAP7_75t_L g868 ( 
.A1(n_661),
.A2(n_685),
.B1(n_494),
.B2(n_644),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_611),
.Y(n_869)
);

OAI21xp33_ASAP7_75t_SL g870 ( 
.A1(n_561),
.A2(n_520),
.B(n_654),
.Y(n_870)
);

BUFx6f_ASAP7_75t_L g871 ( 
.A(n_627),
.Y(n_871)
);

INVxp33_ASAP7_75t_SL g872 ( 
.A(n_630),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_628),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_767),
.B(n_503),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_633),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_634),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_660),
.B(n_734),
.Y(n_877)
);

BUFx6f_ASAP7_75t_L g878 ( 
.A(n_678),
.Y(n_878)
);

INVx2_ASAP7_75t_L g879 ( 
.A(n_637),
.Y(n_879)
);

BUFx4f_ASAP7_75t_L g880 ( 
.A(n_540),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_738),
.B(n_516),
.Y(n_881)
);

AOI22xp33_ASAP7_75t_L g882 ( 
.A1(n_661),
.A2(n_685),
.B1(n_494),
.B2(n_644),
.Y(n_882)
);

INVx2_ASAP7_75t_SL g883 ( 
.A(n_578),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_651),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_653),
.Y(n_885)
);

AOI22xp33_ASAP7_75t_SL g886 ( 
.A1(n_626),
.A2(n_732),
.B1(n_793),
.B2(n_702),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_665),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_730),
.B(n_747),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_646),
.B(n_674),
.Y(n_889)
);

BUFx2_ASAP7_75t_L g890 ( 
.A(n_568),
.Y(n_890)
);

AND2x6_ASAP7_75t_L g891 ( 
.A(n_594),
.B(n_583),
.Y(n_891)
);

AOI22xp33_ASAP7_75t_L g892 ( 
.A1(n_618),
.A2(n_744),
.B1(n_745),
.B2(n_743),
.Y(n_892)
);

AND2x2_ASAP7_75t_L g893 ( 
.A(n_506),
.B(n_771),
.Y(n_893)
);

AND2x6_ASAP7_75t_L g894 ( 
.A(n_581),
.B(n_562),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_676),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_749),
.B(n_764),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_677),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_680),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_691),
.Y(n_899)
);

AOI22xp33_ASAP7_75t_L g900 ( 
.A1(n_618),
.A2(n_743),
.B1(n_667),
.B2(n_681),
.Y(n_900)
);

INVx6_ASAP7_75t_L g901 ( 
.A(n_656),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_692),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_667),
.B(n_681),
.Y(n_903)
);

INVx3_ASAP7_75t_L g904 ( 
.A(n_527),
.Y(n_904)
);

CKINVDCx20_ASAP7_75t_R g905 ( 
.A(n_710),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_768),
.B(n_777),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_700),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_543),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_779),
.B(n_784),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_701),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_703),
.B(n_704),
.Y(n_911)
);

BUFx2_ASAP7_75t_L g912 ( 
.A(n_558),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_706),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_714),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_785),
.B(n_631),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_635),
.B(n_636),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_718),
.Y(n_917)
);

INVx2_ASAP7_75t_SL g918 ( 
.A(n_512),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_703),
.B(n_704),
.Y(n_919)
);

INVx3_ASAP7_75t_L g920 ( 
.A(n_544),
.Y(n_920)
);

BUFx6f_ASAP7_75t_SL g921 ( 
.A(n_656),
.Y(n_921)
);

INVx5_ASAP7_75t_L g922 ( 
.A(n_652),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_679),
.B(n_684),
.Y(n_923)
);

INVx4_ASAP7_75t_L g924 ( 
.A(n_678),
.Y(n_924)
);

BUFx10_ASAP7_75t_L g925 ( 
.A(n_663),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_736),
.B(n_744),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_719),
.Y(n_927)
);

AOI22xp33_ASAP7_75t_L g928 ( 
.A1(n_736),
.A2(n_765),
.B1(n_752),
.B2(n_745),
.Y(n_928)
);

CKINVDCx6p67_ASAP7_75t_R g929 ( 
.A(n_540),
.Y(n_929)
);

AOI22xp33_ASAP7_75t_L g930 ( 
.A1(n_752),
.A2(n_765),
.B1(n_509),
.B2(n_528),
.Y(n_930)
);

INVx2_ASAP7_75t_SL g931 ( 
.A(n_658),
.Y(n_931)
);

BUFx3_ASAP7_75t_L g932 ( 
.A(n_513),
.Y(n_932)
);

AOI22xp33_ASAP7_75t_L g933 ( 
.A1(n_509),
.A2(n_528),
.B1(n_588),
.B2(n_493),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_739),
.Y(n_934)
);

INVx2_ASAP7_75t_SL g935 ( 
.A(n_672),
.Y(n_935)
);

OAI21xp33_ASAP7_75t_L g936 ( 
.A1(n_639),
.A2(n_728),
.B(n_797),
.Y(n_936)
);

BUFx6f_ASAP7_75t_L g937 ( 
.A(n_652),
.Y(n_937)
);

INVx2_ASAP7_75t_SL g938 ( 
.A(n_699),
.Y(n_938)
);

OR2x2_ASAP7_75t_L g939 ( 
.A(n_529),
.B(n_642),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_760),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_SL g941 ( 
.A(n_696),
.B(n_697),
.Y(n_941)
);

BUFx3_ASAP7_75t_L g942 ( 
.A(n_671),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_757),
.B(n_772),
.Y(n_943)
);

AOI22xp33_ASAP7_75t_L g944 ( 
.A1(n_588),
.A2(n_493),
.B1(n_587),
.B2(n_556),
.Y(n_944)
);

INVx2_ASAP7_75t_SL g945 ( 
.A(n_723),
.Y(n_945)
);

BUFx3_ASAP7_75t_L g946 ( 
.A(n_663),
.Y(n_946)
);

AOI22xp33_ASAP7_75t_L g947 ( 
.A1(n_587),
.A2(n_501),
.B1(n_579),
.B2(n_555),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_761),
.Y(n_948)
);

BUFx3_ASAP7_75t_L g949 ( 
.A(n_717),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_518),
.B(n_522),
.Y(n_950)
);

INVx3_ASAP7_75t_L g951 ( 
.A(n_548),
.Y(n_951)
);

INVx3_ASAP7_75t_L g952 ( 
.A(n_572),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_766),
.Y(n_953)
);

AND2x6_ASAP7_75t_L g954 ( 
.A(n_560),
.B(n_557),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_776),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_510),
.B(n_580),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_788),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_515),
.B(n_629),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_789),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_792),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_662),
.B(n_664),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_669),
.B(n_673),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_794),
.Y(n_963)
);

INVx3_ASAP7_75t_L g964 ( 
.A(n_576),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_774),
.B(n_539),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_574),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_606),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_610),
.Y(n_968)
);

NAND3xp33_ASAP7_75t_L g969 ( 
.A(n_686),
.B(n_720),
.C(n_796),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_666),
.Y(n_970)
);

OR2x6_ASAP7_75t_L g971 ( 
.A(n_717),
.B(n_725),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_564),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_708),
.Y(n_973)
);

OAI21xp33_ASAP7_75t_SL g974 ( 
.A1(n_742),
.A2(n_798),
.B(n_565),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_539),
.B(n_579),
.Y(n_975)
);

INVx5_ASAP7_75t_L g976 ( 
.A(n_725),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_566),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_786),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_603),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_549),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_616),
.B(n_783),
.Y(n_981)
);

OR2x2_ASAP7_75t_L g982 ( 
.A(n_687),
.B(n_688),
.Y(n_982)
);

NAND2xp33_ASAP7_75t_L g983 ( 
.A(n_615),
.B(n_547),
.Y(n_983)
);

INVx4_ASAP7_75t_L g984 ( 
.A(n_751),
.Y(n_984)
);

INVx5_ASAP7_75t_L g985 ( 
.A(n_751),
.Y(n_985)
);

INVx3_ASAP7_75t_L g986 ( 
.A(n_563),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_550),
.Y(n_987)
);

NOR2xp33_ASAP7_75t_L g988 ( 
.A(n_695),
.B(n_741),
.Y(n_988)
);

BUFx6f_ASAP7_75t_L g989 ( 
.A(n_753),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_550),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_589),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_707),
.B(n_711),
.Y(n_992)
);

INVx4_ASAP7_75t_L g993 ( 
.A(n_753),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_713),
.B(n_729),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_613),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_614),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_668),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_721),
.B(n_726),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_731),
.B(n_770),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_590),
.Y(n_1000)
);

AOI22xp33_ASAP7_75t_SL g1001 ( 
.A1(n_778),
.A2(n_782),
.B1(n_505),
.B2(n_496),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_525),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_532),
.Y(n_1003)
);

BUFx4f_ASAP7_75t_L g1004 ( 
.A(n_526),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_537),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_546),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_571),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_746),
.B(n_773),
.Y(n_1008)
);

BUFx6f_ASAP7_75t_L g1009 ( 
.A(n_724),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_612),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_SL g1011 ( 
.A(n_758),
.B(n_775),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_526),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_523),
.Y(n_1013)
);

INVxp67_ASAP7_75t_SL g1014 ( 
.A(n_595),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_535),
.Y(n_1015)
);

OAI22xp33_ASAP7_75t_L g1016 ( 
.A1(n_497),
.A2(n_551),
.B1(n_531),
.B2(n_521),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_535),
.Y(n_1017)
);

BUFx3_ASAP7_75t_L g1018 ( 
.A(n_575),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_542),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_542),
.Y(n_1020)
);

AND2x6_ASAP7_75t_L g1021 ( 
.A(n_608),
.B(n_511),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_582),
.Y(n_1022)
);

NAND2xp33_ASAP7_75t_R g1023 ( 
.A(n_495),
.B(n_498),
.Y(n_1023)
);

INVx2_ASAP7_75t_SL g1024 ( 
.A(n_524),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_505),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_519),
.Y(n_1026)
);

INVx1_ASAP7_75t_SL g1027 ( 
.A(n_545),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_514),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_536),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_541),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_507),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_609),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_586),
.B(n_599),
.Y(n_1033)
);

AOI22xp33_ASAP7_75t_L g1034 ( 
.A1(n_661),
.A2(n_685),
.B1(n_399),
.B2(n_596),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_500),
.B(n_624),
.Y(n_1035)
);

INVx3_ASAP7_75t_L g1036 ( 
.A(n_591),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_500),
.B(n_624),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_504),
.Y(n_1038)
);

BUFx3_ASAP7_75t_L g1039 ( 
.A(n_530),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_504),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_586),
.B(n_599),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_586),
.B(n_599),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_504),
.Y(n_1043)
);

BUFx10_ASAP7_75t_L g1044 ( 
.A(n_502),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_504),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_504),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_504),
.Y(n_1047)
);

NOR2x1p5_ASAP7_75t_L g1048 ( 
.A(n_530),
.B(n_456),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_504),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_586),
.B(n_599),
.Y(n_1050)
);

INVx4_ASAP7_75t_L g1051 ( 
.A(n_530),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_504),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_586),
.B(n_599),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_530),
.Y(n_1054)
);

NAND2xp33_ASAP7_75t_SL g1055 ( 
.A(n_552),
.B(n_554),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_500),
.B(n_624),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_504),
.Y(n_1057)
);

INVx5_ASAP7_75t_L g1058 ( 
.A(n_652),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_649),
.B(n_655),
.Y(n_1059)
);

INVx3_ASAP7_75t_L g1060 ( 
.A(n_591),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_504),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_SL g1062 ( 
.A(n_740),
.B(n_367),
.Y(n_1062)
);

AOI22xp33_ASAP7_75t_L g1063 ( 
.A1(n_661),
.A2(n_685),
.B1(n_399),
.B2(n_596),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_586),
.B(n_599),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_508),
.Y(n_1065)
);

INVx3_ASAP7_75t_L g1066 ( 
.A(n_591),
.Y(n_1066)
);

CKINVDCx6p67_ASAP7_75t_R g1067 ( 
.A(n_502),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_504),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_504),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_504),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_500),
.B(n_624),
.Y(n_1071)
);

INVx3_ASAP7_75t_L g1072 ( 
.A(n_591),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_504),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_504),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_640),
.B(n_641),
.Y(n_1075)
);

INVxp67_ASAP7_75t_SL g1076 ( 
.A(n_611),
.Y(n_1076)
);

INVx3_ASAP7_75t_L g1077 ( 
.A(n_591),
.Y(n_1077)
);

AOI22xp33_ASAP7_75t_L g1078 ( 
.A1(n_661),
.A2(n_685),
.B1(n_399),
.B2(n_596),
.Y(n_1078)
);

BUFx3_ASAP7_75t_L g1079 ( 
.A(n_530),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_740),
.Y(n_1080)
);

BUFx2_ASAP7_75t_L g1081 ( 
.A(n_568),
.Y(n_1081)
);

AOI22xp33_ASAP7_75t_L g1082 ( 
.A1(n_661),
.A2(n_685),
.B1(n_399),
.B2(n_596),
.Y(n_1082)
);

BUFx3_ASAP7_75t_L g1083 ( 
.A(n_530),
.Y(n_1083)
);

NOR2x1p5_ASAP7_75t_L g1084 ( 
.A(n_530),
.B(n_456),
.Y(n_1084)
);

INVx2_ASAP7_75t_L g1085 ( 
.A(n_504),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_504),
.Y(n_1086)
);

BUFx10_ASAP7_75t_L g1087 ( 
.A(n_502),
.Y(n_1087)
);

OAI22xp33_ASAP7_75t_L g1088 ( 
.A1(n_643),
.A2(n_698),
.B1(n_675),
.B2(n_796),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_504),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_504),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_504),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_504),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_504),
.Y(n_1093)
);

CKINVDCx6p67_ASAP7_75t_R g1094 ( 
.A(n_502),
.Y(n_1094)
);

INVx3_ASAP7_75t_L g1095 ( 
.A(n_591),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_504),
.Y(n_1096)
);

INVx4_ASAP7_75t_L g1097 ( 
.A(n_530),
.Y(n_1097)
);

BUFx10_ASAP7_75t_L g1098 ( 
.A(n_502),
.Y(n_1098)
);

INVx3_ASAP7_75t_L g1099 ( 
.A(n_591),
.Y(n_1099)
);

OR2x2_ASAP7_75t_L g1100 ( 
.A(n_643),
.B(n_675),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_530),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_586),
.B(n_599),
.Y(n_1102)
);

BUFx4f_ASAP7_75t_L g1103 ( 
.A(n_530),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_504),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_586),
.B(n_599),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_504),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_500),
.B(n_624),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_586),
.B(n_599),
.Y(n_1108)
);

OAI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_643),
.A2(n_698),
.B1(n_675),
.B2(n_796),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_504),
.Y(n_1110)
);

NAND3xp33_ASAP7_75t_L g1111 ( 
.A(n_503),
.B(n_432),
.C(n_376),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_504),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_L g1113 ( 
.A(n_530),
.Y(n_1113)
);

AOI22xp33_ASAP7_75t_L g1114 ( 
.A1(n_661),
.A2(n_685),
.B1(n_399),
.B2(n_596),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_504),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_504),
.Y(n_1116)
);

INVx5_ASAP7_75t_L g1117 ( 
.A(n_652),
.Y(n_1117)
);

NOR3xp33_ASAP7_75t_L g1118 ( 
.A(n_650),
.B(n_432),
.C(n_376),
.Y(n_1118)
);

INVx3_ASAP7_75t_L g1119 ( 
.A(n_591),
.Y(n_1119)
);

INVx2_ASAP7_75t_SL g1120 ( 
.A(n_530),
.Y(n_1120)
);

INVxp33_ASAP7_75t_SL g1121 ( 
.A(n_740),
.Y(n_1121)
);

AO22x2_ASAP7_75t_L g1122 ( 
.A1(n_661),
.A2(n_685),
.B1(n_556),
.B2(n_401),
.Y(n_1122)
);

INVx3_ASAP7_75t_L g1123 ( 
.A(n_591),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_504),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_504),
.Y(n_1125)
);

OR2x2_ASAP7_75t_L g1126 ( 
.A(n_643),
.B(n_675),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_SL g1127 ( 
.A(n_500),
.B(n_624),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_504),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_504),
.Y(n_1129)
);

NAND2xp33_ASAP7_75t_L g1130 ( 
.A(n_593),
.B(n_615),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_504),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_640),
.B(n_641),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_504),
.Y(n_1133)
);

AOI22xp33_ASAP7_75t_L g1134 ( 
.A1(n_661),
.A2(n_685),
.B1(n_399),
.B2(n_596),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_586),
.B(n_599),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_586),
.B(n_599),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_504),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_504),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_504),
.Y(n_1139)
);

OR2x2_ASAP7_75t_L g1140 ( 
.A(n_643),
.B(n_675),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_504),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_504),
.Y(n_1142)
);

AND2x4_ASAP7_75t_L g1143 ( 
.A(n_678),
.B(n_515),
.Y(n_1143)
);

NOR2xp33_ASAP7_75t_L g1144 ( 
.A(n_640),
.B(n_641),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_640),
.B(n_641),
.Y(n_1145)
);

BUFx3_ASAP7_75t_L g1146 ( 
.A(n_530),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_508),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_504),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_504),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_586),
.B(n_599),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_586),
.B(n_599),
.Y(n_1151)
);

BUFx3_ASAP7_75t_L g1152 ( 
.A(n_530),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_508),
.Y(n_1153)
);

AOI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_619),
.A2(n_791),
.B1(n_597),
.B2(n_577),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_504),
.Y(n_1155)
);

INVx3_ASAP7_75t_L g1156 ( 
.A(n_591),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_L g1157 ( 
.A(n_640),
.B(n_641),
.Y(n_1157)
);

BUFx3_ASAP7_75t_L g1158 ( 
.A(n_530),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_504),
.Y(n_1159)
);

CKINVDCx16_ASAP7_75t_R g1160 ( 
.A(n_502),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_504),
.Y(n_1161)
);

INVx2_ASAP7_75t_SL g1162 ( 
.A(n_530),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_500),
.B(n_624),
.Y(n_1163)
);

INVx1_ASAP7_75t_SL g1164 ( 
.A(n_649),
.Y(n_1164)
);

INVx4_ASAP7_75t_L g1165 ( 
.A(n_530),
.Y(n_1165)
);

AOI22xp33_ASAP7_75t_L g1166 ( 
.A1(n_661),
.A2(n_685),
.B1(n_399),
.B2(n_596),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_640),
.B(n_641),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_586),
.B(n_599),
.Y(n_1168)
);

OR2x6_ASAP7_75t_L g1169 ( 
.A(n_540),
.B(n_568),
.Y(n_1169)
);

OAI22xp33_ASAP7_75t_L g1170 ( 
.A1(n_643),
.A2(n_698),
.B1(n_675),
.B2(n_796),
.Y(n_1170)
);

INVx1_ASAP7_75t_SL g1171 ( 
.A(n_649),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_586),
.B(n_599),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_649),
.B(n_655),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_508),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_586),
.B(n_599),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_504),
.Y(n_1176)
);

NAND2xp33_ASAP7_75t_L g1177 ( 
.A(n_593),
.B(n_615),
.Y(n_1177)
);

AOI22xp33_ASAP7_75t_L g1178 ( 
.A1(n_661),
.A2(n_685),
.B1(n_399),
.B2(n_596),
.Y(n_1178)
);

INVx6_ASAP7_75t_L g1179 ( 
.A(n_530),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_500),
.B(n_624),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_500),
.B(n_624),
.Y(n_1181)
);

OR2x6_ASAP7_75t_L g1182 ( 
.A(n_540),
.B(n_568),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_504),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_649),
.B(n_655),
.Y(n_1184)
);

INVx1_ASAP7_75t_SL g1185 ( 
.A(n_649),
.Y(n_1185)
);

HB1xp67_ASAP7_75t_L g1186 ( 
.A(n_530),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_649),
.B(n_655),
.Y(n_1187)
);

INVx4_ASAP7_75t_L g1188 ( 
.A(n_530),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_504),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_504),
.Y(n_1190)
);

OAI22xp33_ASAP7_75t_L g1191 ( 
.A1(n_643),
.A2(n_698),
.B1(n_675),
.B2(n_796),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_649),
.B(n_655),
.Y(n_1192)
);

BUFx2_ASAP7_75t_L g1193 ( 
.A(n_568),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_504),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_504),
.Y(n_1195)
);

BUFx2_ASAP7_75t_L g1196 ( 
.A(n_568),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_504),
.Y(n_1197)
);

INVxp67_ASAP7_75t_L g1198 ( 
.A(n_649),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_504),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_504),
.Y(n_1200)
);

INVx3_ASAP7_75t_L g1201 ( 
.A(n_591),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_504),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_586),
.B(n_599),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_L g1204 ( 
.A(n_640),
.B(n_641),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_504),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_508),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_504),
.Y(n_1207)
);

NOR2xp33_ASAP7_75t_L g1208 ( 
.A(n_640),
.B(n_641),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_508),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_740),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_586),
.B(n_599),
.Y(n_1211)
);

AND2x6_ASAP7_75t_L g1212 ( 
.A(n_585),
.B(n_592),
.Y(n_1212)
);

BUFx2_ASAP7_75t_L g1213 ( 
.A(n_912),
.Y(n_1213)
);

INVx2_ASAP7_75t_SL g1214 ( 
.A(n_1103),
.Y(n_1214)
);

HB1xp67_ASAP7_75t_L g1215 ( 
.A(n_827),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1075),
.A2(n_1144),
.B1(n_1145),
.B2(n_1132),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_801),
.Y(n_1217)
);

AND2x4_ASAP7_75t_L g1218 ( 
.A(n_924),
.B(n_878),
.Y(n_1218)
);

INVxp67_ASAP7_75t_L g1219 ( 
.A(n_861),
.Y(n_1219)
);

AND2x4_ASAP7_75t_L g1220 ( 
.A(n_924),
.B(n_878),
.Y(n_1220)
);

OAI22xp33_ASAP7_75t_SL g1221 ( 
.A1(n_832),
.A2(n_860),
.B1(n_865),
.B2(n_836),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_799),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_878),
.B(n_931),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_800),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_804),
.Y(n_1225)
);

INVx4_ASAP7_75t_L g1226 ( 
.A(n_806),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_811),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_801),
.Y(n_1228)
);

INVx4_ASAP7_75t_L g1229 ( 
.A(n_806),
.Y(n_1229)
);

BUFx2_ASAP7_75t_L g1230 ( 
.A(n_1039),
.Y(n_1230)
);

INVx2_ASAP7_75t_SL g1231 ( 
.A(n_1103),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1075),
.B(n_1132),
.Y(n_1232)
);

BUFx6f_ASAP7_75t_L g1233 ( 
.A(n_806),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_812),
.Y(n_1234)
);

BUFx6f_ASAP7_75t_L g1235 ( 
.A(n_806),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1144),
.B(n_1145),
.Y(n_1236)
);

AND2x4_ASAP7_75t_L g1237 ( 
.A(n_878),
.B(n_935),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_813),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_SL g1239 ( 
.A(n_805),
.B(n_1033),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_823),
.Y(n_1240)
);

AOI21x1_ASAP7_75t_L g1241 ( 
.A1(n_965),
.A2(n_956),
.B(n_1065),
.Y(n_1241)
);

INVxp67_ASAP7_75t_L g1242 ( 
.A(n_1059),
.Y(n_1242)
);

AO22x2_ASAP7_75t_L g1243 ( 
.A1(n_1025),
.A2(n_911),
.B1(n_919),
.B2(n_903),
.Y(n_1243)
);

CKINVDCx20_ASAP7_75t_R g1244 ( 
.A(n_1160),
.Y(n_1244)
);

NOR2xp33_ASAP7_75t_L g1245 ( 
.A(n_1157),
.B(n_1167),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_831),
.Y(n_1246)
);

INVx4_ASAP7_75t_L g1247 ( 
.A(n_843),
.Y(n_1247)
);

BUFx6f_ASAP7_75t_L g1248 ( 
.A(n_843),
.Y(n_1248)
);

HB1xp67_ASAP7_75t_L g1249 ( 
.A(n_1173),
.Y(n_1249)
);

INVxp67_ASAP7_75t_L g1250 ( 
.A(n_1184),
.Y(n_1250)
);

INVx4_ASAP7_75t_L g1251 ( 
.A(n_843),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_834),
.Y(n_1252)
);

AND2x4_ASAP7_75t_L g1253 ( 
.A(n_938),
.B(n_945),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1157),
.B(n_1167),
.Y(n_1254)
);

BUFx6f_ASAP7_75t_L g1255 ( 
.A(n_843),
.Y(n_1255)
);

NOR2xp33_ASAP7_75t_L g1256 ( 
.A(n_1204),
.B(n_1208),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_835),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1147),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_839),
.Y(n_1259)
);

INVx3_ASAP7_75t_L g1260 ( 
.A(n_937),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_1147),
.Y(n_1261)
);

AND2x2_ASAP7_75t_SL g1262 ( 
.A(n_810),
.B(n_868),
.Y(n_1262)
);

OR2x6_ASAP7_75t_L g1263 ( 
.A(n_1169),
.B(n_1182),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1187),
.B(n_1192),
.Y(n_1264)
);

INVxp67_ASAP7_75t_L g1265 ( 
.A(n_846),
.Y(n_1265)
);

AO22x2_ASAP7_75t_L g1266 ( 
.A1(n_926),
.A2(n_1118),
.B1(n_820),
.B2(n_923),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_840),
.Y(n_1267)
);

NOR2xp33_ASAP7_75t_L g1268 ( 
.A(n_1204),
.B(n_1208),
.Y(n_1268)
);

INVx4_ASAP7_75t_SL g1269 ( 
.A(n_894),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_844),
.Y(n_1270)
);

OR2x2_ASAP7_75t_L g1271 ( 
.A(n_848),
.B(n_851),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1153),
.Y(n_1272)
);

AOI22x1_ASAP7_75t_L g1273 ( 
.A1(n_1122),
.A2(n_1000),
.B1(n_1030),
.B2(n_991),
.Y(n_1273)
);

BUFx6f_ASAP7_75t_L g1274 ( 
.A(n_849),
.Y(n_1274)
);

INVx5_ASAP7_75t_L g1275 ( 
.A(n_803),
.Y(n_1275)
);

INVx8_ASAP7_75t_L g1276 ( 
.A(n_976),
.Y(n_1276)
);

AO22x2_ASAP7_75t_L g1277 ( 
.A1(n_1118),
.A2(n_820),
.B1(n_923),
.B2(n_889),
.Y(n_1277)
);

OAI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_824),
.A2(n_826),
.B1(n_1042),
.B2(n_1041),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_L g1279 ( 
.A(n_832),
.B(n_1111),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_L g1280 ( 
.A(n_881),
.B(n_828),
.Y(n_1280)
);

BUFx3_ASAP7_75t_L g1281 ( 
.A(n_932),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_819),
.B(n_1050),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1053),
.B(n_1064),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1040),
.Y(n_1284)
);

NAND2xp33_ASAP7_75t_L g1285 ( 
.A(n_1212),
.B(n_803),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1102),
.B(n_1105),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1164),
.B(n_1171),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1045),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1047),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1153),
.Y(n_1290)
);

HB1xp67_ASAP7_75t_L g1291 ( 
.A(n_1185),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1174),
.Y(n_1292)
);

OR2x2_ASAP7_75t_SL g1293 ( 
.A(n_969),
.B(n_982),
.Y(n_1293)
);

HB1xp67_ASAP7_75t_L g1294 ( 
.A(n_1198),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_893),
.B(n_852),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1174),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1108),
.B(n_1135),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1206),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1049),
.Y(n_1299)
);

OR2x6_ASAP7_75t_L g1300 ( 
.A(n_1169),
.B(n_1182),
.Y(n_1300)
);

BUFx4f_ASAP7_75t_L g1301 ( 
.A(n_829),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_SL g1302 ( 
.A(n_1136),
.B(n_1150),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1206),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1057),
.Y(n_1304)
);

BUFx6f_ASAP7_75t_L g1305 ( 
.A(n_849),
.Y(n_1305)
);

BUFx6f_ASAP7_75t_L g1306 ( 
.A(n_849),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1061),
.Y(n_1307)
);

INVx2_ASAP7_75t_SL g1308 ( 
.A(n_883),
.Y(n_1308)
);

NAND2x1p5_ASAP7_75t_L g1309 ( 
.A(n_815),
.B(n_922),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1068),
.Y(n_1310)
);

NAND3xp33_ASAP7_75t_L g1311 ( 
.A(n_836),
.B(n_865),
.C(n_860),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1069),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1198),
.B(n_1100),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1070),
.Y(n_1314)
);

INVxp67_ASAP7_75t_L g1315 ( 
.A(n_1126),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1151),
.B(n_1168),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1209),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1172),
.B(n_1175),
.Y(n_1318)
);

INVx4_ASAP7_75t_L g1319 ( 
.A(n_849),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1209),
.Y(n_1320)
);

INVxp67_ASAP7_75t_SL g1321 ( 
.A(n_841),
.Y(n_1321)
);

INVx1_ASAP7_75t_SL g1322 ( 
.A(n_814),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1140),
.B(n_837),
.Y(n_1323)
);

BUFx10_ASAP7_75t_L g1324 ( 
.A(n_818),
.Y(n_1324)
);

NOR2xp33_ASAP7_75t_L g1325 ( 
.A(n_807),
.B(n_1088),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1073),
.Y(n_1326)
);

BUFx2_ASAP7_75t_L g1327 ( 
.A(n_1039),
.Y(n_1327)
);

NAND2xp33_ASAP7_75t_L g1328 ( 
.A(n_803),
.B(n_1212),
.Y(n_1328)
);

AND2x4_ASAP7_75t_SL g1329 ( 
.A(n_1044),
.B(n_1087),
.Y(n_1329)
);

BUFx2_ASAP7_75t_L g1330 ( 
.A(n_1079),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1074),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1090),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_877),
.B(n_847),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1091),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1003),
.B(n_1005),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1092),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1104),
.Y(n_1337)
);

HB1xp67_ASAP7_75t_L g1338 ( 
.A(n_990),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1122),
.A2(n_896),
.B1(n_906),
.B2(n_888),
.Y(n_1339)
);

BUFx3_ASAP7_75t_L g1340 ( 
.A(n_932),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_SL g1341 ( 
.A(n_1203),
.B(n_1211),
.Y(n_1341)
);

AOI22xp5_ASAP7_75t_L g1342 ( 
.A1(n_916),
.A2(n_962),
.B1(n_988),
.B2(n_961),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1106),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_830),
.Y(n_1344)
);

INVx3_ASAP7_75t_L g1345 ( 
.A(n_937),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_847),
.B(n_950),
.Y(n_1346)
);

AND2x4_ASAP7_75t_L g1347 ( 
.A(n_1143),
.B(n_942),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_SL g1348 ( 
.A(n_807),
.B(n_1088),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1110),
.Y(n_1349)
);

BUFx6f_ASAP7_75t_L g1350 ( 
.A(n_856),
.Y(n_1350)
);

NAND3x1_ASAP7_75t_L g1351 ( 
.A(n_859),
.B(n_1154),
.C(n_896),
.Y(n_1351)
);

BUFx3_ASAP7_75t_L g1352 ( 
.A(n_942),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_874),
.B(n_1109),
.Y(n_1353)
);

AND2x4_ASAP7_75t_L g1354 ( 
.A(n_1143),
.B(n_1007),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1109),
.B(n_1170),
.Y(n_1355)
);

AND2x4_ASAP7_75t_L g1356 ( 
.A(n_1002),
.B(n_1006),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_SL g1357 ( 
.A1(n_1122),
.A2(n_872),
.B1(n_906),
.B2(n_888),
.Y(n_1357)
);

INVx1_ASAP7_75t_SL g1358 ( 
.A(n_814),
.Y(n_1358)
);

BUFx3_ASAP7_75t_L g1359 ( 
.A(n_1079),
.Y(n_1359)
);

BUFx6f_ASAP7_75t_L g1360 ( 
.A(n_856),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1170),
.B(n_1191),
.Y(n_1361)
);

AND2x4_ASAP7_75t_L g1362 ( 
.A(n_970),
.B(n_973),
.Y(n_1362)
);

INVxp67_ASAP7_75t_L g1363 ( 
.A(n_1186),
.Y(n_1363)
);

INVx3_ASAP7_75t_L g1364 ( 
.A(n_937),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_909),
.A2(n_1063),
.B1(n_1078),
.B2(n_1034),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_918),
.B(n_939),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_897),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_897),
.Y(n_1368)
);

BUFx3_ASAP7_75t_L g1369 ( 
.A(n_1083),
.Y(n_1369)
);

INVx3_ASAP7_75t_L g1370 ( 
.A(n_937),
.Y(n_1370)
);

BUFx6f_ASAP7_75t_L g1371 ( 
.A(n_856),
.Y(n_1371)
);

BUFx3_ASAP7_75t_L g1372 ( 
.A(n_1083),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1115),
.Y(n_1373)
);

BUFx6f_ASAP7_75t_L g1374 ( 
.A(n_856),
.Y(n_1374)
);

INVx3_ASAP7_75t_L g1375 ( 
.A(n_857),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_907),
.Y(n_1376)
);

BUFx6f_ASAP7_75t_L g1377 ( 
.A(n_871),
.Y(n_1377)
);

NAND3x1_ASAP7_75t_L g1378 ( 
.A(n_909),
.B(n_915),
.C(n_916),
.Y(n_1378)
);

BUFx2_ASAP7_75t_L g1379 ( 
.A(n_1146),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_961),
.B(n_962),
.Y(n_1380)
);

BUFx6f_ASAP7_75t_L g1381 ( 
.A(n_871),
.Y(n_1381)
);

BUFx3_ASAP7_75t_L g1382 ( 
.A(n_1146),
.Y(n_1382)
);

BUFx10_ASAP7_75t_L g1383 ( 
.A(n_818),
.Y(n_1383)
);

CKINVDCx8_ASAP7_75t_R g1384 ( 
.A(n_1080),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1116),
.Y(n_1385)
);

AND2x6_ASAP7_75t_L g1386 ( 
.A(n_975),
.B(n_862),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1133),
.Y(n_1387)
);

BUFx6f_ASAP7_75t_L g1388 ( 
.A(n_871),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1137),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_907),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_SL g1391 ( 
.A(n_1191),
.B(n_1016),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1141),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_972),
.B(n_866),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_L g1394 ( 
.A(n_999),
.B(n_1008),
.Y(n_1394)
);

INVx3_ASAP7_75t_L g1395 ( 
.A(n_857),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1142),
.Y(n_1396)
);

AND2x4_ASAP7_75t_L g1397 ( 
.A(n_1152),
.B(n_1158),
.Y(n_1397)
);

BUFx2_ASAP7_75t_L g1398 ( 
.A(n_1152),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1148),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1149),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1034),
.A2(n_1078),
.B1(n_1082),
.B2(n_1063),
.Y(n_1401)
);

BUFx6f_ASAP7_75t_L g1402 ( 
.A(n_871),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_1210),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1155),
.Y(n_1404)
);

AND2x2_ASAP7_75t_L g1405 ( 
.A(n_988),
.B(n_992),
.Y(n_1405)
);

NAND2x1p5_ASAP7_75t_L g1406 ( 
.A(n_815),
.B(n_922),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_992),
.B(n_915),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_913),
.Y(n_1408)
);

BUFx6f_ASAP7_75t_L g1409 ( 
.A(n_1054),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_913),
.Y(n_1410)
);

NAND2x1p5_ASAP7_75t_L g1411 ( 
.A(n_815),
.B(n_922),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_SL g1412 ( 
.A(n_1016),
.B(n_936),
.Y(n_1412)
);

A2O1A1Ixp33_ASAP7_75t_L g1413 ( 
.A1(n_1082),
.A2(n_1134),
.B(n_1166),
.C(n_1114),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1159),
.Y(n_1414)
);

AOI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_994),
.A2(n_1011),
.B1(n_998),
.B2(n_981),
.Y(n_1415)
);

AND2x4_ASAP7_75t_L g1416 ( 
.A(n_1158),
.B(n_1051),
.Y(n_1416)
);

AND2x4_ASAP7_75t_L g1417 ( 
.A(n_1051),
.B(n_1097),
.Y(n_1417)
);

AO22x2_ASAP7_75t_L g1418 ( 
.A1(n_889),
.A2(n_941),
.B1(n_943),
.B2(n_1015),
.Y(n_1418)
);

AND2x4_ASAP7_75t_L g1419 ( 
.A(n_1097),
.B(n_1165),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1161),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1176),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1189),
.Y(n_1422)
);

AOI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_994),
.A2(n_1011),
.B1(n_998),
.B2(n_981),
.Y(n_1423)
);

AOI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_954),
.A2(n_825),
.B1(n_1055),
.B2(n_810),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_809),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1190),
.Y(n_1426)
);

NOR2xp33_ASAP7_75t_L g1427 ( 
.A(n_941),
.B(n_943),
.Y(n_1427)
);

BUFx4f_ASAP7_75t_L g1428 ( 
.A(n_1067),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_822),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_914),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1028),
.B(n_1195),
.Y(n_1431)
);

INVx3_ASAP7_75t_L g1432 ( 
.A(n_815),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1199),
.Y(n_1433)
);

NOR2xp33_ASAP7_75t_SL g1434 ( 
.A(n_1121),
.B(n_1062),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1200),
.Y(n_1435)
);

AOI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_954),
.A2(n_1055),
.B1(n_825),
.B2(n_870),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1202),
.Y(n_1437)
);

NOR2xp33_ASAP7_75t_L g1438 ( 
.A(n_1031),
.B(n_1029),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1207),
.B(n_1024),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_845),
.Y(n_1440)
);

BUFx6f_ASAP7_75t_L g1441 ( 
.A(n_1054),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_914),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_850),
.B(n_853),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_854),
.Y(n_1444)
);

AND2x6_ASAP7_75t_L g1445 ( 
.A(n_869),
.B(n_1013),
.Y(n_1445)
);

INVx2_ASAP7_75t_SL g1446 ( 
.A(n_901),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_855),
.Y(n_1447)
);

AND2x4_ASAP7_75t_L g1448 ( 
.A(n_1165),
.B(n_1188),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_858),
.B(n_1038),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1043),
.Y(n_1450)
);

INVx2_ASAP7_75t_SL g1451 ( 
.A(n_901),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_863),
.Y(n_1452)
);

NOR2xp33_ASAP7_75t_L g1453 ( 
.A(n_1114),
.B(n_1134),
.Y(n_1453)
);

AO22x2_ASAP7_75t_L g1454 ( 
.A1(n_1017),
.A2(n_1020),
.B1(n_1037),
.B2(n_1035),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1046),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1052),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1085),
.Y(n_1457)
);

INVx2_ASAP7_75t_SL g1458 ( 
.A(n_901),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1086),
.Y(n_1459)
);

BUFx6f_ASAP7_75t_L g1460 ( 
.A(n_1054),
.Y(n_1460)
);

NAND3xp33_ASAP7_75t_L g1461 ( 
.A(n_1166),
.B(n_1178),
.C(n_886),
.Y(n_1461)
);

BUFx6f_ASAP7_75t_L g1462 ( 
.A(n_1054),
.Y(n_1462)
);

HB1xp67_ASAP7_75t_L g1463 ( 
.A(n_987),
.Y(n_1463)
);

INVx2_ASAP7_75t_L g1464 ( 
.A(n_1089),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1178),
.B(n_1018),
.Y(n_1465)
);

BUFx4f_ASAP7_75t_L g1466 ( 
.A(n_1094),
.Y(n_1466)
);

BUFx10_ASAP7_75t_L g1467 ( 
.A(n_842),
.Y(n_1467)
);

INVx5_ASAP7_75t_L g1468 ( 
.A(n_803),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1093),
.Y(n_1469)
);

NOR2xp33_ASAP7_75t_L g1470 ( 
.A(n_1018),
.B(n_974),
.Y(n_1470)
);

INVx2_ASAP7_75t_SL g1471 ( 
.A(n_1179),
.Y(n_1471)
);

INVx4_ASAP7_75t_SL g1472 ( 
.A(n_894),
.Y(n_1472)
);

AND2x4_ASAP7_75t_L g1473 ( 
.A(n_1188),
.B(n_978),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1096),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_L g1475 ( 
.A(n_802),
.B(n_1035),
.Y(n_1475)
);

NAND2x1p5_ASAP7_75t_L g1476 ( 
.A(n_922),
.B(n_1058),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1112),
.B(n_1124),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_868),
.B(n_882),
.Y(n_1478)
);

AND2x4_ASAP7_75t_L g1479 ( 
.A(n_986),
.B(n_1101),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1125),
.B(n_1128),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1129),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1131),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1138),
.B(n_1139),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1183),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1194),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1197),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1205),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_864),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1186),
.B(n_968),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_873),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1014),
.A2(n_802),
.B1(n_1181),
.B2(n_1180),
.Y(n_1491)
);

BUFx4f_ASAP7_75t_L g1492 ( 
.A(n_929),
.Y(n_1492)
);

AND3x1_ASAP7_75t_L g1493 ( 
.A(n_882),
.B(n_1019),
.C(n_1012),
.Y(n_1493)
);

AND2x6_ASAP7_75t_L g1494 ( 
.A(n_1013),
.B(n_979),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_875),
.Y(n_1495)
);

AOI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_954),
.A2(n_1037),
.B1(n_1181),
.B2(n_1180),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_876),
.Y(n_1497)
);

OR2x2_ASAP7_75t_SL g1498 ( 
.A(n_1022),
.B(n_1032),
.Y(n_1498)
);

OAI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1014),
.A2(n_1127),
.B1(n_1163),
.B2(n_1107),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_879),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_884),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_885),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_895),
.Y(n_1503)
);

NAND2x1p5_ASAP7_75t_L g1504 ( 
.A(n_1058),
.B(n_1117),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_898),
.Y(n_1505)
);

NAND2x1p5_ASAP7_75t_L g1506 ( 
.A(n_1058),
.B(n_1117),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_887),
.Y(n_1507)
);

BUFx6f_ASAP7_75t_L g1508 ( 
.A(n_1101),
.Y(n_1508)
);

AND2x6_ASAP7_75t_L g1509 ( 
.A(n_995),
.B(n_996),
.Y(n_1509)
);

AND2x6_ASAP7_75t_L g1510 ( 
.A(n_1101),
.B(n_1113),
.Y(n_1510)
);

NOR2xp33_ASAP7_75t_L g1511 ( 
.A(n_1056),
.B(n_1071),
.Y(n_1511)
);

AND2x4_ASAP7_75t_L g1512 ( 
.A(n_986),
.B(n_1101),
.Y(n_1512)
);

OAI22xp5_ASAP7_75t_L g1513 ( 
.A1(n_1056),
.A2(n_1127),
.B1(n_1107),
.B2(n_1163),
.Y(n_1513)
);

CKINVDCx11_ASAP7_75t_R g1514 ( 
.A(n_1044),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_899),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_902),
.Y(n_1516)
);

INVx1_ASAP7_75t_SL g1517 ( 
.A(n_890),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_917),
.Y(n_1518)
);

AO22x2_ASAP7_75t_L g1519 ( 
.A1(n_1071),
.A2(n_1076),
.B1(n_933),
.B2(n_930),
.Y(n_1519)
);

BUFx3_ASAP7_75t_L g1520 ( 
.A(n_1113),
.Y(n_1520)
);

OAI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1023),
.A2(n_1027),
.B1(n_1026),
.B2(n_1004),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_867),
.B(n_1120),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1162),
.B(n_977),
.Y(n_1523)
);

INVx3_ASAP7_75t_L g1524 ( 
.A(n_1058),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_910),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_940),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_L g1527 ( 
.A(n_1113),
.B(n_948),
.Y(n_1527)
);

BUFx6f_ASAP7_75t_L g1528 ( 
.A(n_1113),
.Y(n_1528)
);

AND2x6_ASAP7_75t_L g1529 ( 
.A(n_1010),
.B(n_997),
.Y(n_1529)
);

INVx3_ASAP7_75t_L g1530 ( 
.A(n_1117),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_927),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_934),
.Y(n_1532)
);

BUFx6f_ASAP7_75t_L g1533 ( 
.A(n_1117),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_886),
.A2(n_944),
.B1(n_892),
.B2(n_928),
.Y(n_1534)
);

AND2x4_ASAP7_75t_L g1535 ( 
.A(n_976),
.B(n_985),
.Y(n_1535)
);

BUFx3_ASAP7_75t_L g1536 ( 
.A(n_1179),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_953),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_955),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_957),
.Y(n_1539)
);

BUFx3_ASAP7_75t_L g1540 ( 
.A(n_1179),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_959),
.Y(n_1541)
);

AND2x4_ASAP7_75t_L g1542 ( 
.A(n_976),
.B(n_985),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_904),
.B(n_908),
.Y(n_1543)
);

OAI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_892),
.A2(n_900),
.B1(n_928),
.B2(n_1076),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_960),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_SL g1546 ( 
.A(n_900),
.B(n_944),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_963),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_L g1548 ( 
.A(n_904),
.B(n_908),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_967),
.Y(n_1549)
);

AND2x4_ASAP7_75t_L g1550 ( 
.A(n_976),
.B(n_985),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_920),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_920),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_951),
.B(n_964),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_951),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_952),
.Y(n_1555)
);

AO22x2_ASAP7_75t_L g1556 ( 
.A1(n_933),
.A2(n_930),
.B1(n_1001),
.B2(n_1023),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_952),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_964),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_808),
.Y(n_1559)
);

INVx3_ASAP7_75t_L g1560 ( 
.A(n_894),
.Y(n_1560)
);

BUFx6f_ASAP7_75t_L g1561 ( 
.A(n_894),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_954),
.B(n_894),
.Y(n_1562)
);

NAND2x1p5_ASAP7_75t_L g1563 ( 
.A(n_985),
.B(n_993),
.Y(n_1563)
);

AND2x4_ASAP7_75t_L g1564 ( 
.A(n_966),
.B(n_980),
.Y(n_1564)
);

OR2x6_ASAP7_75t_L g1565 ( 
.A(n_1169),
.B(n_1182),
.Y(n_1565)
);

BUFx6f_ASAP7_75t_L g1566 ( 
.A(n_989),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_954),
.B(n_891),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_808),
.Y(n_1568)
);

INVx3_ASAP7_75t_L g1569 ( 
.A(n_816),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_816),
.Y(n_1570)
);

AND2x4_ASAP7_75t_L g1571 ( 
.A(n_984),
.B(n_993),
.Y(n_1571)
);

AND2x2_ASAP7_75t_SL g1572 ( 
.A(n_947),
.B(n_983),
.Y(n_1572)
);

OR2x6_ASAP7_75t_L g1573 ( 
.A(n_1048),
.B(n_1084),
.Y(n_1573)
);

BUFx3_ASAP7_75t_L g1574 ( 
.A(n_1087),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_821),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_821),
.Y(n_1576)
);

BUFx6f_ASAP7_75t_L g1577 ( 
.A(n_989),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_833),
.Y(n_1578)
);

INVx3_ASAP7_75t_L g1579 ( 
.A(n_833),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_891),
.B(n_1119),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_891),
.B(n_1119),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_838),
.Y(n_1582)
);

OAI221xp5_ASAP7_75t_L g1583 ( 
.A1(n_1001),
.A2(n_1012),
.B1(n_1004),
.B2(n_958),
.C(n_947),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_838),
.Y(n_1584)
);

INVx6_ASAP7_75t_L g1585 ( 
.A(n_1098),
.Y(n_1585)
);

AND2x6_ASAP7_75t_L g1586 ( 
.A(n_989),
.B(n_1009),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1036),
.Y(n_1587)
);

AND2x4_ASAP7_75t_L g1588 ( 
.A(n_984),
.B(n_949),
.Y(n_1588)
);

AND2x6_ASAP7_75t_L g1589 ( 
.A(n_989),
.B(n_1009),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_SL g1590 ( 
.A(n_1009),
.B(n_1066),
.Y(n_1590)
);

BUFx6f_ASAP7_75t_L g1591 ( 
.A(n_803),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1036),
.Y(n_1592)
);

BUFx6f_ASAP7_75t_L g1593 ( 
.A(n_1212),
.Y(n_1593)
);

AO22x2_ASAP7_75t_L g1594 ( 
.A1(n_1021),
.A2(n_983),
.B1(n_949),
.B2(n_946),
.Y(n_1594)
);

AO22x2_ASAP7_75t_L g1595 ( 
.A1(n_1021),
.A2(n_946),
.B1(n_817),
.B2(n_905),
.Y(n_1595)
);

INVx5_ASAP7_75t_L g1596 ( 
.A(n_1212),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1009),
.B(n_1196),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1060),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1060),
.Y(n_1599)
);

OA22x2_ASAP7_75t_L g1600 ( 
.A1(n_971),
.A2(n_1081),
.B1(n_1193),
.B2(n_817),
.Y(n_1600)
);

INVx3_ASAP7_75t_L g1601 ( 
.A(n_1066),
.Y(n_1601)
);

AND2x4_ASAP7_75t_L g1602 ( 
.A(n_971),
.B(n_1095),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1072),
.Y(n_1603)
);

INVx3_ASAP7_75t_L g1604 ( 
.A(n_1072),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1077),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1077),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_971),
.B(n_1156),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1095),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1098),
.B(n_925),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_925),
.B(n_880),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1099),
.Y(n_1611)
);

BUFx6f_ASAP7_75t_L g1612 ( 
.A(n_1212),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_891),
.B(n_1099),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1123),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1123),
.Y(n_1615)
);

BUFx6f_ASAP7_75t_L g1616 ( 
.A(n_1156),
.Y(n_1616)
);

AND2x4_ASAP7_75t_L g1617 ( 
.A(n_1201),
.B(n_1021),
.Y(n_1617)
);

OAI22xp5_ASAP7_75t_L g1618 ( 
.A1(n_1201),
.A2(n_891),
.B1(n_1177),
.B2(n_1130),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1130),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_880),
.B(n_905),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_921),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1177),
.Y(n_1622)
);

NOR2xp33_ASAP7_75t_L g1623 ( 
.A(n_1021),
.B(n_842),
.Y(n_1623)
);

INVx8_ASAP7_75t_L g1624 ( 
.A(n_921),
.Y(n_1624)
);

AND2x4_ASAP7_75t_L g1625 ( 
.A(n_1021),
.B(n_924),
.Y(n_1625)
);

AO22x2_ASAP7_75t_L g1626 ( 
.A1(n_1025),
.A2(n_911),
.B1(n_919),
.B2(n_903),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1075),
.B(n_1132),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_799),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_799),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1075),
.B(n_1132),
.Y(n_1630)
);

INVx8_ASAP7_75t_L g1631 ( 
.A(n_976),
.Y(n_1631)
);

AO22x2_ASAP7_75t_L g1632 ( 
.A1(n_1025),
.A2(n_911),
.B1(n_919),
.B2(n_903),
.Y(n_1632)
);

BUFx3_ASAP7_75t_L g1633 ( 
.A(n_1103),
.Y(n_1633)
);

BUFx3_ASAP7_75t_L g1634 ( 
.A(n_1103),
.Y(n_1634)
);

OAI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1075),
.A2(n_1144),
.B1(n_1145),
.B2(n_1132),
.Y(n_1635)
);

AO22x2_ASAP7_75t_L g1636 ( 
.A1(n_1025),
.A2(n_911),
.B1(n_919),
.B2(n_903),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_801),
.Y(n_1637)
);

INVx8_ASAP7_75t_L g1638 ( 
.A(n_976),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_799),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_799),
.Y(n_1640)
);

BUFx6f_ASAP7_75t_L g1641 ( 
.A(n_806),
.Y(n_1641)
);

OA22x2_ASAP7_75t_L g1642 ( 
.A1(n_1025),
.A2(n_622),
.B1(n_631),
.B2(n_630),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_799),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_L g1644 ( 
.A(n_1075),
.B(n_1132),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_799),
.Y(n_1645)
);

CKINVDCx5p33_ASAP7_75t_R g1646 ( 
.A(n_1080),
.Y(n_1646)
);

NOR2xp33_ASAP7_75t_L g1647 ( 
.A(n_1075),
.B(n_1132),
.Y(n_1647)
);

BUFx6f_ASAP7_75t_L g1648 ( 
.A(n_806),
.Y(n_1648)
);

NOR2xp33_ASAP7_75t_L g1649 ( 
.A(n_1075),
.B(n_1132),
.Y(n_1649)
);

AO22x2_ASAP7_75t_L g1650 ( 
.A1(n_1025),
.A2(n_911),
.B1(n_919),
.B2(n_903),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_799),
.Y(n_1651)
);

AND2x4_ASAP7_75t_L g1652 ( 
.A(n_924),
.B(n_878),
.Y(n_1652)
);

AND2x6_ASAP7_75t_L g1653 ( 
.A(n_1000),
.B(n_937),
.Y(n_1653)
);

OR2x2_ASAP7_75t_SL g1654 ( 
.A(n_1111),
.B(n_969),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_801),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_801),
.Y(n_1656)
);

BUFx3_ASAP7_75t_L g1657 ( 
.A(n_1103),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_799),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_799),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_799),
.Y(n_1660)
);

BUFx3_ASAP7_75t_L g1661 ( 
.A(n_1103),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_799),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_799),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_801),
.Y(n_1664)
);

AND2x4_ASAP7_75t_L g1665 ( 
.A(n_924),
.B(n_878),
.Y(n_1665)
);

OAI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1075),
.A2(n_1144),
.B1(n_1145),
.B2(n_1132),
.Y(n_1666)
);

INVxp67_ASAP7_75t_L g1667 ( 
.A(n_827),
.Y(n_1667)
);

NAND3x1_ASAP7_75t_L g1668 ( 
.A(n_1118),
.B(n_1154),
.C(n_859),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_827),
.B(n_861),
.Y(n_1669)
);

AND2x4_ASAP7_75t_L g1670 ( 
.A(n_924),
.B(n_878),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_SL g1671 ( 
.A(n_805),
.B(n_1033),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1075),
.B(n_1132),
.Y(n_1672)
);

AND2x4_ASAP7_75t_L g1673 ( 
.A(n_924),
.B(n_878),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_799),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_801),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_799),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_799),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_799),
.Y(n_1678)
);

INVx1_ASAP7_75t_SL g1679 ( 
.A(n_912),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_799),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_L g1681 ( 
.A(n_1075),
.B(n_1132),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_799),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_799),
.Y(n_1683)
);

A2O1A1Ixp33_ASAP7_75t_L g1684 ( 
.A1(n_1075),
.A2(n_1144),
.B(n_1145),
.C(n_1132),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1075),
.B(n_1132),
.Y(n_1685)
);

NAND2x1p5_ASAP7_75t_L g1686 ( 
.A(n_815),
.B(n_922),
.Y(n_1686)
);

BUFx3_ASAP7_75t_L g1687 ( 
.A(n_1103),
.Y(n_1687)
);

NOR2xp33_ASAP7_75t_L g1688 ( 
.A(n_1075),
.B(n_1132),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_SL g1689 ( 
.A(n_805),
.B(n_1033),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_799),
.Y(n_1690)
);

AND2x4_ASAP7_75t_L g1691 ( 
.A(n_924),
.B(n_878),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_801),
.Y(n_1692)
);

NOR2xp33_ASAP7_75t_L g1693 ( 
.A(n_1075),
.B(n_1132),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1075),
.B(n_1132),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_799),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_801),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1075),
.B(n_1132),
.Y(n_1697)
);

AO22x2_ASAP7_75t_L g1698 ( 
.A1(n_1025),
.A2(n_911),
.B1(n_919),
.B2(n_903),
.Y(n_1698)
);

INVx2_ASAP7_75t_L g1699 ( 
.A(n_801),
.Y(n_1699)
);

INVx3_ASAP7_75t_L g1700 ( 
.A(n_937),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1075),
.B(n_1132),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_827),
.B(n_861),
.Y(n_1702)
);

AO22x2_ASAP7_75t_L g1703 ( 
.A1(n_1025),
.A2(n_911),
.B1(n_919),
.B2(n_903),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_827),
.B(n_861),
.Y(n_1704)
);

AO22x2_ASAP7_75t_L g1705 ( 
.A1(n_1025),
.A2(n_911),
.B1(n_919),
.B2(n_903),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_799),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1075),
.B(n_1132),
.Y(n_1707)
);

BUFx6f_ASAP7_75t_L g1708 ( 
.A(n_806),
.Y(n_1708)
);

AND2x4_ASAP7_75t_L g1709 ( 
.A(n_924),
.B(n_878),
.Y(n_1709)
);

BUFx6f_ASAP7_75t_L g1710 ( 
.A(n_806),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_801),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_801),
.Y(n_1712)
);

OAI22xp33_ASAP7_75t_L g1713 ( 
.A1(n_824),
.A2(n_826),
.B1(n_1033),
.B2(n_805),
.Y(n_1713)
);

BUFx3_ASAP7_75t_L g1714 ( 
.A(n_1103),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_801),
.Y(n_1715)
);

NOR2xp33_ASAP7_75t_L g1716 ( 
.A(n_1075),
.B(n_1132),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_799),
.Y(n_1717)
);

INVx2_ASAP7_75t_SL g1718 ( 
.A(n_1103),
.Y(n_1718)
);

BUFx6f_ASAP7_75t_L g1719 ( 
.A(n_806),
.Y(n_1719)
);

NOR3xp33_ASAP7_75t_L g1720 ( 
.A(n_1111),
.B(n_1118),
.C(n_432),
.Y(n_1720)
);

BUFx6f_ASAP7_75t_L g1721 ( 
.A(n_806),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_799),
.Y(n_1722)
);

CKINVDCx20_ASAP7_75t_R g1723 ( 
.A(n_1160),
.Y(n_1723)
);

BUFx3_ASAP7_75t_L g1724 ( 
.A(n_1103),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_801),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_801),
.Y(n_1726)
);

BUFx6f_ASAP7_75t_L g1727 ( 
.A(n_806),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_799),
.Y(n_1728)
);

INVx3_ASAP7_75t_L g1729 ( 
.A(n_937),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1075),
.B(n_1132),
.Y(n_1730)
);

INVxp67_ASAP7_75t_L g1731 ( 
.A(n_827),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_799),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_801),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_801),
.Y(n_1734)
);

INVx4_ASAP7_75t_L g1735 ( 
.A(n_806),
.Y(n_1735)
);

BUFx6f_ASAP7_75t_L g1736 ( 
.A(n_806),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_L g1737 ( 
.A(n_1075),
.B(n_1132),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_799),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_799),
.Y(n_1739)
);

OAI22xp5_ASAP7_75t_L g1740 ( 
.A1(n_1075),
.A2(n_1144),
.B1(n_1145),
.B2(n_1132),
.Y(n_1740)
);

CKINVDCx20_ASAP7_75t_R g1741 ( 
.A(n_1160),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_799),
.Y(n_1742)
);

AND2x6_ASAP7_75t_L g1743 ( 
.A(n_1000),
.B(n_937),
.Y(n_1743)
);

CKINVDCx5p33_ASAP7_75t_R g1744 ( 
.A(n_1080),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_799),
.Y(n_1745)
);

INVx4_ASAP7_75t_SL g1746 ( 
.A(n_894),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_799),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_799),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_799),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_827),
.B(n_861),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_801),
.Y(n_1751)
);

AND2x4_ASAP7_75t_L g1752 ( 
.A(n_924),
.B(n_878),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_801),
.Y(n_1753)
);

NOR2xp33_ASAP7_75t_L g1754 ( 
.A(n_1075),
.B(n_1132),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_801),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_801),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1075),
.B(n_1132),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_799),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_827),
.B(n_861),
.Y(n_1759)
);

INVx5_ASAP7_75t_L g1760 ( 
.A(n_803),
.Y(n_1760)
);

BUFx3_ASAP7_75t_L g1761 ( 
.A(n_1103),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_799),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_827),
.B(n_861),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1075),
.B(n_1132),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1075),
.B(n_1132),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1075),
.B(n_1132),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_SL g1767 ( 
.A(n_805),
.B(n_1033),
.Y(n_1767)
);

BUFx6f_ASAP7_75t_L g1768 ( 
.A(n_806),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_799),
.Y(n_1769)
);

CKINVDCx14_ASAP7_75t_R g1770 ( 
.A(n_1080),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_801),
.Y(n_1771)
);

NOR2xp33_ASAP7_75t_L g1772 ( 
.A(n_1075),
.B(n_1132),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_799),
.Y(n_1773)
);

NOR2xp33_ASAP7_75t_L g1774 ( 
.A(n_1075),
.B(n_1132),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_827),
.B(n_861),
.Y(n_1775)
);

INVx1_ASAP7_75t_SL g1776 ( 
.A(n_912),
.Y(n_1776)
);

NOR2xp33_ASAP7_75t_L g1777 ( 
.A(n_1075),
.B(n_1132),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_799),
.Y(n_1778)
);

AND2x6_ASAP7_75t_L g1779 ( 
.A(n_1000),
.B(n_937),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_801),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_801),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_799),
.Y(n_1782)
);

AOI22xp5_ASAP7_75t_L g1783 ( 
.A1(n_1118),
.A2(n_619),
.B1(n_791),
.B2(n_916),
.Y(n_1783)
);

AND2x4_ASAP7_75t_L g1784 ( 
.A(n_924),
.B(n_878),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_799),
.Y(n_1785)
);

INVx3_ASAP7_75t_L g1786 ( 
.A(n_937),
.Y(n_1786)
);

NOR2xp33_ASAP7_75t_L g1787 ( 
.A(n_1075),
.B(n_1132),
.Y(n_1787)
);

INVx2_ASAP7_75t_SL g1788 ( 
.A(n_1103),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_801),
.Y(n_1789)
);

BUFx3_ASAP7_75t_L g1790 ( 
.A(n_1103),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_SL g1791 ( 
.A(n_805),
.B(n_1033),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_801),
.Y(n_1792)
);

BUFx6f_ASAP7_75t_L g1793 ( 
.A(n_806),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_799),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_801),
.Y(n_1795)
);

OR2x6_ASAP7_75t_L g1796 ( 
.A(n_1169),
.B(n_1182),
.Y(n_1796)
);

AND2x4_ASAP7_75t_L g1797 ( 
.A(n_924),
.B(n_878),
.Y(n_1797)
);

AND2x6_ASAP7_75t_L g1798 ( 
.A(n_1000),
.B(n_937),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_799),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_801),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_801),
.Y(n_1801)
);

BUFx6f_ASAP7_75t_L g1802 ( 
.A(n_806),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_801),
.Y(n_1803)
);

INVx2_ASAP7_75t_L g1804 ( 
.A(n_801),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_799),
.Y(n_1805)
);

BUFx6f_ASAP7_75t_L g1806 ( 
.A(n_806),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_827),
.B(n_861),
.Y(n_1807)
);

BUFx6f_ASAP7_75t_L g1808 ( 
.A(n_806),
.Y(n_1808)
);

OR2x2_ASAP7_75t_L g1809 ( 
.A(n_846),
.B(n_848),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_799),
.Y(n_1810)
);

CKINVDCx5p33_ASAP7_75t_R g1811 ( 
.A(n_1080),
.Y(n_1811)
);

AND2x6_ASAP7_75t_L g1812 ( 
.A(n_1000),
.B(n_937),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_799),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_801),
.Y(n_1814)
);

AO22x2_ASAP7_75t_L g1815 ( 
.A1(n_1025),
.A2(n_911),
.B1(n_919),
.B2(n_903),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_799),
.Y(n_1816)
);

NOR2xp33_ASAP7_75t_L g1817 ( 
.A(n_1245),
.B(n_1256),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1367),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1367),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_SL g1820 ( 
.A(n_1342),
.B(n_1434),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_L g1821 ( 
.A(n_1394),
.B(n_1245),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1394),
.B(n_1256),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1268),
.B(n_1644),
.Y(n_1823)
);

INVx5_ASAP7_75t_L g1824 ( 
.A(n_1591),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1217),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1268),
.B(n_1644),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1368),
.Y(n_1827)
);

A2O1A1Ixp33_ASAP7_75t_L g1828 ( 
.A1(n_1787),
.A2(n_1649),
.B(n_1681),
.C(n_1647),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1647),
.B(n_1649),
.Y(n_1829)
);

OAI22xp5_ASAP7_75t_SL g1830 ( 
.A1(n_1401),
.A2(n_1365),
.B1(n_1461),
.B2(n_1783),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_SL g1831 ( 
.A(n_1380),
.B(n_1405),
.Y(n_1831)
);

NOR3x1_ASAP7_75t_L g1832 ( 
.A(n_1583),
.B(n_1635),
.C(n_1216),
.Y(n_1832)
);

O2A1O1Ixp33_ASAP7_75t_L g1833 ( 
.A1(n_1684),
.A2(n_1221),
.B(n_1740),
.C(n_1666),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1681),
.B(n_1688),
.Y(n_1834)
);

BUFx6f_ASAP7_75t_L g1835 ( 
.A(n_1591),
.Y(n_1835)
);

AOI22xp5_ASAP7_75t_L g1836 ( 
.A1(n_1688),
.A2(n_1693),
.B1(n_1737),
.B2(n_1716),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1368),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1693),
.B(n_1716),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1217),
.Y(n_1839)
);

AOI22xp33_ASAP7_75t_L g1840 ( 
.A1(n_1720),
.A2(n_1453),
.B1(n_1311),
.B2(n_1412),
.Y(n_1840)
);

AOI22xp5_ASAP7_75t_L g1841 ( 
.A1(n_1737),
.A2(n_1772),
.B1(n_1774),
.B2(n_1754),
.Y(n_1841)
);

OR2x2_ASAP7_75t_L g1842 ( 
.A(n_1407),
.B(n_1293),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1754),
.B(n_1772),
.Y(n_1843)
);

NOR2x2_ASAP7_75t_L g1844 ( 
.A(n_1263),
.B(n_1300),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1774),
.B(n_1777),
.Y(n_1845)
);

AOI22xp5_ASAP7_75t_L g1846 ( 
.A1(n_1777),
.A2(n_1787),
.B1(n_1378),
.B2(n_1279),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1684),
.B(n_1232),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1376),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1236),
.B(n_1254),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1228),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1376),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1627),
.B(n_1630),
.Y(n_1852)
);

AOI22xp33_ASAP7_75t_L g1853 ( 
.A1(n_1720),
.A2(n_1453),
.B1(n_1412),
.B2(n_1279),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1672),
.B(n_1685),
.Y(n_1854)
);

INVx2_ASAP7_75t_SL g1855 ( 
.A(n_1359),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1390),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1694),
.B(n_1697),
.Y(n_1857)
);

NAND3xp33_ASAP7_75t_L g1858 ( 
.A(n_1339),
.B(n_1423),
.C(n_1415),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_SL g1859 ( 
.A(n_1333),
.B(n_1323),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1390),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1701),
.B(n_1707),
.Y(n_1861)
);

OR2x2_ASAP7_75t_L g1862 ( 
.A(n_1339),
.B(n_1654),
.Y(n_1862)
);

NOR2xp33_ASAP7_75t_L g1863 ( 
.A(n_1730),
.B(n_1757),
.Y(n_1863)
);

OAI22x1_ASAP7_75t_SL g1864 ( 
.A1(n_1403),
.A2(n_1811),
.B1(n_1744),
.B2(n_1646),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_L g1865 ( 
.A(n_1764),
.B(n_1765),
.Y(n_1865)
);

OAI22xp5_ASAP7_75t_SL g1866 ( 
.A1(n_1401),
.A2(n_1365),
.B1(n_1357),
.B2(n_1262),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1228),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_SL g1868 ( 
.A(n_1766),
.B(n_1280),
.Y(n_1868)
);

AND2x2_ASAP7_75t_SL g1869 ( 
.A(n_1572),
.B(n_1325),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1408),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1321),
.B(n_1283),
.Y(n_1871)
);

NOR2xp33_ASAP7_75t_L g1872 ( 
.A(n_1470),
.B(n_1280),
.Y(n_1872)
);

NOR2xp33_ASAP7_75t_SL g1873 ( 
.A(n_1384),
.B(n_1413),
.Y(n_1873)
);

NAND3xp33_ASAP7_75t_SL g1874 ( 
.A(n_1357),
.B(n_1391),
.C(n_1353),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1321),
.B(n_1286),
.Y(n_1875)
);

NOR2xp33_ASAP7_75t_L g1876 ( 
.A(n_1470),
.B(n_1282),
.Y(n_1876)
);

NOR2xp33_ASAP7_75t_L g1877 ( 
.A(n_1265),
.B(n_1809),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1572),
.B(n_1295),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1297),
.B(n_1316),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1264),
.B(n_1669),
.Y(n_1880)
);

CKINVDCx5p33_ASAP7_75t_R g1881 ( 
.A(n_1452),
.Y(n_1881)
);

NOR2xp33_ASAP7_75t_L g1882 ( 
.A(n_1265),
.B(n_1271),
.Y(n_1882)
);

NOR2xp33_ASAP7_75t_L g1883 ( 
.A(n_1315),
.B(n_1679),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1318),
.B(n_1393),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1258),
.Y(n_1885)
);

NOR2xp33_ASAP7_75t_L g1886 ( 
.A(n_1315),
.B(n_1776),
.Y(n_1886)
);

CKINVDCx20_ASAP7_75t_R g1887 ( 
.A(n_1244),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1702),
.B(n_1704),
.Y(n_1888)
);

AOI22xp5_ASAP7_75t_L g1889 ( 
.A1(n_1325),
.A2(n_1391),
.B1(n_1351),
.B2(n_1668),
.Y(n_1889)
);

INVx3_ASAP7_75t_L g1890 ( 
.A(n_1591),
.Y(n_1890)
);

BUFx12f_ASAP7_75t_L g1891 ( 
.A(n_1514),
.Y(n_1891)
);

AND2x4_ASAP7_75t_L g1892 ( 
.A(n_1269),
.B(n_1472),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1278),
.B(n_1713),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1278),
.B(n_1713),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1239),
.B(n_1302),
.Y(n_1895)
);

INVx5_ASAP7_75t_L g1896 ( 
.A(n_1593),
.Y(n_1896)
);

OAI21xp5_ASAP7_75t_L g1897 ( 
.A1(n_1475),
.A2(n_1511),
.B(n_1427),
.Y(n_1897)
);

CKINVDCx5p33_ASAP7_75t_R g1898 ( 
.A(n_1770),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_SL g1899 ( 
.A(n_1750),
.B(n_1759),
.Y(n_1899)
);

BUFx2_ASAP7_75t_L g1900 ( 
.A(n_1213),
.Y(n_1900)
);

INVx3_ASAP7_75t_L g1901 ( 
.A(n_1593),
.Y(n_1901)
);

AND2x4_ASAP7_75t_L g1902 ( 
.A(n_1269),
.B(n_1472),
.Y(n_1902)
);

NOR2xp33_ASAP7_75t_L g1903 ( 
.A(n_1219),
.B(n_1242),
.Y(n_1903)
);

INVx4_ASAP7_75t_L g1904 ( 
.A(n_1269),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1408),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1239),
.B(n_1302),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1341),
.B(n_1671),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_SL g1908 ( 
.A(n_1763),
.B(n_1775),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1341),
.B(n_1671),
.Y(n_1909)
);

OR2x6_ASAP7_75t_L g1910 ( 
.A(n_1567),
.B(n_1593),
.Y(n_1910)
);

INVxp33_ASAP7_75t_L g1911 ( 
.A(n_1291),
.Y(n_1911)
);

AOI22xp33_ASAP7_75t_L g1912 ( 
.A1(n_1348),
.A2(n_1262),
.B1(n_1642),
.B2(n_1427),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1807),
.B(n_1689),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1689),
.B(n_1767),
.Y(n_1914)
);

AOI22xp33_ASAP7_75t_L g1915 ( 
.A1(n_1348),
.A2(n_1642),
.B1(n_1355),
.B2(n_1361),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_SL g1916 ( 
.A(n_1366),
.B(n_1287),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1258),
.Y(n_1917)
);

NOR2xp33_ASAP7_75t_L g1918 ( 
.A(n_1219),
.B(n_1242),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1767),
.B(n_1791),
.Y(n_1919)
);

INVx2_ASAP7_75t_L g1920 ( 
.A(n_1261),
.Y(n_1920)
);

AOI22xp33_ASAP7_75t_L g1921 ( 
.A1(n_1465),
.A2(n_1277),
.B1(n_1511),
.B2(n_1475),
.Y(n_1921)
);

O2A1O1Ixp5_ASAP7_75t_L g1922 ( 
.A1(n_1513),
.A2(n_1499),
.B(n_1491),
.C(n_1413),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1261),
.Y(n_1923)
);

AND2x4_ASAP7_75t_L g1924 ( 
.A(n_1472),
.B(n_1746),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_SL g1925 ( 
.A(n_1250),
.B(n_1667),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1272),
.Y(n_1926)
);

NOR2xp33_ASAP7_75t_L g1927 ( 
.A(n_1250),
.B(n_1667),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1791),
.B(n_1438),
.Y(n_1928)
);

OR2x2_ASAP7_75t_L g1929 ( 
.A(n_1478),
.B(n_1534),
.Y(n_1929)
);

AOI22xp33_ASAP7_75t_L g1930 ( 
.A1(n_1277),
.A2(n_1356),
.B1(n_1249),
.B2(n_1215),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_SL g1931 ( 
.A(n_1731),
.B(n_1335),
.Y(n_1931)
);

AND2x2_ASAP7_75t_SL g1932 ( 
.A(n_1285),
.B(n_1328),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1438),
.B(n_1273),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1534),
.B(n_1619),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1622),
.B(n_1277),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1546),
.B(n_1266),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1410),
.Y(n_1937)
);

NOR2xp33_ASAP7_75t_SL g1938 ( 
.A(n_1322),
.B(n_1358),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_L g1939 ( 
.A(n_1546),
.B(n_1266),
.Y(n_1939)
);

OR2x2_ASAP7_75t_L g1940 ( 
.A(n_1544),
.B(n_1215),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_L g1941 ( 
.A(n_1266),
.B(n_1496),
.Y(n_1941)
);

OAI22xp5_ASAP7_75t_L g1942 ( 
.A1(n_1556),
.A2(n_1594),
.B1(n_1519),
.B2(n_1431),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1418),
.B(n_1519),
.Y(n_1943)
);

INVx2_ASAP7_75t_SL g1944 ( 
.A(n_1275),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1410),
.Y(n_1945)
);

OAI21xp5_ASAP7_75t_L g1946 ( 
.A1(n_1436),
.A2(n_1241),
.B(n_1618),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1418),
.B(n_1519),
.Y(n_1947)
);

NAND2xp5_ASAP7_75t_L g1948 ( 
.A(n_1418),
.B(n_1731),
.Y(n_1948)
);

INVx8_ASAP7_75t_L g1949 ( 
.A(n_1510),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_L g1950 ( 
.A(n_1249),
.B(n_1243),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1243),
.B(n_1626),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_SL g1952 ( 
.A(n_1335),
.B(n_1346),
.Y(n_1952)
);

NAND2x1p5_ASAP7_75t_L g1953 ( 
.A(n_1275),
.B(n_1468),
.Y(n_1953)
);

BUFx6f_ASAP7_75t_SL g1954 ( 
.A(n_1535),
.Y(n_1954)
);

HB1xp67_ASAP7_75t_L g1955 ( 
.A(n_1291),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1430),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1272),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1243),
.B(n_1626),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1626),
.B(n_1632),
.Y(n_1959)
);

NOR2xp33_ASAP7_75t_L g1960 ( 
.A(n_1521),
.B(n_1313),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1632),
.B(n_1636),
.Y(n_1961)
);

NOR2xp33_ASAP7_75t_L g1962 ( 
.A(n_1521),
.B(n_1439),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1632),
.B(n_1636),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1636),
.B(n_1650),
.Y(n_1964)
);

NOR2x2_ASAP7_75t_L g1965 ( 
.A(n_1263),
.B(n_1300),
.Y(n_1965)
);

AOI22xp33_ASAP7_75t_L g1966 ( 
.A1(n_1356),
.A2(n_1556),
.B1(n_1354),
.B2(n_1617),
.Y(n_1966)
);

BUFx3_ASAP7_75t_L g1967 ( 
.A(n_1276),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1430),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1442),
.Y(n_1969)
);

AOI21xp5_ASAP7_75t_L g1970 ( 
.A1(n_1285),
.A2(n_1328),
.B(n_1580),
.Y(n_1970)
);

AOI22xp5_ASAP7_75t_L g1971 ( 
.A1(n_1594),
.A2(n_1556),
.B1(n_1623),
.B2(n_1625),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1650),
.B(n_1698),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1650),
.B(n_1698),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1698),
.B(n_1703),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1442),
.Y(n_1975)
);

AOI22xp33_ASAP7_75t_L g1976 ( 
.A1(n_1354),
.A2(n_1617),
.B1(n_1386),
.B2(n_1253),
.Y(n_1976)
);

AOI22xp33_ASAP7_75t_SL g1977 ( 
.A1(n_1595),
.A2(n_1600),
.B1(n_1623),
.B2(n_1594),
.Y(n_1977)
);

NAND3xp33_ASAP7_75t_L g1978 ( 
.A(n_1424),
.B(n_1294),
.C(n_1493),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_SL g1979 ( 
.A(n_1535),
.B(n_1542),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_SL g1980 ( 
.A(n_1542),
.B(n_1550),
.Y(n_1980)
);

BUFx3_ASAP7_75t_L g1981 ( 
.A(n_1276),
.Y(n_1981)
);

NAND2x1_ASAP7_75t_L g1982 ( 
.A(n_1653),
.B(n_1743),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1296),
.Y(n_1983)
);

AOI22xp33_ASAP7_75t_L g1984 ( 
.A1(n_1386),
.A2(n_1253),
.B1(n_1595),
.B2(n_1600),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1703),
.B(n_1705),
.Y(n_1985)
);

HB1xp67_ASAP7_75t_L g1986 ( 
.A(n_1489),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_SL g1987 ( 
.A(n_1550),
.B(n_1347),
.Y(n_1987)
);

OAI22xp5_ASAP7_75t_L g1988 ( 
.A1(n_1498),
.A2(n_1703),
.B1(n_1815),
.B2(n_1705),
.Y(n_1988)
);

OR2x2_ASAP7_75t_L g1989 ( 
.A(n_1463),
.B(n_1581),
.Y(n_1989)
);

NOR2xp33_ASAP7_75t_L g1990 ( 
.A(n_1294),
.B(n_1517),
.Y(n_1990)
);

NAND3xp33_ASAP7_75t_L g1991 ( 
.A(n_1440),
.B(n_1450),
.C(n_1447),
.Y(n_1991)
);

INVx8_ASAP7_75t_L g1992 ( 
.A(n_1510),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_SL g1993 ( 
.A(n_1347),
.B(n_1564),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1296),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1298),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1705),
.B(n_1815),
.Y(n_1996)
);

AOI22xp5_ASAP7_75t_L g1997 ( 
.A1(n_1625),
.A2(n_1815),
.B1(n_1386),
.B2(n_1595),
.Y(n_1997)
);

NOR2xp33_ASAP7_75t_L g1998 ( 
.A(n_1363),
.B(n_1308),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1454),
.B(n_1386),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1298),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1454),
.B(n_1386),
.Y(n_2001)
);

NAND2xp5_ASAP7_75t_L g2002 ( 
.A(n_1454),
.B(n_1509),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1303),
.Y(n_2003)
);

AOI22xp33_ASAP7_75t_SL g2004 ( 
.A1(n_1770),
.A2(n_1620),
.B1(n_1624),
.B2(n_1509),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_L g2005 ( 
.A(n_1509),
.B(n_1444),
.Y(n_2005)
);

NAND3xp33_ASAP7_75t_L g2006 ( 
.A(n_1455),
.B(n_1457),
.C(n_1456),
.Y(n_2006)
);

NOR2xp33_ASAP7_75t_SL g2007 ( 
.A(n_1301),
.B(n_1428),
.Y(n_2007)
);

NOR2xp33_ASAP7_75t_L g2008 ( 
.A(n_1363),
.B(n_1443),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1509),
.B(n_1444),
.Y(n_2009)
);

NAND2xp33_ASAP7_75t_L g2010 ( 
.A(n_1509),
.B(n_1533),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1303),
.Y(n_2011)
);

INVx2_ASAP7_75t_SL g2012 ( 
.A(n_1359),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1317),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1317),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1459),
.B(n_1464),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1459),
.B(n_1464),
.Y(n_2016)
);

NOR2xp33_ASAP7_75t_SL g2017 ( 
.A(n_1301),
.B(n_1428),
.Y(n_2017)
);

OAI22xp5_ASAP7_75t_L g2018 ( 
.A1(n_1222),
.A2(n_1224),
.B1(n_1227),
.B2(n_1225),
.Y(n_2018)
);

AOI22xp33_ASAP7_75t_L g2019 ( 
.A1(n_1564),
.A2(n_1445),
.B1(n_1429),
.B2(n_1425),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1481),
.B(n_1482),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1320),
.Y(n_2021)
);

A2O1A1Ixp33_ASAP7_75t_L g2022 ( 
.A1(n_1527),
.A2(n_1548),
.B(n_1477),
.C(n_1480),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1481),
.B(n_1482),
.Y(n_2023)
);

NOR2xp33_ASAP7_75t_L g2024 ( 
.A(n_1449),
.B(n_1483),
.Y(n_2024)
);

AOI22xp5_ASAP7_75t_L g2025 ( 
.A1(n_1469),
.A2(n_1474),
.B1(n_1486),
.B2(n_1484),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1637),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_1637),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_SL g2028 ( 
.A(n_1416),
.B(n_1397),
.Y(n_2028)
);

HB1xp67_ASAP7_75t_L g2029 ( 
.A(n_1281),
.Y(n_2029)
);

NAND2xp5_ASAP7_75t_L g2030 ( 
.A(n_1485),
.B(n_1375),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_SL g2031 ( 
.A(n_1416),
.B(n_1397),
.Y(n_2031)
);

NOR2xp33_ASAP7_75t_L g2032 ( 
.A(n_1375),
.B(n_1395),
.Y(n_2032)
);

NOR2xp33_ASAP7_75t_L g2033 ( 
.A(n_1395),
.B(n_1487),
.Y(n_2033)
);

NOR3xp33_ASAP7_75t_L g2034 ( 
.A(n_1597),
.B(n_1621),
.C(n_1562),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1485),
.B(n_1445),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1655),
.Y(n_2036)
);

AOI22xp33_ASAP7_75t_L g2037 ( 
.A1(n_1445),
.A2(n_1237),
.B1(n_1223),
.B2(n_1362),
.Y(n_2037)
);

NOR3xp33_ASAP7_75t_L g2038 ( 
.A(n_1597),
.B(n_1621),
.C(n_1610),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_SL g2039 ( 
.A(n_1362),
.B(n_1417),
.Y(n_2039)
);

AND2x6_ASAP7_75t_SL g2040 ( 
.A(n_1573),
.B(n_1263),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1655),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1656),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_SL g2043 ( 
.A(n_1417),
.B(n_1419),
.Y(n_2043)
);

NOR3xp33_ASAP7_75t_L g2044 ( 
.A(n_1214),
.B(n_1718),
.C(n_1231),
.Y(n_2044)
);

NOR2xp33_ASAP7_75t_SL g2045 ( 
.A(n_1466),
.B(n_1492),
.Y(n_2045)
);

AOI22xp5_ASAP7_75t_L g2046 ( 
.A1(n_1494),
.A2(n_1238),
.B1(n_1240),
.B2(n_1234),
.Y(n_2046)
);

NOR2xp33_ASAP7_75t_L g2047 ( 
.A(n_1523),
.B(n_1223),
.Y(n_2047)
);

NOR2xp67_ASAP7_75t_L g2048 ( 
.A(n_1432),
.B(n_1524),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1656),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1344),
.B(n_1494),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_SL g2051 ( 
.A(n_1419),
.B(n_1448),
.Y(n_2051)
);

INVx2_ASAP7_75t_L g2052 ( 
.A(n_1664),
.Y(n_2052)
);

AOI22xp33_ASAP7_75t_L g2053 ( 
.A1(n_1237),
.A2(n_1602),
.B1(n_1607),
.B2(n_1494),
.Y(n_2053)
);

INVx2_ASAP7_75t_L g2054 ( 
.A(n_1664),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_1344),
.B(n_1488),
.Y(n_2055)
);

AOI22xp33_ASAP7_75t_L g2056 ( 
.A1(n_1602),
.A2(n_1607),
.B1(n_1494),
.B2(n_1252),
.Y(n_2056)
);

INVx8_ASAP7_75t_L g2057 ( 
.A(n_1510),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1675),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1675),
.Y(n_2059)
);

O2A1O1Ixp33_ASAP7_75t_L g2060 ( 
.A1(n_1463),
.A2(n_1338),
.B(n_1549),
.C(n_1257),
.Y(n_2060)
);

NAND2x1_ASAP7_75t_L g2061 ( 
.A(n_1653),
.B(n_1743),
.Y(n_2061)
);

AOI22xp5_ASAP7_75t_L g2062 ( 
.A1(n_1494),
.A2(n_1259),
.B1(n_1267),
.B2(n_1246),
.Y(n_2062)
);

AOI22xp33_ASAP7_75t_L g2063 ( 
.A1(n_1270),
.A2(n_1288),
.B1(n_1289),
.B2(n_1284),
.Y(n_2063)
);

AOI22xp5_ASAP7_75t_L g2064 ( 
.A1(n_1299),
.A2(n_1304),
.B1(n_1310),
.B2(n_1307),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1692),
.Y(n_2065)
);

AOI22xp33_ASAP7_75t_L g2066 ( 
.A1(n_1312),
.A2(n_1314),
.B1(n_1331),
.B2(n_1326),
.Y(n_2066)
);

NOR2xp33_ASAP7_75t_L g2067 ( 
.A(n_1332),
.B(n_1816),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1548),
.B(n_1334),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_1336),
.B(n_1337),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_1343),
.B(n_1349),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_SL g2071 ( 
.A(n_1448),
.B(n_1633),
.Y(n_2071)
);

AND2x4_ASAP7_75t_L g2072 ( 
.A(n_1746),
.B(n_1561),
.Y(n_2072)
);

NOR2xp33_ASAP7_75t_SL g2073 ( 
.A(n_1466),
.B(n_1492),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_1373),
.B(n_1385),
.Y(n_2074)
);

INVx2_ASAP7_75t_SL g2075 ( 
.A(n_1275),
.Y(n_2075)
);

AOI22xp33_ASAP7_75t_L g2076 ( 
.A1(n_1387),
.A2(n_1392),
.B1(n_1396),
.B2(n_1389),
.Y(n_2076)
);

INVx3_ASAP7_75t_L g2077 ( 
.A(n_1593),
.Y(n_2077)
);

AOI22xp5_ASAP7_75t_L g2078 ( 
.A1(n_1399),
.A2(n_1404),
.B1(n_1414),
.B2(n_1400),
.Y(n_2078)
);

AND2x6_ASAP7_75t_SL g2079 ( 
.A(n_1573),
.B(n_1300),
.Y(n_2079)
);

INVx2_ASAP7_75t_SL g2080 ( 
.A(n_1369),
.Y(n_2080)
);

INVx2_ASAP7_75t_SL g2081 ( 
.A(n_1369),
.Y(n_2081)
);

AOI22xp33_ASAP7_75t_L g2082 ( 
.A1(n_1420),
.A2(n_1421),
.B1(n_1426),
.B2(n_1422),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_1433),
.B(n_1435),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1692),
.Y(n_2084)
);

HB1xp67_ASAP7_75t_L g2085 ( 
.A(n_1281),
.Y(n_2085)
);

NOR2xp33_ASAP7_75t_L g2086 ( 
.A(n_1437),
.B(n_1628),
.Y(n_2086)
);

CKINVDCx5p33_ASAP7_75t_R g2087 ( 
.A(n_1514),
.Y(n_2087)
);

NAND2x1_ASAP7_75t_L g2088 ( 
.A(n_1653),
.B(n_1743),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_1629),
.B(n_1639),
.Y(n_2089)
);

OR2x2_ASAP7_75t_L g2090 ( 
.A(n_1613),
.B(n_1338),
.Y(n_2090)
);

NOR3x1_ASAP7_75t_L g2091 ( 
.A(n_1788),
.B(n_1451),
.C(n_1446),
.Y(n_2091)
);

AOI22xp5_ASAP7_75t_L g2092 ( 
.A1(n_1640),
.A2(n_1645),
.B1(n_1651),
.B2(n_1643),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_1658),
.B(n_1659),
.Y(n_2093)
);

BUFx6f_ASAP7_75t_L g2094 ( 
.A(n_1612),
.Y(n_2094)
);

NOR2xp33_ASAP7_75t_L g2095 ( 
.A(n_1660),
.B(n_1662),
.Y(n_2095)
);

AOI22xp33_ASAP7_75t_L g2096 ( 
.A1(n_1663),
.A2(n_1676),
.B1(n_1677),
.B2(n_1674),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_L g2097 ( 
.A(n_1678),
.B(n_1680),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_SL g2098 ( 
.A(n_1633),
.B(n_1634),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_1682),
.B(n_1683),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_L g2100 ( 
.A(n_1690),
.B(n_1695),
.Y(n_2100)
);

NOR2xp33_ASAP7_75t_L g2101 ( 
.A(n_1706),
.B(n_1717),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_SL g2102 ( 
.A(n_1634),
.B(n_1657),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_1722),
.B(n_1728),
.Y(n_2103)
);

OAI22xp5_ASAP7_75t_L g2104 ( 
.A1(n_1732),
.A2(n_1739),
.B1(n_1742),
.B2(n_1738),
.Y(n_2104)
);

INVx4_ASAP7_75t_L g2105 ( 
.A(n_1746),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1745),
.B(n_1747),
.Y(n_2106)
);

INVx2_ASAP7_75t_L g2107 ( 
.A(n_1696),
.Y(n_2107)
);

BUFx3_ASAP7_75t_L g2108 ( 
.A(n_1276),
.Y(n_2108)
);

AND2x6_ASAP7_75t_SL g2109 ( 
.A(n_1573),
.B(n_1565),
.Y(n_2109)
);

BUFx2_ASAP7_75t_L g2110 ( 
.A(n_1230),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_SL g2111 ( 
.A(n_1657),
.B(n_1661),
.Y(n_2111)
);

NOR3xp33_ASAP7_75t_SL g2112 ( 
.A(n_1590),
.B(n_1527),
.C(n_1501),
.Y(n_2112)
);

HB1xp67_ASAP7_75t_L g2113 ( 
.A(n_1340),
.Y(n_2113)
);

NOR2xp33_ASAP7_75t_L g2114 ( 
.A(n_1748),
.B(n_1749),
.Y(n_2114)
);

AOI22xp5_ASAP7_75t_L g2115 ( 
.A1(n_1758),
.A2(n_1769),
.B1(n_1773),
.B2(n_1762),
.Y(n_2115)
);

OAI22xp33_ASAP7_75t_L g2116 ( 
.A1(n_1565),
.A2(n_1796),
.B1(n_1687),
.B2(n_1714),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_1778),
.B(n_1782),
.Y(n_2117)
);

INVx8_ASAP7_75t_L g2118 ( 
.A(n_1510),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_1785),
.B(n_1794),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_1799),
.B(n_1805),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1699),
.Y(n_2121)
);

OAI22xp5_ASAP7_75t_L g2122 ( 
.A1(n_1810),
.A2(n_1813),
.B1(n_1468),
.B2(n_1596),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_1488),
.B(n_1495),
.Y(n_2123)
);

NAND2xp5_ASAP7_75t_L g2124 ( 
.A(n_1495),
.B(n_1497),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1711),
.Y(n_2125)
);

BUFx3_ASAP7_75t_L g2126 ( 
.A(n_1631),
.Y(n_2126)
);

NAND3xp33_ASAP7_75t_SL g2127 ( 
.A(n_1543),
.B(n_1553),
.C(n_1503),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1712),
.Y(n_2128)
);

INVxp67_ASAP7_75t_L g2129 ( 
.A(n_1340),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_SL g2130 ( 
.A(n_1661),
.B(n_1687),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1712),
.Y(n_2131)
);

NOR2xp67_ASAP7_75t_L g2132 ( 
.A(n_1432),
.B(n_1524),
.Y(n_2132)
);

NAND2xp33_ASAP7_75t_L g2133 ( 
.A(n_1533),
.B(n_1561),
.Y(n_2133)
);

AOI221xp5_ASAP7_75t_L g2134 ( 
.A1(n_1490),
.A2(n_1516),
.B1(n_1515),
.B2(n_1525),
.C(n_1505),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_1497),
.B(n_1500),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_SL g2136 ( 
.A(n_1714),
.B(n_1724),
.Y(n_2136)
);

AOI22xp33_ASAP7_75t_L g2137 ( 
.A1(n_1500),
.A2(n_1502),
.B1(n_1507),
.B2(n_1518),
.Y(n_2137)
);

AOI22xp33_ASAP7_75t_L g2138 ( 
.A1(n_1502),
.A2(n_1518),
.B1(n_1507),
.B2(n_1539),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_1538),
.B(n_1539),
.Y(n_2139)
);

AOI22xp33_ASAP7_75t_L g2140 ( 
.A1(n_1538),
.A2(n_1541),
.B1(n_1531),
.B2(n_1532),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_L g2141 ( 
.A(n_1715),
.B(n_1725),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_SL g2142 ( 
.A(n_1724),
.B(n_1761),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_1715),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_L g2144 ( 
.A(n_1725),
.B(n_1726),
.Y(n_2144)
);

BUFx3_ASAP7_75t_L g2145 ( 
.A(n_1631),
.Y(n_2145)
);

AOI21xp5_ASAP7_75t_L g2146 ( 
.A1(n_1275),
.A2(n_1596),
.B(n_1468),
.Y(n_2146)
);

NOR2xp33_ASAP7_75t_L g2147 ( 
.A(n_1352),
.B(n_1526),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_1726),
.B(n_1733),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_1733),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_1734),
.B(n_1751),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_SL g2151 ( 
.A(n_1761),
.B(n_1790),
.Y(n_2151)
);

HB1xp67_ASAP7_75t_L g2152 ( 
.A(n_1352),
.Y(n_2152)
);

AND2x2_ASAP7_75t_L g2153 ( 
.A(n_1559),
.B(n_1582),
.Y(n_2153)
);

NOR2xp33_ASAP7_75t_L g2154 ( 
.A(n_1327),
.B(n_1330),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_1751),
.B(n_1753),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1753),
.Y(n_2156)
);

OR2x2_ASAP7_75t_L g2157 ( 
.A(n_1565),
.B(n_1796),
.Y(n_2157)
);

NOR2xp33_ASAP7_75t_L g2158 ( 
.A(n_1379),
.B(n_1398),
.Y(n_2158)
);

INVx2_ASAP7_75t_SL g2159 ( 
.A(n_1468),
.Y(n_2159)
);

BUFx6f_ASAP7_75t_L g2160 ( 
.A(n_1612),
.Y(n_2160)
);

NAND2xp5_ASAP7_75t_SL g2161 ( 
.A(n_1790),
.B(n_1566),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_1755),
.B(n_1756),
.Y(n_2162)
);

NOR2xp67_ASAP7_75t_SL g2163 ( 
.A(n_1596),
.B(n_1760),
.Y(n_2163)
);

AOI22xp5_ASAP7_75t_L g2164 ( 
.A1(n_1537),
.A2(n_1545),
.B1(n_1547),
.B2(n_1529),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_1755),
.B(n_1756),
.Y(n_2165)
);

AOI21xp5_ASAP7_75t_L g2166 ( 
.A1(n_1596),
.A2(n_1760),
.B(n_1771),
.Y(n_2166)
);

HB1xp67_ASAP7_75t_L g2167 ( 
.A(n_1372),
.Y(n_2167)
);

NOR3xp33_ASAP7_75t_SL g2168 ( 
.A(n_1590),
.B(n_1552),
.C(n_1551),
.Y(n_2168)
);

NOR2xp33_ASAP7_75t_L g2169 ( 
.A(n_1522),
.B(n_1554),
.Y(n_2169)
);

NAND2xp5_ASAP7_75t_L g2170 ( 
.A(n_1780),
.B(n_1781),
.Y(n_2170)
);

CKINVDCx16_ASAP7_75t_R g2171 ( 
.A(n_1244),
.Y(n_2171)
);

INVx2_ASAP7_75t_SL g2172 ( 
.A(n_1760),
.Y(n_2172)
);

NOR2xp33_ASAP7_75t_L g2173 ( 
.A(n_1555),
.B(n_1557),
.Y(n_2173)
);

NOR2xp33_ASAP7_75t_L g2174 ( 
.A(n_1558),
.B(n_1372),
.Y(n_2174)
);

AND2x2_ASAP7_75t_L g2175 ( 
.A(n_1559),
.B(n_1582),
.Y(n_2175)
);

NOR2x1p5_ASAP7_75t_L g2176 ( 
.A(n_1574),
.B(n_1560),
.Y(n_2176)
);

NAND2xp5_ASAP7_75t_L g2177 ( 
.A(n_1780),
.B(n_1781),
.Y(n_2177)
);

INVx3_ASAP7_75t_L g2178 ( 
.A(n_1612),
.Y(n_2178)
);

INVx2_ASAP7_75t_SL g2179 ( 
.A(n_1760),
.Y(n_2179)
);

INVx2_ASAP7_75t_L g2180 ( 
.A(n_1789),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_L g2181 ( 
.A(n_1789),
.B(n_1792),
.Y(n_2181)
);

OR2x2_ASAP7_75t_L g2182 ( 
.A(n_1796),
.B(n_1587),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_1792),
.B(n_1795),
.Y(n_2183)
);

OR2x6_ASAP7_75t_L g2184 ( 
.A(n_1612),
.B(n_1561),
.Y(n_2184)
);

NOR2xp33_ASAP7_75t_L g2185 ( 
.A(n_1382),
.B(n_1473),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_SL g2186 ( 
.A(n_1566),
.B(n_1577),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_L g2187 ( 
.A(n_1795),
.B(n_1800),
.Y(n_2187)
);

OAI22xp5_ASAP7_75t_L g2188 ( 
.A1(n_1561),
.A2(n_1560),
.B1(n_1804),
.B2(n_1803),
.Y(n_2188)
);

OAI21xp5_ASAP7_75t_L g2189 ( 
.A1(n_1800),
.A2(n_1803),
.B(n_1801),
.Y(n_2189)
);

INVxp67_ASAP7_75t_SL g2190 ( 
.A(n_1233),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_1804),
.B(n_1814),
.Y(n_2191)
);

AOI22xp5_ASAP7_75t_L g2192 ( 
.A1(n_1529),
.A2(n_1743),
.B1(n_1653),
.B2(n_1812),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_1814),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_1290),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_SL g2195 ( 
.A(n_1566),
.B(n_1577),
.Y(n_2195)
);

BUFx6f_ASAP7_75t_L g2196 ( 
.A(n_1533),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_1587),
.B(n_1592),
.Y(n_2197)
);

AND2x4_ASAP7_75t_L g2198 ( 
.A(n_1218),
.B(n_1220),
.Y(n_2198)
);

CKINVDCx5p33_ASAP7_75t_R g2199 ( 
.A(n_1723),
.Y(n_2199)
);

NAND2xp5_ASAP7_75t_L g2200 ( 
.A(n_1592),
.B(n_1598),
.Y(n_2200)
);

INVx2_ASAP7_75t_SL g2201 ( 
.A(n_1616),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_L g2202 ( 
.A(n_1598),
.B(n_1611),
.Y(n_2202)
);

AOI22xp33_ASAP7_75t_L g2203 ( 
.A1(n_1606),
.A2(n_1611),
.B1(n_1614),
.B2(n_1529),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1292),
.Y(n_2204)
);

NAND2xp5_ASAP7_75t_L g2205 ( 
.A(n_1614),
.B(n_1653),
.Y(n_2205)
);

AND2x2_ASAP7_75t_L g2206 ( 
.A(n_1569),
.B(n_1579),
.Y(n_2206)
);

AOI22xp5_ASAP7_75t_L g2207 ( 
.A1(n_1529),
.A2(n_1812),
.B1(n_1798),
.B2(n_1779),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_1743),
.B(n_1779),
.Y(n_2208)
);

NOR2xp33_ASAP7_75t_L g2209 ( 
.A(n_1382),
.B(n_1473),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_1779),
.B(n_1798),
.Y(n_2210)
);

AND2x2_ASAP7_75t_L g2211 ( 
.A(n_1569),
.B(n_1579),
.Y(n_2211)
);

NAND2x1p5_ASAP7_75t_L g2212 ( 
.A(n_1533),
.B(n_1530),
.Y(n_2212)
);

NAND2xp5_ASAP7_75t_SL g2213 ( 
.A(n_1566),
.B(n_1577),
.Y(n_2213)
);

BUFx5_ASAP7_75t_L g2214 ( 
.A(n_1779),
.Y(n_2214)
);

INVx2_ASAP7_75t_L g2215 ( 
.A(n_1601),
.Y(n_2215)
);

AND2x6_ASAP7_75t_SL g2216 ( 
.A(n_1609),
.B(n_1571),
.Y(n_2216)
);

OAI22xp5_ASAP7_75t_L g2217 ( 
.A1(n_1601),
.A2(n_1604),
.B1(n_1577),
.B2(n_1615),
.Y(n_2217)
);

OR2x6_ASAP7_75t_L g2218 ( 
.A(n_1631),
.B(n_1638),
.Y(n_2218)
);

INVx2_ASAP7_75t_SL g2219 ( 
.A(n_1536),
.Y(n_2219)
);

INVx2_ASAP7_75t_L g2220 ( 
.A(n_1604),
.Y(n_2220)
);

INVx3_ASAP7_75t_L g2221 ( 
.A(n_1779),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_1798),
.B(n_1812),
.Y(n_2222)
);

OR2x2_ASAP7_75t_L g2223 ( 
.A(n_1568),
.B(n_1570),
.Y(n_2223)
);

BUFx12f_ASAP7_75t_SL g2224 ( 
.A(n_1233),
.Y(n_2224)
);

INVx2_ASAP7_75t_L g2225 ( 
.A(n_1530),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_SL g2226 ( 
.A(n_1588),
.B(n_1571),
.Y(n_2226)
);

INVx2_ASAP7_75t_SL g2227 ( 
.A(n_1536),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_1798),
.B(n_1812),
.Y(n_2228)
);

INVx2_ASAP7_75t_L g2229 ( 
.A(n_1575),
.Y(n_2229)
);

AOI22xp33_ASAP7_75t_L g2230 ( 
.A1(n_1529),
.A2(n_1218),
.B1(n_1220),
.B2(n_1797),
.Y(n_2230)
);

AOI22xp33_ASAP7_75t_L g2231 ( 
.A1(n_1652),
.A2(n_1665),
.B1(n_1670),
.B2(n_1797),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_1798),
.Y(n_2232)
);

NAND3xp33_ASAP7_75t_SL g2233 ( 
.A(n_1563),
.B(n_1723),
.C(n_1741),
.Y(n_2233)
);

NAND2xp5_ASAP7_75t_L g2234 ( 
.A(n_1812),
.B(n_1479),
.Y(n_2234)
);

NOR2xp67_ASAP7_75t_L g2235 ( 
.A(n_1260),
.B(n_1345),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_1576),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_SL g2237 ( 
.A(n_1588),
.B(n_1479),
.Y(n_2237)
);

INVx6_ASAP7_75t_L g2238 ( 
.A(n_1638),
.Y(n_2238)
);

AOI22xp33_ASAP7_75t_L g2239 ( 
.A1(n_1652),
.A2(n_1665),
.B1(n_1784),
.B2(n_1752),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_L g2240 ( 
.A(n_1512),
.B(n_1578),
.Y(n_2240)
);

NOR2xp33_ASAP7_75t_SL g2241 ( 
.A(n_1638),
.B(n_1624),
.Y(n_2241)
);

AOI21xp5_ASAP7_75t_L g2242 ( 
.A1(n_1309),
.A2(n_1406),
.B(n_1504),
.Y(n_2242)
);

BUFx2_ASAP7_75t_L g2243 ( 
.A(n_1510),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_1512),
.B(n_1584),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_1599),
.Y(n_2245)
);

AND2x2_ASAP7_75t_L g2246 ( 
.A(n_1603),
.B(n_1605),
.Y(n_2246)
);

NOR2xp33_ASAP7_75t_L g2247 ( 
.A(n_1458),
.B(n_1563),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_SL g2248 ( 
.A(n_1670),
.B(n_1673),
.Y(n_2248)
);

BUFx6f_ASAP7_75t_L g2249 ( 
.A(n_1233),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_L g2250 ( 
.A(n_1608),
.B(n_1260),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_SL g2251 ( 
.A(n_1673),
.B(n_1691),
.Y(n_2251)
);

AO221x1_ASAP7_75t_L g2252 ( 
.A1(n_1616),
.A2(n_1808),
.B1(n_1806),
.B2(n_1233),
.C(n_1235),
.Y(n_2252)
);

OAI22xp33_ASAP7_75t_L g2253 ( 
.A1(n_1624),
.A2(n_1741),
.B1(n_1585),
.B2(n_1574),
.Y(n_2253)
);

INVx3_ASAP7_75t_L g2254 ( 
.A(n_1309),
.Y(n_2254)
);

AND2x4_ASAP7_75t_L g2255 ( 
.A(n_1691),
.B(n_1709),
.Y(n_2255)
);

INVx8_ASAP7_75t_L g2256 ( 
.A(n_1586),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_1345),
.B(n_1364),
.Y(n_2257)
);

AND2x4_ASAP7_75t_L g2258 ( 
.A(n_1709),
.B(n_1784),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_1364),
.B(n_1700),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_1370),
.B(n_1700),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_1406),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_1370),
.B(n_1729),
.Y(n_2262)
);

INVx4_ASAP7_75t_L g2263 ( 
.A(n_1235),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_1411),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_1729),
.B(n_1786),
.Y(n_2265)
);

INVxp67_ASAP7_75t_L g2266 ( 
.A(n_1586),
.Y(n_2266)
);

O2A1O1Ixp33_ASAP7_75t_L g2267 ( 
.A1(n_1520),
.A2(n_1786),
.B(n_1752),
.C(n_1471),
.Y(n_2267)
);

NOR2xp33_ASAP7_75t_L g2268 ( 
.A(n_1540),
.B(n_1585),
.Y(n_2268)
);

AOI221xp5_ASAP7_75t_L g2269 ( 
.A1(n_1540),
.A2(n_1329),
.B1(n_1616),
.B2(n_1520),
.C(n_1247),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_L g2270 ( 
.A(n_1616),
.B(n_1460),
.Y(n_2270)
);

INVxp67_ASAP7_75t_L g2271 ( 
.A(n_1586),
.Y(n_2271)
);

NAND2xp33_ASAP7_75t_L g2272 ( 
.A(n_1586),
.B(n_1589),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_L g2273 ( 
.A(n_1235),
.B(n_1462),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_1411),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_SL g2275 ( 
.A(n_1467),
.B(n_1460),
.Y(n_2275)
);

INVx3_ASAP7_75t_L g2276 ( 
.A(n_1476),
.Y(n_2276)
);

NOR2xp33_ASAP7_75t_L g2277 ( 
.A(n_1585),
.B(n_1226),
.Y(n_2277)
);

INVx1_ASAP7_75t_SL g2278 ( 
.A(n_1235),
.Y(n_2278)
);

AND2x6_ASAP7_75t_SL g2279 ( 
.A(n_1324),
.B(n_1383),
.Y(n_2279)
);

INVx2_ASAP7_75t_SL g2280 ( 
.A(n_1248),
.Y(n_2280)
);

INVx2_ASAP7_75t_SL g2281 ( 
.A(n_1248),
.Y(n_2281)
);

INVx5_ASAP7_75t_L g2282 ( 
.A(n_1248),
.Y(n_2282)
);

NOR2xp33_ASAP7_75t_SL g2283 ( 
.A(n_1586),
.B(n_1589),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_1248),
.B(n_1462),
.Y(n_2284)
);

NAND2xp5_ASAP7_75t_L g2285 ( 
.A(n_1255),
.B(n_1462),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_1255),
.B(n_1462),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_L g2287 ( 
.A(n_1255),
.B(n_1808),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_1255),
.B(n_1808),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_L g2289 ( 
.A(n_1274),
.B(n_1808),
.Y(n_2289)
);

NAND2xp5_ASAP7_75t_L g2290 ( 
.A(n_1274),
.B(n_1806),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_1274),
.B(n_1806),
.Y(n_2291)
);

NOR2xp33_ASAP7_75t_SL g2292 ( 
.A(n_1589),
.B(n_1467),
.Y(n_2292)
);

A2O1A1Ixp33_ASAP7_75t_L g2293 ( 
.A1(n_1329),
.A2(n_1460),
.B(n_1802),
.C(n_1793),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_1274),
.B(n_1806),
.Y(n_2294)
);

NAND2xp5_ASAP7_75t_L g2295 ( 
.A(n_1305),
.B(n_1802),
.Y(n_2295)
);

INVx2_ASAP7_75t_L g2296 ( 
.A(n_1476),
.Y(n_2296)
);

AOI22xp5_ASAP7_75t_L g2297 ( 
.A1(n_1589),
.A2(n_1226),
.B1(n_1229),
.B2(n_1247),
.Y(n_2297)
);

OAI22xp5_ASAP7_75t_L g2298 ( 
.A1(n_1305),
.A2(n_1802),
.B1(n_1793),
.B2(n_1306),
.Y(n_2298)
);

AOI22xp5_ASAP7_75t_L g2299 ( 
.A1(n_1589),
.A2(n_1229),
.B1(n_1251),
.B2(n_1735),
.Y(n_2299)
);

AOI221xp5_ASAP7_75t_L g2300 ( 
.A1(n_1251),
.A2(n_1735),
.B1(n_1319),
.B2(n_1306),
.C(n_1508),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_L g2301 ( 
.A(n_1305),
.B(n_1306),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_1305),
.B(n_1306),
.Y(n_2302)
);

AOI22xp33_ASAP7_75t_SL g2303 ( 
.A1(n_1324),
.A2(n_1383),
.B1(n_1350),
.B2(n_1360),
.Y(n_2303)
);

AOI22xp33_ASAP7_75t_L g2304 ( 
.A1(n_1319),
.A2(n_1350),
.B1(n_1360),
.B2(n_1371),
.Y(n_2304)
);

OAI21xp5_ASAP7_75t_L g2305 ( 
.A1(n_1504),
.A2(n_1686),
.B(n_1506),
.Y(n_2305)
);

OAI22xp5_ASAP7_75t_L g2306 ( 
.A1(n_1350),
.A2(n_1360),
.B1(n_1371),
.B2(n_1374),
.Y(n_2306)
);

AOI22xp33_ASAP7_75t_L g2307 ( 
.A1(n_1371),
.A2(n_1374),
.B1(n_1377),
.B2(n_1381),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_1506),
.Y(n_2308)
);

INVx2_ASAP7_75t_SL g2309 ( 
.A(n_1371),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_1374),
.B(n_1377),
.Y(n_2310)
);

XOR2x2_ASAP7_75t_L g2311 ( 
.A(n_1686),
.B(n_1802),
.Y(n_2311)
);

OAI22xp5_ASAP7_75t_L g2312 ( 
.A1(n_1374),
.A2(n_1377),
.B1(n_1381),
.B2(n_1388),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_L g2313 ( 
.A(n_1377),
.B(n_1381),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_SL g2314 ( 
.A(n_1381),
.B(n_1388),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_1388),
.B(n_1402),
.Y(n_2315)
);

NOR2xp33_ASAP7_75t_L g2316 ( 
.A(n_1388),
.B(n_1402),
.Y(n_2316)
);

NOR2xp33_ASAP7_75t_L g2317 ( 
.A(n_1402),
.B(n_1409),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_1402),
.Y(n_2318)
);

AND2x2_ASAP7_75t_L g2319 ( 
.A(n_1409),
.B(n_1441),
.Y(n_2319)
);

INVx2_ASAP7_75t_SL g2320 ( 
.A(n_1409),
.Y(n_2320)
);

AOI22xp33_ASAP7_75t_L g2321 ( 
.A1(n_1409),
.A2(n_1441),
.B1(n_1460),
.B2(n_1508),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_1441),
.B(n_1508),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_1441),
.B(n_1508),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_L g2324 ( 
.A(n_1528),
.B(n_1641),
.Y(n_2324)
);

INVx2_ASAP7_75t_SL g2325 ( 
.A(n_1793),
.Y(n_2325)
);

INVx2_ASAP7_75t_L g2326 ( 
.A(n_1528),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_1528),
.B(n_1641),
.Y(n_2327)
);

INVx2_ASAP7_75t_L g2328 ( 
.A(n_1528),
.Y(n_2328)
);

OAI22xp5_ASAP7_75t_L g2329 ( 
.A1(n_1641),
.A2(n_1648),
.B1(n_1708),
.B2(n_1710),
.Y(n_2329)
);

AND2x2_ASAP7_75t_L g2330 ( 
.A(n_1641),
.B(n_1648),
.Y(n_2330)
);

NOR2xp33_ASAP7_75t_L g2331 ( 
.A(n_1648),
.B(n_1708),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_L g2332 ( 
.A(n_1648),
.B(n_1708),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_1710),
.B(n_1719),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_L g2334 ( 
.A(n_1710),
.B(n_1719),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_1719),
.B(n_1721),
.Y(n_2335)
);

NOR2xp33_ASAP7_75t_L g2336 ( 
.A(n_1719),
.B(n_1721),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_1721),
.B(n_1727),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_1721),
.Y(n_2338)
);

NOR2xp33_ASAP7_75t_L g2339 ( 
.A(n_1727),
.B(n_1736),
.Y(n_2339)
);

BUFx4_ASAP7_75t_L g2340 ( 
.A(n_1727),
.Y(n_2340)
);

NOR2x1p5_ASAP7_75t_L g2341 ( 
.A(n_1727),
.B(n_1736),
.Y(n_2341)
);

BUFx3_ASAP7_75t_L g2342 ( 
.A(n_1736),
.Y(n_2342)
);

AOI21xp5_ASAP7_75t_L g2343 ( 
.A1(n_1793),
.A2(n_1736),
.B(n_1768),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_1768),
.Y(n_2344)
);

INVx2_ASAP7_75t_SL g2345 ( 
.A(n_1768),
.Y(n_2345)
);

NOR2x1p5_ASAP7_75t_L g2346 ( 
.A(n_1768),
.B(n_829),
.Y(n_2346)
);

NOR2xp33_ASAP7_75t_L g2347 ( 
.A(n_1245),
.B(n_1256),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_1367),
.Y(n_2348)
);

NAND2xp33_ASAP7_75t_L g2349 ( 
.A(n_1378),
.B(n_1342),
.Y(n_2349)
);

OR2x2_ASAP7_75t_L g2350 ( 
.A(n_1342),
.B(n_1380),
.Y(n_2350)
);

AOI22xp5_ASAP7_75t_L g2351 ( 
.A1(n_1342),
.A2(n_1256),
.B1(n_1268),
.B2(n_1245),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_1217),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2354)
);

AOI22xp33_ASAP7_75t_L g2355 ( 
.A1(n_1461),
.A2(n_1118),
.B1(n_1122),
.B2(n_1720),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_L g2356 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2356)
);

AND2x2_ASAP7_75t_L g2357 ( 
.A(n_1380),
.B(n_1405),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_SL g2358 ( 
.A(n_1342),
.B(n_1434),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_SL g2359 ( 
.A(n_1342),
.B(n_1434),
.Y(n_2359)
);

NOR2xp33_ASAP7_75t_L g2360 ( 
.A(n_1245),
.B(n_1256),
.Y(n_2360)
);

AOI22xp5_ASAP7_75t_L g2361 ( 
.A1(n_1342),
.A2(n_1256),
.B1(n_1268),
.B2(n_1245),
.Y(n_2361)
);

AND2x2_ASAP7_75t_L g2362 ( 
.A(n_1380),
.B(n_1405),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_1217),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2364)
);

INVx2_ASAP7_75t_SL g2365 ( 
.A(n_1275),
.Y(n_2365)
);

HB1xp67_ASAP7_75t_L g2366 ( 
.A(n_1213),
.Y(n_2366)
);

INVx5_ASAP7_75t_L g2367 ( 
.A(n_1591),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_1217),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_1367),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_1367),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_L g2372 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2372)
);

AND2x6_ASAP7_75t_SL g2373 ( 
.A(n_1573),
.B(n_1623),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_L g2374 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2374)
);

AOI22xp33_ASAP7_75t_L g2375 ( 
.A1(n_1461),
.A2(n_1118),
.B1(n_1122),
.B2(n_1720),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_SL g2376 ( 
.A(n_1342),
.B(n_1434),
.Y(n_2376)
);

AND2x2_ASAP7_75t_L g2377 ( 
.A(n_1380),
.B(n_1405),
.Y(n_2377)
);

NAND2xp5_ASAP7_75t_L g2378 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2378)
);

AOI22xp5_ASAP7_75t_L g2379 ( 
.A1(n_1342),
.A2(n_1256),
.B1(n_1268),
.B2(n_1245),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2380)
);

AOI22xp33_ASAP7_75t_L g2381 ( 
.A1(n_1461),
.A2(n_1118),
.B1(n_1122),
.B2(n_1720),
.Y(n_2381)
);

NAND2xp5_ASAP7_75t_SL g2382 ( 
.A(n_1342),
.B(n_1434),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_1367),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_SL g2384 ( 
.A(n_1342),
.B(n_1434),
.Y(n_2384)
);

AND2x6_ASAP7_75t_SL g2385 ( 
.A(n_1573),
.B(n_1623),
.Y(n_2385)
);

INVx2_ASAP7_75t_L g2386 ( 
.A(n_1217),
.Y(n_2386)
);

AND2x4_ASAP7_75t_L g2387 ( 
.A(n_1269),
.B(n_1472),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_SL g2388 ( 
.A(n_1342),
.B(n_1434),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_SL g2389 ( 
.A(n_1342),
.B(n_1434),
.Y(n_2389)
);

INVx2_ASAP7_75t_L g2390 ( 
.A(n_1217),
.Y(n_2390)
);

INVx8_ASAP7_75t_L g2391 ( 
.A(n_1510),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_L g2392 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2392)
);

INVx2_ASAP7_75t_L g2393 ( 
.A(n_1217),
.Y(n_2393)
);

NAND2xp5_ASAP7_75t_L g2394 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2394)
);

AOI22xp5_ASAP7_75t_L g2395 ( 
.A1(n_1342),
.A2(n_1256),
.B1(n_1268),
.B2(n_1245),
.Y(n_2395)
);

AOI22xp5_ASAP7_75t_L g2396 ( 
.A1(n_1342),
.A2(n_1256),
.B1(n_1268),
.B2(n_1245),
.Y(n_2396)
);

A2O1A1Ixp33_ASAP7_75t_L g2397 ( 
.A1(n_1342),
.A2(n_1256),
.B(n_1268),
.C(n_1245),
.Y(n_2397)
);

BUFx3_ASAP7_75t_L g2398 ( 
.A(n_1276),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_SL g2399 ( 
.A(n_1342),
.B(n_1434),
.Y(n_2399)
);

INVxp67_ASAP7_75t_L g2400 ( 
.A(n_1213),
.Y(n_2400)
);

O2A1O1Ixp5_ASAP7_75t_L g2401 ( 
.A1(n_1391),
.A2(n_1412),
.B(n_1348),
.C(n_860),
.Y(n_2401)
);

INVx4_ASAP7_75t_L g2402 ( 
.A(n_1269),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2403)
);

NOR2xp33_ASAP7_75t_L g2404 ( 
.A(n_1245),
.B(n_1256),
.Y(n_2404)
);

AND2x4_ASAP7_75t_SL g2405 ( 
.A(n_1561),
.B(n_1591),
.Y(n_2405)
);

BUFx12f_ASAP7_75t_L g2406 ( 
.A(n_1514),
.Y(n_2406)
);

AOI22xp5_ASAP7_75t_L g2407 ( 
.A1(n_1342),
.A2(n_1256),
.B1(n_1268),
.B2(n_1245),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_SL g2408 ( 
.A(n_1342),
.B(n_1434),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_1367),
.Y(n_2409)
);

OR2x2_ASAP7_75t_L g2410 ( 
.A(n_1342),
.B(n_1380),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_1367),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_1217),
.Y(n_2412)
);

AOI22xp33_ASAP7_75t_L g2413 ( 
.A1(n_1461),
.A2(n_1118),
.B1(n_1122),
.B2(n_1720),
.Y(n_2413)
);

NAND2xp5_ASAP7_75t_L g2414 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2414)
);

AOI22xp5_ASAP7_75t_L g2415 ( 
.A1(n_1342),
.A2(n_1256),
.B1(n_1268),
.B2(n_1245),
.Y(n_2415)
);

INVxp33_ASAP7_75t_L g2416 ( 
.A(n_1213),
.Y(n_2416)
);

OR2x2_ASAP7_75t_L g2417 ( 
.A(n_1342),
.B(n_1380),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_L g2418 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_1367),
.Y(n_2419)
);

INVxp67_ASAP7_75t_L g2420 ( 
.A(n_1213),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_SL g2421 ( 
.A(n_1342),
.B(n_1434),
.Y(n_2421)
);

INVx3_ASAP7_75t_L g2422 ( 
.A(n_1591),
.Y(n_2422)
);

NOR2xp33_ASAP7_75t_L g2423 ( 
.A(n_1245),
.B(n_1256),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_L g2424 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2424)
);

NAND2xp5_ASAP7_75t_L g2425 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2425)
);

AND2x4_ASAP7_75t_L g2426 ( 
.A(n_1269),
.B(n_1472),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_SL g2427 ( 
.A(n_1342),
.B(n_1434),
.Y(n_2427)
);

AOI22xp33_ASAP7_75t_L g2428 ( 
.A1(n_1461),
.A2(n_1118),
.B1(n_1122),
.B2(n_1720),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_1367),
.Y(n_2429)
);

NAND2xp5_ASAP7_75t_L g2430 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2432)
);

CKINVDCx5p33_ASAP7_75t_R g2433 ( 
.A(n_1403),
.Y(n_2433)
);

CKINVDCx20_ASAP7_75t_R g2434 ( 
.A(n_1244),
.Y(n_2434)
);

OAI22xp5_ASAP7_75t_L g2435 ( 
.A1(n_1342),
.A2(n_1256),
.B1(n_1268),
.B2(n_1245),
.Y(n_2435)
);

CKINVDCx5p33_ASAP7_75t_R g2436 ( 
.A(n_1403),
.Y(n_2436)
);

BUFx3_ASAP7_75t_L g2437 ( 
.A(n_1276),
.Y(n_2437)
);

AOI22xp33_ASAP7_75t_L g2438 ( 
.A1(n_1461),
.A2(n_1118),
.B1(n_1122),
.B2(n_1720),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_L g2439 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2439)
);

OAI21xp5_ASAP7_75t_L g2440 ( 
.A1(n_1415),
.A2(n_1423),
.B(n_1394),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_1367),
.Y(n_2441)
);

NOR2xp33_ASAP7_75t_L g2442 ( 
.A(n_1245),
.B(n_1256),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_L g2443 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2443)
);

AOI22xp5_ASAP7_75t_L g2444 ( 
.A1(n_1342),
.A2(n_1256),
.B1(n_1268),
.B2(n_1245),
.Y(n_2444)
);

NAND3xp33_ASAP7_75t_L g2445 ( 
.A(n_1720),
.B(n_1118),
.C(n_1111),
.Y(n_2445)
);

NOR3xp33_ASAP7_75t_SL g2446 ( 
.A(n_1521),
.B(n_1023),
.C(n_1583),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_L g2447 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_L g2448 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2448)
);

HB1xp67_ASAP7_75t_L g2449 ( 
.A(n_1213),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_L g2450 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2450)
);

NOR2xp33_ASAP7_75t_L g2451 ( 
.A(n_1245),
.B(n_1256),
.Y(n_2451)
);

NAND2xp5_ASAP7_75t_L g2452 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2452)
);

AND2x4_ASAP7_75t_L g2453 ( 
.A(n_1269),
.B(n_1472),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_L g2454 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2454)
);

NAND2xp5_ASAP7_75t_L g2455 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2455)
);

NOR2xp33_ASAP7_75t_L g2456 ( 
.A(n_1245),
.B(n_1256),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_1367),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_1367),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_L g2459 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2460)
);

INVx1_ASAP7_75t_L g2461 ( 
.A(n_1367),
.Y(n_2461)
);

NOR2xp67_ASAP7_75t_L g2462 ( 
.A(n_1311),
.B(n_1342),
.Y(n_2462)
);

NAND2xp5_ASAP7_75t_L g2463 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2463)
);

NAND2xp5_ASAP7_75t_L g2464 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2464)
);

NAND2xp5_ASAP7_75t_L g2465 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_L g2467 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2467)
);

NOR3xp33_ASAP7_75t_L g2468 ( 
.A(n_1216),
.B(n_1111),
.C(n_1635),
.Y(n_2468)
);

NAND2xp5_ASAP7_75t_SL g2469 ( 
.A(n_1342),
.B(n_1434),
.Y(n_2469)
);

NAND2xp5_ASAP7_75t_L g2470 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2470)
);

AND2x2_ASAP7_75t_L g2471 ( 
.A(n_1380),
.B(n_1405),
.Y(n_2471)
);

INVxp67_ASAP7_75t_L g2472 ( 
.A(n_1213),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_1367),
.Y(n_2473)
);

AOI21xp5_ASAP7_75t_L g2474 ( 
.A1(n_1412),
.A2(n_1321),
.B(n_1394),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_1367),
.Y(n_2475)
);

INVx4_ASAP7_75t_L g2476 ( 
.A(n_1269),
.Y(n_2476)
);

NAND2xp5_ASAP7_75t_SL g2477 ( 
.A(n_1342),
.B(n_1434),
.Y(n_2477)
);

O2A1O1Ixp33_ASAP7_75t_L g2478 ( 
.A1(n_1684),
.A2(n_1221),
.B(n_1635),
.C(n_1216),
.Y(n_2478)
);

NAND2xp5_ASAP7_75t_L g2479 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2479)
);

INVx3_ASAP7_75t_L g2480 ( 
.A(n_1591),
.Y(n_2480)
);

INVx4_ASAP7_75t_L g2481 ( 
.A(n_1269),
.Y(n_2481)
);

AND2x2_ASAP7_75t_L g2482 ( 
.A(n_1380),
.B(n_1405),
.Y(n_2482)
);

OR2x6_ASAP7_75t_L g2483 ( 
.A(n_1391),
.B(n_1567),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_1367),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_1367),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_L g2486 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2486)
);

INVx3_ASAP7_75t_L g2487 ( 
.A(n_1591),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_L g2488 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_L g2489 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2489)
);

NAND2xp5_ASAP7_75t_L g2490 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2490)
);

NAND2xp5_ASAP7_75t_SL g2491 ( 
.A(n_1342),
.B(n_1434),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_1367),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_L g2493 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_L g2494 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2494)
);

OR2x2_ASAP7_75t_L g2495 ( 
.A(n_1342),
.B(n_1380),
.Y(n_2495)
);

NAND3xp33_ASAP7_75t_L g2496 ( 
.A(n_1720),
.B(n_1118),
.C(n_1111),
.Y(n_2496)
);

BUFx6f_ASAP7_75t_L g2497 ( 
.A(n_1591),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_L g2498 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2498)
);

INVx1_ASAP7_75t_L g2499 ( 
.A(n_1367),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_L g2500 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2500)
);

INVx8_ASAP7_75t_L g2501 ( 
.A(n_1510),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_1367),
.Y(n_2502)
);

NAND2xp5_ASAP7_75t_SL g2503 ( 
.A(n_1342),
.B(n_1434),
.Y(n_2503)
);

NOR2xp33_ASAP7_75t_L g2504 ( 
.A(n_1245),
.B(n_1256),
.Y(n_2504)
);

BUFx3_ASAP7_75t_L g2505 ( 
.A(n_1276),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_1367),
.Y(n_2506)
);

NAND2xp5_ASAP7_75t_L g2507 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_1367),
.Y(n_2508)
);

NOR2x2_ASAP7_75t_L g2509 ( 
.A(n_1263),
.B(n_1025),
.Y(n_2509)
);

AOI22xp5_ASAP7_75t_L g2510 ( 
.A1(n_1342),
.A2(n_1256),
.B1(n_1268),
.B2(n_1245),
.Y(n_2510)
);

AND2x6_ASAP7_75t_SL g2511 ( 
.A(n_1573),
.B(n_1623),
.Y(n_2511)
);

NAND2xp5_ASAP7_75t_L g2512 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2512)
);

BUFx3_ASAP7_75t_L g2513 ( 
.A(n_1276),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_L g2514 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2514)
);

AOI221xp5_ASAP7_75t_L g2515 ( 
.A1(n_1216),
.A2(n_1666),
.B1(n_1740),
.B2(n_1635),
.C(n_1221),
.Y(n_2515)
);

NAND2xp5_ASAP7_75t_L g2516 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2516)
);

CKINVDCx5p33_ASAP7_75t_R g2517 ( 
.A(n_1403),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_L g2518 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2518)
);

NAND2xp5_ASAP7_75t_L g2519 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2519)
);

AOI21xp5_ASAP7_75t_L g2520 ( 
.A1(n_1412),
.A2(n_1321),
.B(n_1394),
.Y(n_2520)
);

INVx2_ASAP7_75t_SL g2521 ( 
.A(n_1275),
.Y(n_2521)
);

INVx2_ASAP7_75t_SL g2522 ( 
.A(n_1275),
.Y(n_2522)
);

CKINVDCx5p33_ASAP7_75t_R g2523 ( 
.A(n_1403),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_1367),
.Y(n_2524)
);

NOR2xp33_ASAP7_75t_L g2525 ( 
.A(n_1245),
.B(n_1256),
.Y(n_2525)
);

NAND2xp5_ASAP7_75t_L g2526 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2526)
);

INVxp67_ASAP7_75t_SL g2527 ( 
.A(n_1321),
.Y(n_2527)
);

NOR3xp33_ASAP7_75t_L g2528 ( 
.A(n_1216),
.B(n_1111),
.C(n_1635),
.Y(n_2528)
);

OAI221xp5_ASAP7_75t_L g2529 ( 
.A1(n_1342),
.A2(n_1783),
.B1(n_1063),
.B2(n_1082),
.C(n_1078),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_SL g2530 ( 
.A(n_1342),
.B(n_1434),
.Y(n_2530)
);

INVx2_ASAP7_75t_SL g2531 ( 
.A(n_1359),
.Y(n_2531)
);

OA22x2_ASAP7_75t_L g2532 ( 
.A1(n_1783),
.A2(n_1342),
.B1(n_1025),
.B2(n_1154),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_1367),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2534)
);

NAND2xp5_ASAP7_75t_L g2535 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2535)
);

AOI22xp5_ASAP7_75t_L g2536 ( 
.A1(n_1342),
.A2(n_1256),
.B1(n_1268),
.B2(n_1245),
.Y(n_2536)
);

NAND2xp5_ASAP7_75t_L g2537 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2537)
);

OAI21xp5_ASAP7_75t_L g2538 ( 
.A1(n_1415),
.A2(n_1423),
.B(n_1394),
.Y(n_2538)
);

AND2x2_ASAP7_75t_L g2539 ( 
.A(n_1380),
.B(n_1405),
.Y(n_2539)
);

INVx2_ASAP7_75t_SL g2540 ( 
.A(n_1359),
.Y(n_2540)
);

NAND2xp33_ASAP7_75t_L g2541 ( 
.A(n_1378),
.B(n_1342),
.Y(n_2541)
);

NAND2xp5_ASAP7_75t_L g2542 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_L g2543 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_L g2544 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2544)
);

NOR3xp33_ASAP7_75t_L g2545 ( 
.A(n_1216),
.B(n_1111),
.C(n_1635),
.Y(n_2545)
);

NOR3xp33_ASAP7_75t_L g2546 ( 
.A(n_1216),
.B(n_1111),
.C(n_1635),
.Y(n_2546)
);

NAND2xp5_ASAP7_75t_L g2547 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2547)
);

AND2x4_ASAP7_75t_L g2548 ( 
.A(n_1269),
.B(n_1472),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_SL g2549 ( 
.A(n_1342),
.B(n_1434),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_1367),
.Y(n_2550)
);

NOR3xp33_ASAP7_75t_L g2551 ( 
.A(n_1216),
.B(n_1111),
.C(n_1635),
.Y(n_2551)
);

INVxp67_ASAP7_75t_L g2552 ( 
.A(n_1213),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_SL g2553 ( 
.A(n_1342),
.B(n_1434),
.Y(n_2553)
);

INVx1_ASAP7_75t_SL g2554 ( 
.A(n_1679),
.Y(n_2554)
);

NAND2xp5_ASAP7_75t_L g2555 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_SL g2556 ( 
.A(n_1342),
.B(n_1434),
.Y(n_2556)
);

NAND2xp5_ASAP7_75t_SL g2557 ( 
.A(n_1342),
.B(n_1434),
.Y(n_2557)
);

AOI22xp5_ASAP7_75t_L g2558 ( 
.A1(n_1342),
.A2(n_1256),
.B1(n_1268),
.B2(n_1245),
.Y(n_2558)
);

AND2x2_ASAP7_75t_L g2559 ( 
.A(n_1380),
.B(n_1405),
.Y(n_2559)
);

INVx2_ASAP7_75t_L g2560 ( 
.A(n_1217),
.Y(n_2560)
);

AOI22xp5_ASAP7_75t_L g2561 ( 
.A1(n_1342),
.A2(n_1256),
.B1(n_1268),
.B2(n_1245),
.Y(n_2561)
);

INVx2_ASAP7_75t_L g2562 ( 
.A(n_1217),
.Y(n_2562)
);

AOI22xp33_ASAP7_75t_L g2563 ( 
.A1(n_1461),
.A2(n_1118),
.B1(n_1122),
.B2(n_1720),
.Y(n_2563)
);

INVx2_ASAP7_75t_L g2564 ( 
.A(n_1217),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_L g2565 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2565)
);

NAND2xp5_ASAP7_75t_L g2566 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2566)
);

NOR2xp33_ASAP7_75t_L g2567 ( 
.A(n_1245),
.B(n_1256),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_1367),
.Y(n_2568)
);

INVx3_ASAP7_75t_L g2569 ( 
.A(n_1591),
.Y(n_2569)
);

NOR2xp33_ASAP7_75t_R g2570 ( 
.A(n_1403),
.B(n_740),
.Y(n_2570)
);

NOR2xp33_ASAP7_75t_L g2571 ( 
.A(n_1245),
.B(n_1256),
.Y(n_2571)
);

NAND2xp5_ASAP7_75t_L g2572 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2572)
);

NAND2xp5_ASAP7_75t_SL g2573 ( 
.A(n_1342),
.B(n_1434),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_SL g2574 ( 
.A(n_1342),
.B(n_1434),
.Y(n_2574)
);

HB1xp67_ASAP7_75t_L g2575 ( 
.A(n_1213),
.Y(n_2575)
);

NAND2xp5_ASAP7_75t_L g2576 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2576)
);

INVx5_ASAP7_75t_L g2577 ( 
.A(n_1591),
.Y(n_2577)
);

AOI22xp5_ASAP7_75t_L g2578 ( 
.A1(n_1342),
.A2(n_1256),
.B1(n_1268),
.B2(n_1245),
.Y(n_2578)
);

NAND2xp33_ASAP7_75t_L g2579 ( 
.A(n_1378),
.B(n_1342),
.Y(n_2579)
);

INVx4_ASAP7_75t_L g2580 ( 
.A(n_1269),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_1367),
.Y(n_2581)
);

INVx2_ASAP7_75t_L g2582 ( 
.A(n_1217),
.Y(n_2582)
);

NAND2xp5_ASAP7_75t_L g2583 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2583)
);

AOI22xp33_ASAP7_75t_L g2584 ( 
.A1(n_1461),
.A2(n_1118),
.B1(n_1122),
.B2(n_1720),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_L g2585 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2585)
);

NAND2x1_ASAP7_75t_L g2586 ( 
.A(n_1653),
.B(n_1743),
.Y(n_2586)
);

AND2x4_ASAP7_75t_L g2587 ( 
.A(n_1269),
.B(n_1472),
.Y(n_2587)
);

OAI22xp5_ASAP7_75t_L g2588 ( 
.A1(n_1342),
.A2(n_1256),
.B1(n_1268),
.B2(n_1245),
.Y(n_2588)
);

NAND2xp5_ASAP7_75t_SL g2589 ( 
.A(n_1342),
.B(n_1434),
.Y(n_2589)
);

NAND2xp5_ASAP7_75t_L g2590 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2590)
);

NAND2xp5_ASAP7_75t_L g2591 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2591)
);

NOR2xp33_ASAP7_75t_L g2592 ( 
.A(n_1245),
.B(n_1256),
.Y(n_2592)
);

AND2x6_ASAP7_75t_L g2593 ( 
.A(n_1436),
.B(n_1591),
.Y(n_2593)
);

NAND2xp5_ASAP7_75t_L g2594 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2594)
);

NAND2xp5_ASAP7_75t_SL g2595 ( 
.A(n_1342),
.B(n_1434),
.Y(n_2595)
);

NOR2x1p5_ASAP7_75t_L g2596 ( 
.A(n_1461),
.B(n_829),
.Y(n_2596)
);

NAND2xp5_ASAP7_75t_L g2597 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2597)
);

NAND2xp5_ASAP7_75t_L g2598 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2598)
);

AOI22xp33_ASAP7_75t_SL g2599 ( 
.A1(n_1461),
.A2(n_626),
.B1(n_702),
.B2(n_623),
.Y(n_2599)
);

NOR2xp33_ASAP7_75t_L g2600 ( 
.A(n_1245),
.B(n_1256),
.Y(n_2600)
);

NOR2x2_ASAP7_75t_L g2601 ( 
.A(n_1263),
.B(n_1025),
.Y(n_2601)
);

NAND2xp5_ASAP7_75t_L g2602 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2602)
);

AND2x2_ASAP7_75t_L g2603 ( 
.A(n_1380),
.B(n_1405),
.Y(n_2603)
);

INVx1_ASAP7_75t_SL g2604 ( 
.A(n_1679),
.Y(n_2604)
);

NAND2x1p5_ASAP7_75t_L g2605 ( 
.A(n_1275),
.B(n_1468),
.Y(n_2605)
);

NAND2xp5_ASAP7_75t_SL g2606 ( 
.A(n_1342),
.B(n_1434),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_1367),
.Y(n_2607)
);

NOR2xp33_ASAP7_75t_L g2608 ( 
.A(n_1245),
.B(n_1256),
.Y(n_2608)
);

NOR3xp33_ASAP7_75t_L g2609 ( 
.A(n_1216),
.B(n_1111),
.C(n_1635),
.Y(n_2609)
);

NAND2xp5_ASAP7_75t_L g2610 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2610)
);

INVx1_ASAP7_75t_L g2611 ( 
.A(n_1367),
.Y(n_2611)
);

NAND2xp5_ASAP7_75t_L g2612 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2612)
);

INVx2_ASAP7_75t_SL g2613 ( 
.A(n_1359),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_SL g2614 ( 
.A(n_1342),
.B(n_1434),
.Y(n_2614)
);

NOR2xp67_ASAP7_75t_L g2615 ( 
.A(n_1311),
.B(n_1342),
.Y(n_2615)
);

AOI21xp5_ASAP7_75t_L g2616 ( 
.A1(n_1412),
.A2(n_1321),
.B(n_1394),
.Y(n_2616)
);

AOI22xp33_ASAP7_75t_L g2617 ( 
.A1(n_1461),
.A2(n_1118),
.B1(n_1122),
.B2(n_1720),
.Y(n_2617)
);

NAND2xp5_ASAP7_75t_L g2618 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2618)
);

AOI22xp5_ASAP7_75t_L g2619 ( 
.A1(n_1342),
.A2(n_1256),
.B1(n_1268),
.B2(n_1245),
.Y(n_2619)
);

NAND2xp5_ASAP7_75t_L g2620 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2620)
);

NOR2xp33_ASAP7_75t_L g2621 ( 
.A(n_1245),
.B(n_1256),
.Y(n_2621)
);

NOR2xp67_ASAP7_75t_L g2622 ( 
.A(n_1311),
.B(n_1342),
.Y(n_2622)
);

NOR2xp33_ASAP7_75t_L g2623 ( 
.A(n_1245),
.B(n_1256),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_L g2624 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2624)
);

NAND2xp5_ASAP7_75t_L g2625 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2625)
);

NAND2xp33_ASAP7_75t_L g2626 ( 
.A(n_1378),
.B(n_1342),
.Y(n_2626)
);

INVx2_ASAP7_75t_SL g2627 ( 
.A(n_1275),
.Y(n_2627)
);

NAND2xp5_ASAP7_75t_L g2628 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2628)
);

NOR2x2_ASAP7_75t_L g2629 ( 
.A(n_1263),
.B(n_1025),
.Y(n_2629)
);

NOR3xp33_ASAP7_75t_L g2630 ( 
.A(n_1216),
.B(n_1111),
.C(n_1635),
.Y(n_2630)
);

NOR3x1_ASAP7_75t_L g2631 ( 
.A(n_1461),
.B(n_1111),
.C(n_410),
.Y(n_2631)
);

AOI22xp33_ASAP7_75t_L g2632 ( 
.A1(n_1461),
.A2(n_1118),
.B1(n_1122),
.B2(n_1720),
.Y(n_2632)
);

NAND2xp5_ASAP7_75t_L g2633 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2633)
);

NAND2xp33_ASAP7_75t_L g2634 ( 
.A(n_1378),
.B(n_1342),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_1367),
.Y(n_2635)
);

AOI21xp5_ASAP7_75t_L g2636 ( 
.A1(n_1412),
.A2(n_1321),
.B(n_1394),
.Y(n_2636)
);

INVxp33_ASAP7_75t_L g2637 ( 
.A(n_1213),
.Y(n_2637)
);

NAND3xp33_ASAP7_75t_L g2638 ( 
.A(n_1720),
.B(n_1118),
.C(n_1111),
.Y(n_2638)
);

NAND2xp5_ASAP7_75t_L g2639 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2639)
);

NAND2xp5_ASAP7_75t_SL g2640 ( 
.A(n_1342),
.B(n_1434),
.Y(n_2640)
);

NAND2x1p5_ASAP7_75t_L g2641 ( 
.A(n_1275),
.B(n_1468),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_1367),
.Y(n_2642)
);

AND2x2_ASAP7_75t_L g2643 ( 
.A(n_1380),
.B(n_1405),
.Y(n_2643)
);

A2O1A1Ixp33_ASAP7_75t_L g2644 ( 
.A1(n_1342),
.A2(n_1256),
.B(n_1268),
.C(n_1245),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_L g2645 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2645)
);

BUFx6f_ASAP7_75t_SL g2646 ( 
.A(n_1535),
.Y(n_2646)
);

INVx2_ASAP7_75t_L g2647 ( 
.A(n_1217),
.Y(n_2647)
);

NOR2xp33_ASAP7_75t_L g2648 ( 
.A(n_1245),
.B(n_1256),
.Y(n_2648)
);

INVx1_ASAP7_75t_SL g2649 ( 
.A(n_1679),
.Y(n_2649)
);

NAND2xp5_ASAP7_75t_L g2650 ( 
.A(n_1394),
.B(n_1245),
.Y(n_2650)
);

NOR2xp33_ASAP7_75t_L g2651 ( 
.A(n_1245),
.B(n_1256),
.Y(n_2651)
);

BUFx8_ASAP7_75t_L g2652 ( 
.A(n_1954),
.Y(n_2652)
);

AOI22xp5_ASAP7_75t_L g2653 ( 
.A1(n_2462),
.A2(n_2622),
.B1(n_2615),
.B2(n_2588),
.Y(n_2653)
);

CKINVDCx5p33_ASAP7_75t_R g2654 ( 
.A(n_2570),
.Y(n_2654)
);

NAND2xp5_ASAP7_75t_L g2655 ( 
.A(n_2440),
.B(n_2538),
.Y(n_2655)
);

BUFx3_ASAP7_75t_L g2656 ( 
.A(n_2593),
.Y(n_2656)
);

HB1xp67_ASAP7_75t_L g2657 ( 
.A(n_1989),
.Y(n_2657)
);

INVx2_ASAP7_75t_SL g2658 ( 
.A(n_2252),
.Y(n_2658)
);

BUFx4f_ASAP7_75t_L g2659 ( 
.A(n_2256),
.Y(n_2659)
);

BUFx4f_ASAP7_75t_L g2660 ( 
.A(n_2256),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_1895),
.Y(n_2661)
);

BUFx6f_ASAP7_75t_L g2662 ( 
.A(n_1932),
.Y(n_2662)
);

INVx2_ASAP7_75t_L g2663 ( 
.A(n_1895),
.Y(n_2663)
);

INVx2_ASAP7_75t_L g2664 ( 
.A(n_1906),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_1906),
.Y(n_2665)
);

NAND2xp5_ASAP7_75t_L g2666 ( 
.A(n_2440),
.B(n_2538),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_1907),
.Y(n_2667)
);

NOR2xp33_ASAP7_75t_L g2668 ( 
.A(n_1872),
.B(n_1817),
.Y(n_2668)
);

AOI22xp33_ASAP7_75t_L g2669 ( 
.A1(n_2468),
.A2(n_2528),
.B1(n_2546),
.B2(n_2545),
.Y(n_2669)
);

BUFx8_ASAP7_75t_SL g2670 ( 
.A(n_1891),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_1907),
.Y(n_2671)
);

INVx4_ASAP7_75t_L g2672 ( 
.A(n_2214),
.Y(n_2672)
);

HB1xp67_ASAP7_75t_L g2673 ( 
.A(n_1989),
.Y(n_2673)
);

HB1xp67_ASAP7_75t_L g2674 ( 
.A(n_2090),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_1909),
.Y(n_2675)
);

BUFx6f_ASAP7_75t_L g2676 ( 
.A(n_1932),
.Y(n_2676)
);

BUFx6f_ASAP7_75t_L g2677 ( 
.A(n_1932),
.Y(n_2677)
);

NAND2xp5_ASAP7_75t_L g2678 ( 
.A(n_1847),
.B(n_2474),
.Y(n_2678)
);

BUFx2_ASAP7_75t_L g2679 ( 
.A(n_1946),
.Y(n_2679)
);

BUFx2_ASAP7_75t_L g2680 ( 
.A(n_1946),
.Y(n_2680)
);

NAND2xp5_ASAP7_75t_L g2681 ( 
.A(n_1847),
.B(n_2474),
.Y(n_2681)
);

OR2x4_ASAP7_75t_L g2682 ( 
.A(n_1876),
.B(n_1874),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_1909),
.Y(n_2683)
);

INVx5_ASAP7_75t_L g2684 ( 
.A(n_2256),
.Y(n_2684)
);

INVx1_ASAP7_75t_SL g2685 ( 
.A(n_1950),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_1914),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_1914),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_1919),
.Y(n_2688)
);

NOR2xp33_ASAP7_75t_L g2689 ( 
.A(n_2347),
.B(n_2360),
.Y(n_2689)
);

INVx2_ASAP7_75t_L g2690 ( 
.A(n_1919),
.Y(n_2690)
);

INVx2_ASAP7_75t_L g2691 ( 
.A(n_1935),
.Y(n_2691)
);

BUFx3_ASAP7_75t_L g2692 ( 
.A(n_2593),
.Y(n_2692)
);

INVx2_ASAP7_75t_L g2693 ( 
.A(n_1935),
.Y(n_2693)
);

HB1xp67_ASAP7_75t_L g2694 ( 
.A(n_2090),
.Y(n_2694)
);

INVx2_ASAP7_75t_L g2695 ( 
.A(n_1825),
.Y(n_2695)
);

AOI22xp33_ASAP7_75t_L g2696 ( 
.A1(n_2551),
.A2(n_2609),
.B1(n_2630),
.B2(n_1830),
.Y(n_2696)
);

INVx2_ASAP7_75t_SL g2697 ( 
.A(n_2252),
.Y(n_2697)
);

INVx2_ASAP7_75t_SL g2698 ( 
.A(n_1982),
.Y(n_2698)
);

A2O1A1Ixp33_ASAP7_75t_L g2699 ( 
.A1(n_1922),
.A2(n_2397),
.B(n_2644),
.C(n_1897),
.Y(n_2699)
);

NAND2xp5_ASAP7_75t_L g2700 ( 
.A(n_2520),
.B(n_2636),
.Y(n_2700)
);

AOI22xp33_ASAP7_75t_L g2701 ( 
.A1(n_1830),
.A2(n_2588),
.B1(n_2435),
.B2(n_2529),
.Y(n_2701)
);

INVx2_ASAP7_75t_L g2702 ( 
.A(n_1825),
.Y(n_2702)
);

INVx2_ASAP7_75t_L g2703 ( 
.A(n_1825),
.Y(n_2703)
);

OR2x2_ASAP7_75t_L g2704 ( 
.A(n_1941),
.B(n_1951),
.Y(n_2704)
);

NAND2xp5_ASAP7_75t_SL g2705 ( 
.A(n_2351),
.B(n_2361),
.Y(n_2705)
);

NAND2xp5_ASAP7_75t_L g2706 ( 
.A(n_2520),
.B(n_2616),
.Y(n_2706)
);

AOI22xp5_ASAP7_75t_L g2707 ( 
.A1(n_2462),
.A2(n_2622),
.B1(n_2615),
.B2(n_2435),
.Y(n_2707)
);

BUFx4f_ASAP7_75t_L g2708 ( 
.A(n_2256),
.Y(n_2708)
);

OR2x2_ASAP7_75t_L g2709 ( 
.A(n_1941),
.B(n_1958),
.Y(n_2709)
);

NAND2xp5_ASAP7_75t_L g2710 ( 
.A(n_2616),
.B(n_2636),
.Y(n_2710)
);

AND2x6_ASAP7_75t_SL g2711 ( 
.A(n_2404),
.B(n_2423),
.Y(n_2711)
);

BUFx6f_ASAP7_75t_L g2712 ( 
.A(n_1982),
.Y(n_2712)
);

AND3x1_ASAP7_75t_SL g2713 ( 
.A(n_2529),
.B(n_2596),
.C(n_2515),
.Y(n_2713)
);

AND2x4_ASAP7_75t_L g2714 ( 
.A(n_2483),
.B(n_1910),
.Y(n_2714)
);

NAND2xp5_ASAP7_75t_SL g2715 ( 
.A(n_2351),
.B(n_2361),
.Y(n_2715)
);

AOI22xp5_ASAP7_75t_L g2716 ( 
.A1(n_2349),
.A2(n_2579),
.B1(n_2626),
.B2(n_2541),
.Y(n_2716)
);

CKINVDCx5p33_ASAP7_75t_R g2717 ( 
.A(n_2433),
.Y(n_2717)
);

BUFx6f_ASAP7_75t_L g2718 ( 
.A(n_2061),
.Y(n_2718)
);

NOR2xp33_ASAP7_75t_L g2719 ( 
.A(n_2442),
.B(n_2451),
.Y(n_2719)
);

NAND2xp5_ASAP7_75t_SL g2720 ( 
.A(n_2379),
.B(n_2395),
.Y(n_2720)
);

CKINVDCx5p33_ASAP7_75t_R g2721 ( 
.A(n_2436),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_L g2722 ( 
.A(n_1897),
.B(n_1869),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_1959),
.Y(n_2723)
);

AND2x4_ASAP7_75t_L g2724 ( 
.A(n_2483),
.B(n_1910),
.Y(n_2724)
);

INVx2_ASAP7_75t_L g2725 ( 
.A(n_1839),
.Y(n_2725)
);

INVx2_ASAP7_75t_L g2726 ( 
.A(n_1850),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_L g2727 ( 
.A(n_1869),
.B(n_1853),
.Y(n_2727)
);

INVx1_ASAP7_75t_SL g2728 ( 
.A(n_1950),
.Y(n_2728)
);

INVx2_ASAP7_75t_SL g2729 ( 
.A(n_2088),
.Y(n_2729)
);

AO21x2_ASAP7_75t_L g2730 ( 
.A1(n_1893),
.A2(n_1894),
.B(n_1858),
.Y(n_2730)
);

AND2x2_ASAP7_75t_L g2731 ( 
.A(n_1869),
.B(n_1921),
.Y(n_2731)
);

AND3x1_ASAP7_75t_SL g2732 ( 
.A(n_2596),
.B(n_2515),
.C(n_2599),
.Y(n_2732)
);

AOI22xp5_ASAP7_75t_L g2733 ( 
.A1(n_2634),
.A2(n_2379),
.B1(n_2396),
.B2(n_2395),
.Y(n_2733)
);

INVx3_ASAP7_75t_L g2734 ( 
.A(n_2061),
.Y(n_2734)
);

NAND2xp5_ASAP7_75t_L g2735 ( 
.A(n_1840),
.B(n_1915),
.Y(n_2735)
);

INVx2_ASAP7_75t_L g2736 ( 
.A(n_1850),
.Y(n_2736)
);

NAND2xp5_ASAP7_75t_L g2737 ( 
.A(n_2645),
.B(n_2650),
.Y(n_2737)
);

O2A1O1Ixp33_ASAP7_75t_L g2738 ( 
.A1(n_1828),
.A2(n_1893),
.B(n_1894),
.C(n_1833),
.Y(n_2738)
);

AOI22xp5_ASAP7_75t_L g2739 ( 
.A1(n_2396),
.A2(n_2415),
.B1(n_2444),
.B2(n_2407),
.Y(n_2739)
);

INVx2_ASAP7_75t_SL g2740 ( 
.A(n_2088),
.Y(n_2740)
);

BUFx2_ASAP7_75t_L g2741 ( 
.A(n_1961),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_1961),
.Y(n_2742)
);

INVx2_ASAP7_75t_L g2743 ( 
.A(n_1850),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_1963),
.Y(n_2744)
);

BUFx3_ASAP7_75t_L g2745 ( 
.A(n_2593),
.Y(n_2745)
);

BUFx2_ASAP7_75t_L g2746 ( 
.A(n_1963),
.Y(n_2746)
);

NOR2x1p5_ASAP7_75t_L g2747 ( 
.A(n_2586),
.B(n_1874),
.Y(n_2747)
);

BUFx4f_ASAP7_75t_L g2748 ( 
.A(n_2256),
.Y(n_2748)
);

NOR2xp33_ASAP7_75t_R g2749 ( 
.A(n_2517),
.B(n_2523),
.Y(n_2749)
);

INVx2_ASAP7_75t_L g2750 ( 
.A(n_1867),
.Y(n_2750)
);

INVx5_ASAP7_75t_L g2751 ( 
.A(n_1949),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_L g2752 ( 
.A(n_2639),
.B(n_2645),
.Y(n_2752)
);

CKINVDCx20_ASAP7_75t_R g2753 ( 
.A(n_1887),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_1964),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_1964),
.Y(n_2755)
);

BUFx8_ASAP7_75t_L g2756 ( 
.A(n_1954),
.Y(n_2756)
);

AO22x1_ASAP7_75t_L g2757 ( 
.A1(n_1832),
.A2(n_2527),
.B1(n_2631),
.B2(n_2456),
.Y(n_2757)
);

INVxp67_ASAP7_75t_L g2758 ( 
.A(n_1871),
.Y(n_2758)
);

INVx2_ASAP7_75t_SL g2759 ( 
.A(n_2586),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_L g2760 ( 
.A(n_2650),
.B(n_1821),
.Y(n_2760)
);

INVx2_ASAP7_75t_L g2761 ( 
.A(n_1867),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_1821),
.B(n_1822),
.Y(n_2762)
);

AOI21xp5_ASAP7_75t_L g2763 ( 
.A1(n_1871),
.A2(n_1875),
.B(n_1879),
.Y(n_2763)
);

AND2x4_ASAP7_75t_L g2764 ( 
.A(n_2483),
.B(n_1910),
.Y(n_2764)
);

NOR2xp33_ASAP7_75t_L g2765 ( 
.A(n_2504),
.B(n_2525),
.Y(n_2765)
);

AND3x1_ASAP7_75t_L g2766 ( 
.A(n_2446),
.B(n_2415),
.C(n_2407),
.Y(n_2766)
);

A2O1A1Ixp33_ASAP7_75t_L g2767 ( 
.A1(n_1833),
.A2(n_2478),
.B(n_2510),
.C(n_2444),
.Y(n_2767)
);

BUFx3_ASAP7_75t_L g2768 ( 
.A(n_2593),
.Y(n_2768)
);

BUFx6f_ASAP7_75t_L g2769 ( 
.A(n_2593),
.Y(n_2769)
);

NAND2xp5_ASAP7_75t_L g2770 ( 
.A(n_2639),
.B(n_1822),
.Y(n_2770)
);

AOI22xp33_ASAP7_75t_L g2771 ( 
.A1(n_2567),
.A2(n_2592),
.B1(n_2600),
.B2(n_2571),
.Y(n_2771)
);

CKINVDCx5p33_ASAP7_75t_R g2772 ( 
.A(n_1864),
.Y(n_2772)
);

AOI22xp5_ASAP7_75t_L g2773 ( 
.A1(n_2510),
.A2(n_2558),
.B1(n_2561),
.B2(n_2536),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_1972),
.Y(n_2774)
);

NAND3xp33_ASAP7_75t_L g2775 ( 
.A(n_2445),
.B(n_2638),
.C(n_2496),
.Y(n_2775)
);

INVx2_ASAP7_75t_SL g2776 ( 
.A(n_2214),
.Y(n_2776)
);

INVx1_ASAP7_75t_L g2777 ( 
.A(n_1972),
.Y(n_2777)
);

NAND2xp5_ASAP7_75t_L g2778 ( 
.A(n_2352),
.B(n_2354),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_1973),
.Y(n_2779)
);

BUFx3_ASAP7_75t_L g2780 ( 
.A(n_2593),
.Y(n_2780)
);

BUFx6f_ASAP7_75t_L g2781 ( 
.A(n_2593),
.Y(n_2781)
);

CKINVDCx5p33_ASAP7_75t_R g2782 ( 
.A(n_1864),
.Y(n_2782)
);

BUFx6f_ASAP7_75t_L g2783 ( 
.A(n_2593),
.Y(n_2783)
);

BUFx12f_ASAP7_75t_L g2784 ( 
.A(n_1881),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_1973),
.Y(n_2785)
);

OR2x2_ASAP7_75t_L g2786 ( 
.A(n_1974),
.B(n_1985),
.Y(n_2786)
);

AOI21xp5_ASAP7_75t_L g2787 ( 
.A1(n_1875),
.A2(n_1879),
.B(n_1884),
.Y(n_2787)
);

INVx4_ASAP7_75t_L g2788 ( 
.A(n_2214),
.Y(n_2788)
);

BUFx2_ASAP7_75t_L g2789 ( 
.A(n_2483),
.Y(n_2789)
);

BUFx3_ASAP7_75t_L g2790 ( 
.A(n_2483),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_1974),
.Y(n_2791)
);

INVx3_ASAP7_75t_L g2792 ( 
.A(n_2214),
.Y(n_2792)
);

AND2x4_ASAP7_75t_L g2793 ( 
.A(n_1910),
.B(n_1970),
.Y(n_2793)
);

BUFx3_ASAP7_75t_L g2794 ( 
.A(n_2214),
.Y(n_2794)
);

NAND2xp5_ASAP7_75t_SL g2795 ( 
.A(n_2536),
.B(n_2558),
.Y(n_2795)
);

NAND2xp5_ASAP7_75t_L g2796 ( 
.A(n_2352),
.B(n_2354),
.Y(n_2796)
);

AND2x4_ASAP7_75t_L g2797 ( 
.A(n_1910),
.B(n_1970),
.Y(n_2797)
);

BUFx3_ASAP7_75t_L g2798 ( 
.A(n_2214),
.Y(n_2798)
);

INVx2_ASAP7_75t_L g2799 ( 
.A(n_1885),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_1985),
.Y(n_2800)
);

INVx1_ASAP7_75t_SL g2801 ( 
.A(n_1948),
.Y(n_2801)
);

INVx2_ASAP7_75t_L g2802 ( 
.A(n_1885),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_1996),
.Y(n_2803)
);

NOR2xp33_ASAP7_75t_L g2804 ( 
.A(n_2608),
.B(n_2621),
.Y(n_2804)
);

BUFx3_ASAP7_75t_L g2805 ( 
.A(n_2214),
.Y(n_2805)
);

NAND2xp5_ASAP7_75t_L g2806 ( 
.A(n_2356),
.B(n_2633),
.Y(n_2806)
);

AO22x1_ASAP7_75t_L g2807 ( 
.A1(n_1832),
.A2(n_2631),
.B1(n_2648),
.B2(n_2623),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_SL g2808 ( 
.A(n_2561),
.B(n_2578),
.Y(n_2808)
);

NOR2x1_ASAP7_75t_R g2809 ( 
.A(n_1891),
.B(n_2406),
.Y(n_2809)
);

NAND2xp5_ASAP7_75t_L g2810 ( 
.A(n_2356),
.B(n_2364),
.Y(n_2810)
);

HB1xp67_ASAP7_75t_L g2811 ( 
.A(n_1955),
.Y(n_2811)
);

BUFx3_ASAP7_75t_L g2812 ( 
.A(n_2214),
.Y(n_2812)
);

BUFx6f_ASAP7_75t_L g2813 ( 
.A(n_2208),
.Y(n_2813)
);

INVx2_ASAP7_75t_SL g2814 ( 
.A(n_2214),
.Y(n_2814)
);

AOI22xp5_ASAP7_75t_L g2815 ( 
.A1(n_2578),
.A2(n_2619),
.B1(n_1866),
.B2(n_1889),
.Y(n_2815)
);

BUFx2_ASAP7_75t_L g2816 ( 
.A(n_1999),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_1996),
.Y(n_2817)
);

AOI22xp33_ASAP7_75t_L g2818 ( 
.A1(n_2651),
.A2(n_1866),
.B1(n_2619),
.B2(n_1858),
.Y(n_2818)
);

NAND2xp5_ASAP7_75t_L g2819 ( 
.A(n_2364),
.B(n_2369),
.Y(n_2819)
);

AOI22xp5_ASAP7_75t_SL g2820 ( 
.A1(n_2532),
.A2(n_1988),
.B1(n_1962),
.B2(n_1826),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_1943),
.Y(n_2821)
);

BUFx3_ASAP7_75t_L g2822 ( 
.A(n_2214),
.Y(n_2822)
);

BUFx6f_ASAP7_75t_L g2823 ( 
.A(n_2208),
.Y(n_2823)
);

INVx2_ASAP7_75t_SL g2824 ( 
.A(n_2221),
.Y(n_2824)
);

AOI22xp33_ASAP7_75t_L g2825 ( 
.A1(n_2445),
.A2(n_2496),
.B1(n_2638),
.B2(n_2632),
.Y(n_2825)
);

INVxp67_ASAP7_75t_L g2826 ( 
.A(n_1948),
.Y(n_2826)
);

INVx2_ASAP7_75t_L g2827 ( 
.A(n_1917),
.Y(n_2827)
);

NAND2xp5_ASAP7_75t_L g2828 ( 
.A(n_2369),
.B(n_2372),
.Y(n_2828)
);

INVx2_ASAP7_75t_L g2829 ( 
.A(n_1917),
.Y(n_2829)
);

INVx2_ASAP7_75t_L g2830 ( 
.A(n_1917),
.Y(n_2830)
);

INVx2_ASAP7_75t_SL g2831 ( 
.A(n_2221),
.Y(n_2831)
);

INVx2_ASAP7_75t_L g2832 ( 
.A(n_1920),
.Y(n_2832)
);

AND2x2_ASAP7_75t_L g2833 ( 
.A(n_1936),
.B(n_1939),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_1943),
.Y(n_2834)
);

AND2x2_ASAP7_75t_L g2835 ( 
.A(n_1936),
.B(n_1939),
.Y(n_2835)
);

AND2x4_ASAP7_75t_L g2836 ( 
.A(n_1892),
.B(n_1902),
.Y(n_2836)
);

NAND2xp5_ASAP7_75t_L g2837 ( 
.A(n_2372),
.B(n_2374),
.Y(n_2837)
);

INVx2_ASAP7_75t_L g2838 ( 
.A(n_1920),
.Y(n_2838)
);

NAND2xp5_ASAP7_75t_L g2839 ( 
.A(n_2374),
.B(n_2378),
.Y(n_2839)
);

INVx3_ASAP7_75t_L g2840 ( 
.A(n_2221),
.Y(n_2840)
);

NAND2x1p5_ASAP7_75t_L g2841 ( 
.A(n_2192),
.B(n_2207),
.Y(n_2841)
);

AND2x4_ASAP7_75t_L g2842 ( 
.A(n_1892),
.B(n_1902),
.Y(n_2842)
);

INVx2_ASAP7_75t_L g2843 ( 
.A(n_1920),
.Y(n_2843)
);

NAND2xp5_ASAP7_75t_L g2844 ( 
.A(n_2378),
.B(n_2380),
.Y(n_2844)
);

BUFx2_ASAP7_75t_L g2845 ( 
.A(n_1999),
.Y(n_2845)
);

INVx2_ASAP7_75t_L g2846 ( 
.A(n_1923),
.Y(n_2846)
);

AND2x4_ASAP7_75t_L g2847 ( 
.A(n_1892),
.B(n_1902),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_1947),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_1947),
.Y(n_2849)
);

INVx2_ASAP7_75t_L g2850 ( 
.A(n_1923),
.Y(n_2850)
);

NAND2xp5_ASAP7_75t_L g2851 ( 
.A(n_2625),
.B(n_2628),
.Y(n_2851)
);

INVx2_ASAP7_75t_L g2852 ( 
.A(n_1923),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2001),
.Y(n_2853)
);

BUFx12f_ASAP7_75t_L g2854 ( 
.A(n_2279),
.Y(n_2854)
);

INVx3_ASAP7_75t_L g2855 ( 
.A(n_2221),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_L g2856 ( 
.A(n_2628),
.B(n_2633),
.Y(n_2856)
);

HB1xp67_ASAP7_75t_L g2857 ( 
.A(n_2188),
.Y(n_2857)
);

INVx2_ASAP7_75t_L g2858 ( 
.A(n_1926),
.Y(n_2858)
);

INVx4_ASAP7_75t_L g2859 ( 
.A(n_1949),
.Y(n_2859)
);

NOR2xp33_ASAP7_75t_L g2860 ( 
.A(n_1836),
.B(n_1841),
.Y(n_2860)
);

HB1xp67_ASAP7_75t_L g2861 ( 
.A(n_2188),
.Y(n_2861)
);

AND2x4_ASAP7_75t_L g2862 ( 
.A(n_1892),
.B(n_1902),
.Y(n_2862)
);

INVx2_ASAP7_75t_L g2863 ( 
.A(n_1926),
.Y(n_2863)
);

NAND2xp5_ASAP7_75t_SL g2864 ( 
.A(n_1846),
.B(n_2380),
.Y(n_2864)
);

INVx2_ASAP7_75t_SL g2865 ( 
.A(n_2232),
.Y(n_2865)
);

NAND2xp5_ASAP7_75t_L g2866 ( 
.A(n_2392),
.B(n_2394),
.Y(n_2866)
);

INVxp33_ASAP7_75t_L g2867 ( 
.A(n_1883),
.Y(n_2867)
);

NAND2xp5_ASAP7_75t_SL g2868 ( 
.A(n_1846),
.B(n_2392),
.Y(n_2868)
);

BUFx6f_ASAP7_75t_L g2869 ( 
.A(n_2210),
.Y(n_2869)
);

OR2x2_ASAP7_75t_L g2870 ( 
.A(n_1862),
.B(n_2001),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2189),
.Y(n_2871)
);

INVx2_ASAP7_75t_SL g2872 ( 
.A(n_2232),
.Y(n_2872)
);

INVx1_ASAP7_75t_L g2873 ( 
.A(n_2189),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_L g2874 ( 
.A(n_2394),
.B(n_2403),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_1926),
.Y(n_2875)
);

INVx6_ASAP7_75t_L g2876 ( 
.A(n_1904),
.Y(n_2876)
);

NOR2xp33_ASAP7_75t_L g2877 ( 
.A(n_1836),
.B(n_1841),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_1957),
.Y(n_2878)
);

HB1xp67_ASAP7_75t_L g2879 ( 
.A(n_2050),
.Y(n_2879)
);

INVxp67_ASAP7_75t_L g2880 ( 
.A(n_1940),
.Y(n_2880)
);

INVx5_ASAP7_75t_L g2881 ( 
.A(n_1949),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_L g2882 ( 
.A(n_2625),
.B(n_2403),
.Y(n_2882)
);

INVx2_ASAP7_75t_L g2883 ( 
.A(n_1957),
.Y(n_2883)
);

HB1xp67_ASAP7_75t_L g2884 ( 
.A(n_2050),
.Y(n_2884)
);

AND2x4_ASAP7_75t_L g2885 ( 
.A(n_1924),
.B(n_2387),
.Y(n_2885)
);

BUFx3_ASAP7_75t_L g2886 ( 
.A(n_2311),
.Y(n_2886)
);

INVx2_ASAP7_75t_L g2887 ( 
.A(n_2000),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2414),
.B(n_2418),
.Y(n_2888)
);

INVx3_ASAP7_75t_L g2889 ( 
.A(n_1835),
.Y(n_2889)
);

AOI22xp33_ASAP7_75t_L g2890 ( 
.A1(n_2355),
.A2(n_2375),
.B1(n_2413),
.B2(n_2381),
.Y(n_2890)
);

BUFx2_ASAP7_75t_L g2891 ( 
.A(n_2002),
.Y(n_2891)
);

NAND2xp5_ASAP7_75t_SL g2892 ( 
.A(n_2414),
.B(n_2418),
.Y(n_2892)
);

INVx2_ASAP7_75t_L g2893 ( 
.A(n_2000),
.Y(n_2893)
);

HB1xp67_ASAP7_75t_L g2894 ( 
.A(n_1940),
.Y(n_2894)
);

NAND2xp5_ASAP7_75t_L g2895 ( 
.A(n_2424),
.B(n_2425),
.Y(n_2895)
);

AOI22xp33_ASAP7_75t_L g2896 ( 
.A1(n_2428),
.A2(n_2438),
.B1(n_2584),
.B2(n_2563),
.Y(n_2896)
);

BUFx3_ASAP7_75t_L g2897 ( 
.A(n_2311),
.Y(n_2897)
);

BUFx2_ASAP7_75t_L g2898 ( 
.A(n_2002),
.Y(n_2898)
);

NAND2xp5_ASAP7_75t_L g2899 ( 
.A(n_2424),
.B(n_2425),
.Y(n_2899)
);

INVx2_ASAP7_75t_L g2900 ( 
.A(n_2014),
.Y(n_2900)
);

BUFx6f_ASAP7_75t_L g2901 ( 
.A(n_2210),
.Y(n_2901)
);

BUFx2_ASAP7_75t_L g2902 ( 
.A(n_1997),
.Y(n_2902)
);

INVx5_ASAP7_75t_L g2903 ( 
.A(n_1949),
.Y(n_2903)
);

INVx2_ASAP7_75t_SL g2904 ( 
.A(n_1944),
.Y(n_2904)
);

BUFx6f_ASAP7_75t_L g2905 ( 
.A(n_2222),
.Y(n_2905)
);

NAND2xp5_ASAP7_75t_L g2906 ( 
.A(n_2430),
.B(n_2431),
.Y(n_2906)
);

AOI22xp33_ASAP7_75t_L g2907 ( 
.A1(n_2617),
.A2(n_1862),
.B1(n_2553),
.B2(n_2503),
.Y(n_2907)
);

INVx3_ASAP7_75t_L g2908 ( 
.A(n_1835),
.Y(n_2908)
);

BUFx3_ASAP7_75t_L g2909 ( 
.A(n_2311),
.Y(n_2909)
);

NAND2xp5_ASAP7_75t_SL g2910 ( 
.A(n_2430),
.B(n_2431),
.Y(n_2910)
);

OR2x2_ASAP7_75t_SL g2911 ( 
.A(n_2350),
.B(n_2410),
.Y(n_2911)
);

BUFx2_ASAP7_75t_L g2912 ( 
.A(n_1997),
.Y(n_2912)
);

AND2x4_ASAP7_75t_L g2913 ( 
.A(n_1924),
.B(n_2387),
.Y(n_2913)
);

INVx2_ASAP7_75t_SL g2914 ( 
.A(n_1944),
.Y(n_2914)
);

INVx4_ASAP7_75t_L g2915 ( 
.A(n_1949),
.Y(n_2915)
);

INVx3_ASAP7_75t_L g2916 ( 
.A(n_1835),
.Y(n_2916)
);

BUFx6f_ASAP7_75t_L g2917 ( 
.A(n_2222),
.Y(n_2917)
);

CKINVDCx5p33_ASAP7_75t_R g2918 ( 
.A(n_1891),
.Y(n_2918)
);

HB1xp67_ASAP7_75t_L g2919 ( 
.A(n_1986),
.Y(n_2919)
);

INVx2_ASAP7_75t_L g2920 ( 
.A(n_2027),
.Y(n_2920)
);

INVx5_ASAP7_75t_L g2921 ( 
.A(n_1992),
.Y(n_2921)
);

AND2x4_ASAP7_75t_L g2922 ( 
.A(n_1924),
.B(n_2387),
.Y(n_2922)
);

NOR2xp33_ASAP7_75t_L g2923 ( 
.A(n_1823),
.B(n_1826),
.Y(n_2923)
);

INVx1_ASAP7_75t_SL g2924 ( 
.A(n_2350),
.Y(n_2924)
);

INVx1_ASAP7_75t_SL g2925 ( 
.A(n_2410),
.Y(n_2925)
);

INVx2_ASAP7_75t_L g2926 ( 
.A(n_2052),
.Y(n_2926)
);

INVx4_ASAP7_75t_L g2927 ( 
.A(n_1992),
.Y(n_2927)
);

BUFx3_ASAP7_75t_L g2928 ( 
.A(n_1971),
.Y(n_2928)
);

CKINVDCx5p33_ASAP7_75t_R g2929 ( 
.A(n_2406),
.Y(n_2929)
);

INVx2_ASAP7_75t_L g2930 ( 
.A(n_2054),
.Y(n_2930)
);

AOI22xp5_ASAP7_75t_L g2931 ( 
.A1(n_1889),
.A2(n_1912),
.B1(n_1863),
.B2(n_1831),
.Y(n_2931)
);

INVx3_ASAP7_75t_L g2932 ( 
.A(n_1835),
.Y(n_2932)
);

INVx1_ASAP7_75t_SL g2933 ( 
.A(n_2417),
.Y(n_2933)
);

BUFx2_ASAP7_75t_L g2934 ( 
.A(n_2046),
.Y(n_2934)
);

NAND3xp33_ASAP7_75t_SL g2935 ( 
.A(n_2401),
.B(n_2478),
.C(n_2358),
.Y(n_2935)
);

AND2x6_ASAP7_75t_SL g2936 ( 
.A(n_2618),
.B(n_2620),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_L g2937 ( 
.A(n_2618),
.B(n_2620),
.Y(n_2937)
);

AND2x4_ASAP7_75t_L g2938 ( 
.A(n_1924),
.B(n_2387),
.Y(n_2938)
);

O2A1O1Ixp33_ASAP7_75t_L g2939 ( 
.A1(n_2432),
.A2(n_2443),
.B(n_2447),
.C(n_2439),
.Y(n_2939)
);

INVx2_ASAP7_75t_SL g2940 ( 
.A(n_1944),
.Y(n_2940)
);

AOI22xp5_ASAP7_75t_L g2941 ( 
.A1(n_2532),
.A2(n_1820),
.B1(n_2376),
.B2(n_2359),
.Y(n_2941)
);

AOI22xp5_ASAP7_75t_L g2942 ( 
.A1(n_2532),
.A2(n_2382),
.B1(n_2388),
.B2(n_2384),
.Y(n_2942)
);

INVx4_ASAP7_75t_L g2943 ( 
.A(n_1992),
.Y(n_2943)
);

AOI22xp33_ASAP7_75t_L g2944 ( 
.A1(n_2469),
.A2(n_2556),
.B1(n_2399),
.B2(n_2408),
.Y(n_2944)
);

AND2x4_ASAP7_75t_L g2945 ( 
.A(n_2426),
.B(n_2453),
.Y(n_2945)
);

NAND2xp5_ASAP7_75t_L g2946 ( 
.A(n_2624),
.B(n_2432),
.Y(n_2946)
);

CKINVDCx20_ASAP7_75t_R g2947 ( 
.A(n_2434),
.Y(n_2947)
);

INVx5_ASAP7_75t_L g2948 ( 
.A(n_1992),
.Y(n_2948)
);

INVx2_ASAP7_75t_L g2949 ( 
.A(n_2107),
.Y(n_2949)
);

NAND2xp5_ASAP7_75t_L g2950 ( 
.A(n_2439),
.B(n_2443),
.Y(n_2950)
);

BUFx6f_ASAP7_75t_L g2951 ( 
.A(n_2228),
.Y(n_2951)
);

INVx1_ASAP7_75t_SL g2952 ( 
.A(n_2417),
.Y(n_2952)
);

NAND2xp5_ASAP7_75t_L g2953 ( 
.A(n_2447),
.B(n_2448),
.Y(n_2953)
);

INVx2_ASAP7_75t_SL g2954 ( 
.A(n_2075),
.Y(n_2954)
);

BUFx2_ASAP7_75t_L g2955 ( 
.A(n_2046),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_L g2956 ( 
.A(n_2448),
.B(n_2450),
.Y(n_2956)
);

INVx2_ASAP7_75t_SL g2957 ( 
.A(n_2075),
.Y(n_2957)
);

INVx2_ASAP7_75t_L g2958 ( 
.A(n_2131),
.Y(n_2958)
);

OAI22xp33_ASAP7_75t_L g2959 ( 
.A1(n_1823),
.A2(n_1834),
.B1(n_1838),
.B2(n_1829),
.Y(n_2959)
);

AOI22xp5_ASAP7_75t_L g2960 ( 
.A1(n_2389),
.A2(n_2421),
.B1(n_2477),
.B2(n_2427),
.Y(n_2960)
);

INVx5_ASAP7_75t_L g2961 ( 
.A(n_1992),
.Y(n_2961)
);

NAND2xp5_ASAP7_75t_L g2962 ( 
.A(n_2450),
.B(n_2452),
.Y(n_2962)
);

AOI22xp33_ASAP7_75t_L g2963 ( 
.A1(n_2530),
.A2(n_2549),
.B1(n_2557),
.B2(n_2491),
.Y(n_2963)
);

BUFx8_ASAP7_75t_L g2964 ( 
.A(n_1954),
.Y(n_2964)
);

BUFx5_ASAP7_75t_L g2965 ( 
.A(n_1878),
.Y(n_2965)
);

INVx3_ASAP7_75t_L g2966 ( 
.A(n_1835),
.Y(n_2966)
);

INVx2_ASAP7_75t_L g2967 ( 
.A(n_2149),
.Y(n_2967)
);

NOR2xp67_ASAP7_75t_L g2968 ( 
.A(n_2146),
.B(n_2192),
.Y(n_2968)
);

INVx2_ASAP7_75t_SL g2969 ( 
.A(n_2075),
.Y(n_2969)
);

AND2x4_ASAP7_75t_L g2970 ( 
.A(n_2426),
.B(n_2453),
.Y(n_2970)
);

AND2x2_ASAP7_75t_SL g2971 ( 
.A(n_2207),
.B(n_2010),
.Y(n_2971)
);

NAND2xp5_ASAP7_75t_L g2972 ( 
.A(n_2452),
.B(n_2454),
.Y(n_2972)
);

AND2x4_ASAP7_75t_L g2973 ( 
.A(n_2426),
.B(n_2453),
.Y(n_2973)
);

AND2x4_ASAP7_75t_L g2974 ( 
.A(n_2426),
.B(n_2453),
.Y(n_2974)
);

INVx4_ASAP7_75t_L g2975 ( 
.A(n_2057),
.Y(n_2975)
);

BUFx3_ASAP7_75t_L g2976 ( 
.A(n_1971),
.Y(n_2976)
);

INVx3_ASAP7_75t_L g2977 ( 
.A(n_1835),
.Y(n_2977)
);

NAND2xp5_ASAP7_75t_L g2978 ( 
.A(n_2454),
.B(n_2455),
.Y(n_2978)
);

BUFx6f_ASAP7_75t_L g2979 ( 
.A(n_2228),
.Y(n_2979)
);

AND2x6_ASAP7_75t_L g2980 ( 
.A(n_2548),
.B(n_2587),
.Y(n_2980)
);

AND3x2_ASAP7_75t_SL g2981 ( 
.A(n_1988),
.B(n_1977),
.C(n_1942),
.Y(n_2981)
);

INVx5_ASAP7_75t_L g2982 ( 
.A(n_2057),
.Y(n_2982)
);

BUFx3_ASAP7_75t_L g2983 ( 
.A(n_2062),
.Y(n_2983)
);

CKINVDCx5p33_ASAP7_75t_R g2984 ( 
.A(n_2406),
.Y(n_2984)
);

NAND2xp5_ASAP7_75t_L g2985 ( 
.A(n_2455),
.B(n_2459),
.Y(n_2985)
);

BUFx12f_ASAP7_75t_L g2986 ( 
.A(n_2279),
.Y(n_2986)
);

NAND2xp5_ASAP7_75t_L g2987 ( 
.A(n_2459),
.B(n_2460),
.Y(n_2987)
);

INVx2_ASAP7_75t_SL g2988 ( 
.A(n_2159),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_L g2989 ( 
.A(n_2460),
.B(n_2463),
.Y(n_2989)
);

BUFx2_ASAP7_75t_L g2990 ( 
.A(n_2062),
.Y(n_2990)
);

NAND2xp5_ASAP7_75t_L g2991 ( 
.A(n_2624),
.B(n_2463),
.Y(n_2991)
);

BUFx3_ASAP7_75t_L g2992 ( 
.A(n_2057),
.Y(n_2992)
);

INVx1_ASAP7_75t_SL g2993 ( 
.A(n_2495),
.Y(n_2993)
);

NAND2xp5_ASAP7_75t_SL g2994 ( 
.A(n_2464),
.B(n_2465),
.Y(n_2994)
);

INVx3_ASAP7_75t_L g2995 ( 
.A(n_2094),
.Y(n_2995)
);

NAND2xp5_ASAP7_75t_L g2996 ( 
.A(n_2464),
.B(n_2465),
.Y(n_2996)
);

NOR2xp33_ASAP7_75t_L g2997 ( 
.A(n_1829),
.B(n_1834),
.Y(n_2997)
);

OR2x2_ASAP7_75t_L g2998 ( 
.A(n_1942),
.B(n_2495),
.Y(n_2998)
);

CKINVDCx5p33_ASAP7_75t_R g2999 ( 
.A(n_2087),
.Y(n_2999)
);

NAND2xp5_ASAP7_75t_L g3000 ( 
.A(n_2466),
.B(n_2467),
.Y(n_3000)
);

BUFx2_ASAP7_75t_L g3001 ( 
.A(n_2005),
.Y(n_3001)
);

INVx2_ASAP7_75t_SL g3002 ( 
.A(n_2159),
.Y(n_3002)
);

BUFx6f_ASAP7_75t_L g3003 ( 
.A(n_2057),
.Y(n_3003)
);

INVx2_ASAP7_75t_L g3004 ( 
.A(n_2180),
.Y(n_3004)
);

BUFx3_ASAP7_75t_L g3005 ( 
.A(n_2057),
.Y(n_3005)
);

INVx2_ASAP7_75t_L g3006 ( 
.A(n_2180),
.Y(n_3006)
);

INVx2_ASAP7_75t_SL g3007 ( 
.A(n_2159),
.Y(n_3007)
);

OAI22xp5_ASAP7_75t_L g3008 ( 
.A1(n_2466),
.A2(n_2470),
.B1(n_2479),
.B2(n_2467),
.Y(n_3008)
);

AND2x4_ASAP7_75t_L g3009 ( 
.A(n_2548),
.B(n_2587),
.Y(n_3009)
);

CKINVDCx5p33_ASAP7_75t_R g3010 ( 
.A(n_2199),
.Y(n_3010)
);

NAND2xp5_ASAP7_75t_SL g3011 ( 
.A(n_2470),
.B(n_2479),
.Y(n_3011)
);

OR2x2_ASAP7_75t_L g3012 ( 
.A(n_2486),
.B(n_2488),
.Y(n_3012)
);

BUFx6f_ASAP7_75t_SL g3013 ( 
.A(n_2548),
.Y(n_3013)
);

AND2x4_ASAP7_75t_L g3014 ( 
.A(n_2548),
.B(n_2587),
.Y(n_3014)
);

CKINVDCx5p33_ASAP7_75t_R g3015 ( 
.A(n_1898),
.Y(n_3015)
);

INVxp67_ASAP7_75t_L g3016 ( 
.A(n_1933),
.Y(n_3016)
);

BUFx3_ASAP7_75t_L g3017 ( 
.A(n_2118),
.Y(n_3017)
);

AND2x4_ASAP7_75t_L g3018 ( 
.A(n_2587),
.B(n_2072),
.Y(n_3018)
);

INVxp67_ASAP7_75t_SL g3019 ( 
.A(n_2060),
.Y(n_3019)
);

INVx2_ASAP7_75t_L g3020 ( 
.A(n_2353),
.Y(n_3020)
);

BUFx6f_ASAP7_75t_L g3021 ( 
.A(n_2118),
.Y(n_3021)
);

INVx2_ASAP7_75t_L g3022 ( 
.A(n_2363),
.Y(n_3022)
);

BUFx3_ASAP7_75t_L g3023 ( 
.A(n_2118),
.Y(n_3023)
);

INVx2_ASAP7_75t_L g3024 ( 
.A(n_2368),
.Y(n_3024)
);

CKINVDCx14_ASAP7_75t_R g3025 ( 
.A(n_2233),
.Y(n_3025)
);

INVx3_ASAP7_75t_L g3026 ( 
.A(n_2094),
.Y(n_3026)
);

NAND2xp5_ASAP7_75t_L g3027 ( 
.A(n_2486),
.B(n_2488),
.Y(n_3027)
);

CKINVDCx8_ASAP7_75t_R g3028 ( 
.A(n_2216),
.Y(n_3028)
);

NAND2xp5_ASAP7_75t_SL g3029 ( 
.A(n_2489),
.B(n_2490),
.Y(n_3029)
);

NAND2x1p5_ASAP7_75t_L g3030 ( 
.A(n_2163),
.B(n_2164),
.Y(n_3030)
);

NAND2xp5_ASAP7_75t_L g3031 ( 
.A(n_2489),
.B(n_2490),
.Y(n_3031)
);

NOR2x1p5_ASAP7_75t_L g3032 ( 
.A(n_1842),
.B(n_2493),
.Y(n_3032)
);

BUFx4f_ASAP7_75t_L g3033 ( 
.A(n_2118),
.Y(n_3033)
);

AOI22xp5_ASAP7_75t_L g3034 ( 
.A1(n_2573),
.A2(n_2589),
.B1(n_2595),
.B2(n_2574),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_L g3035 ( 
.A(n_2493),
.B(n_2494),
.Y(n_3035)
);

BUFx6f_ASAP7_75t_L g3036 ( 
.A(n_2118),
.Y(n_3036)
);

OR2x2_ASAP7_75t_SL g3037 ( 
.A(n_1842),
.B(n_1978),
.Y(n_3037)
);

BUFx2_ASAP7_75t_L g3038 ( 
.A(n_2164),
.Y(n_3038)
);

CKINVDCx5p33_ASAP7_75t_R g3039 ( 
.A(n_2171),
.Y(n_3039)
);

INVx2_ASAP7_75t_SL g3040 ( 
.A(n_2172),
.Y(n_3040)
);

NAND2xp5_ASAP7_75t_L g3041 ( 
.A(n_2494),
.B(n_2498),
.Y(n_3041)
);

AOI22xp33_ASAP7_75t_L g3042 ( 
.A1(n_2606),
.A2(n_2640),
.B1(n_2614),
.B2(n_2500),
.Y(n_3042)
);

NOR2x1_ASAP7_75t_L g3043 ( 
.A(n_1933),
.B(n_1928),
.Y(n_3043)
);

INVx5_ASAP7_75t_L g3044 ( 
.A(n_2391),
.Y(n_3044)
);

AO22x1_ASAP7_75t_L g3045 ( 
.A1(n_2038),
.A2(n_2122),
.B1(n_2500),
.B2(n_2498),
.Y(n_3045)
);

INVx2_ASAP7_75t_L g3046 ( 
.A(n_2386),
.Y(n_3046)
);

AND2x4_ASAP7_75t_L g3047 ( 
.A(n_2072),
.B(n_2184),
.Y(n_3047)
);

BUFx6f_ASAP7_75t_L g3048 ( 
.A(n_2391),
.Y(n_3048)
);

NAND2xp5_ASAP7_75t_SL g3049 ( 
.A(n_2507),
.B(n_2512),
.Y(n_3049)
);

AOI22xp33_ASAP7_75t_L g3050 ( 
.A1(n_2507),
.A2(n_2514),
.B1(n_2516),
.B2(n_2512),
.Y(n_3050)
);

BUFx3_ASAP7_75t_L g3051 ( 
.A(n_2391),
.Y(n_3051)
);

INVx2_ASAP7_75t_SL g3052 ( 
.A(n_2172),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_L g3053 ( 
.A(n_2514),
.B(n_2612),
.Y(n_3053)
);

INVx3_ASAP7_75t_L g3054 ( 
.A(n_2094),
.Y(n_3054)
);

INVx1_ASAP7_75t_SL g3055 ( 
.A(n_1913),
.Y(n_3055)
);

O2A1O1Ixp5_ASAP7_75t_L g3056 ( 
.A1(n_1928),
.A2(n_2122),
.B(n_2518),
.C(n_2516),
.Y(n_3056)
);

INVx2_ASAP7_75t_L g3057 ( 
.A(n_2390),
.Y(n_3057)
);

INVx3_ASAP7_75t_L g3058 ( 
.A(n_2094),
.Y(n_3058)
);

AOI22xp33_ASAP7_75t_L g3059 ( 
.A1(n_2518),
.A2(n_2526),
.B1(n_2534),
.B2(n_2519),
.Y(n_3059)
);

INVx2_ASAP7_75t_L g3060 ( 
.A(n_2390),
.Y(n_3060)
);

NOR2x1p5_ASAP7_75t_L g3061 ( 
.A(n_2519),
.B(n_2526),
.Y(n_3061)
);

NOR2xp33_ASAP7_75t_L g3062 ( 
.A(n_1838),
.B(n_1843),
.Y(n_3062)
);

AND2x2_ASAP7_75t_L g3063 ( 
.A(n_1878),
.B(n_1929),
.Y(n_3063)
);

AOI22xp5_ASAP7_75t_L g3064 ( 
.A1(n_2534),
.A2(n_2535),
.B1(n_2542),
.B2(n_2537),
.Y(n_3064)
);

AND2x4_ASAP7_75t_L g3065 ( 
.A(n_2072),
.B(n_2184),
.Y(n_3065)
);

INVx2_ASAP7_75t_L g3066 ( 
.A(n_2393),
.Y(n_3066)
);

INVx4_ASAP7_75t_L g3067 ( 
.A(n_2391),
.Y(n_3067)
);

INVxp67_ASAP7_75t_L g3068 ( 
.A(n_1978),
.Y(n_3068)
);

CKINVDCx16_ASAP7_75t_R g3069 ( 
.A(n_2171),
.Y(n_3069)
);

BUFx2_ASAP7_75t_L g3070 ( 
.A(n_2005),
.Y(n_3070)
);

NAND2xp5_ASAP7_75t_L g3071 ( 
.A(n_2535),
.B(n_2537),
.Y(n_3071)
);

INVx4_ASAP7_75t_L g3072 ( 
.A(n_2391),
.Y(n_3072)
);

BUFx2_ASAP7_75t_L g3073 ( 
.A(n_2009),
.Y(n_3073)
);

CKINVDCx5p33_ASAP7_75t_R g3074 ( 
.A(n_2373),
.Y(n_3074)
);

BUFx6f_ASAP7_75t_L g3075 ( 
.A(n_2501),
.Y(n_3075)
);

BUFx6f_ASAP7_75t_L g3076 ( 
.A(n_2501),
.Y(n_3076)
);

NAND2xp5_ASAP7_75t_L g3077 ( 
.A(n_2542),
.B(n_2543),
.Y(n_3077)
);

AND2x4_ASAP7_75t_L g3078 ( 
.A(n_2072),
.B(n_2184),
.Y(n_3078)
);

INVx3_ASAP7_75t_L g3079 ( 
.A(n_2094),
.Y(n_3079)
);

INVx5_ASAP7_75t_L g3080 ( 
.A(n_2501),
.Y(n_3080)
);

NOR2xp33_ASAP7_75t_L g3081 ( 
.A(n_1843),
.B(n_1845),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_L g3082 ( 
.A(n_2543),
.B(n_2544),
.Y(n_3082)
);

BUFx3_ASAP7_75t_L g3083 ( 
.A(n_2501),
.Y(n_3083)
);

INVx2_ASAP7_75t_L g3084 ( 
.A(n_2412),
.Y(n_3084)
);

NAND2x1p5_ASAP7_75t_L g3085 ( 
.A(n_2163),
.B(n_1904),
.Y(n_3085)
);

OR2x6_ASAP7_75t_SL g3086 ( 
.A(n_2544),
.B(n_2547),
.Y(n_3086)
);

CKINVDCx20_ASAP7_75t_R g3087 ( 
.A(n_1900),
.Y(n_3087)
);

INVx1_ASAP7_75t_SL g3088 ( 
.A(n_1913),
.Y(n_3088)
);

INVx2_ASAP7_75t_SL g3089 ( 
.A(n_2172),
.Y(n_3089)
);

HB1xp67_ASAP7_75t_L g3090 ( 
.A(n_2035),
.Y(n_3090)
);

INVx2_ASAP7_75t_SL g3091 ( 
.A(n_2179),
.Y(n_3091)
);

INVx5_ASAP7_75t_L g3092 ( 
.A(n_2501),
.Y(n_3092)
);

NAND2xp5_ASAP7_75t_L g3093 ( 
.A(n_2547),
.B(n_2555),
.Y(n_3093)
);

INVx5_ASAP7_75t_L g3094 ( 
.A(n_1904),
.Y(n_3094)
);

BUFx4f_ASAP7_75t_L g3095 ( 
.A(n_1953),
.Y(n_3095)
);

INVx3_ASAP7_75t_L g3096 ( 
.A(n_2094),
.Y(n_3096)
);

AND2x4_ASAP7_75t_SL g3097 ( 
.A(n_1904),
.B(n_2105),
.Y(n_3097)
);

BUFx4f_ASAP7_75t_L g3098 ( 
.A(n_1953),
.Y(n_3098)
);

AOI22xp5_ASAP7_75t_L g3099 ( 
.A1(n_2555),
.A2(n_2566),
.B1(n_2572),
.B2(n_2565),
.Y(n_3099)
);

AOI22xp5_ASAP7_75t_SL g3100 ( 
.A1(n_1845),
.A2(n_2565),
.B1(n_2572),
.B2(n_2566),
.Y(n_3100)
);

BUFx4f_ASAP7_75t_L g3101 ( 
.A(n_1953),
.Y(n_3101)
);

AND2x4_ASAP7_75t_L g3102 ( 
.A(n_2184),
.B(n_1824),
.Y(n_3102)
);

NOR2xp33_ASAP7_75t_L g3103 ( 
.A(n_2576),
.B(n_2583),
.Y(n_3103)
);

AND2x2_ASAP7_75t_L g3104 ( 
.A(n_1929),
.B(n_2357),
.Y(n_3104)
);

AND2x4_ASAP7_75t_L g3105 ( 
.A(n_2184),
.B(n_1824),
.Y(n_3105)
);

NOR2x1p5_ASAP7_75t_L g3106 ( 
.A(n_2576),
.B(n_2583),
.Y(n_3106)
);

INVx3_ASAP7_75t_L g3107 ( 
.A(n_2160),
.Y(n_3107)
);

AND2x6_ASAP7_75t_L g3108 ( 
.A(n_2160),
.B(n_2497),
.Y(n_3108)
);

NAND2xp5_ASAP7_75t_L g3109 ( 
.A(n_2585),
.B(n_2590),
.Y(n_3109)
);

NAND2xp5_ASAP7_75t_L g3110 ( 
.A(n_2585),
.B(n_2590),
.Y(n_3110)
);

AND2x4_ASAP7_75t_L g3111 ( 
.A(n_1824),
.B(n_1896),
.Y(n_3111)
);

BUFx3_ASAP7_75t_L g3112 ( 
.A(n_2605),
.Y(n_3112)
);

NAND2x1p5_ASAP7_75t_L g3113 ( 
.A(n_2105),
.B(n_2402),
.Y(n_3113)
);

AND2x2_ASAP7_75t_L g3114 ( 
.A(n_2357),
.B(n_2362),
.Y(n_3114)
);

NAND2xp5_ASAP7_75t_SL g3115 ( 
.A(n_2591),
.B(n_2594),
.Y(n_3115)
);

OR2x6_ASAP7_75t_L g3116 ( 
.A(n_2146),
.B(n_2166),
.Y(n_3116)
);

OR2x2_ASAP7_75t_L g3117 ( 
.A(n_2591),
.B(n_2594),
.Y(n_3117)
);

INVxp67_ASAP7_75t_SL g3118 ( 
.A(n_2060),
.Y(n_3118)
);

NAND2xp5_ASAP7_75t_L g3119 ( 
.A(n_2597),
.B(n_2598),
.Y(n_3119)
);

BUFx6f_ASAP7_75t_L g3120 ( 
.A(n_2605),
.Y(n_3120)
);

INVx5_ASAP7_75t_L g3121 ( 
.A(n_2105),
.Y(n_3121)
);

INVx5_ASAP7_75t_L g3122 ( 
.A(n_2105),
.Y(n_3122)
);

BUFx2_ASAP7_75t_L g3123 ( 
.A(n_1844),
.Y(n_3123)
);

BUFx2_ASAP7_75t_L g3124 ( 
.A(n_1965),
.Y(n_3124)
);

CKINVDCx5p33_ASAP7_75t_R g3125 ( 
.A(n_2373),
.Y(n_3125)
);

NAND2xp5_ASAP7_75t_L g3126 ( 
.A(n_2597),
.B(n_2598),
.Y(n_3126)
);

INVx1_ASAP7_75t_SL g3127 ( 
.A(n_2009),
.Y(n_3127)
);

INVxp67_ASAP7_75t_SL g3128 ( 
.A(n_2340),
.Y(n_3128)
);

BUFx3_ASAP7_75t_L g3129 ( 
.A(n_2605),
.Y(n_3129)
);

INVx5_ASAP7_75t_L g3130 ( 
.A(n_2402),
.Y(n_3130)
);

INVx3_ASAP7_75t_L g3131 ( 
.A(n_2160),
.Y(n_3131)
);

INVx2_ASAP7_75t_SL g3132 ( 
.A(n_2179),
.Y(n_3132)
);

NAND2xp5_ASAP7_75t_L g3133 ( 
.A(n_2602),
.B(n_2610),
.Y(n_3133)
);

OR2x6_ASAP7_75t_L g3134 ( 
.A(n_2166),
.B(n_2641),
.Y(n_3134)
);

AND2x2_ASAP7_75t_L g3135 ( 
.A(n_2362),
.B(n_2377),
.Y(n_3135)
);

NAND2xp5_ASAP7_75t_L g3136 ( 
.A(n_2602),
.B(n_2610),
.Y(n_3136)
);

AND2x2_ASAP7_75t_L g3137 ( 
.A(n_2377),
.B(n_2471),
.Y(n_3137)
);

NAND2xp33_ASAP7_75t_L g3138 ( 
.A(n_1884),
.B(n_2612),
.Y(n_3138)
);

INVx2_ASAP7_75t_SL g3139 ( 
.A(n_2179),
.Y(n_3139)
);

INVx3_ASAP7_75t_L g3140 ( 
.A(n_2160),
.Y(n_3140)
);

BUFx2_ASAP7_75t_L g3141 ( 
.A(n_2157),
.Y(n_3141)
);

INVx2_ASAP7_75t_SL g3142 ( 
.A(n_2365),
.Y(n_3142)
);

BUFx8_ASAP7_75t_SL g3143 ( 
.A(n_2340),
.Y(n_3143)
);

NAND2xp5_ASAP7_75t_SL g3144 ( 
.A(n_1873),
.B(n_1868),
.Y(n_3144)
);

NAND2x1p5_ASAP7_75t_L g3145 ( 
.A(n_2402),
.B(n_2476),
.Y(n_3145)
);

NAND2xp5_ASAP7_75t_L g3146 ( 
.A(n_1934),
.B(n_1849),
.Y(n_3146)
);

BUFx3_ASAP7_75t_L g3147 ( 
.A(n_2641),
.Y(n_3147)
);

BUFx6f_ASAP7_75t_L g3148 ( 
.A(n_2641),
.Y(n_3148)
);

NAND2xp5_ASAP7_75t_SL g3149 ( 
.A(n_1873),
.B(n_2112),
.Y(n_3149)
);

INVxp67_ASAP7_75t_L g3150 ( 
.A(n_2035),
.Y(n_3150)
);

NAND2xp5_ASAP7_75t_SL g3151 ( 
.A(n_1849),
.B(n_1852),
.Y(n_3151)
);

NAND2xp5_ASAP7_75t_L g3152 ( 
.A(n_1934),
.B(n_1852),
.Y(n_3152)
);

NAND2x1p5_ASAP7_75t_L g3153 ( 
.A(n_2402),
.B(n_2476),
.Y(n_3153)
);

INVx1_ASAP7_75t_SL g3154 ( 
.A(n_2182),
.Y(n_3154)
);

NOR2x1_ASAP7_75t_L g3155 ( 
.A(n_2127),
.B(n_2272),
.Y(n_3155)
);

NAND2xp5_ASAP7_75t_L g3156 ( 
.A(n_1854),
.B(n_1857),
.Y(n_3156)
);

AND2x2_ASAP7_75t_L g3157 ( 
.A(n_2471),
.B(n_2482),
.Y(n_3157)
);

BUFx4f_ASAP7_75t_L g3158 ( 
.A(n_2160),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_L g3159 ( 
.A(n_1854),
.B(n_1857),
.Y(n_3159)
);

NAND2xp33_ASAP7_75t_L g3160 ( 
.A(n_1824),
.B(n_1896),
.Y(n_3160)
);

INVx4_ASAP7_75t_L g3161 ( 
.A(n_1824),
.Y(n_3161)
);

INVx3_ASAP7_75t_L g3162 ( 
.A(n_2160),
.Y(n_3162)
);

BUFx3_ASAP7_75t_L g3163 ( 
.A(n_2243),
.Y(n_3163)
);

BUFx3_ASAP7_75t_L g3164 ( 
.A(n_2243),
.Y(n_3164)
);

INVx6_ASAP7_75t_L g3165 ( 
.A(n_2476),
.Y(n_3165)
);

INVx3_ASAP7_75t_L g3166 ( 
.A(n_2497),
.Y(n_3166)
);

BUFx6f_ASAP7_75t_L g3167 ( 
.A(n_2497),
.Y(n_3167)
);

CKINVDCx5p33_ASAP7_75t_R g3168 ( 
.A(n_2385),
.Y(n_3168)
);

AND2x4_ASAP7_75t_SL g3169 ( 
.A(n_2476),
.B(n_2481),
.Y(n_3169)
);

BUFx3_ASAP7_75t_L g3170 ( 
.A(n_2157),
.Y(n_3170)
);

BUFx2_ASAP7_75t_L g3171 ( 
.A(n_2205),
.Y(n_3171)
);

INVx3_ASAP7_75t_L g3172 ( 
.A(n_2497),
.Y(n_3172)
);

AOI22xp5_ASAP7_75t_L g3173 ( 
.A1(n_2482),
.A2(n_2539),
.B1(n_2603),
.B2(n_2559),
.Y(n_3173)
);

NOR2x1_ASAP7_75t_L g3174 ( 
.A(n_2127),
.B(n_2205),
.Y(n_3174)
);

AND3x1_ASAP7_75t_SL g3175 ( 
.A(n_2346),
.B(n_2176),
.C(n_2269),
.Y(n_3175)
);

NOR2xp33_ASAP7_75t_L g3176 ( 
.A(n_1861),
.B(n_1865),
.Y(n_3176)
);

BUFx3_ASAP7_75t_L g3177 ( 
.A(n_2497),
.Y(n_3177)
);

AOI22xp5_ASAP7_75t_L g3178 ( 
.A1(n_2539),
.A2(n_2559),
.B1(n_2643),
.B2(n_2603),
.Y(n_3178)
);

BUFx4f_ASAP7_75t_L g3179 ( 
.A(n_2365),
.Y(n_3179)
);

BUFx2_ASAP7_75t_L g3180 ( 
.A(n_2509),
.Y(n_3180)
);

INVx2_ASAP7_75t_SL g3181 ( 
.A(n_2365),
.Y(n_3181)
);

BUFx12f_ASAP7_75t_L g3182 ( 
.A(n_2385),
.Y(n_3182)
);

BUFx3_ASAP7_75t_L g3183 ( 
.A(n_1824),
.Y(n_3183)
);

NAND2xp5_ASAP7_75t_SL g3184 ( 
.A(n_1861),
.B(n_1865),
.Y(n_3184)
);

NAND2xp5_ASAP7_75t_SL g3185 ( 
.A(n_2034),
.B(n_2643),
.Y(n_3185)
);

NAND2xp5_ASAP7_75t_L g3186 ( 
.A(n_2560),
.B(n_2562),
.Y(n_3186)
);

AND2x2_ASAP7_75t_L g3187 ( 
.A(n_1930),
.B(n_1966),
.Y(n_3187)
);

AND2x2_ASAP7_75t_SL g3188 ( 
.A(n_2283),
.B(n_2481),
.Y(n_3188)
);

HB1xp67_ASAP7_75t_L g3189 ( 
.A(n_2182),
.Y(n_3189)
);

AOI21xp5_ASAP7_75t_L g3190 ( 
.A1(n_2022),
.A2(n_2283),
.B(n_2133),
.Y(n_3190)
);

NAND2x1p5_ASAP7_75t_L g3191 ( 
.A(n_2481),
.B(n_2580),
.Y(n_3191)
);

OR2x6_ASAP7_75t_L g3192 ( 
.A(n_2521),
.B(n_2522),
.Y(n_3192)
);

INVxp67_ASAP7_75t_SL g3193 ( 
.A(n_2267),
.Y(n_3193)
);

AND2x4_ASAP7_75t_L g3194 ( 
.A(n_1824),
.B(n_1896),
.Y(n_3194)
);

INVxp67_ASAP7_75t_L g3195 ( 
.A(n_2068),
.Y(n_3195)
);

INVxp67_ASAP7_75t_L g3196 ( 
.A(n_2068),
.Y(n_3196)
);

BUFx6f_ASAP7_75t_L g3197 ( 
.A(n_1896),
.Y(n_3197)
);

BUFx6f_ASAP7_75t_L g3198 ( 
.A(n_1896),
.Y(n_3198)
);

OR2x2_ASAP7_75t_SL g3199 ( 
.A(n_2233),
.B(n_1991),
.Y(n_3199)
);

AND2x4_ASAP7_75t_L g3200 ( 
.A(n_1896),
.B(n_2367),
.Y(n_3200)
);

INVx2_ASAP7_75t_SL g3201 ( 
.A(n_2521),
.Y(n_3201)
);

NOR2xp33_ASAP7_75t_L g3202 ( 
.A(n_1960),
.B(n_1859),
.Y(n_3202)
);

NAND2xp5_ASAP7_75t_L g3203 ( 
.A(n_2564),
.B(n_2582),
.Y(n_3203)
);

OAI22xp33_ASAP7_75t_L g3204 ( 
.A1(n_2064),
.A2(n_2078),
.B1(n_2115),
.B2(n_2092),
.Y(n_3204)
);

CKINVDCx5p33_ASAP7_75t_R g3205 ( 
.A(n_2511),
.Y(n_3205)
);

AOI22xp5_ASAP7_75t_L g3206 ( 
.A1(n_1877),
.A2(n_1882),
.B1(n_1908),
.B2(n_1899),
.Y(n_3206)
);

AND2x4_ASAP7_75t_L g3207 ( 
.A(n_1896),
.B(n_2367),
.Y(n_3207)
);

NOR2xp33_ASAP7_75t_R g3208 ( 
.A(n_2045),
.B(n_2073),
.Y(n_3208)
);

CKINVDCx5p33_ASAP7_75t_R g3209 ( 
.A(n_2511),
.Y(n_3209)
);

A2O1A1Ixp33_ASAP7_75t_L g3210 ( 
.A1(n_2024),
.A2(n_2086),
.B(n_2095),
.C(n_2067),
.Y(n_3210)
);

BUFx3_ASAP7_75t_L g3211 ( 
.A(n_2367),
.Y(n_3211)
);

HB1xp67_ASAP7_75t_L g3212 ( 
.A(n_2298),
.Y(n_3212)
);

BUFx3_ASAP7_75t_L g3213 ( 
.A(n_2367),
.Y(n_3213)
);

AOI22xp5_ASAP7_75t_L g3214 ( 
.A1(n_2116),
.A2(n_1984),
.B1(n_1888),
.B2(n_1880),
.Y(n_3214)
);

CKINVDCx5p33_ASAP7_75t_R g3215 ( 
.A(n_1900),
.Y(n_3215)
);

INVx3_ASAP7_75t_SL g3216 ( 
.A(n_2481),
.Y(n_3216)
);

AND2x4_ASAP7_75t_L g3217 ( 
.A(n_2367),
.B(n_2577),
.Y(n_3217)
);

BUFx3_ASAP7_75t_L g3218 ( 
.A(n_2367),
.Y(n_3218)
);

NAND2xp5_ASAP7_75t_L g3219 ( 
.A(n_2647),
.B(n_1818),
.Y(n_3219)
);

NAND2xp5_ASAP7_75t_L g3220 ( 
.A(n_1818),
.B(n_1819),
.Y(n_3220)
);

NOR2xp67_ASAP7_75t_L g3221 ( 
.A(n_2521),
.B(n_2522),
.Y(n_3221)
);

BUFx3_ASAP7_75t_L g3222 ( 
.A(n_2367),
.Y(n_3222)
);

AOI22xp5_ASAP7_75t_L g3223 ( 
.A1(n_1880),
.A2(n_1888),
.B1(n_1918),
.B2(n_1903),
.Y(n_3223)
);

INVx1_ASAP7_75t_L g3224 ( 
.A(n_1819),
.Y(n_3224)
);

BUFx2_ASAP7_75t_L g3225 ( 
.A(n_2601),
.Y(n_3225)
);

CKINVDCx5p33_ASAP7_75t_R g3226 ( 
.A(n_2040),
.Y(n_3226)
);

HB1xp67_ASAP7_75t_L g3227 ( 
.A(n_2298),
.Y(n_3227)
);

INVx1_ASAP7_75t_SL g3228 ( 
.A(n_2629),
.Y(n_3228)
);

OAI22xp5_ASAP7_75t_SL g3229 ( 
.A1(n_2004),
.A2(n_1976),
.B1(n_1927),
.B2(n_1990),
.Y(n_3229)
);

NOR2x1_ASAP7_75t_L g3230 ( 
.A(n_2580),
.B(n_1991),
.Y(n_3230)
);

OR2x6_ASAP7_75t_L g3231 ( 
.A(n_2522),
.B(n_2627),
.Y(n_3231)
);

INVxp67_ASAP7_75t_L g3232 ( 
.A(n_2101),
.Y(n_3232)
);

INVx1_ASAP7_75t_L g3233 ( 
.A(n_1827),
.Y(n_3233)
);

INVx2_ASAP7_75t_L g3234 ( 
.A(n_1827),
.Y(n_3234)
);

CKINVDCx5p33_ASAP7_75t_R g3235 ( 
.A(n_2040),
.Y(n_3235)
);

NOR2xp33_ASAP7_75t_L g3236 ( 
.A(n_1911),
.B(n_1916),
.Y(n_3236)
);

BUFx3_ASAP7_75t_L g3237 ( 
.A(n_2577),
.Y(n_3237)
);

INVx2_ASAP7_75t_L g3238 ( 
.A(n_1837),
.Y(n_3238)
);

AOI22xp5_ASAP7_75t_L g3239 ( 
.A1(n_1925),
.A2(n_2006),
.B1(n_2008),
.B2(n_2025),
.Y(n_3239)
);

INVx2_ASAP7_75t_L g3240 ( 
.A(n_1837),
.Y(n_3240)
);

BUFx6f_ASAP7_75t_L g3241 ( 
.A(n_2577),
.Y(n_3241)
);

AOI22xp33_ASAP7_75t_L g3242 ( 
.A1(n_1931),
.A2(n_2114),
.B1(n_1952),
.B2(n_2006),
.Y(n_3242)
);

INVx5_ASAP7_75t_L g3243 ( 
.A(n_2580),
.Y(n_3243)
);

INVx1_ASAP7_75t_L g3244 ( 
.A(n_1848),
.Y(n_3244)
);

BUFx2_ASAP7_75t_L g3245 ( 
.A(n_2216),
.Y(n_3245)
);

AND2x4_ASAP7_75t_L g3246 ( 
.A(n_2577),
.B(n_2580),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_1848),
.Y(n_3247)
);

NAND2xp5_ASAP7_75t_L g3248 ( 
.A(n_1851),
.B(n_1856),
.Y(n_3248)
);

AND2x4_ASAP7_75t_L g3249 ( 
.A(n_2577),
.B(n_2627),
.Y(n_3249)
);

HB1xp67_ASAP7_75t_L g3250 ( 
.A(n_2306),
.Y(n_3250)
);

NAND2xp5_ASAP7_75t_L g3251 ( 
.A(n_1851),
.B(n_1856),
.Y(n_3251)
);

INVx1_ASAP7_75t_L g3252 ( 
.A(n_1860),
.Y(n_3252)
);

INVx1_ASAP7_75t_L g3253 ( 
.A(n_1860),
.Y(n_3253)
);

INVx2_ASAP7_75t_L g3254 ( 
.A(n_1870),
.Y(n_3254)
);

AND2x4_ASAP7_75t_L g3255 ( 
.A(n_2577),
.B(n_2627),
.Y(n_3255)
);

INVx1_ASAP7_75t_L g3256 ( 
.A(n_1870),
.Y(n_3256)
);

CKINVDCx5p33_ASAP7_75t_R g3257 ( 
.A(n_2079),
.Y(n_3257)
);

HB1xp67_ASAP7_75t_L g3258 ( 
.A(n_2306),
.Y(n_3258)
);

INVx2_ASAP7_75t_L g3259 ( 
.A(n_1905),
.Y(n_3259)
);

BUFx2_ASAP7_75t_L g3260 ( 
.A(n_2079),
.Y(n_3260)
);

NAND2xp5_ASAP7_75t_L g3261 ( 
.A(n_1905),
.B(n_1937),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_1937),
.Y(n_3262)
);

NAND2xp5_ASAP7_75t_L g3263 ( 
.A(n_1945),
.B(n_1956),
.Y(n_3263)
);

NAND2xp5_ASAP7_75t_SL g3264 ( 
.A(n_2025),
.B(n_2056),
.Y(n_3264)
);

HB1xp67_ASAP7_75t_L g3265 ( 
.A(n_2312),
.Y(n_3265)
);

HB1xp67_ASAP7_75t_L g3266 ( 
.A(n_2312),
.Y(n_3266)
);

NAND2x1p5_ASAP7_75t_L g3267 ( 
.A(n_2577),
.B(n_1890),
.Y(n_3267)
);

INVx2_ASAP7_75t_L g3268 ( 
.A(n_1945),
.Y(n_3268)
);

AND2x4_ASAP7_75t_L g3269 ( 
.A(n_1901),
.B(n_2077),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_1956),
.Y(n_3270)
);

AOI22xp5_ASAP7_75t_L g3271 ( 
.A1(n_2047),
.A2(n_1938),
.B1(n_2104),
.B2(n_2018),
.Y(n_3271)
);

AND2x2_ASAP7_75t_SL g3272 ( 
.A(n_2405),
.B(n_2292),
.Y(n_3272)
);

AND2x4_ASAP7_75t_L g3273 ( 
.A(n_1901),
.B(n_2077),
.Y(n_3273)
);

INVx2_ASAP7_75t_L g3274 ( 
.A(n_1968),
.Y(n_3274)
);

BUFx4f_ASAP7_75t_L g3275 ( 
.A(n_2218),
.Y(n_3275)
);

BUFx12f_ASAP7_75t_L g3276 ( 
.A(n_2109),
.Y(n_3276)
);

AND2x2_ASAP7_75t_L g3277 ( 
.A(n_2055),
.B(n_1968),
.Y(n_3277)
);

INVx2_ASAP7_75t_SL g3278 ( 
.A(n_2282),
.Y(n_3278)
);

AOI22xp5_ASAP7_75t_L g3279 ( 
.A1(n_1938),
.A2(n_2104),
.B1(n_2018),
.B2(n_2053),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_1969),
.Y(n_3280)
);

AOI22xp33_ASAP7_75t_L g3281 ( 
.A1(n_2134),
.A2(n_2070),
.B1(n_2074),
.B2(n_2069),
.Y(n_3281)
);

NAND2xp5_ASAP7_75t_SL g3282 ( 
.A(n_2019),
.B(n_2269),
.Y(n_3282)
);

INVx1_ASAP7_75t_L g3283 ( 
.A(n_1969),
.Y(n_3283)
);

INVxp67_ASAP7_75t_L g3284 ( 
.A(n_2069),
.Y(n_3284)
);

INVx1_ASAP7_75t_L g3285 ( 
.A(n_1975),
.Y(n_3285)
);

BUFx3_ASAP7_75t_L g3286 ( 
.A(n_2405),
.Y(n_3286)
);

BUFx3_ASAP7_75t_L g3287 ( 
.A(n_2405),
.Y(n_3287)
);

NOR2xp33_ASAP7_75t_L g3288 ( 
.A(n_2554),
.B(n_2604),
.Y(n_3288)
);

NAND2xp5_ASAP7_75t_L g3289 ( 
.A(n_1975),
.B(n_1983),
.Y(n_3289)
);

INVx2_ASAP7_75t_L g3290 ( 
.A(n_1983),
.Y(n_3290)
);

NAND2xp5_ASAP7_75t_L g3291 ( 
.A(n_1994),
.B(n_1995),
.Y(n_3291)
);

AO22x1_ASAP7_75t_L g3292 ( 
.A1(n_2305),
.A2(n_2091),
.B1(n_2234),
.B2(n_2044),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_L g3293 ( 
.A(n_1994),
.B(n_1995),
.Y(n_3293)
);

INVxp67_ASAP7_75t_L g3294 ( 
.A(n_2070),
.Y(n_3294)
);

AND2x2_ASAP7_75t_L g3295 ( 
.A(n_2055),
.B(n_2003),
.Y(n_3295)
);

CKINVDCx5p33_ASAP7_75t_R g3296 ( 
.A(n_2109),
.Y(n_3296)
);

INVx2_ASAP7_75t_L g3297 ( 
.A(n_2003),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_2011),
.Y(n_3298)
);

INVxp67_ASAP7_75t_SL g3299 ( 
.A(n_2267),
.Y(n_3299)
);

INVx1_ASAP7_75t_L g3300 ( 
.A(n_2011),
.Y(n_3300)
);

INVx1_ASAP7_75t_L g3301 ( 
.A(n_2013),
.Y(n_3301)
);

INVx2_ASAP7_75t_L g3302 ( 
.A(n_2013),
.Y(n_3302)
);

HB1xp67_ASAP7_75t_L g3303 ( 
.A(n_2329),
.Y(n_3303)
);

AOI22xp33_ASAP7_75t_L g3304 ( 
.A1(n_2134),
.A2(n_2083),
.B1(n_2089),
.B2(n_2074),
.Y(n_3304)
);

INVx1_ASAP7_75t_L g3305 ( 
.A(n_2021),
.Y(n_3305)
);

INVx2_ASAP7_75t_L g3306 ( 
.A(n_2021),
.Y(n_3306)
);

NAND2xp5_ASAP7_75t_SL g3307 ( 
.A(n_2168),
.B(n_2300),
.Y(n_3307)
);

INVx1_ASAP7_75t_L g3308 ( 
.A(n_2026),
.Y(n_3308)
);

BUFx8_ASAP7_75t_L g3309 ( 
.A(n_1954),
.Y(n_3309)
);

NOR2xp33_ASAP7_75t_L g3310 ( 
.A(n_2554),
.B(n_2604),
.Y(n_3310)
);

INVx5_ASAP7_75t_L g3311 ( 
.A(n_2218),
.Y(n_3311)
);

INVx2_ASAP7_75t_L g3312 ( 
.A(n_2026),
.Y(n_3312)
);

INVx2_ASAP7_75t_L g3313 ( 
.A(n_2036),
.Y(n_3313)
);

NAND2xp5_ASAP7_75t_SL g3314 ( 
.A(n_2300),
.B(n_2292),
.Y(n_3314)
);

INVx2_ASAP7_75t_SL g3315 ( 
.A(n_2282),
.Y(n_3315)
);

INVx2_ASAP7_75t_L g3316 ( 
.A(n_2036),
.Y(n_3316)
);

OR2x2_ASAP7_75t_SL g3317 ( 
.A(n_2234),
.B(n_2238),
.Y(n_3317)
);

NAND2xp5_ASAP7_75t_L g3318 ( 
.A(n_2041),
.B(n_2042),
.Y(n_3318)
);

INVx1_ASAP7_75t_L g3319 ( 
.A(n_2041),
.Y(n_3319)
);

NOR2xp33_ASAP7_75t_L g3320 ( 
.A(n_2649),
.B(n_2416),
.Y(n_3320)
);

NAND2xp5_ASAP7_75t_L g3321 ( 
.A(n_2042),
.B(n_2049),
.Y(n_3321)
);

INVx2_ASAP7_75t_L g3322 ( 
.A(n_2049),
.Y(n_3322)
);

INVxp67_ASAP7_75t_L g3323 ( 
.A(n_2083),
.Y(n_3323)
);

INVx1_ASAP7_75t_L g3324 ( 
.A(n_2058),
.Y(n_3324)
);

NAND2xp5_ASAP7_75t_L g3325 ( 
.A(n_2058),
.B(n_2059),
.Y(n_3325)
);

AND2x4_ASAP7_75t_L g3326 ( 
.A(n_2178),
.B(n_2422),
.Y(n_3326)
);

NAND2xp5_ASAP7_75t_L g3327 ( 
.A(n_2059),
.B(n_2065),
.Y(n_3327)
);

NAND2xp5_ASAP7_75t_L g3328 ( 
.A(n_2065),
.B(n_2084),
.Y(n_3328)
);

NAND2xp5_ASAP7_75t_L g3329 ( 
.A(n_2084),
.B(n_2121),
.Y(n_3329)
);

AND2x2_ASAP7_75t_L g3330 ( 
.A(n_2121),
.B(n_2125),
.Y(n_3330)
);

NAND2xp5_ASAP7_75t_L g3331 ( 
.A(n_2125),
.B(n_2128),
.Y(n_3331)
);

INVx1_ASAP7_75t_L g3332 ( 
.A(n_2128),
.Y(n_3332)
);

BUFx6f_ASAP7_75t_L g3333 ( 
.A(n_2249),
.Y(n_3333)
);

NAND2xp5_ASAP7_75t_L g3334 ( 
.A(n_2143),
.B(n_2156),
.Y(n_3334)
);

NAND2xp5_ASAP7_75t_L g3335 ( 
.A(n_2143),
.B(n_2156),
.Y(n_3335)
);

AND2x4_ASAP7_75t_L g3336 ( 
.A(n_2178),
.B(n_2422),
.Y(n_3336)
);

OR2x6_ASAP7_75t_L g3337 ( 
.A(n_2242),
.B(n_2305),
.Y(n_3337)
);

BUFx6f_ASAP7_75t_L g3338 ( 
.A(n_2249),
.Y(n_3338)
);

INVx2_ASAP7_75t_L g3339 ( 
.A(n_2193),
.Y(n_3339)
);

INVx1_ASAP7_75t_L g3340 ( 
.A(n_2193),
.Y(n_3340)
);

AND2x4_ASAP7_75t_L g3341 ( 
.A(n_2178),
.B(n_2422),
.Y(n_3341)
);

NAND2xp5_ASAP7_75t_L g3342 ( 
.A(n_2348),
.B(n_2370),
.Y(n_3342)
);

INVx1_ASAP7_75t_L g3343 ( 
.A(n_2348),
.Y(n_3343)
);

BUFx2_ASAP7_75t_L g3344 ( 
.A(n_2110),
.Y(n_3344)
);

BUFx3_ASAP7_75t_L g3345 ( 
.A(n_2282),
.Y(n_3345)
);

INVx1_ASAP7_75t_L g3346 ( 
.A(n_2370),
.Y(n_3346)
);

INVx2_ASAP7_75t_L g3347 ( 
.A(n_2371),
.Y(n_3347)
);

AO221x1_ASAP7_75t_L g3348 ( 
.A1(n_2329),
.A2(n_2253),
.B1(n_2217),
.B2(n_2271),
.C(n_2266),
.Y(n_3348)
);

INVx2_ASAP7_75t_L g3349 ( 
.A(n_2371),
.Y(n_3349)
);

NAND2xp5_ASAP7_75t_L g3350 ( 
.A(n_2383),
.B(n_2409),
.Y(n_3350)
);

NAND2xp5_ASAP7_75t_L g3351 ( 
.A(n_2383),
.B(n_2409),
.Y(n_3351)
);

INVx1_ASAP7_75t_L g3352 ( 
.A(n_2411),
.Y(n_3352)
);

BUFx6f_ASAP7_75t_SL g3353 ( 
.A(n_2218),
.Y(n_3353)
);

INVx2_ASAP7_75t_L g3354 ( 
.A(n_2411),
.Y(n_3354)
);

INVx1_ASAP7_75t_L g3355 ( 
.A(n_2419),
.Y(n_3355)
);

OR2x6_ASAP7_75t_L g3356 ( 
.A(n_2242),
.B(n_2218),
.Y(n_3356)
);

NAND2x1p5_ASAP7_75t_L g3357 ( 
.A(n_2480),
.B(n_2487),
.Y(n_3357)
);

AOI22xp33_ASAP7_75t_L g3358 ( 
.A1(n_2089),
.A2(n_2097),
.B1(n_2099),
.B2(n_2093),
.Y(n_3358)
);

OAI21xp5_ASAP7_75t_L g3359 ( 
.A1(n_2141),
.A2(n_2148),
.B(n_2144),
.Y(n_3359)
);

NOR2xp33_ASAP7_75t_L g3360 ( 
.A(n_2649),
.B(n_2637),
.Y(n_3360)
);

NAND2xp5_ASAP7_75t_L g3361 ( 
.A(n_2429),
.B(n_2441),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_2441),
.Y(n_3362)
);

NAND2x1p5_ASAP7_75t_L g3363 ( 
.A(n_2480),
.B(n_2487),
.Y(n_3363)
);

OR2x2_ASAP7_75t_L g3364 ( 
.A(n_2217),
.B(n_2030),
.Y(n_3364)
);

INVx1_ASAP7_75t_L g3365 ( 
.A(n_2457),
.Y(n_3365)
);

OR2x6_ASAP7_75t_L g3366 ( 
.A(n_2218),
.B(n_2480),
.Y(n_3366)
);

INVx4_ASAP7_75t_L g3367 ( 
.A(n_2282),
.Y(n_3367)
);

INVx1_ASAP7_75t_L g3368 ( 
.A(n_2458),
.Y(n_3368)
);

HB1xp67_ASAP7_75t_L g3369 ( 
.A(n_2458),
.Y(n_3369)
);

INVx2_ASAP7_75t_SL g3370 ( 
.A(n_2282),
.Y(n_3370)
);

INVxp67_ASAP7_75t_L g3371 ( 
.A(n_2093),
.Y(n_3371)
);

INVx2_ASAP7_75t_L g3372 ( 
.A(n_2461),
.Y(n_3372)
);

INVx1_ASAP7_75t_L g3373 ( 
.A(n_2461),
.Y(n_3373)
);

BUFx5_ASAP7_75t_L g3374 ( 
.A(n_2198),
.Y(n_3374)
);

BUFx3_ASAP7_75t_L g3375 ( 
.A(n_2282),
.Y(n_3375)
);

NAND2xp5_ASAP7_75t_L g3376 ( 
.A(n_2473),
.B(n_2475),
.Y(n_3376)
);

INVx1_ASAP7_75t_L g3377 ( 
.A(n_2473),
.Y(n_3377)
);

INVx2_ASAP7_75t_L g3378 ( 
.A(n_2475),
.Y(n_3378)
);

INVx1_ASAP7_75t_L g3379 ( 
.A(n_2484),
.Y(n_3379)
);

BUFx3_ASAP7_75t_L g3380 ( 
.A(n_2282),
.Y(n_3380)
);

INVx1_ASAP7_75t_SL g3381 ( 
.A(n_2030),
.Y(n_3381)
);

INVx1_ASAP7_75t_L g3382 ( 
.A(n_2484),
.Y(n_3382)
);

INVxp67_ASAP7_75t_L g3383 ( 
.A(n_2097),
.Y(n_3383)
);

AOI22xp5_ASAP7_75t_L g3384 ( 
.A1(n_2064),
.A2(n_2078),
.B1(n_2115),
.B2(n_2092),
.Y(n_3384)
);

INVx2_ASAP7_75t_SL g3385 ( 
.A(n_2296),
.Y(n_3385)
);

INVx2_ASAP7_75t_L g3386 ( 
.A(n_2485),
.Y(n_3386)
);

INVx2_ASAP7_75t_L g3387 ( 
.A(n_2485),
.Y(n_3387)
);

INVx2_ASAP7_75t_SL g3388 ( 
.A(n_2296),
.Y(n_3388)
);

OAI21x1_ASAP7_75t_L g3389 ( 
.A1(n_2343),
.A2(n_2144),
.B(n_2141),
.Y(n_3389)
);

OR2x6_ASAP7_75t_L g3390 ( 
.A(n_2569),
.B(n_2296),
.Y(n_3390)
);

INVx2_ASAP7_75t_L g3391 ( 
.A(n_2492),
.Y(n_3391)
);

NAND2xp5_ASAP7_75t_SL g3392 ( 
.A(n_2033),
.B(n_2203),
.Y(n_3392)
);

INVx1_ASAP7_75t_L g3393 ( 
.A(n_2492),
.Y(n_3393)
);

NAND2xp5_ASAP7_75t_L g3394 ( 
.A(n_2499),
.B(n_2502),
.Y(n_3394)
);

OR2x6_ASAP7_75t_L g3395 ( 
.A(n_2569),
.B(n_2308),
.Y(n_3395)
);

INVx2_ASAP7_75t_SL g3396 ( 
.A(n_2308),
.Y(n_3396)
);

HB1xp67_ASAP7_75t_L g3397 ( 
.A(n_2499),
.Y(n_3397)
);

AND2x2_ASAP7_75t_SL g3398 ( 
.A(n_2241),
.B(n_2230),
.Y(n_3398)
);

INVx3_ASAP7_75t_L g3399 ( 
.A(n_2196),
.Y(n_3399)
);

AOI22xp33_ASAP7_75t_SL g3400 ( 
.A1(n_2007),
.A2(n_2017),
.B1(n_2073),
.B2(n_2045),
.Y(n_3400)
);

OAI22xp33_ASAP7_75t_L g3401 ( 
.A1(n_2099),
.A2(n_2103),
.B1(n_2106),
.B2(n_2100),
.Y(n_3401)
);

INVx3_ASAP7_75t_L g3402 ( 
.A(n_2196),
.Y(n_3402)
);

INVx2_ASAP7_75t_L g3403 ( 
.A(n_2502),
.Y(n_3403)
);

AND2x4_ASAP7_75t_SL g3404 ( 
.A(n_2308),
.B(n_2254),
.Y(n_3404)
);

NAND2xp5_ASAP7_75t_L g3405 ( 
.A(n_2506),
.B(n_2508),
.Y(n_3405)
);

INVxp67_ASAP7_75t_SL g3406 ( 
.A(n_2100),
.Y(n_3406)
);

BUFx6f_ASAP7_75t_L g3407 ( 
.A(n_2196),
.Y(n_3407)
);

HB1xp67_ASAP7_75t_L g3408 ( 
.A(n_2506),
.Y(n_3408)
);

AOI22xp5_ASAP7_75t_L g3409 ( 
.A1(n_2169),
.A2(n_2140),
.B1(n_2037),
.B2(n_2147),
.Y(n_3409)
);

INVx1_ASAP7_75t_L g3410 ( 
.A(n_2508),
.Y(n_3410)
);

BUFx6f_ASAP7_75t_L g3411 ( 
.A(n_2196),
.Y(n_3411)
);

BUFx2_ASAP7_75t_L g3412 ( 
.A(n_2110),
.Y(n_3412)
);

INVx1_ASAP7_75t_L g3413 ( 
.A(n_2524),
.Y(n_3413)
);

NAND2xp5_ASAP7_75t_L g3414 ( 
.A(n_2524),
.B(n_2533),
.Y(n_3414)
);

INVx3_ASAP7_75t_L g3415 ( 
.A(n_2196),
.Y(n_3415)
);

NAND2xp5_ASAP7_75t_SL g3416 ( 
.A(n_2293),
.B(n_2103),
.Y(n_3416)
);

INVx4_ASAP7_75t_L g3417 ( 
.A(n_2646),
.Y(n_3417)
);

INVx1_ASAP7_75t_L g3418 ( 
.A(n_2533),
.Y(n_3418)
);

NAND2xp5_ASAP7_75t_SL g3419 ( 
.A(n_2106),
.B(n_2117),
.Y(n_3419)
);

INVx2_ASAP7_75t_L g3420 ( 
.A(n_2550),
.Y(n_3420)
);

BUFx6f_ASAP7_75t_L g3421 ( 
.A(n_2196),
.Y(n_3421)
);

INVx2_ASAP7_75t_L g3422 ( 
.A(n_2550),
.Y(n_3422)
);

BUFx6f_ASAP7_75t_L g3423 ( 
.A(n_2342),
.Y(n_3423)
);

INVxp67_ASAP7_75t_L g3424 ( 
.A(n_2117),
.Y(n_3424)
);

INVx3_ASAP7_75t_L g3425 ( 
.A(n_2263),
.Y(n_3425)
);

BUFx6f_ASAP7_75t_L g3426 ( 
.A(n_2342),
.Y(n_3426)
);

INVx2_ASAP7_75t_SL g3427 ( 
.A(n_2254),
.Y(n_3427)
);

INVx2_ASAP7_75t_SL g3428 ( 
.A(n_2254),
.Y(n_3428)
);

NAND2xp5_ASAP7_75t_L g3429 ( 
.A(n_2568),
.B(n_2581),
.Y(n_3429)
);

INVxp67_ASAP7_75t_SL g3430 ( 
.A(n_2119),
.Y(n_3430)
);

INVx1_ASAP7_75t_L g3431 ( 
.A(n_2568),
.Y(n_3431)
);

INVx1_ASAP7_75t_L g3432 ( 
.A(n_2581),
.Y(n_3432)
);

BUFx6f_ASAP7_75t_L g3433 ( 
.A(n_2342),
.Y(n_3433)
);

BUFx4f_ASAP7_75t_L g3434 ( 
.A(n_2238),
.Y(n_3434)
);

A2O1A1Ixp33_ASAP7_75t_L g3435 ( 
.A1(n_2119),
.A2(n_2120),
.B(n_2063),
.C(n_2076),
.Y(n_3435)
);

BUFx8_ASAP7_75t_L g3436 ( 
.A(n_2646),
.Y(n_3436)
);

INVx1_ASAP7_75t_L g3437 ( 
.A(n_2607),
.Y(n_3437)
);

NAND2xp5_ASAP7_75t_L g3438 ( 
.A(n_2607),
.B(n_2611),
.Y(n_3438)
);

NAND2xp5_ASAP7_75t_L g3439 ( 
.A(n_2611),
.B(n_2635),
.Y(n_3439)
);

AND2x2_ASAP7_75t_L g3440 ( 
.A(n_2635),
.B(n_2642),
.Y(n_3440)
);

INVx5_ASAP7_75t_L g3441 ( 
.A(n_2238),
.Y(n_3441)
);

BUFx3_ASAP7_75t_L g3442 ( 
.A(n_2238),
.Y(n_3442)
);

NAND2xp5_ASAP7_75t_L g3443 ( 
.A(n_2642),
.B(n_2148),
.Y(n_3443)
);

INVx1_ASAP7_75t_L g3444 ( 
.A(n_2150),
.Y(n_3444)
);

NAND2xp5_ASAP7_75t_L g3445 ( 
.A(n_2150),
.B(n_2155),
.Y(n_3445)
);

NOR2xp33_ASAP7_75t_L g3446 ( 
.A(n_2400),
.B(n_2420),
.Y(n_3446)
);

NAND2xp5_ASAP7_75t_L g3447 ( 
.A(n_2155),
.B(n_2162),
.Y(n_3447)
);

HB1xp67_ASAP7_75t_L g3448 ( 
.A(n_2229),
.Y(n_3448)
);

INVx1_ASAP7_75t_L g3449 ( 
.A(n_2162),
.Y(n_3449)
);

NAND2xp5_ASAP7_75t_L g3450 ( 
.A(n_2165),
.B(n_2170),
.Y(n_3450)
);

INVx2_ASAP7_75t_L g3451 ( 
.A(n_2165),
.Y(n_3451)
);

INVx2_ASAP7_75t_SL g3452 ( 
.A(n_2254),
.Y(n_3452)
);

NOR2xp33_ASAP7_75t_L g3453 ( 
.A(n_2472),
.B(n_2552),
.Y(n_3453)
);

OR2x2_ASAP7_75t_SL g3454 ( 
.A(n_2238),
.B(n_2240),
.Y(n_3454)
);

INVx2_ASAP7_75t_SL g3455 ( 
.A(n_2276),
.Y(n_3455)
);

INVx2_ASAP7_75t_L g3456 ( 
.A(n_2170),
.Y(n_3456)
);

AO22x1_ASAP7_75t_L g3457 ( 
.A1(n_2091),
.A2(n_2190),
.B1(n_2261),
.B2(n_2264),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_2177),
.Y(n_3458)
);

HB1xp67_ASAP7_75t_L g3459 ( 
.A(n_2229),
.Y(n_3459)
);

OAI22xp5_ASAP7_75t_L g3460 ( 
.A1(n_2120),
.A2(n_2096),
.B1(n_2066),
.B2(n_2082),
.Y(n_3460)
);

HB1xp67_ASAP7_75t_L g3461 ( 
.A(n_2229),
.Y(n_3461)
);

AND2x4_ASAP7_75t_L g3462 ( 
.A(n_2198),
.B(n_2255),
.Y(n_3462)
);

NAND2xp5_ASAP7_75t_L g3463 ( 
.A(n_2177),
.B(n_2181),
.Y(n_3463)
);

INVx1_ASAP7_75t_L g3464 ( 
.A(n_2181),
.Y(n_3464)
);

INVx1_ASAP7_75t_L g3465 ( 
.A(n_2183),
.Y(n_3465)
);

AOI22xp5_ASAP7_75t_L g3466 ( 
.A1(n_2241),
.A2(n_2071),
.B1(n_2646),
.B2(n_2258),
.Y(n_3466)
);

NAND2xp5_ASAP7_75t_L g3467 ( 
.A(n_2183),
.B(n_2187),
.Y(n_3467)
);

CKINVDCx5p33_ASAP7_75t_R g3468 ( 
.A(n_2366),
.Y(n_3468)
);

INVx4_ASAP7_75t_L g3469 ( 
.A(n_2646),
.Y(n_3469)
);

AND3x1_ASAP7_75t_L g3470 ( 
.A(n_2007),
.B(n_2017),
.C(n_2247),
.Y(n_3470)
);

INVx2_ASAP7_75t_L g3471 ( 
.A(n_2187),
.Y(n_3471)
);

INVx1_ASAP7_75t_L g3472 ( 
.A(n_2191),
.Y(n_3472)
);

INVxp67_ASAP7_75t_L g3473 ( 
.A(n_2245),
.Y(n_3473)
);

NAND2xp5_ASAP7_75t_L g3474 ( 
.A(n_3406),
.B(n_2015),
.Y(n_3474)
);

HB1xp67_ASAP7_75t_L g3475 ( 
.A(n_3344),
.Y(n_3475)
);

OR2x2_ASAP7_75t_L g3476 ( 
.A(n_2704),
.B(n_2245),
.Y(n_3476)
);

OAI21xp33_ASAP7_75t_SL g3477 ( 
.A1(n_3188),
.A2(n_2195),
.B(n_2186),
.Y(n_3477)
);

AOI22xp33_ASAP7_75t_L g3478 ( 
.A1(n_2669),
.A2(n_1993),
.B1(n_1886),
.B2(n_2449),
.Y(n_3478)
);

BUFx6f_ASAP7_75t_L g3479 ( 
.A(n_3356),
.Y(n_3479)
);

O2A1O1Ixp33_ASAP7_75t_SL g3480 ( 
.A1(n_3210),
.A2(n_2275),
.B(n_2161),
.C(n_2111),
.Y(n_3480)
);

O2A1O1Ixp33_ASAP7_75t_L g3481 ( 
.A1(n_3210),
.A2(n_2136),
.B(n_2098),
.C(n_2142),
.Y(n_3481)
);

AOI21xp5_ASAP7_75t_L g3482 ( 
.A1(n_2700),
.A2(n_2710),
.B(n_2706),
.Y(n_3482)
);

AOI21xp5_ASAP7_75t_L g3483 ( 
.A1(n_2700),
.A2(n_2343),
.B(n_2191),
.Y(n_3483)
);

AOI21xp5_ASAP7_75t_L g3484 ( 
.A1(n_2700),
.A2(n_2213),
.B(n_2248),
.Y(n_3484)
);

NAND2xp5_ASAP7_75t_L g3485 ( 
.A(n_3406),
.B(n_2015),
.Y(n_3485)
);

INVx1_ASAP7_75t_L g3486 ( 
.A(n_2691),
.Y(n_3486)
);

OAI22xp5_ASAP7_75t_L g3487 ( 
.A1(n_2771),
.A2(n_2303),
.B1(n_2138),
.B2(n_2137),
.Y(n_3487)
);

O2A1O1Ixp33_ASAP7_75t_L g3488 ( 
.A1(n_2668),
.A2(n_2151),
.B(n_2130),
.C(n_2102),
.Y(n_3488)
);

AOI21xp5_ASAP7_75t_L g3489 ( 
.A1(n_2706),
.A2(n_2251),
.B(n_2051),
.Y(n_3489)
);

NAND2xp5_ASAP7_75t_SL g3490 ( 
.A(n_2960),
.B(n_2198),
.Y(n_3490)
);

CKINVDCx11_ASAP7_75t_R g3491 ( 
.A(n_2753),
.Y(n_3491)
);

AOI21xp5_ASAP7_75t_L g3492 ( 
.A1(n_2706),
.A2(n_2043),
.B(n_2123),
.Y(n_3492)
);

NAND2xp5_ASAP7_75t_L g3493 ( 
.A(n_3406),
.B(n_2016),
.Y(n_3493)
);

INVx2_ASAP7_75t_SL g3494 ( 
.A(n_3311),
.Y(n_3494)
);

AOI22x1_ASAP7_75t_L g3495 ( 
.A1(n_2820),
.A2(n_2176),
.B1(n_2341),
.B2(n_2245),
.Y(n_3495)
);

OR2x2_ASAP7_75t_L g3496 ( 
.A(n_2704),
.B(n_2194),
.Y(n_3496)
);

BUFx3_ASAP7_75t_L g3497 ( 
.A(n_2652),
.Y(n_3497)
);

AO22x1_ASAP7_75t_L g3498 ( 
.A1(n_3128),
.A2(n_2277),
.B1(n_1967),
.B2(n_2505),
.Y(n_3498)
);

NOR2xp67_ASAP7_75t_L g3499 ( 
.A(n_2775),
.B(n_2276),
.Y(n_3499)
);

INVx2_ASAP7_75t_L g3500 ( 
.A(n_2663),
.Y(n_3500)
);

BUFx8_ASAP7_75t_SL g3501 ( 
.A(n_2753),
.Y(n_3501)
);

NOR2xp67_ASAP7_75t_L g3502 ( 
.A(n_2775),
.B(n_2276),
.Y(n_3502)
);

BUFx3_ASAP7_75t_L g3503 ( 
.A(n_2652),
.Y(n_3503)
);

OAI21xp5_ASAP7_75t_L g3504 ( 
.A1(n_2669),
.A2(n_2032),
.B(n_2240),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_L g3505 ( 
.A(n_3430),
.B(n_2016),
.Y(n_3505)
);

NAND2xp5_ASAP7_75t_SL g3506 ( 
.A(n_2960),
.B(n_2198),
.Y(n_3506)
);

INVx2_ASAP7_75t_SL g3507 ( 
.A(n_3311),
.Y(n_3507)
);

OAI22xp5_ASAP7_75t_L g3508 ( 
.A1(n_2771),
.A2(n_2236),
.B1(n_2223),
.B2(n_2023),
.Y(n_3508)
);

OAI22xp5_ASAP7_75t_L g3509 ( 
.A1(n_2668),
.A2(n_2236),
.B1(n_2223),
.B2(n_2023),
.Y(n_3509)
);

O2A1O1Ixp33_ASAP7_75t_L g3510 ( 
.A1(n_2767),
.A2(n_2575),
.B(n_2039),
.C(n_2226),
.Y(n_3510)
);

NOR2xp33_ASAP7_75t_L g3511 ( 
.A(n_2867),
.B(n_2129),
.Y(n_3511)
);

NAND2xp5_ASAP7_75t_L g3512 ( 
.A(n_3430),
.B(n_2020),
.Y(n_3512)
);

INVx3_ASAP7_75t_SL g3513 ( 
.A(n_2654),
.Y(n_3513)
);

INVx2_ASAP7_75t_L g3514 ( 
.A(n_2663),
.Y(n_3514)
);

AOI33xp33_ASAP7_75t_L g3515 ( 
.A1(n_2696),
.A2(n_1855),
.A3(n_2540),
.B1(n_2531),
.B2(n_2613),
.B3(n_2081),
.Y(n_3515)
);

AOI21xp5_ASAP7_75t_L g3516 ( 
.A1(n_2710),
.A2(n_2124),
.B(n_2123),
.Y(n_3516)
);

NAND2xp5_ASAP7_75t_L g3517 ( 
.A(n_3430),
.B(n_2020),
.Y(n_3517)
);

AOI21xp5_ASAP7_75t_L g3518 ( 
.A1(n_2710),
.A2(n_2135),
.B(n_2124),
.Y(n_3518)
);

BUFx2_ASAP7_75t_L g3519 ( 
.A(n_2789),
.Y(n_3519)
);

INVxp67_ASAP7_75t_L g3520 ( 
.A(n_2811),
.Y(n_3520)
);

INVx1_ASAP7_75t_L g3521 ( 
.A(n_2691),
.Y(n_3521)
);

NAND2xp5_ASAP7_75t_L g3522 ( 
.A(n_2758),
.B(n_2135),
.Y(n_3522)
);

NAND2xp5_ASAP7_75t_L g3523 ( 
.A(n_2758),
.B(n_2139),
.Y(n_3523)
);

NOR2x1p5_ASAP7_75t_SL g3524 ( 
.A(n_2871),
.B(n_2225),
.Y(n_3524)
);

HB1xp67_ASAP7_75t_L g3525 ( 
.A(n_2894),
.Y(n_3525)
);

NAND2xp5_ASAP7_75t_L g3526 ( 
.A(n_2758),
.B(n_2139),
.Y(n_3526)
);

AND2x2_ASAP7_75t_L g3527 ( 
.A(n_3063),
.B(n_2153),
.Y(n_3527)
);

NOR2xp33_ASAP7_75t_L g3528 ( 
.A(n_2867),
.B(n_2154),
.Y(n_3528)
);

CKINVDCx20_ASAP7_75t_R g3529 ( 
.A(n_2947),
.Y(n_3529)
);

BUFx3_ASAP7_75t_L g3530 ( 
.A(n_2652),
.Y(n_3530)
);

HB1xp67_ASAP7_75t_L g3531 ( 
.A(n_3344),
.Y(n_3531)
);

NAND2xp5_ASAP7_75t_L g3532 ( 
.A(n_2787),
.B(n_2153),
.Y(n_3532)
);

A2O1A1Ixp33_ASAP7_75t_L g3533 ( 
.A1(n_2716),
.A2(n_2174),
.B(n_2185),
.C(n_2209),
.Y(n_3533)
);

NOR2xp67_ASAP7_75t_SL g3534 ( 
.A(n_3028),
.B(n_1967),
.Y(n_3534)
);

AND2x4_ASAP7_75t_SL g3535 ( 
.A(n_2769),
.B(n_2297),
.Y(n_3535)
);

OAI22xp5_ASAP7_75t_L g3536 ( 
.A1(n_2815),
.A2(n_2173),
.B1(n_2244),
.B2(n_2194),
.Y(n_3536)
);

NAND2xp5_ASAP7_75t_SL g3537 ( 
.A(n_2960),
.B(n_2255),
.Y(n_3537)
);

INVx2_ASAP7_75t_L g3538 ( 
.A(n_2663),
.Y(n_3538)
);

INVx1_ASAP7_75t_L g3539 ( 
.A(n_2691),
.Y(n_3539)
);

NAND2xp5_ASAP7_75t_L g3540 ( 
.A(n_2787),
.B(n_2175),
.Y(n_3540)
);

AOI22xp5_ASAP7_75t_L g3541 ( 
.A1(n_3034),
.A2(n_2255),
.B1(n_2258),
.B2(n_2237),
.Y(n_3541)
);

OAI22xp5_ASAP7_75t_L g3542 ( 
.A1(n_2815),
.A2(n_2244),
.B1(n_2204),
.B2(n_2239),
.Y(n_3542)
);

NAND2xp5_ASAP7_75t_L g3543 ( 
.A(n_2939),
.B(n_2175),
.Y(n_3543)
);

NAND2xp5_ASAP7_75t_L g3544 ( 
.A(n_2939),
.B(n_2204),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_2691),
.Y(n_3545)
);

OAI22xp5_ASAP7_75t_L g3546 ( 
.A1(n_2815),
.A2(n_2231),
.B1(n_2321),
.B2(n_2307),
.Y(n_3546)
);

AOI21xp5_ASAP7_75t_L g3547 ( 
.A1(n_2763),
.A2(n_2314),
.B(n_2200),
.Y(n_3547)
);

NOR2xp33_ASAP7_75t_L g3548 ( 
.A(n_2689),
.B(n_2158),
.Y(n_3548)
);

OAI21xp5_ASAP7_75t_L g3549 ( 
.A1(n_2696),
.A2(n_2250),
.B(n_2197),
.Y(n_3549)
);

OAI22xp5_ASAP7_75t_L g3550 ( 
.A1(n_2689),
.A2(n_2304),
.B1(n_1998),
.B2(n_2346),
.Y(n_3550)
);

NOR2xp33_ASAP7_75t_SL g3551 ( 
.A(n_3143),
.B(n_2224),
.Y(n_3551)
);

AOI21xp5_ASAP7_75t_L g3552 ( 
.A1(n_2763),
.A2(n_2666),
.B(n_2655),
.Y(n_3552)
);

NOR2xp33_ASAP7_75t_L g3553 ( 
.A(n_2719),
.B(n_2029),
.Y(n_3553)
);

AOI22x1_ASAP7_75t_L g3554 ( 
.A1(n_2820),
.A2(n_2341),
.B1(n_2212),
.B2(n_2220),
.Y(n_3554)
);

A2O1A1Ixp33_ASAP7_75t_L g3555 ( 
.A1(n_2716),
.A2(n_1987),
.B(n_1980),
.C(n_1979),
.Y(n_3555)
);

AOI21xp5_ASAP7_75t_L g3556 ( 
.A1(n_2763),
.A2(n_2202),
.B(n_2200),
.Y(n_3556)
);

INVx2_ASAP7_75t_SL g3557 ( 
.A(n_3311),
.Y(n_3557)
);

NAND2xp5_ASAP7_75t_L g3558 ( 
.A(n_2939),
.B(n_3195),
.Y(n_3558)
);

INVx2_ASAP7_75t_L g3559 ( 
.A(n_2663),
.Y(n_3559)
);

BUFx4f_ASAP7_75t_L g3560 ( 
.A(n_3188),
.Y(n_3560)
);

INVx2_ASAP7_75t_L g3561 ( 
.A(n_2663),
.Y(n_3561)
);

NAND2xp5_ASAP7_75t_SL g3562 ( 
.A(n_3034),
.B(n_2255),
.Y(n_3562)
);

AOI21xp5_ASAP7_75t_L g3563 ( 
.A1(n_2655),
.A2(n_2197),
.B(n_2202),
.Y(n_3563)
);

AND2x2_ASAP7_75t_SL g3564 ( 
.A(n_2679),
.B(n_2258),
.Y(n_3564)
);

OAI22xp5_ASAP7_75t_L g3565 ( 
.A1(n_2719),
.A2(n_1855),
.B1(n_2540),
.B2(n_2531),
.Y(n_3565)
);

OAI22xp5_ASAP7_75t_L g3566 ( 
.A1(n_2765),
.A2(n_2804),
.B1(n_2701),
.B2(n_2818),
.Y(n_3566)
);

AND2x2_ASAP7_75t_L g3567 ( 
.A(n_3063),
.B(n_2318),
.Y(n_3567)
);

OAI21xp5_ASAP7_75t_L g3568 ( 
.A1(n_2775),
.A2(n_2250),
.B(n_2299),
.Y(n_3568)
);

NAND2xp5_ASAP7_75t_L g3569 ( 
.A(n_3195),
.B(n_2215),
.Y(n_3569)
);

AO21x1_ASAP7_75t_L g3570 ( 
.A1(n_3019),
.A2(n_2265),
.B(n_2262),
.Y(n_3570)
);

NAND2xp5_ASAP7_75t_L g3571 ( 
.A(n_3196),
.B(n_3195),
.Y(n_3571)
);

OR2x6_ASAP7_75t_SL g3572 ( 
.A(n_2666),
.B(n_2261),
.Y(n_3572)
);

OAI22xp5_ASAP7_75t_L g3573 ( 
.A1(n_2765),
.A2(n_2613),
.B1(n_2081),
.B2(n_2012),
.Y(n_3573)
);

NAND2xp5_ASAP7_75t_SL g3574 ( 
.A(n_3034),
.B(n_2258),
.Y(n_3574)
);

NOR2xp33_ASAP7_75t_L g3575 ( 
.A(n_2804),
.B(n_2085),
.Y(n_3575)
);

INVx2_ASAP7_75t_L g3576 ( 
.A(n_2664),
.Y(n_3576)
);

NAND3xp33_ASAP7_75t_L g3577 ( 
.A(n_2944),
.B(n_2963),
.C(n_2825),
.Y(n_3577)
);

NAND2xp5_ASAP7_75t_SL g3578 ( 
.A(n_2944),
.B(n_2012),
.Y(n_3578)
);

BUFx6f_ASAP7_75t_L g3579 ( 
.A(n_3356),
.Y(n_3579)
);

OAI22xp5_ASAP7_75t_SL g3580 ( 
.A1(n_2818),
.A2(n_2080),
.B1(n_2152),
.B2(n_2113),
.Y(n_3580)
);

INVx2_ASAP7_75t_L g3581 ( 
.A(n_2664),
.Y(n_3581)
);

NOR2xp33_ASAP7_75t_SL g3582 ( 
.A(n_3143),
.B(n_2224),
.Y(n_3582)
);

OAI22xp5_ASAP7_75t_L g3583 ( 
.A1(n_2701),
.A2(n_2080),
.B1(n_2297),
.B2(n_2299),
.Y(n_3583)
);

NAND2xp5_ASAP7_75t_SL g3584 ( 
.A(n_2963),
.B(n_2206),
.Y(n_3584)
);

O2A1O1Ixp5_ASAP7_75t_L g3585 ( 
.A1(n_3149),
.A2(n_2705),
.B(n_2720),
.C(n_2715),
.Y(n_3585)
);

INVx6_ASAP7_75t_L g3586 ( 
.A(n_2652),
.Y(n_3586)
);

OAI21x1_ASAP7_75t_L g3587 ( 
.A1(n_3190),
.A2(n_2220),
.B(n_2215),
.Y(n_3587)
);

AND2x2_ASAP7_75t_L g3588 ( 
.A(n_3063),
.B(n_2833),
.Y(n_3588)
);

NAND2xp5_ASAP7_75t_SL g3589 ( 
.A(n_3042),
.B(n_2206),
.Y(n_3589)
);

NAND2xp5_ASAP7_75t_SL g3590 ( 
.A(n_3042),
.B(n_2211),
.Y(n_3590)
);

AND2x2_ASAP7_75t_SL g3591 ( 
.A(n_2679),
.B(n_2680),
.Y(n_3591)
);

AOI21xp5_ASAP7_75t_L g3592 ( 
.A1(n_2666),
.A2(n_2028),
.B(n_2031),
.Y(n_3592)
);

NAND2xp5_ASAP7_75t_L g3593 ( 
.A(n_3196),
.B(n_2225),
.Y(n_3593)
);

AOI22xp5_ASAP7_75t_L g3594 ( 
.A1(n_2941),
.A2(n_2246),
.B1(n_2268),
.B2(n_2211),
.Y(n_3594)
);

NAND2xp5_ASAP7_75t_L g3595 ( 
.A(n_3196),
.B(n_2959),
.Y(n_3595)
);

AOI21xp5_ASAP7_75t_L g3596 ( 
.A1(n_3160),
.A2(n_2270),
.B(n_2048),
.Y(n_3596)
);

NOR2xp33_ASAP7_75t_L g3597 ( 
.A(n_2711),
.B(n_2167),
.Y(n_3597)
);

AND2x6_ASAP7_75t_L g3598 ( 
.A(n_2769),
.B(n_2276),
.Y(n_3598)
);

AOI21xp5_ASAP7_75t_L g3599 ( 
.A1(n_3160),
.A2(n_2681),
.B(n_2678),
.Y(n_3599)
);

AOI22xp33_ASAP7_75t_L g3600 ( 
.A1(n_2705),
.A2(n_2720),
.B1(n_2795),
.B2(n_2715),
.Y(n_3600)
);

A2O1A1Ixp33_ASAP7_75t_L g3601 ( 
.A1(n_2716),
.A2(n_1967),
.B(n_1981),
.C(n_2505),
.Y(n_3601)
);

O2A1O1Ixp33_ASAP7_75t_L g3602 ( 
.A1(n_2767),
.A2(n_2265),
.B(n_2257),
.C(n_2262),
.Y(n_3602)
);

AND2x2_ASAP7_75t_L g3603 ( 
.A(n_3063),
.B(n_2318),
.Y(n_3603)
);

AOI21xp5_ASAP7_75t_L g3604 ( 
.A1(n_2678),
.A2(n_2270),
.B(n_2048),
.Y(n_3604)
);

OAI22xp5_ASAP7_75t_L g3605 ( 
.A1(n_2890),
.A2(n_2896),
.B1(n_2739),
.B2(n_2773),
.Y(n_3605)
);

INVx2_ASAP7_75t_L g3606 ( 
.A(n_2664),
.Y(n_3606)
);

AOI21xp5_ASAP7_75t_L g3607 ( 
.A1(n_2678),
.A2(n_2132),
.B(n_2225),
.Y(n_3607)
);

OR2x2_ASAP7_75t_L g3608 ( 
.A(n_2704),
.B(n_2257),
.Y(n_3608)
);

INVx2_ASAP7_75t_L g3609 ( 
.A(n_2664),
.Y(n_3609)
);

NOR2xp33_ASAP7_75t_SL g3610 ( 
.A(n_3434),
.B(n_2224),
.Y(n_3610)
);

INVx1_ASAP7_75t_L g3611 ( 
.A(n_2693),
.Y(n_3611)
);

BUFx6f_ASAP7_75t_L g3612 ( 
.A(n_3356),
.Y(n_3612)
);

INVx2_ASAP7_75t_L g3613 ( 
.A(n_2664),
.Y(n_3613)
);

INVx1_ASAP7_75t_L g3614 ( 
.A(n_2693),
.Y(n_3614)
);

CKINVDCx5p33_ASAP7_75t_R g3615 ( 
.A(n_2749),
.Y(n_3615)
);

AND2x2_ASAP7_75t_L g3616 ( 
.A(n_2833),
.B(n_2318),
.Y(n_3616)
);

CKINVDCx16_ASAP7_75t_R g3617 ( 
.A(n_2749),
.Y(n_3617)
);

INVx3_ASAP7_75t_L g3618 ( 
.A(n_2712),
.Y(n_3618)
);

O2A1O1Ixp33_ASAP7_75t_L g3619 ( 
.A1(n_3149),
.A2(n_2260),
.B(n_2259),
.C(n_2246),
.Y(n_3619)
);

BUFx3_ASAP7_75t_L g3620 ( 
.A(n_2652),
.Y(n_3620)
);

AOI22xp5_ASAP7_75t_L g3621 ( 
.A1(n_2941),
.A2(n_2219),
.B1(n_2227),
.B2(n_2274),
.Y(n_3621)
);

OAI21xp33_ASAP7_75t_L g3622 ( 
.A1(n_2825),
.A2(n_1981),
.B(n_2108),
.Y(n_3622)
);

NOR2xp33_ASAP7_75t_L g3623 ( 
.A(n_2711),
.B(n_3202),
.Y(n_3623)
);

AOI21xp5_ASAP7_75t_L g3624 ( 
.A1(n_2681),
.A2(n_3190),
.B(n_3401),
.Y(n_3624)
);

NAND2xp5_ASAP7_75t_SL g3625 ( 
.A(n_2942),
.B(n_2274),
.Y(n_3625)
);

OR2x6_ASAP7_75t_L g3626 ( 
.A(n_3356),
.B(n_2212),
.Y(n_3626)
);

NOR2xp33_ASAP7_75t_L g3627 ( 
.A(n_2711),
.B(n_3202),
.Y(n_3627)
);

HB1xp67_ASAP7_75t_L g3628 ( 
.A(n_3344),
.Y(n_3628)
);

NAND2xp5_ASAP7_75t_L g3629 ( 
.A(n_2959),
.B(n_2328),
.Y(n_3629)
);

OR2x6_ASAP7_75t_L g3630 ( 
.A(n_3356),
.B(n_2212),
.Y(n_3630)
);

NOR2xp33_ASAP7_75t_L g3631 ( 
.A(n_3320),
.B(n_2260),
.Y(n_3631)
);

NAND2xp5_ASAP7_75t_L g3632 ( 
.A(n_3176),
.B(n_2328),
.Y(n_3632)
);

NAND2xp5_ASAP7_75t_L g3633 ( 
.A(n_3176),
.B(n_2328),
.Y(n_3633)
);

NAND2xp5_ASAP7_75t_SL g3634 ( 
.A(n_2942),
.B(n_2264),
.Y(n_3634)
);

NOR2x1_ASAP7_75t_L g3635 ( 
.A(n_3401),
.B(n_2513),
.Y(n_3635)
);

AOI33xp33_ASAP7_75t_L g3636 ( 
.A1(n_2907),
.A2(n_2338),
.A3(n_2278),
.B1(n_2201),
.B2(n_2319),
.B3(n_2330),
.Y(n_3636)
);

AOI21xp5_ASAP7_75t_L g3637 ( 
.A1(n_3190),
.A2(n_2201),
.B(n_2331),
.Y(n_3637)
);

AOI21xp5_ASAP7_75t_L g3638 ( 
.A1(n_2699),
.A2(n_2336),
.B(n_2317),
.Y(n_3638)
);

BUFx6f_ASAP7_75t_L g3639 ( 
.A(n_3356),
.Y(n_3639)
);

NAND2xp5_ASAP7_75t_SL g3640 ( 
.A(n_2942),
.B(n_1981),
.Y(n_3640)
);

INVx2_ASAP7_75t_L g3641 ( 
.A(n_2690),
.Y(n_3641)
);

NAND2xp5_ASAP7_75t_SL g3642 ( 
.A(n_3239),
.B(n_2108),
.Y(n_3642)
);

OAI22xp5_ASAP7_75t_L g3643 ( 
.A1(n_2890),
.A2(n_2108),
.B1(n_2126),
.B2(n_2145),
.Y(n_3643)
);

INVx2_ASAP7_75t_L g3644 ( 
.A(n_2690),
.Y(n_3644)
);

NOR3xp33_ASAP7_75t_L g3645 ( 
.A(n_2807),
.B(n_2259),
.C(n_2294),
.Y(n_3645)
);

AOI21xp5_ASAP7_75t_L g3646 ( 
.A1(n_2699),
.A2(n_2339),
.B(n_2316),
.Y(n_3646)
);

NAND2x1p5_ASAP7_75t_L g3647 ( 
.A(n_3311),
.B(n_2126),
.Y(n_3647)
);

INVx2_ASAP7_75t_L g3648 ( 
.A(n_2690),
.Y(n_3648)
);

NAND2xp5_ASAP7_75t_SL g3649 ( 
.A(n_3239),
.B(n_2126),
.Y(n_3649)
);

OAI21xp33_ASAP7_75t_SL g3650 ( 
.A1(n_3188),
.A2(n_2309),
.B(n_2320),
.Y(n_3650)
);

NAND2xp5_ASAP7_75t_L g3651 ( 
.A(n_3016),
.B(n_2344),
.Y(n_3651)
);

INVx2_ASAP7_75t_L g3652 ( 
.A(n_2690),
.Y(n_3652)
);

O2A1O1Ixp33_ASAP7_75t_SL g3653 ( 
.A1(n_3314),
.A2(n_2315),
.B(n_2334),
.C(n_2273),
.Y(n_3653)
);

NAND2xp5_ASAP7_75t_L g3654 ( 
.A(n_3016),
.B(n_2344),
.Y(n_3654)
);

NAND2xp5_ASAP7_75t_SL g3655 ( 
.A(n_3239),
.B(n_2145),
.Y(n_3655)
);

NAND2xp5_ASAP7_75t_L g3656 ( 
.A(n_3016),
.B(n_2344),
.Y(n_3656)
);

INVx2_ASAP7_75t_SL g3657 ( 
.A(n_3311),
.Y(n_3657)
);

AOI21xp5_ASAP7_75t_L g3658 ( 
.A1(n_3138),
.A2(n_2313),
.B(n_2335),
.Y(n_3658)
);

AOI22xp5_ASAP7_75t_L g3659 ( 
.A1(n_2732),
.A2(n_2235),
.B1(n_2145),
.B2(n_2505),
.Y(n_3659)
);

OAI21xp5_ASAP7_75t_L g3660 ( 
.A1(n_2653),
.A2(n_2313),
.B(n_2273),
.Y(n_3660)
);

NAND3xp33_ASAP7_75t_L g3661 ( 
.A(n_2907),
.B(n_2513),
.C(n_2437),
.Y(n_3661)
);

NOR3xp33_ASAP7_75t_L g3662 ( 
.A(n_2807),
.B(n_2315),
.C(n_2337),
.Y(n_3662)
);

AOI21xp5_ASAP7_75t_L g3663 ( 
.A1(n_3138),
.A2(n_2302),
.B(n_2334),
.Y(n_3663)
);

NAND2xp5_ASAP7_75t_L g3664 ( 
.A(n_3146),
.B(n_2326),
.Y(n_3664)
);

O2A1O1Ixp5_ASAP7_75t_L g3665 ( 
.A1(n_2795),
.A2(n_2808),
.B(n_3056),
.C(n_3307),
.Y(n_3665)
);

AND2x2_ASAP7_75t_L g3666 ( 
.A(n_2833),
.B(n_2326),
.Y(n_3666)
);

HB1xp67_ASAP7_75t_L g3667 ( 
.A(n_2894),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_SL g3668 ( 
.A(n_3400),
.B(n_2437),
.Y(n_3668)
);

NAND2xp5_ASAP7_75t_L g3669 ( 
.A(n_3146),
.B(n_2326),
.Y(n_3669)
);

BUFx6f_ASAP7_75t_L g3670 ( 
.A(n_3356),
.Y(n_3670)
);

AOI22xp33_ASAP7_75t_L g3671 ( 
.A1(n_2808),
.A2(n_2513),
.B1(n_2437),
.B2(n_2398),
.Y(n_3671)
);

AOI21xp5_ASAP7_75t_L g3672 ( 
.A1(n_3337),
.A2(n_2294),
.B(n_2332),
.Y(n_3672)
);

INVx1_ASAP7_75t_L g3673 ( 
.A(n_2693),
.Y(n_3673)
);

NAND2xp5_ASAP7_75t_L g3674 ( 
.A(n_3146),
.B(n_2330),
.Y(n_3674)
);

AOI21xp5_ASAP7_75t_L g3675 ( 
.A1(n_3337),
.A2(n_2295),
.B(n_2332),
.Y(n_3675)
);

AND2x4_ASAP7_75t_L g3676 ( 
.A(n_2714),
.B(n_2398),
.Y(n_3676)
);

AOI22xp33_ASAP7_75t_L g3677 ( 
.A1(n_2860),
.A2(n_2398),
.B1(n_2319),
.B2(n_2235),
.Y(n_3677)
);

AOI21xp5_ASAP7_75t_L g3678 ( 
.A1(n_3337),
.A2(n_2302),
.B(n_2327),
.Y(n_3678)
);

NAND2xp5_ASAP7_75t_L g3679 ( 
.A(n_3152),
.B(n_2278),
.Y(n_3679)
);

NAND2xp5_ASAP7_75t_L g3680 ( 
.A(n_3152),
.B(n_2301),
.Y(n_3680)
);

NOR2xp33_ASAP7_75t_L g3681 ( 
.A(n_3320),
.B(n_2301),
.Y(n_3681)
);

AOI21xp5_ASAP7_75t_L g3682 ( 
.A1(n_3337),
.A2(n_2337),
.B(n_2335),
.Y(n_3682)
);

NOR2xp33_ASAP7_75t_L g3683 ( 
.A(n_3360),
.B(n_2295),
.Y(n_3683)
);

AOI21xp5_ASAP7_75t_L g3684 ( 
.A1(n_3337),
.A2(n_2291),
.B(n_2333),
.Y(n_3684)
);

BUFx6f_ASAP7_75t_L g3685 ( 
.A(n_3356),
.Y(n_3685)
);

NOR2xp33_ASAP7_75t_L g3686 ( 
.A(n_3360),
.B(n_2291),
.Y(n_3686)
);

OAI21xp33_ASAP7_75t_L g3687 ( 
.A1(n_2733),
.A2(n_2896),
.B(n_2877),
.Y(n_3687)
);

AOI21xp5_ASAP7_75t_L g3688 ( 
.A1(n_3337),
.A2(n_2333),
.B(n_2324),
.Y(n_3688)
);

AOI21xp5_ASAP7_75t_L g3689 ( 
.A1(n_3337),
.A2(n_2290),
.B(n_2324),
.Y(n_3689)
);

INVx2_ASAP7_75t_L g3690 ( 
.A(n_3268),
.Y(n_3690)
);

INVx1_ASAP7_75t_L g3691 ( 
.A(n_2693),
.Y(n_3691)
);

NAND2xp5_ASAP7_75t_L g3692 ( 
.A(n_3152),
.B(n_2290),
.Y(n_3692)
);

BUFx6f_ASAP7_75t_L g3693 ( 
.A(n_3356),
.Y(n_3693)
);

NAND2xp5_ASAP7_75t_L g3694 ( 
.A(n_2661),
.B(n_2289),
.Y(n_3694)
);

NOR2xp33_ASAP7_75t_L g3695 ( 
.A(n_2947),
.B(n_2289),
.Y(n_3695)
);

CKINVDCx14_ASAP7_75t_R g3696 ( 
.A(n_2717),
.Y(n_3696)
);

AOI22x1_ASAP7_75t_L g3697 ( 
.A1(n_2820),
.A2(n_3100),
.B1(n_3118),
.B2(n_3019),
.Y(n_3697)
);

AO21x1_ASAP7_75t_L g3698 ( 
.A1(n_3019),
.A2(n_2323),
.B(n_2322),
.Y(n_3698)
);

AO32x1_ASAP7_75t_L g3699 ( 
.A1(n_2658),
.A2(n_2280),
.A3(n_2320),
.B1(n_2309),
.B2(n_2345),
.Y(n_3699)
);

NAND2xp5_ASAP7_75t_SL g3700 ( 
.A(n_3400),
.B(n_2323),
.Y(n_3700)
);

NAND2x1p5_ASAP7_75t_L g3701 ( 
.A(n_3311),
.B(n_2280),
.Y(n_3701)
);

BUFx2_ASAP7_75t_L g3702 ( 
.A(n_2789),
.Y(n_3702)
);

OR2x6_ASAP7_75t_L g3703 ( 
.A(n_3337),
.B(n_2280),
.Y(n_3703)
);

BUFx3_ASAP7_75t_L g3704 ( 
.A(n_2652),
.Y(n_3704)
);

INVx1_ASAP7_75t_L g3705 ( 
.A(n_2693),
.Y(n_3705)
);

AOI21xp5_ASAP7_75t_L g3706 ( 
.A1(n_3314),
.A2(n_2287),
.B(n_2284),
.Y(n_3706)
);

NAND2xp5_ASAP7_75t_L g3707 ( 
.A(n_2661),
.B(n_2287),
.Y(n_3707)
);

NAND2xp5_ASAP7_75t_SL g3708 ( 
.A(n_3400),
.B(n_2288),
.Y(n_3708)
);

AOI21xp5_ASAP7_75t_L g3709 ( 
.A1(n_3116),
.A2(n_2310),
.B(n_2285),
.Y(n_3709)
);

O2A1O1Ixp5_ASAP7_75t_L g3710 ( 
.A1(n_3056),
.A2(n_2285),
.B(n_2286),
.C(n_2322),
.Y(n_3710)
);

INVx1_ASAP7_75t_SL g3711 ( 
.A(n_3412),
.Y(n_3711)
);

A2O1A1Ixp33_ASAP7_75t_L g3712 ( 
.A1(n_2733),
.A2(n_2320),
.B(n_2281),
.C(n_2325),
.Y(n_3712)
);

O2A1O1Ixp33_ASAP7_75t_L g3713 ( 
.A1(n_3144),
.A2(n_2286),
.B(n_2281),
.C(n_2325),
.Y(n_3713)
);

NOR2xp33_ASAP7_75t_L g3714 ( 
.A(n_3468),
.B(n_2345),
.Y(n_3714)
);

BUFx6f_ASAP7_75t_L g3715 ( 
.A(n_2769),
.Y(n_3715)
);

AOI21x1_ASAP7_75t_L g3716 ( 
.A1(n_2757),
.A2(n_3457),
.B(n_3045),
.Y(n_3716)
);

NAND2xp5_ASAP7_75t_L g3717 ( 
.A(n_2665),
.B(n_2667),
.Y(n_3717)
);

INVx6_ASAP7_75t_L g3718 ( 
.A(n_2652),
.Y(n_3718)
);

NOR2xp33_ASAP7_75t_L g3719 ( 
.A(n_3468),
.B(n_3010),
.Y(n_3719)
);

INVx2_ASAP7_75t_SL g3720 ( 
.A(n_3311),
.Y(n_3720)
);

INVx3_ASAP7_75t_L g3721 ( 
.A(n_2712),
.Y(n_3721)
);

INVx1_ASAP7_75t_SL g3722 ( 
.A(n_3412),
.Y(n_3722)
);

BUFx2_ASAP7_75t_L g3723 ( 
.A(n_2789),
.Y(n_3723)
);

AOI21x1_ASAP7_75t_L g3724 ( 
.A1(n_2757),
.A2(n_3457),
.B(n_3045),
.Y(n_3724)
);

O2A1O1Ixp5_ASAP7_75t_L g3725 ( 
.A1(n_3056),
.A2(n_3307),
.B(n_2807),
.C(n_3045),
.Y(n_3725)
);

AND2x2_ASAP7_75t_L g3726 ( 
.A(n_2835),
.B(n_3055),
.Y(n_3726)
);

AO32x2_ASAP7_75t_L g3727 ( 
.A1(n_2658),
.A2(n_2697),
.A3(n_3008),
.B1(n_3229),
.B2(n_2872),
.Y(n_3727)
);

AO32x2_ASAP7_75t_L g3728 ( 
.A1(n_2658),
.A2(n_2697),
.A3(n_3008),
.B1(n_3229),
.B2(n_2872),
.Y(n_3728)
);

OAI22xp5_ASAP7_75t_L g3729 ( 
.A1(n_2739),
.A2(n_2773),
.B1(n_3384),
.B2(n_3232),
.Y(n_3729)
);

NAND2xp5_ASAP7_75t_SL g3730 ( 
.A(n_3206),
.B(n_2931),
.Y(n_3730)
);

NAND2x1p5_ASAP7_75t_L g3731 ( 
.A(n_3311),
.B(n_3155),
.Y(n_3731)
);

NAND2xp5_ASAP7_75t_L g3732 ( 
.A(n_2667),
.B(n_2671),
.Y(n_3732)
);

BUFx4f_ASAP7_75t_L g3733 ( 
.A(n_3188),
.Y(n_3733)
);

NAND2xp5_ASAP7_75t_SL g3734 ( 
.A(n_3206),
.B(n_2931),
.Y(n_3734)
);

NAND2xp5_ASAP7_75t_L g3735 ( 
.A(n_2671),
.B(n_2675),
.Y(n_3735)
);

AOI21xp5_ASAP7_75t_L g3736 ( 
.A1(n_3116),
.A2(n_2680),
.B(n_2679),
.Y(n_3736)
);

AOI22xp33_ASAP7_75t_L g3737 ( 
.A1(n_2860),
.A2(n_2877),
.B1(n_3229),
.B2(n_2935),
.Y(n_3737)
);

AND2x4_ASAP7_75t_L g3738 ( 
.A(n_2714),
.B(n_2724),
.Y(n_3738)
);

BUFx2_ASAP7_75t_L g3739 ( 
.A(n_2657),
.Y(n_3739)
);

AO21x1_ASAP7_75t_L g3740 ( 
.A1(n_3118),
.A2(n_3204),
.B(n_2738),
.Y(n_3740)
);

AOI21xp5_ASAP7_75t_L g3741 ( 
.A1(n_3116),
.A2(n_2680),
.B(n_3179),
.Y(n_3741)
);

NOR2xp33_ASAP7_75t_L g3742 ( 
.A(n_3010),
.B(n_3114),
.Y(n_3742)
);

O2A1O1Ixp33_ASAP7_75t_L g3743 ( 
.A1(n_3144),
.A2(n_2935),
.B(n_3184),
.C(n_3151),
.Y(n_3743)
);

INVx4_ASAP7_75t_L g3744 ( 
.A(n_3441),
.Y(n_3744)
);

O2A1O1Ixp5_ASAP7_75t_L g3745 ( 
.A1(n_3118),
.A2(n_2757),
.B(n_3416),
.C(n_2868),
.Y(n_3745)
);

NAND2xp5_ASAP7_75t_SL g3746 ( 
.A(n_3242),
.B(n_2653),
.Y(n_3746)
);

NAND2xp5_ASAP7_75t_L g3747 ( 
.A(n_2671),
.B(n_2675),
.Y(n_3747)
);

AOI21xp5_ASAP7_75t_L g3748 ( 
.A1(n_3116),
.A2(n_3179),
.B(n_3230),
.Y(n_3748)
);

AO32x2_ASAP7_75t_L g3749 ( 
.A1(n_2658),
.A2(n_2697),
.A3(n_3008),
.B1(n_2872),
.B2(n_2865),
.Y(n_3749)
);

BUFx6f_ASAP7_75t_L g3750 ( 
.A(n_2769),
.Y(n_3750)
);

NAND2xp5_ASAP7_75t_L g3751 ( 
.A(n_2675),
.B(n_2683),
.Y(n_3751)
);

AOI21xp5_ASAP7_75t_L g3752 ( 
.A1(n_3116),
.A2(n_3179),
.B(n_3230),
.Y(n_3752)
);

CKINVDCx5p33_ASAP7_75t_R g3753 ( 
.A(n_2717),
.Y(n_3753)
);

INVx1_ASAP7_75t_SL g3754 ( 
.A(n_3412),
.Y(n_3754)
);

AOI21xp5_ASAP7_75t_L g3755 ( 
.A1(n_3116),
.A2(n_3179),
.B(n_3230),
.Y(n_3755)
);

AOI22xp5_ASAP7_75t_L g3756 ( 
.A1(n_2732),
.A2(n_2766),
.B1(n_2733),
.B2(n_2739),
.Y(n_3756)
);

OAI22xp5_ASAP7_75t_L g3757 ( 
.A1(n_2773),
.A2(n_3384),
.B1(n_3232),
.B2(n_2766),
.Y(n_3757)
);

BUFx6f_ASAP7_75t_L g3758 ( 
.A(n_2769),
.Y(n_3758)
);

O2A1O1Ixp33_ASAP7_75t_L g3759 ( 
.A1(n_2935),
.A2(n_3151),
.B(n_3184),
.C(n_3068),
.Y(n_3759)
);

NAND2x1p5_ASAP7_75t_L g3760 ( 
.A(n_3311),
.B(n_3155),
.Y(n_3760)
);

O2A1O1Ixp33_ASAP7_75t_SL g3761 ( 
.A1(n_3128),
.A2(n_3232),
.B(n_3435),
.C(n_3416),
.Y(n_3761)
);

AOI22xp5_ASAP7_75t_L g3762 ( 
.A1(n_2766),
.A2(n_2713),
.B1(n_2707),
.B2(n_2653),
.Y(n_3762)
);

OR2x2_ASAP7_75t_L g3763 ( 
.A(n_2704),
.B(n_2709),
.Y(n_3763)
);

NAND2xp5_ASAP7_75t_SL g3764 ( 
.A(n_3242),
.B(n_2707),
.Y(n_3764)
);

AOI21xp5_ASAP7_75t_L g3765 ( 
.A1(n_3116),
.A2(n_3179),
.B(n_2682),
.Y(n_3765)
);

AOI21xp5_ASAP7_75t_L g3766 ( 
.A1(n_3116),
.A2(n_3179),
.B(n_2682),
.Y(n_3766)
);

AOI21xp5_ASAP7_75t_L g3767 ( 
.A1(n_3179),
.A2(n_2682),
.B(n_3204),
.Y(n_3767)
);

AOI21xp5_ASAP7_75t_L g3768 ( 
.A1(n_2682),
.A2(n_3158),
.B(n_3134),
.Y(n_3768)
);

NAND2xp5_ASAP7_75t_L g3769 ( 
.A(n_2683),
.B(n_2686),
.Y(n_3769)
);

NAND3xp33_ASAP7_75t_L g3770 ( 
.A(n_2707),
.B(n_3068),
.C(n_2738),
.Y(n_3770)
);

OAI22xp5_ASAP7_75t_L g3771 ( 
.A1(n_3384),
.A2(n_2897),
.B1(n_2909),
.B2(n_2886),
.Y(n_3771)
);

NAND2xp5_ASAP7_75t_L g3772 ( 
.A(n_2683),
.B(n_2686),
.Y(n_3772)
);

NOR2xp33_ASAP7_75t_L g3773 ( 
.A(n_3114),
.B(n_3135),
.Y(n_3773)
);

INVx2_ASAP7_75t_SL g3774 ( 
.A(n_3311),
.Y(n_3774)
);

NAND2xp5_ASAP7_75t_L g3775 ( 
.A(n_2686),
.B(n_2687),
.Y(n_3775)
);

NAND2xp5_ASAP7_75t_SL g3776 ( 
.A(n_3470),
.B(n_3409),
.Y(n_3776)
);

NAND2xp5_ASAP7_75t_L g3777 ( 
.A(n_2687),
.B(n_2688),
.Y(n_3777)
);

NOR2xp33_ASAP7_75t_L g3778 ( 
.A(n_3114),
.B(n_3135),
.Y(n_3778)
);

OA22x2_ASAP7_75t_L g3779 ( 
.A1(n_3348),
.A2(n_3271),
.B1(n_3214),
.B2(n_3279),
.Y(n_3779)
);

AO21x1_ASAP7_75t_L g3780 ( 
.A1(n_2738),
.A2(n_2868),
.B(n_2864),
.Y(n_3780)
);

HB1xp67_ASAP7_75t_L g3781 ( 
.A(n_2919),
.Y(n_3781)
);

OAI21xp5_ASAP7_75t_L g3782 ( 
.A1(n_3068),
.A2(n_2864),
.B(n_3174),
.Y(n_3782)
);

A2O1A1Ixp33_ASAP7_75t_L g3783 ( 
.A1(n_3100),
.A2(n_3279),
.B(n_2983),
.C(n_3103),
.Y(n_3783)
);

INVx2_ASAP7_75t_L g3784 ( 
.A(n_3386),
.Y(n_3784)
);

AOI22xp33_ASAP7_75t_L g3785 ( 
.A1(n_3032),
.A2(n_3025),
.B1(n_2983),
.B2(n_2928),
.Y(n_3785)
);

A2O1A1Ixp33_ASAP7_75t_L g3786 ( 
.A1(n_3100),
.A2(n_3279),
.B(n_2983),
.C(n_3103),
.Y(n_3786)
);

BUFx2_ASAP7_75t_L g3787 ( 
.A(n_2657),
.Y(n_3787)
);

NOR2xp33_ASAP7_75t_L g3788 ( 
.A(n_3114),
.B(n_3135),
.Y(n_3788)
);

NOR2xp33_ASAP7_75t_L g3789 ( 
.A(n_3135),
.B(n_3137),
.Y(n_3789)
);

INVx2_ASAP7_75t_L g3790 ( 
.A(n_3238),
.Y(n_3790)
);

NAND2xp5_ASAP7_75t_SL g3791 ( 
.A(n_3064),
.B(n_3099),
.Y(n_3791)
);

INVx3_ASAP7_75t_L g3792 ( 
.A(n_2712),
.Y(n_3792)
);

AOI21xp5_ASAP7_75t_L g3793 ( 
.A1(n_2682),
.A2(n_3158),
.B(n_3134),
.Y(n_3793)
);

NAND2xp5_ASAP7_75t_L g3794 ( 
.A(n_2687),
.B(n_2688),
.Y(n_3794)
);

AOI21xp5_ASAP7_75t_L g3795 ( 
.A1(n_3158),
.A2(n_3134),
.B(n_3434),
.Y(n_3795)
);

OAI21xp5_ASAP7_75t_L g3796 ( 
.A1(n_3174),
.A2(n_3043),
.B(n_3435),
.Y(n_3796)
);

AND2x2_ASAP7_75t_L g3797 ( 
.A(n_2835),
.B(n_3055),
.Y(n_3797)
);

BUFx2_ASAP7_75t_L g3798 ( 
.A(n_2673),
.Y(n_3798)
);

AND2x2_ASAP7_75t_L g3799 ( 
.A(n_3055),
.B(n_3088),
.Y(n_3799)
);

NAND2xp5_ASAP7_75t_SL g3800 ( 
.A(n_3064),
.B(n_3099),
.Y(n_3800)
);

CKINVDCx6p67_ASAP7_75t_R g3801 ( 
.A(n_2784),
.Y(n_3801)
);

NOR2xp33_ASAP7_75t_SL g3802 ( 
.A(n_3434),
.B(n_3128),
.Y(n_3802)
);

BUFx6f_ASAP7_75t_L g3803 ( 
.A(n_2769),
.Y(n_3803)
);

INVx1_ASAP7_75t_SL g3804 ( 
.A(n_3154),
.Y(n_3804)
);

AOI21xp5_ASAP7_75t_L g3805 ( 
.A1(n_3158),
.A2(n_3134),
.B(n_3434),
.Y(n_3805)
);

NAND2xp5_ASAP7_75t_L g3806 ( 
.A(n_2688),
.B(n_3284),
.Y(n_3806)
);

NOR3xp33_ASAP7_75t_L g3807 ( 
.A(n_3292),
.B(n_3185),
.C(n_3264),
.Y(n_3807)
);

AOI21xp5_ASAP7_75t_L g3808 ( 
.A1(n_3158),
.A2(n_3134),
.B(n_3434),
.Y(n_3808)
);

AOI22xp33_ASAP7_75t_L g3809 ( 
.A1(n_3032),
.A2(n_3025),
.B1(n_2983),
.B2(n_2976),
.Y(n_3809)
);

NOR2x1_ASAP7_75t_R g3810 ( 
.A(n_2654),
.B(n_2854),
.Y(n_3810)
);

NOR2xp33_ASAP7_75t_L g3811 ( 
.A(n_3137),
.B(n_3157),
.Y(n_3811)
);

NAND2xp5_ASAP7_75t_SL g3812 ( 
.A(n_3064),
.B(n_3099),
.Y(n_3812)
);

NAND2xp5_ASAP7_75t_SL g3813 ( 
.A(n_3208),
.B(n_3358),
.Y(n_3813)
);

NAND2xp5_ASAP7_75t_L g3814 ( 
.A(n_3284),
.B(n_3294),
.Y(n_3814)
);

NOR2xp33_ASAP7_75t_L g3815 ( 
.A(n_3137),
.B(n_3157),
.Y(n_3815)
);

AOI21xp5_ASAP7_75t_L g3816 ( 
.A1(n_3158),
.A2(n_3134),
.B(n_3434),
.Y(n_3816)
);

INVx2_ASAP7_75t_L g3817 ( 
.A(n_3234),
.Y(n_3817)
);

CKINVDCx5p33_ASAP7_75t_R g3818 ( 
.A(n_2721),
.Y(n_3818)
);

NAND2xp33_ASAP7_75t_L g3819 ( 
.A(n_3208),
.B(n_3074),
.Y(n_3819)
);

NOR2xp33_ASAP7_75t_SL g3820 ( 
.A(n_3434),
.B(n_3028),
.Y(n_3820)
);

BUFx6f_ASAP7_75t_L g3821 ( 
.A(n_2769),
.Y(n_3821)
);

OAI22xp5_ASAP7_75t_L g3822 ( 
.A1(n_2886),
.A2(n_2897),
.B1(n_2909),
.B2(n_3050),
.Y(n_3822)
);

NOR2xp33_ASAP7_75t_L g3823 ( 
.A(n_3137),
.B(n_3157),
.Y(n_3823)
);

AOI21xp5_ASAP7_75t_L g3824 ( 
.A1(n_3134),
.A2(n_3299),
.B(n_3193),
.Y(n_3824)
);

O2A1O1Ixp33_ASAP7_75t_L g3825 ( 
.A1(n_2892),
.A2(n_2994),
.B(n_3011),
.C(n_2910),
.Y(n_3825)
);

NAND2xp5_ASAP7_75t_SL g3826 ( 
.A(n_3358),
.B(n_3271),
.Y(n_3826)
);

AOI21xp5_ASAP7_75t_L g3827 ( 
.A1(n_3134),
.A2(n_3299),
.B(n_3193),
.Y(n_3827)
);

OAI21xp5_ASAP7_75t_L g3828 ( 
.A1(n_3174),
.A2(n_3043),
.B(n_3392),
.Y(n_3828)
);

NAND2xp5_ASAP7_75t_L g3829 ( 
.A(n_3284),
.B(n_3294),
.Y(n_3829)
);

OAI21x1_ASAP7_75t_L g3830 ( 
.A1(n_3389),
.A2(n_3155),
.B(n_2792),
.Y(n_3830)
);

OR2x6_ASAP7_75t_SL g3831 ( 
.A(n_2998),
.B(n_2722),
.Y(n_3831)
);

BUFx2_ASAP7_75t_L g3832 ( 
.A(n_2673),
.Y(n_3832)
);

OAI22xp5_ASAP7_75t_L g3833 ( 
.A1(n_2886),
.A2(n_2897),
.B1(n_2909),
.B2(n_3050),
.Y(n_3833)
);

O2A1O1Ixp33_ASAP7_75t_L g3834 ( 
.A1(n_2892),
.A2(n_2994),
.B(n_3011),
.C(n_2910),
.Y(n_3834)
);

NAND2xp5_ASAP7_75t_L g3835 ( 
.A(n_3294),
.B(n_3323),
.Y(n_3835)
);

AOI221xp5_ASAP7_75t_L g3836 ( 
.A1(n_2735),
.A2(n_3304),
.B1(n_3281),
.B2(n_3460),
.C(n_2997),
.Y(n_3836)
);

INVx2_ASAP7_75t_L g3837 ( 
.A(n_3254),
.Y(n_3837)
);

AOI21xp5_ASAP7_75t_L g3838 ( 
.A1(n_3193),
.A2(n_3299),
.B(n_3419),
.Y(n_3838)
);

NAND2xp5_ASAP7_75t_SL g3839 ( 
.A(n_3271),
.B(n_3156),
.Y(n_3839)
);

OAI22xp5_ASAP7_75t_L g3840 ( 
.A1(n_2886),
.A2(n_2897),
.B1(n_2909),
.B2(n_3059),
.Y(n_3840)
);

NAND2xp5_ASAP7_75t_SL g3841 ( 
.A(n_3156),
.B(n_3159),
.Y(n_3841)
);

NAND2xp5_ASAP7_75t_L g3842 ( 
.A(n_3323),
.B(n_3371),
.Y(n_3842)
);

O2A1O1Ixp33_ASAP7_75t_SL g3843 ( 
.A1(n_3282),
.A2(n_3159),
.B(n_3156),
.C(n_2735),
.Y(n_3843)
);

BUFx10_ASAP7_75t_L g3844 ( 
.A(n_3097),
.Y(n_3844)
);

NAND2xp5_ASAP7_75t_L g3845 ( 
.A(n_3323),
.B(n_3371),
.Y(n_3845)
);

OAI22xp5_ASAP7_75t_L g3846 ( 
.A1(n_2886),
.A2(n_2897),
.B1(n_2909),
.B2(n_3059),
.Y(n_3846)
);

AO32x2_ASAP7_75t_L g3847 ( 
.A1(n_2697),
.A2(n_2872),
.A3(n_2865),
.B1(n_3388),
.B2(n_3385),
.Y(n_3847)
);

NAND2xp5_ASAP7_75t_L g3848 ( 
.A(n_3371),
.B(n_3383),
.Y(n_3848)
);

NAND2xp5_ASAP7_75t_SL g3849 ( 
.A(n_3159),
.B(n_3223),
.Y(n_3849)
);

AOI22xp5_ASAP7_75t_L g3850 ( 
.A1(n_2713),
.A2(n_2923),
.B1(n_3062),
.B2(n_2997),
.Y(n_3850)
);

O2A1O1Ixp33_ASAP7_75t_L g3851 ( 
.A1(n_3029),
.A2(n_3115),
.B(n_3049),
.C(n_3185),
.Y(n_3851)
);

NAND2xp5_ASAP7_75t_SL g3852 ( 
.A(n_3223),
.B(n_3281),
.Y(n_3852)
);

NOR2xp33_ASAP7_75t_L g3853 ( 
.A(n_3157),
.B(n_3087),
.Y(n_3853)
);

O2A1O1Ixp33_ASAP7_75t_L g3854 ( 
.A1(n_3029),
.A2(n_3115),
.B(n_3049),
.C(n_3264),
.Y(n_3854)
);

BUFx6f_ASAP7_75t_L g3855 ( 
.A(n_2769),
.Y(n_3855)
);

AOI21xp5_ASAP7_75t_L g3856 ( 
.A1(n_3419),
.A2(n_3098),
.B(n_3095),
.Y(n_3856)
);

AND2x2_ASAP7_75t_L g3857 ( 
.A(n_3088),
.B(n_2891),
.Y(n_3857)
);

NAND2xp5_ASAP7_75t_SL g3858 ( 
.A(n_3223),
.B(n_3304),
.Y(n_3858)
);

NAND2xp5_ASAP7_75t_L g3859 ( 
.A(n_3383),
.B(n_3424),
.Y(n_3859)
);

NOR2x1_ASAP7_75t_SL g3860 ( 
.A(n_2769),
.B(n_2781),
.Y(n_3860)
);

AND2x2_ASAP7_75t_L g3861 ( 
.A(n_3088),
.B(n_2891),
.Y(n_3861)
);

INVx2_ASAP7_75t_L g3862 ( 
.A(n_3290),
.Y(n_3862)
);

NAND2xp5_ASAP7_75t_L g3863 ( 
.A(n_3383),
.B(n_3424),
.Y(n_3863)
);

BUFx2_ASAP7_75t_L g3864 ( 
.A(n_3141),
.Y(n_3864)
);

AOI21xp33_ASAP7_75t_L g3865 ( 
.A1(n_2735),
.A2(n_2730),
.B(n_2727),
.Y(n_3865)
);

OAI21xp5_ASAP7_75t_L g3866 ( 
.A1(n_3043),
.A2(n_3392),
.B(n_3282),
.Y(n_3866)
);

INVx2_ASAP7_75t_L g3867 ( 
.A(n_3234),
.Y(n_3867)
);

OAI21xp5_ASAP7_75t_L g3868 ( 
.A1(n_3460),
.A2(n_2727),
.B(n_2923),
.Y(n_3868)
);

INVx2_ASAP7_75t_L g3869 ( 
.A(n_3274),
.Y(n_3869)
);

NAND2xp5_ASAP7_75t_L g3870 ( 
.A(n_2924),
.B(n_2925),
.Y(n_3870)
);

NAND2xp5_ASAP7_75t_L g3871 ( 
.A(n_2924),
.B(n_2925),
.Y(n_3871)
);

AOI22xp33_ASAP7_75t_L g3872 ( 
.A1(n_3032),
.A2(n_2983),
.B1(n_2976),
.B2(n_2928),
.Y(n_3872)
);

OR2x6_ASAP7_75t_L g3873 ( 
.A(n_2793),
.B(n_2797),
.Y(n_3873)
);

AOI21xp5_ASAP7_75t_L g3874 ( 
.A1(n_3095),
.A2(n_3101),
.B(n_3098),
.Y(n_3874)
);

OAI21xp5_ASAP7_75t_L g3875 ( 
.A1(n_3460),
.A2(n_2727),
.B(n_3062),
.Y(n_3875)
);

INVx6_ASAP7_75t_L g3876 ( 
.A(n_2756),
.Y(n_3876)
);

INVx2_ASAP7_75t_L g3877 ( 
.A(n_3354),
.Y(n_3877)
);

O2A1O1Ixp33_ASAP7_75t_L g3878 ( 
.A1(n_2737),
.A2(n_2752),
.B(n_2762),
.C(n_2760),
.Y(n_3878)
);

NOR2xp33_ASAP7_75t_L g3879 ( 
.A(n_3087),
.B(n_2721),
.Y(n_3879)
);

INVx2_ASAP7_75t_L g3880 ( 
.A(n_3234),
.Y(n_3880)
);

BUFx6f_ASAP7_75t_L g3881 ( 
.A(n_2769),
.Y(n_3881)
);

NOR2xp33_ASAP7_75t_L g3882 ( 
.A(n_3081),
.B(n_3215),
.Y(n_3882)
);

BUFx8_ASAP7_75t_SL g3883 ( 
.A(n_2670),
.Y(n_3883)
);

AOI21x1_ASAP7_75t_L g3884 ( 
.A1(n_3457),
.A2(n_3292),
.B(n_3221),
.Y(n_3884)
);

NAND2xp5_ASAP7_75t_L g3885 ( 
.A(n_2925),
.B(n_2933),
.Y(n_3885)
);

O2A1O1Ixp33_ASAP7_75t_L g3886 ( 
.A1(n_2737),
.A2(n_2752),
.B(n_2762),
.C(n_2760),
.Y(n_3886)
);

AOI21xp5_ASAP7_75t_L g3887 ( 
.A1(n_3095),
.A2(n_3101),
.B(n_3098),
.Y(n_3887)
);

AOI21xp5_ASAP7_75t_L g3888 ( 
.A1(n_3095),
.A2(n_3101),
.B(n_3098),
.Y(n_3888)
);

O2A1O1Ixp33_ASAP7_75t_L g3889 ( 
.A1(n_2737),
.A2(n_2752),
.B(n_2762),
.C(n_2760),
.Y(n_3889)
);

INVxp67_ASAP7_75t_L g3890 ( 
.A(n_2811),
.Y(n_3890)
);

AOI21xp5_ASAP7_75t_L g3891 ( 
.A1(n_3095),
.A2(n_3101),
.B(n_3098),
.Y(n_3891)
);

OAI21x1_ASAP7_75t_L g3892 ( 
.A1(n_3389),
.A2(n_2792),
.B(n_2734),
.Y(n_3892)
);

AOI21xp5_ASAP7_75t_L g3893 ( 
.A1(n_3101),
.A2(n_3188),
.B(n_3275),
.Y(n_3893)
);

NAND2xp5_ASAP7_75t_L g3894 ( 
.A(n_2933),
.B(n_2952),
.Y(n_3894)
);

OAI22xp5_ASAP7_75t_L g3895 ( 
.A1(n_3081),
.A2(n_2778),
.B1(n_2796),
.B2(n_2770),
.Y(n_3895)
);

NAND2xp5_ASAP7_75t_L g3896 ( 
.A(n_2933),
.B(n_2952),
.Y(n_3896)
);

NAND2xp5_ASAP7_75t_L g3897 ( 
.A(n_2952),
.B(n_2993),
.Y(n_3897)
);

NAND2x1p5_ASAP7_75t_L g3898 ( 
.A(n_3311),
.B(n_3094),
.Y(n_3898)
);

INVx1_ASAP7_75t_L g3899 ( 
.A(n_2723),
.Y(n_3899)
);

OR2x6_ASAP7_75t_L g3900 ( 
.A(n_2793),
.B(n_2797),
.Y(n_3900)
);

NOR2xp33_ASAP7_75t_L g3901 ( 
.A(n_3215),
.B(n_3069),
.Y(n_3901)
);

NAND2xp5_ASAP7_75t_SL g3902 ( 
.A(n_3209),
.B(n_3074),
.Y(n_3902)
);

OAI22xp5_ASAP7_75t_L g3903 ( 
.A1(n_2770),
.A2(n_2796),
.B1(n_2806),
.B2(n_2778),
.Y(n_3903)
);

BUFx6f_ASAP7_75t_L g3904 ( 
.A(n_2781),
.Y(n_3904)
);

OAI21xp5_ASAP7_75t_L g3905 ( 
.A1(n_3150),
.A2(n_2968),
.B(n_2778),
.Y(n_3905)
);

NAND2xp5_ASAP7_75t_L g3906 ( 
.A(n_2993),
.B(n_3012),
.Y(n_3906)
);

INVx2_ASAP7_75t_L g3907 ( 
.A(n_3274),
.Y(n_3907)
);

INVx1_ASAP7_75t_L g3908 ( 
.A(n_2723),
.Y(n_3908)
);

BUFx6f_ASAP7_75t_L g3909 ( 
.A(n_2781),
.Y(n_3909)
);

NAND2xp5_ASAP7_75t_L g3910 ( 
.A(n_2993),
.B(n_3012),
.Y(n_3910)
);

BUFx3_ASAP7_75t_L g3911 ( 
.A(n_2756),
.Y(n_3911)
);

OAI22xp5_ASAP7_75t_L g3912 ( 
.A1(n_2770),
.A2(n_2806),
.B1(n_2810),
.B2(n_2796),
.Y(n_3912)
);

OR2x6_ASAP7_75t_SL g3913 ( 
.A(n_2998),
.B(n_2722),
.Y(n_3913)
);

OAI21x1_ASAP7_75t_L g3914 ( 
.A1(n_3389),
.A2(n_2792),
.B(n_2734),
.Y(n_3914)
);

NAND2xp5_ASAP7_75t_L g3915 ( 
.A(n_3012),
.B(n_3117),
.Y(n_3915)
);

AOI21xp5_ASAP7_75t_L g3916 ( 
.A1(n_3275),
.A2(n_3030),
.B(n_2814),
.Y(n_3916)
);

NAND2xp5_ASAP7_75t_SL g3917 ( 
.A(n_3125),
.B(n_3168),
.Y(n_3917)
);

INVx2_ASAP7_75t_L g3918 ( 
.A(n_3238),
.Y(n_3918)
);

AND2x4_ASAP7_75t_L g3919 ( 
.A(n_2714),
.B(n_2724),
.Y(n_3919)
);

CKINVDCx20_ASAP7_75t_R g3920 ( 
.A(n_2670),
.Y(n_3920)
);

INVx1_ASAP7_75t_L g3921 ( 
.A(n_2723),
.Y(n_3921)
);

AOI22xp5_ASAP7_75t_L g3922 ( 
.A1(n_3061),
.A2(n_3106),
.B1(n_3214),
.B2(n_3228),
.Y(n_3922)
);

INVx1_ASAP7_75t_L g3923 ( 
.A(n_2742),
.Y(n_3923)
);

NAND3xp33_ASAP7_75t_L g3924 ( 
.A(n_3236),
.B(n_3214),
.C(n_3288),
.Y(n_3924)
);

A2O1A1Ixp33_ASAP7_75t_SL g3925 ( 
.A1(n_3236),
.A2(n_2734),
.B(n_3425),
.C(n_3466),
.Y(n_3925)
);

AOI22xp5_ASAP7_75t_L g3926 ( 
.A1(n_3061),
.A2(n_3106),
.B1(n_3228),
.B2(n_2810),
.Y(n_3926)
);

NAND2xp5_ASAP7_75t_L g3927 ( 
.A(n_3012),
.B(n_3117),
.Y(n_3927)
);

AOI21xp5_ASAP7_75t_L g3928 ( 
.A1(n_3275),
.A2(n_3030),
.B(n_2814),
.Y(n_3928)
);

AOI21xp5_ASAP7_75t_L g3929 ( 
.A1(n_3275),
.A2(n_3030),
.B(n_2814),
.Y(n_3929)
);

NAND2xp5_ASAP7_75t_L g3930 ( 
.A(n_3117),
.B(n_2730),
.Y(n_3930)
);

AOI21x1_ASAP7_75t_L g3931 ( 
.A1(n_3292),
.A2(n_3221),
.B(n_2968),
.Y(n_3931)
);

O2A1O1Ixp33_ASAP7_75t_SL g3932 ( 
.A1(n_3228),
.A2(n_2810),
.B(n_2819),
.C(n_2806),
.Y(n_3932)
);

INVx3_ASAP7_75t_L g3933 ( 
.A(n_2712),
.Y(n_3933)
);

INVx2_ASAP7_75t_L g3934 ( 
.A(n_3240),
.Y(n_3934)
);

NAND3xp33_ASAP7_75t_L g3935 ( 
.A(n_3288),
.B(n_3310),
.C(n_3178),
.Y(n_3935)
);

A2O1A1Ixp33_ASAP7_75t_L g3936 ( 
.A1(n_2656),
.A2(n_2745),
.B(n_2768),
.C(n_2692),
.Y(n_3936)
);

INVx2_ASAP7_75t_L g3937 ( 
.A(n_3240),
.Y(n_3937)
);

INVxp67_ASAP7_75t_L g3938 ( 
.A(n_2919),
.Y(n_3938)
);

AND2x2_ASAP7_75t_SL g3939 ( 
.A(n_2934),
.B(n_3272),
.Y(n_3939)
);

AOI21xp5_ASAP7_75t_L g3940 ( 
.A1(n_3275),
.A2(n_3030),
.B(n_2814),
.Y(n_3940)
);

NAND2xp5_ASAP7_75t_L g3941 ( 
.A(n_2730),
.B(n_2819),
.Y(n_3941)
);

BUFx6f_ASAP7_75t_L g3942 ( 
.A(n_2781),
.Y(n_3942)
);

A2O1A1Ixp33_ASAP7_75t_L g3943 ( 
.A1(n_2656),
.A2(n_2745),
.B(n_2768),
.C(n_2692),
.Y(n_3943)
);

INVx4_ASAP7_75t_L g3944 ( 
.A(n_3441),
.Y(n_3944)
);

INVx2_ASAP7_75t_L g3945 ( 
.A(n_3259),
.Y(n_3945)
);

INVx1_ASAP7_75t_L g3946 ( 
.A(n_2742),
.Y(n_3946)
);

AOI21xp5_ASAP7_75t_L g3947 ( 
.A1(n_3275),
.A2(n_3030),
.B(n_2776),
.Y(n_3947)
);

NAND3xp33_ASAP7_75t_L g3948 ( 
.A(n_3310),
.B(n_3178),
.C(n_3173),
.Y(n_3948)
);

NAND2x2_ASAP7_75t_L g3949 ( 
.A(n_3061),
.B(n_3106),
.Y(n_3949)
);

AND2x4_ASAP7_75t_L g3950 ( 
.A(n_2714),
.B(n_2724),
.Y(n_3950)
);

NAND2xp5_ASAP7_75t_L g3951 ( 
.A(n_2730),
.B(n_2819),
.Y(n_3951)
);

AOI21xp5_ASAP7_75t_L g3952 ( 
.A1(n_3275),
.A2(n_3030),
.B(n_2776),
.Y(n_3952)
);

NAND2xp5_ASAP7_75t_SL g3953 ( 
.A(n_3125),
.B(n_3168),
.Y(n_3953)
);

AOI22xp5_ASAP7_75t_L g3954 ( 
.A1(n_2828),
.A2(n_2839),
.B1(n_2844),
.B2(n_2837),
.Y(n_3954)
);

NAND3xp33_ASAP7_75t_L g3955 ( 
.A(n_3173),
.B(n_3178),
.C(n_2837),
.Y(n_3955)
);

AOI21xp5_ASAP7_75t_L g3956 ( 
.A1(n_2776),
.A2(n_3272),
.B(n_3085),
.Y(n_3956)
);

INVxp67_ASAP7_75t_L g3957 ( 
.A(n_3189),
.Y(n_3957)
);

NAND3xp33_ASAP7_75t_SL g3958 ( 
.A(n_3205),
.B(n_3209),
.C(n_3028),
.Y(n_3958)
);

OAI21x1_ASAP7_75t_L g3959 ( 
.A1(n_3389),
.A2(n_2792),
.B(n_2734),
.Y(n_3959)
);

NOR2xp33_ASAP7_75t_L g3960 ( 
.A(n_3069),
.B(n_3039),
.Y(n_3960)
);

NOR2xp33_ASAP7_75t_L g3961 ( 
.A(n_3069),
.B(n_3039),
.Y(n_3961)
);

AO21x1_ASAP7_75t_L g3962 ( 
.A1(n_2722),
.A2(n_2744),
.B(n_2742),
.Y(n_3962)
);

INVx1_ASAP7_75t_L g3963 ( 
.A(n_2744),
.Y(n_3963)
);

INVx1_ASAP7_75t_L g3964 ( 
.A(n_2744),
.Y(n_3964)
);

INVx1_ASAP7_75t_SL g3965 ( 
.A(n_3154),
.Y(n_3965)
);

AOI21xp5_ASAP7_75t_L g3966 ( 
.A1(n_2776),
.A2(n_3272),
.B(n_3085),
.Y(n_3966)
);

AOI21x1_ASAP7_75t_L g3967 ( 
.A1(n_3221),
.A2(n_2968),
.B(n_3192),
.Y(n_3967)
);

INVx1_ASAP7_75t_L g3968 ( 
.A(n_2754),
.Y(n_3968)
);

NAND2xp5_ASAP7_75t_L g3969 ( 
.A(n_2730),
.B(n_2828),
.Y(n_3969)
);

INVx1_ASAP7_75t_L g3970 ( 
.A(n_2754),
.Y(n_3970)
);

NAND2xp5_ASAP7_75t_SL g3971 ( 
.A(n_3205),
.B(n_3028),
.Y(n_3971)
);

NOR2xp33_ASAP7_75t_L g3972 ( 
.A(n_3446),
.B(n_3453),
.Y(n_3972)
);

NOR2xp33_ASAP7_75t_SL g3973 ( 
.A(n_2809),
.B(n_3441),
.Y(n_3973)
);

NOR2xp33_ASAP7_75t_L g3974 ( 
.A(n_3446),
.B(n_3453),
.Y(n_3974)
);

NAND2xp5_ASAP7_75t_L g3975 ( 
.A(n_2828),
.B(n_2837),
.Y(n_3975)
);

NOR2xp33_ASAP7_75t_L g3976 ( 
.A(n_3173),
.B(n_3180),
.Y(n_3976)
);

AOI21xp5_ASAP7_75t_L g3977 ( 
.A1(n_3272),
.A2(n_3085),
.B(n_2797),
.Y(n_3977)
);

O2A1O1Ixp5_ASAP7_75t_L g3978 ( 
.A1(n_2793),
.A2(n_2797),
.B(n_2788),
.C(n_2672),
.Y(n_3978)
);

INVx1_ASAP7_75t_L g3979 ( 
.A(n_2754),
.Y(n_3979)
);

NAND2xp5_ASAP7_75t_L g3980 ( 
.A(n_2839),
.B(n_2844),
.Y(n_3980)
);

NOR2xp33_ASAP7_75t_SL g3981 ( 
.A(n_2809),
.B(n_3441),
.Y(n_3981)
);

AOI21xp5_ASAP7_75t_L g3982 ( 
.A1(n_3272),
.A2(n_3085),
.B(n_2797),
.Y(n_3982)
);

NAND2xp5_ASAP7_75t_SL g3983 ( 
.A(n_3245),
.B(n_3466),
.Y(n_3983)
);

NAND2xp5_ASAP7_75t_L g3984 ( 
.A(n_2839),
.B(n_2844),
.Y(n_3984)
);

OR2x6_ASAP7_75t_SL g3985 ( 
.A(n_2998),
.B(n_2709),
.Y(n_3985)
);

INVx1_ASAP7_75t_L g3986 ( 
.A(n_2755),
.Y(n_3986)
);

NAND3xp33_ASAP7_75t_SL g3987 ( 
.A(n_3226),
.B(n_3257),
.C(n_3235),
.Y(n_3987)
);

INVx2_ASAP7_75t_SL g3988 ( 
.A(n_2714),
.Y(n_3988)
);

INVx1_ASAP7_75t_L g3989 ( 
.A(n_2755),
.Y(n_3989)
);

OAI21xp5_ASAP7_75t_L g3990 ( 
.A1(n_3150),
.A2(n_2856),
.B(n_2851),
.Y(n_3990)
);

CKINVDCx6p67_ASAP7_75t_R g3991 ( 
.A(n_2784),
.Y(n_3991)
);

INVx1_ASAP7_75t_L g3992 ( 
.A(n_2755),
.Y(n_3992)
);

AOI21xp5_ASAP7_75t_L g3993 ( 
.A1(n_3085),
.A2(n_2797),
.B(n_2793),
.Y(n_3993)
);

NAND2xp5_ASAP7_75t_L g3994 ( 
.A(n_2851),
.B(n_2856),
.Y(n_3994)
);

NAND2xp5_ASAP7_75t_L g3995 ( 
.A(n_2851),
.B(n_2856),
.Y(n_3995)
);

NAND2xp5_ASAP7_75t_L g3996 ( 
.A(n_2866),
.B(n_2874),
.Y(n_3996)
);

NAND2xp5_ASAP7_75t_SL g3997 ( 
.A(n_3245),
.B(n_3466),
.Y(n_3997)
);

AND2x2_ASAP7_75t_L g3998 ( 
.A(n_2898),
.B(n_3104),
.Y(n_3998)
);

AND2x2_ASAP7_75t_L g3999 ( 
.A(n_2898),
.B(n_3104),
.Y(n_3999)
);

A2O1A1Ixp33_ASAP7_75t_L g4000 ( 
.A1(n_2656),
.A2(n_2745),
.B(n_2768),
.C(n_2692),
.Y(n_4000)
);

NAND2xp5_ASAP7_75t_SL g4001 ( 
.A(n_3245),
.B(n_3398),
.Y(n_4001)
);

NAND2xp5_ASAP7_75t_L g4002 ( 
.A(n_2866),
.B(n_2874),
.Y(n_4002)
);

INVx1_ASAP7_75t_SL g4003 ( 
.A(n_3154),
.Y(n_4003)
);

AOI21xp33_ASAP7_75t_L g4004 ( 
.A1(n_2955),
.A2(n_2990),
.B(n_2934),
.Y(n_4004)
);

AOI21x1_ASAP7_75t_L g4005 ( 
.A1(n_3192),
.A2(n_3231),
.B(n_2873),
.Y(n_4005)
);

OAI22xp5_ASAP7_75t_L g4006 ( 
.A1(n_2866),
.A2(n_2874),
.B1(n_2888),
.B2(n_2882),
.Y(n_4006)
);

CKINVDCx10_ASAP7_75t_R g4007 ( 
.A(n_3013),
.Y(n_4007)
);

OAI22xp5_ASAP7_75t_L g4008 ( 
.A1(n_2882),
.A2(n_2888),
.B1(n_2899),
.B2(n_2895),
.Y(n_4008)
);

NAND2xp5_ASAP7_75t_L g4009 ( 
.A(n_2882),
.B(n_2888),
.Y(n_4009)
);

A2O1A1Ixp33_ASAP7_75t_SL g4010 ( 
.A1(n_2734),
.A2(n_3425),
.B(n_2826),
.C(n_3402),
.Y(n_4010)
);

AND2x2_ASAP7_75t_L g4011 ( 
.A(n_3104),
.B(n_2853),
.Y(n_4011)
);

AOI21xp5_ASAP7_75t_L g4012 ( 
.A1(n_3085),
.A2(n_2797),
.B(n_2793),
.Y(n_4012)
);

AOI21xp5_ASAP7_75t_L g4013 ( 
.A1(n_2793),
.A2(n_2971),
.B(n_2660),
.Y(n_4013)
);

INVx1_ASAP7_75t_L g4014 ( 
.A(n_2774),
.Y(n_4014)
);

NAND3xp33_ASAP7_75t_L g4015 ( 
.A(n_2895),
.B(n_2906),
.C(n_2899),
.Y(n_4015)
);

NOR2xp33_ASAP7_75t_L g4016 ( 
.A(n_3180),
.B(n_3225),
.Y(n_4016)
);

AOI21x1_ASAP7_75t_L g4017 ( 
.A1(n_3192),
.A2(n_3231),
.B(n_2873),
.Y(n_4017)
);

AND2x6_ASAP7_75t_SL g4018 ( 
.A(n_2809),
.B(n_3366),
.Y(n_4018)
);

NOR2xp33_ASAP7_75t_L g4019 ( 
.A(n_3180),
.B(n_3225),
.Y(n_4019)
);

O2A1O1Ixp33_ASAP7_75t_L g4020 ( 
.A1(n_2895),
.A2(n_2906),
.B(n_2937),
.C(n_2899),
.Y(n_4020)
);

NAND2xp5_ASAP7_75t_L g4021 ( 
.A(n_2906),
.B(n_2937),
.Y(n_4021)
);

NAND2xp5_ASAP7_75t_L g4022 ( 
.A(n_2937),
.B(n_2946),
.Y(n_4022)
);

OAI22x1_ASAP7_75t_L g4023 ( 
.A1(n_2902),
.A2(n_2912),
.B1(n_2934),
.B2(n_2955),
.Y(n_4023)
);

AOI21xp5_ASAP7_75t_L g4024 ( 
.A1(n_2793),
.A2(n_2971),
.B(n_2660),
.Y(n_4024)
);

A2O1A1Ixp33_ASAP7_75t_L g4025 ( 
.A1(n_2656),
.A2(n_2745),
.B(n_2768),
.C(n_2692),
.Y(n_4025)
);

NAND2xp5_ASAP7_75t_L g4026 ( 
.A(n_2946),
.B(n_2950),
.Y(n_4026)
);

BUFx12f_ASAP7_75t_L g4027 ( 
.A(n_2918),
.Y(n_4027)
);

AOI21xp5_ASAP7_75t_L g4028 ( 
.A1(n_2971),
.A2(n_2659),
.B(n_2660),
.Y(n_4028)
);

OAI22xp5_ASAP7_75t_L g4029 ( 
.A1(n_2946),
.A2(n_2953),
.B1(n_2956),
.B2(n_2950),
.Y(n_4029)
);

NAND2xp5_ASAP7_75t_L g4030 ( 
.A(n_2950),
.B(n_2953),
.Y(n_4030)
);

NAND2x1p5_ASAP7_75t_L g4031 ( 
.A(n_3094),
.B(n_3121),
.Y(n_4031)
);

AOI21xp5_ASAP7_75t_L g4032 ( 
.A1(n_2971),
.A2(n_2659),
.B(n_2660),
.Y(n_4032)
);

OAI21xp33_ASAP7_75t_L g4033 ( 
.A1(n_2731),
.A2(n_2956),
.B(n_2953),
.Y(n_4033)
);

O2A1O1Ixp33_ASAP7_75t_L g4034 ( 
.A1(n_2956),
.A2(n_2972),
.B(n_2978),
.C(n_2962),
.Y(n_4034)
);

OAI21xp5_ASAP7_75t_L g4035 ( 
.A1(n_3150),
.A2(n_2972),
.B(n_2962),
.Y(n_4035)
);

INVx2_ASAP7_75t_L g4036 ( 
.A(n_3238),
.Y(n_4036)
);

INVx2_ASAP7_75t_L g4037 ( 
.A(n_3238),
.Y(n_4037)
);

OAI21xp5_ASAP7_75t_L g4038 ( 
.A1(n_2962),
.A2(n_2978),
.B(n_2972),
.Y(n_4038)
);

NAND2xp5_ASAP7_75t_SL g4039 ( 
.A(n_3245),
.B(n_3398),
.Y(n_4039)
);

AND2x2_ASAP7_75t_L g4040 ( 
.A(n_3104),
.B(n_2853),
.Y(n_4040)
);

NAND2xp5_ASAP7_75t_L g4041 ( 
.A(n_2978),
.B(n_2985),
.Y(n_4041)
);

O2A1O1Ixp5_ASAP7_75t_L g4042 ( 
.A1(n_2672),
.A2(n_2788),
.B(n_2777),
.C(n_2779),
.Y(n_4042)
);

NAND2xp5_ASAP7_75t_L g4043 ( 
.A(n_2985),
.B(n_2987),
.Y(n_4043)
);

NOR2xp33_ASAP7_75t_SL g4044 ( 
.A(n_3441),
.B(n_3417),
.Y(n_4044)
);

AND2x2_ASAP7_75t_L g4045 ( 
.A(n_2853),
.B(n_2816),
.Y(n_4045)
);

AOI21xp5_ASAP7_75t_L g4046 ( 
.A1(n_2971),
.A2(n_2659),
.B(n_2660),
.Y(n_4046)
);

AOI21xp5_ASAP7_75t_L g4047 ( 
.A1(n_2659),
.A2(n_2708),
.B(n_2660),
.Y(n_4047)
);

O2A1O1Ixp33_ASAP7_75t_SL g4048 ( 
.A1(n_2985),
.A2(n_2987),
.B(n_2991),
.C(n_2989),
.Y(n_4048)
);

AND2x4_ASAP7_75t_L g4049 ( 
.A(n_2714),
.B(n_2724),
.Y(n_4049)
);

AND2x4_ASAP7_75t_L g4050 ( 
.A(n_2724),
.B(n_2764),
.Y(n_4050)
);

O2A1O1Ixp5_ASAP7_75t_L g4051 ( 
.A1(n_2672),
.A2(n_2788),
.B(n_2777),
.C(n_2779),
.Y(n_4051)
);

AOI21xp5_ASAP7_75t_L g4052 ( 
.A1(n_2659),
.A2(n_2708),
.B(n_2660),
.Y(n_4052)
);

NOR2xp33_ASAP7_75t_SL g4053 ( 
.A(n_3441),
.B(n_3417),
.Y(n_4053)
);

NAND2xp5_ASAP7_75t_SL g4054 ( 
.A(n_3398),
.B(n_3226),
.Y(n_4054)
);

BUFx2_ASAP7_75t_L g4055 ( 
.A(n_3141),
.Y(n_4055)
);

NAND3xp33_ASAP7_75t_L g4056 ( 
.A(n_2987),
.B(n_2991),
.C(n_2989),
.Y(n_4056)
);

AOI21x1_ASAP7_75t_L g4057 ( 
.A1(n_3192),
.A2(n_3231),
.B(n_2873),
.Y(n_4057)
);

NOR2xp33_ASAP7_75t_L g4058 ( 
.A(n_3225),
.B(n_3170),
.Y(n_4058)
);

NAND2xp5_ASAP7_75t_SL g4059 ( 
.A(n_3398),
.B(n_3235),
.Y(n_4059)
);

OAI22xp5_ASAP7_75t_L g4060 ( 
.A1(n_2989),
.A2(n_2996),
.B1(n_3000),
.B2(n_2991),
.Y(n_4060)
);

NAND2xp5_ASAP7_75t_L g4061 ( 
.A(n_2996),
.B(n_3000),
.Y(n_4061)
);

AOI22xp5_ASAP7_75t_L g4062 ( 
.A1(n_2996),
.A2(n_3000),
.B1(n_3031),
.B2(n_3027),
.Y(n_4062)
);

OA22x2_ASAP7_75t_L g4063 ( 
.A1(n_3348),
.A2(n_3124),
.B1(n_3123),
.B2(n_2912),
.Y(n_4063)
);

O2A1O1Ixp33_ASAP7_75t_SL g4064 ( 
.A1(n_3027),
.A2(n_3031),
.B(n_3041),
.C(n_3035),
.Y(n_4064)
);

AOI22xp5_ASAP7_75t_L g4065 ( 
.A1(n_3027),
.A2(n_3031),
.B1(n_3041),
.B2(n_3035),
.Y(n_4065)
);

NOR2xp33_ASAP7_75t_L g4066 ( 
.A(n_3170),
.B(n_3015),
.Y(n_4066)
);

NAND2xp5_ASAP7_75t_L g4067 ( 
.A(n_3035),
.B(n_3041),
.Y(n_4067)
);

O2A1O1Ixp33_ASAP7_75t_L g4068 ( 
.A1(n_3053),
.A2(n_3077),
.B(n_3082),
.C(n_3071),
.Y(n_4068)
);

NAND2xp5_ASAP7_75t_L g4069 ( 
.A(n_3053),
.B(n_3071),
.Y(n_4069)
);

NAND2xp5_ASAP7_75t_L g4070 ( 
.A(n_3053),
.B(n_3071),
.Y(n_4070)
);

INVx1_ASAP7_75t_L g4071 ( 
.A(n_2774),
.Y(n_4071)
);

OR2x2_ASAP7_75t_L g4072 ( 
.A(n_2709),
.B(n_2801),
.Y(n_4072)
);

NOR2xp67_ASAP7_75t_L g4073 ( 
.A(n_2826),
.B(n_3417),
.Y(n_4073)
);

OAI22xp5_ASAP7_75t_L g4074 ( 
.A1(n_3077),
.A2(n_3093),
.B1(n_3109),
.B2(n_3082),
.Y(n_4074)
);

AOI21xp5_ASAP7_75t_L g4075 ( 
.A1(n_2659),
.A2(n_2748),
.B(n_2708),
.Y(n_4075)
);

NOR2xp33_ASAP7_75t_L g4076 ( 
.A(n_3170),
.B(n_3015),
.Y(n_4076)
);

OAI22xp5_ASAP7_75t_L g4077 ( 
.A1(n_3077),
.A2(n_3093),
.B1(n_3109),
.B2(n_3082),
.Y(n_4077)
);

BUFx4f_ASAP7_75t_SL g4078 ( 
.A(n_2784),
.Y(n_4078)
);

AOI21xp5_ASAP7_75t_L g4079 ( 
.A1(n_2708),
.A2(n_3033),
.B(n_2748),
.Y(n_4079)
);

AOI22x1_ASAP7_75t_L g4080 ( 
.A1(n_2747),
.A2(n_2990),
.B1(n_2955),
.B2(n_3038),
.Y(n_4080)
);

NOR2xp33_ASAP7_75t_L g4081 ( 
.A(n_3170),
.B(n_3123),
.Y(n_4081)
);

NAND2xp5_ASAP7_75t_L g4082 ( 
.A(n_3093),
.B(n_3109),
.Y(n_4082)
);

CKINVDCx5p33_ASAP7_75t_R g4083 ( 
.A(n_2784),
.Y(n_4083)
);

NAND2xp5_ASAP7_75t_SL g4084 ( 
.A(n_3398),
.B(n_3257),
.Y(n_4084)
);

A2O1A1Ixp33_ASAP7_75t_L g4085 ( 
.A1(n_2780),
.A2(n_2934),
.B(n_2976),
.C(n_2928),
.Y(n_4085)
);

NAND2xp5_ASAP7_75t_SL g4086 ( 
.A(n_3296),
.B(n_3110),
.Y(n_4086)
);

NAND2xp5_ASAP7_75t_L g4087 ( 
.A(n_3110),
.B(n_3119),
.Y(n_4087)
);

INVx1_ASAP7_75t_L g4088 ( 
.A(n_2785),
.Y(n_4088)
);

OAI22xp5_ASAP7_75t_L g4089 ( 
.A1(n_3110),
.A2(n_3126),
.B1(n_3133),
.B2(n_3119),
.Y(n_4089)
);

INVx2_ASAP7_75t_L g4090 ( 
.A(n_3234),
.Y(n_4090)
);

AOI21xp5_ASAP7_75t_L g4091 ( 
.A1(n_2708),
.A2(n_3033),
.B(n_2748),
.Y(n_4091)
);

HB1xp67_ASAP7_75t_L g4092 ( 
.A(n_3189),
.Y(n_4092)
);

O2A1O1Ixp33_ASAP7_75t_SL g4093 ( 
.A1(n_3119),
.A2(n_3126),
.B(n_3136),
.C(n_3133),
.Y(n_4093)
);

BUFx4f_ASAP7_75t_L g4094 ( 
.A(n_3216),
.Y(n_4094)
);

NAND2xp5_ASAP7_75t_L g4095 ( 
.A(n_3126),
.B(n_3133),
.Y(n_4095)
);

INVx11_ASAP7_75t_L g4096 ( 
.A(n_2980),
.Y(n_4096)
);

NOR2xp33_ASAP7_75t_L g4097 ( 
.A(n_3170),
.B(n_3123),
.Y(n_4097)
);

OAI21x1_ASAP7_75t_L g4098 ( 
.A1(n_2792),
.A2(n_2734),
.B(n_3267),
.Y(n_4098)
);

NOR2xp33_ASAP7_75t_SL g4099 ( 
.A(n_3441),
.B(n_3417),
.Y(n_4099)
);

AOI21xp5_ASAP7_75t_L g4100 ( 
.A1(n_2748),
.A2(n_3033),
.B(n_3359),
.Y(n_4100)
);

OAI22xp5_ASAP7_75t_L g4101 ( 
.A1(n_3136),
.A2(n_2780),
.B1(n_3038),
.B2(n_2990),
.Y(n_4101)
);

NAND2xp5_ASAP7_75t_L g4102 ( 
.A(n_3136),
.B(n_3381),
.Y(n_4102)
);

OAI22xp5_ASAP7_75t_SL g4103 ( 
.A1(n_2772),
.A2(n_2782),
.B1(n_3296),
.B2(n_3199),
.Y(n_4103)
);

AOI21xp5_ASAP7_75t_L g4104 ( 
.A1(n_3033),
.A2(n_3359),
.B(n_3194),
.Y(n_4104)
);

OAI21xp5_ASAP7_75t_L g4105 ( 
.A1(n_2826),
.A2(n_2880),
.B(n_3038),
.Y(n_4105)
);

NAND2xp5_ASAP7_75t_L g4106 ( 
.A(n_3381),
.B(n_2674),
.Y(n_4106)
);

NOR2xp33_ASAP7_75t_L g4107 ( 
.A(n_3123),
.B(n_3124),
.Y(n_4107)
);

BUFx3_ASAP7_75t_L g4108 ( 
.A(n_2756),
.Y(n_4108)
);

NOR2xp33_ASAP7_75t_L g4109 ( 
.A(n_3124),
.B(n_3182),
.Y(n_4109)
);

BUFx12f_ASAP7_75t_L g4110 ( 
.A(n_2918),
.Y(n_4110)
);

NOR3xp33_ASAP7_75t_L g4111 ( 
.A(n_3260),
.B(n_3124),
.C(n_3417),
.Y(n_4111)
);

OAI22xp5_ASAP7_75t_L g4112 ( 
.A1(n_2780),
.A2(n_3038),
.B1(n_2976),
.B2(n_2928),
.Y(n_4112)
);

AOI22x1_ASAP7_75t_L g4113 ( 
.A1(n_2747),
.A2(n_2841),
.B1(n_3216),
.B2(n_3260),
.Y(n_4113)
);

AOI21xp5_ASAP7_75t_L g4114 ( 
.A1(n_3033),
.A2(n_3194),
.B(n_3111),
.Y(n_4114)
);

AOI21xp5_ASAP7_75t_L g4115 ( 
.A1(n_3111),
.A2(n_3200),
.B(n_3194),
.Y(n_4115)
);

A2O1A1Ixp33_ASAP7_75t_L g4116 ( 
.A1(n_2780),
.A2(n_2928),
.B(n_2976),
.C(n_2731),
.Y(n_4116)
);

NAND2xp5_ASAP7_75t_L g4117 ( 
.A(n_3381),
.B(n_2674),
.Y(n_4117)
);

OAI21xp33_ASAP7_75t_SL g4118 ( 
.A1(n_3348),
.A2(n_2747),
.B(n_2865),
.Y(n_4118)
);

NAND2xp5_ASAP7_75t_SL g4119 ( 
.A(n_3260),
.B(n_3182),
.Y(n_4119)
);

NAND2xp5_ASAP7_75t_SL g4120 ( 
.A(n_3260),
.B(n_3182),
.Y(n_4120)
);

NAND2xp5_ASAP7_75t_SL g4121 ( 
.A(n_3182),
.B(n_3374),
.Y(n_4121)
);

NOR2x1p5_ASAP7_75t_L g4122 ( 
.A(n_3182),
.B(n_3276),
.Y(n_4122)
);

OAI22xp5_ASAP7_75t_L g4123 ( 
.A1(n_2780),
.A2(n_3037),
.B1(n_2783),
.B2(n_2781),
.Y(n_4123)
);

AOI21xp5_ASAP7_75t_L g4124 ( 
.A1(n_3111),
.A2(n_3200),
.B(n_3194),
.Y(n_4124)
);

BUFx6f_ASAP7_75t_L g4125 ( 
.A(n_2781),
.Y(n_4125)
);

AOI21xp5_ASAP7_75t_L g4126 ( 
.A1(n_3111),
.A2(n_3200),
.B(n_3194),
.Y(n_4126)
);

BUFx3_ASAP7_75t_L g4127 ( 
.A(n_2756),
.Y(n_4127)
);

NAND2xp5_ASAP7_75t_L g4128 ( 
.A(n_2694),
.B(n_2880),
.Y(n_4128)
);

NAND2xp5_ASAP7_75t_SL g4129 ( 
.A(n_3374),
.B(n_3462),
.Y(n_4129)
);

AOI21xp5_ASAP7_75t_L g4130 ( 
.A1(n_3111),
.A2(n_3207),
.B(n_3200),
.Y(n_4130)
);

BUFx12f_ASAP7_75t_L g4131 ( 
.A(n_2929),
.Y(n_4131)
);

OR2x2_ASAP7_75t_L g4132 ( 
.A(n_2801),
.B(n_2786),
.Y(n_4132)
);

NOR2xp33_ASAP7_75t_L g4133 ( 
.A(n_2784),
.B(n_3462),
.Y(n_4133)
);

NAND2xp5_ASAP7_75t_SL g4134 ( 
.A(n_3374),
.B(n_3462),
.Y(n_4134)
);

INVx3_ASAP7_75t_SL g4135 ( 
.A(n_2929),
.Y(n_4135)
);

INVx1_ASAP7_75t_L g4136 ( 
.A(n_2785),
.Y(n_4136)
);

INVx3_ASAP7_75t_L g4137 ( 
.A(n_2712),
.Y(n_4137)
);

BUFx12f_ASAP7_75t_L g4138 ( 
.A(n_2984),
.Y(n_4138)
);

NAND2xp5_ASAP7_75t_L g4139 ( 
.A(n_3127),
.B(n_3444),
.Y(n_4139)
);

INVx2_ASAP7_75t_L g4140 ( 
.A(n_3259),
.Y(n_4140)
);

NOR2xp33_ASAP7_75t_L g4141 ( 
.A(n_3462),
.B(n_2772),
.Y(n_4141)
);

O2A1O1Ixp33_ASAP7_75t_SL g4142 ( 
.A1(n_2865),
.A2(n_3315),
.B(n_3370),
.C(n_3278),
.Y(n_4142)
);

NAND2xp5_ASAP7_75t_L g4143 ( 
.A(n_3127),
.B(n_3444),
.Y(n_4143)
);

NAND2xp5_ASAP7_75t_L g4144 ( 
.A(n_3444),
.B(n_3449),
.Y(n_4144)
);

NAND2xp5_ASAP7_75t_SL g4145 ( 
.A(n_3374),
.B(n_3462),
.Y(n_4145)
);

OAI21xp33_ASAP7_75t_L g4146 ( 
.A1(n_2731),
.A2(n_3187),
.B(n_2998),
.Y(n_4146)
);

O2A1O1Ixp5_ASAP7_75t_SL g4147 ( 
.A1(n_2785),
.A2(n_2791),
.B(n_2803),
.C(n_2800),
.Y(n_4147)
);

INVx2_ASAP7_75t_L g4148 ( 
.A(n_3297),
.Y(n_4148)
);

AOI21x1_ASAP7_75t_L g4149 ( 
.A1(n_3192),
.A2(n_3231),
.B(n_2871),
.Y(n_4149)
);

NAND2xp5_ASAP7_75t_L g4150 ( 
.A(n_3449),
.B(n_3458),
.Y(n_4150)
);

AOI21xp5_ASAP7_75t_L g4151 ( 
.A1(n_3200),
.A2(n_3217),
.B(n_3207),
.Y(n_4151)
);

INVx8_ASAP7_75t_L g4152 ( 
.A(n_2980),
.Y(n_4152)
);

NAND2xp5_ASAP7_75t_L g4153 ( 
.A(n_3449),
.B(n_3458),
.Y(n_4153)
);

BUFx12f_ASAP7_75t_L g4154 ( 
.A(n_2984),
.Y(n_4154)
);

INVx3_ASAP7_75t_L g4155 ( 
.A(n_2712),
.Y(n_4155)
);

AOI21xp5_ASAP7_75t_L g4156 ( 
.A1(n_3207),
.A2(n_3217),
.B(n_3121),
.Y(n_4156)
);

INVx1_ASAP7_75t_SL g4157 ( 
.A(n_3277),
.Y(n_4157)
);

NAND2xp5_ASAP7_75t_L g4158 ( 
.A(n_3458),
.B(n_3464),
.Y(n_4158)
);

BUFx2_ASAP7_75t_L g4159 ( 
.A(n_3171),
.Y(n_4159)
);

A2O1A1Ixp33_ASAP7_75t_L g4160 ( 
.A1(n_2731),
.A2(n_2783),
.B(n_2781),
.C(n_3187),
.Y(n_4160)
);

NOR3xp33_ASAP7_75t_L g4161 ( 
.A(n_3417),
.B(n_3469),
.C(n_3187),
.Y(n_4161)
);

NAND2xp5_ASAP7_75t_L g4162 ( 
.A(n_3464),
.B(n_3465),
.Y(n_4162)
);

INVx1_ASAP7_75t_L g4163 ( 
.A(n_2791),
.Y(n_4163)
);

O2A1O1Ixp33_ASAP7_75t_L g4164 ( 
.A1(n_2857),
.A2(n_2861),
.B(n_3227),
.C(n_3212),
.Y(n_4164)
);

INVx2_ASAP7_75t_L g4165 ( 
.A(n_3302),
.Y(n_4165)
);

NAND2xp5_ASAP7_75t_SL g4166 ( 
.A(n_3374),
.B(n_3462),
.Y(n_4166)
);

NAND2xp5_ASAP7_75t_L g4167 ( 
.A(n_3464),
.B(n_3465),
.Y(n_4167)
);

BUFx2_ASAP7_75t_L g4168 ( 
.A(n_3171),
.Y(n_4168)
);

AND2x4_ASAP7_75t_SL g4169 ( 
.A(n_2783),
.B(n_3417),
.Y(n_4169)
);

AOI21xp5_ASAP7_75t_L g4170 ( 
.A1(n_3207),
.A2(n_3217),
.B(n_3121),
.Y(n_4170)
);

AOI21xp5_ASAP7_75t_L g4171 ( 
.A1(n_3207),
.A2(n_3217),
.B(n_3121),
.Y(n_4171)
);

A2O1A1Ixp33_ASAP7_75t_L g4172 ( 
.A1(n_2783),
.A2(n_3187),
.B(n_2902),
.C(n_2912),
.Y(n_4172)
);

NAND2xp5_ASAP7_75t_L g4173 ( 
.A(n_3465),
.B(n_3472),
.Y(n_4173)
);

AOI21x1_ASAP7_75t_L g4174 ( 
.A1(n_3192),
.A2(n_3231),
.B(n_2871),
.Y(n_4174)
);

NAND2xp5_ASAP7_75t_L g4175 ( 
.A(n_3472),
.B(n_2821),
.Y(n_4175)
);

NAND2xp5_ASAP7_75t_L g4176 ( 
.A(n_3472),
.B(n_2821),
.Y(n_4176)
);

NAND2xp5_ASAP7_75t_L g4177 ( 
.A(n_2821),
.B(n_2834),
.Y(n_4177)
);

AOI221xp5_ASAP7_75t_L g4178 ( 
.A1(n_2834),
.A2(n_2849),
.B1(n_2848),
.B2(n_2902),
.C(n_2791),
.Y(n_4178)
);

BUFx3_ASAP7_75t_L g4179 ( 
.A(n_2756),
.Y(n_4179)
);

NOR2xp33_ASAP7_75t_L g4180 ( 
.A(n_3462),
.B(n_2782),
.Y(n_4180)
);

NAND2xp5_ASAP7_75t_L g4181 ( 
.A(n_2834),
.B(n_2848),
.Y(n_4181)
);

INVx2_ASAP7_75t_L g4182 ( 
.A(n_3302),
.Y(n_4182)
);

AOI21xp5_ASAP7_75t_L g4183 ( 
.A1(n_3207),
.A2(n_3217),
.B(n_3121),
.Y(n_4183)
);

INVx1_ASAP7_75t_L g4184 ( 
.A(n_2800),
.Y(n_4184)
);

INVx1_ASAP7_75t_L g4185 ( 
.A(n_2800),
.Y(n_4185)
);

AOI21xp5_ASAP7_75t_L g4186 ( 
.A1(n_3094),
.A2(n_3122),
.B(n_3121),
.Y(n_4186)
);

AOI21xp5_ASAP7_75t_L g4187 ( 
.A1(n_3094),
.A2(n_3122),
.B(n_3121),
.Y(n_4187)
);

BUFx2_ASAP7_75t_L g4188 ( 
.A(n_3171),
.Y(n_4188)
);

NAND2xp5_ASAP7_75t_L g4189 ( 
.A(n_2848),
.B(n_2849),
.Y(n_4189)
);

INVx1_ASAP7_75t_L g4190 ( 
.A(n_2803),
.Y(n_4190)
);

NAND2xp5_ASAP7_75t_L g4191 ( 
.A(n_2849),
.B(n_3456),
.Y(n_4191)
);

NAND2xp5_ASAP7_75t_L g4192 ( 
.A(n_3456),
.B(n_3471),
.Y(n_4192)
);

INVx8_ASAP7_75t_L g4193 ( 
.A(n_2980),
.Y(n_4193)
);

OAI22xp5_ASAP7_75t_L g4194 ( 
.A1(n_2783),
.A2(n_2870),
.B1(n_3199),
.B2(n_3086),
.Y(n_4194)
);

NOR2xp33_ASAP7_75t_SL g4195 ( 
.A(n_3441),
.B(n_3469),
.Y(n_4195)
);

AOI21xp5_ASAP7_75t_L g4196 ( 
.A1(n_3094),
.A2(n_3122),
.B(n_3121),
.Y(n_4196)
);

NAND2xp5_ASAP7_75t_L g4197 ( 
.A(n_3451),
.B(n_3456),
.Y(n_4197)
);

A2O1A1Ixp33_ASAP7_75t_SL g4198 ( 
.A1(n_2734),
.A2(n_3425),
.B(n_3402),
.C(n_3415),
.Y(n_4198)
);

OR2x6_ASAP7_75t_SL g4199 ( 
.A(n_2786),
.B(n_2803),
.Y(n_4199)
);

AND2x2_ASAP7_75t_L g4200 ( 
.A(n_2816),
.B(n_2845),
.Y(n_4200)
);

AOI21xp5_ASAP7_75t_L g4201 ( 
.A1(n_3094),
.A2(n_3130),
.B(n_3122),
.Y(n_4201)
);

O2A1O1Ixp5_ASAP7_75t_L g4202 ( 
.A1(n_2672),
.A2(n_2788),
.B(n_2817),
.C(n_2764),
.Y(n_4202)
);

AOI21xp5_ASAP7_75t_L g4203 ( 
.A1(n_3094),
.A2(n_3130),
.B(n_3122),
.Y(n_4203)
);

NAND2xp5_ASAP7_75t_L g4204 ( 
.A(n_3451),
.B(n_3471),
.Y(n_4204)
);

OAI21x1_ASAP7_75t_L g4205 ( 
.A1(n_2792),
.A2(n_3267),
.B(n_2841),
.Y(n_4205)
);

INVx1_ASAP7_75t_L g4206 ( 
.A(n_2817),
.Y(n_4206)
);

INVx1_ASAP7_75t_L g4207 ( 
.A(n_2817),
.Y(n_4207)
);

NAND2xp5_ASAP7_75t_L g4208 ( 
.A(n_3451),
.B(n_3456),
.Y(n_4208)
);

NAND2xp5_ASAP7_75t_L g4209 ( 
.A(n_3451),
.B(n_3456),
.Y(n_4209)
);

NAND2xp5_ASAP7_75t_L g4210 ( 
.A(n_3451),
.B(n_3471),
.Y(n_4210)
);

NOR2xp33_ASAP7_75t_L g4211 ( 
.A(n_3276),
.B(n_2999),
.Y(n_4211)
);

AND2x2_ASAP7_75t_L g4212 ( 
.A(n_2816),
.B(n_2845),
.Y(n_4212)
);

NAND2xp5_ASAP7_75t_SL g4213 ( 
.A(n_3374),
.B(n_2965),
.Y(n_4213)
);

INVxp67_ASAP7_75t_L g4214 ( 
.A(n_3448),
.Y(n_4214)
);

NAND2xp5_ASAP7_75t_L g4215 ( 
.A(n_3471),
.B(n_2879),
.Y(n_4215)
);

NOR2xp67_ASAP7_75t_R g4216 ( 
.A(n_3276),
.B(n_2684),
.Y(n_4216)
);

NAND3xp33_ASAP7_75t_L g4217 ( 
.A(n_3090),
.B(n_2884),
.C(n_2879),
.Y(n_4217)
);

BUFx6f_ASAP7_75t_L g4218 ( 
.A(n_2712),
.Y(n_4218)
);

NAND2xp5_ASAP7_75t_SL g4219 ( 
.A(n_3374),
.B(n_2965),
.Y(n_4219)
);

INVx4_ASAP7_75t_L g4220 ( 
.A(n_3441),
.Y(n_4220)
);

NAND2xp5_ASAP7_75t_L g4221 ( 
.A(n_3471),
.B(n_2884),
.Y(n_4221)
);

NOR2xp33_ASAP7_75t_R g4222 ( 
.A(n_2999),
.B(n_2854),
.Y(n_4222)
);

NAND2xp5_ASAP7_75t_SL g4223 ( 
.A(n_3374),
.B(n_2965),
.Y(n_4223)
);

AOI21xp5_ASAP7_75t_L g4224 ( 
.A1(n_3094),
.A2(n_3130),
.B(n_3122),
.Y(n_4224)
);

INVx1_ASAP7_75t_L g4225 ( 
.A(n_2741),
.Y(n_4225)
);

BUFx6f_ASAP7_75t_L g4226 ( 
.A(n_2712),
.Y(n_4226)
);

O2A1O1Ixp33_ASAP7_75t_SL g4227 ( 
.A1(n_3278),
.A2(n_3370),
.B(n_3315),
.C(n_2831),
.Y(n_4227)
);

INVxp67_ASAP7_75t_L g4228 ( 
.A(n_3448),
.Y(n_4228)
);

AOI21xp5_ASAP7_75t_L g4229 ( 
.A1(n_3094),
.A2(n_3130),
.B(n_3122),
.Y(n_4229)
);

NOR2xp33_ASAP7_75t_L g4230 ( 
.A(n_3276),
.B(n_2813),
.Y(n_4230)
);

NAND3xp33_ASAP7_75t_SL g4231 ( 
.A(n_3113),
.B(n_3153),
.C(n_3145),
.Y(n_4231)
);

NAND2xp5_ASAP7_75t_SL g4232 ( 
.A(n_3374),
.B(n_2965),
.Y(n_4232)
);

BUFx6f_ASAP7_75t_L g4233 ( 
.A(n_2712),
.Y(n_4233)
);

INVx1_ASAP7_75t_L g4234 ( 
.A(n_2741),
.Y(n_4234)
);

OR2x6_ASAP7_75t_L g4235 ( 
.A(n_2724),
.B(n_2764),
.Y(n_4235)
);

BUFx3_ASAP7_75t_L g4236 ( 
.A(n_2756),
.Y(n_4236)
);

NAND2xp5_ASAP7_75t_SL g4237 ( 
.A(n_3374),
.B(n_2965),
.Y(n_4237)
);

HB1xp67_ASAP7_75t_L g4238 ( 
.A(n_3001),
.Y(n_4238)
);

INVx3_ASAP7_75t_L g4239 ( 
.A(n_2712),
.Y(n_4239)
);

BUFx8_ASAP7_75t_L g4240 ( 
.A(n_3013),
.Y(n_4240)
);

BUFx6f_ASAP7_75t_L g4241 ( 
.A(n_2718),
.Y(n_4241)
);

NAND2x1p5_ASAP7_75t_L g4242 ( 
.A(n_3122),
.B(n_3130),
.Y(n_4242)
);

NOR2xp33_ASAP7_75t_L g4243 ( 
.A(n_3276),
.B(n_2813),
.Y(n_4243)
);

O2A1O1Ixp33_ASAP7_75t_L g4244 ( 
.A1(n_2857),
.A2(n_2861),
.B(n_3227),
.C(n_3212),
.Y(n_4244)
);

NOR2xp33_ASAP7_75t_L g4245 ( 
.A(n_2813),
.B(n_2823),
.Y(n_4245)
);

OAI21xp5_ASAP7_75t_L g4246 ( 
.A1(n_3364),
.A2(n_3090),
.B(n_2685),
.Y(n_4246)
);

OAI22x1_ASAP7_75t_L g4247 ( 
.A1(n_2741),
.A2(n_2746),
.B1(n_2685),
.B2(n_2728),
.Y(n_4247)
);

BUFx6f_ASAP7_75t_L g4248 ( 
.A(n_2718),
.Y(n_4248)
);

A2O1A1Ixp33_ASAP7_75t_SL g4249 ( 
.A1(n_3425),
.A2(n_3402),
.B(n_3415),
.C(n_3399),
.Y(n_4249)
);

AOI21xp5_ASAP7_75t_L g4250 ( 
.A1(n_3130),
.A2(n_3243),
.B(n_3441),
.Y(n_4250)
);

NAND2x1p5_ASAP7_75t_L g4251 ( 
.A(n_3130),
.B(n_3243),
.Y(n_4251)
);

NAND2xp5_ASAP7_75t_SL g4252 ( 
.A(n_3374),
.B(n_2965),
.Y(n_4252)
);

AND2x2_ASAP7_75t_SL g4253 ( 
.A(n_2724),
.B(n_2764),
.Y(n_4253)
);

OAI21xp33_ASAP7_75t_L g4254 ( 
.A1(n_2685),
.A2(n_2728),
.B(n_3364),
.Y(n_4254)
);

AOI21xp5_ASAP7_75t_L g4255 ( 
.A1(n_3130),
.A2(n_3243),
.B(n_3441),
.Y(n_4255)
);

INVx3_ASAP7_75t_L g4256 ( 
.A(n_2718),
.Y(n_4256)
);

NOR2xp67_ASAP7_75t_L g4257 ( 
.A(n_3469),
.B(n_2698),
.Y(n_4257)
);

NAND2xp5_ASAP7_75t_L g4258 ( 
.A(n_3277),
.B(n_3295),
.Y(n_4258)
);

O2A1O1Ixp33_ASAP7_75t_L g4259 ( 
.A1(n_3250),
.A2(n_3258),
.B(n_3266),
.C(n_3265),
.Y(n_4259)
);

NAND2xp5_ASAP7_75t_L g4260 ( 
.A(n_3277),
.B(n_3295),
.Y(n_4260)
);

O2A1O1Ixp33_ASAP7_75t_L g4261 ( 
.A1(n_3250),
.A2(n_3258),
.B(n_3266),
.C(n_3265),
.Y(n_4261)
);

AOI21xp5_ASAP7_75t_L g4262 ( 
.A1(n_3130),
.A2(n_3243),
.B(n_3198),
.Y(n_4262)
);

AOI22xp5_ASAP7_75t_L g4263 ( 
.A1(n_3175),
.A2(n_2986),
.B1(n_2854),
.B2(n_3001),
.Y(n_4263)
);

AOI21x1_ASAP7_75t_L g4264 ( 
.A1(n_3192),
.A2(n_3231),
.B(n_3369),
.Y(n_4264)
);

NAND2xp5_ASAP7_75t_L g4265 ( 
.A(n_3277),
.B(n_3295),
.Y(n_4265)
);

A2O1A1Ixp33_ASAP7_75t_L g4266 ( 
.A1(n_2790),
.A2(n_2764),
.B(n_3199),
.C(n_3169),
.Y(n_4266)
);

AOI22x1_ASAP7_75t_L g4267 ( 
.A1(n_2841),
.A2(n_3216),
.B1(n_3145),
.B2(n_3153),
.Y(n_4267)
);

OA21x2_ASAP7_75t_L g4268 ( 
.A1(n_2741),
.A2(n_2746),
.B(n_3070),
.Y(n_4268)
);

INVx3_ASAP7_75t_L g4269 ( 
.A(n_2718),
.Y(n_4269)
);

NOR2xp33_ASAP7_75t_L g4270 ( 
.A(n_2813),
.B(n_2823),
.Y(n_4270)
);

OAI22xp5_ASAP7_75t_L g4271 ( 
.A1(n_3086),
.A2(n_2786),
.B1(n_3473),
.B2(n_2676),
.Y(n_4271)
);

INVx1_ASAP7_75t_L g4272 ( 
.A(n_2746),
.Y(n_4272)
);

NOR2xp33_ASAP7_75t_L g4273 ( 
.A(n_2813),
.B(n_2823),
.Y(n_4273)
);

OR2x6_ASAP7_75t_SL g4274 ( 
.A(n_2786),
.B(n_3364),
.Y(n_4274)
);

AND2x2_ASAP7_75t_L g4275 ( 
.A(n_3070),
.B(n_3073),
.Y(n_4275)
);

NAND2xp5_ASAP7_75t_SL g4276 ( 
.A(n_3374),
.B(n_2965),
.Y(n_4276)
);

OAI22xp5_ASAP7_75t_L g4277 ( 
.A1(n_3086),
.A2(n_3473),
.B1(n_2676),
.B2(n_2677),
.Y(n_4277)
);

O2A1O1Ixp33_ASAP7_75t_L g4278 ( 
.A1(n_3303),
.A2(n_3364),
.B(n_2728),
.C(n_3443),
.Y(n_4278)
);

BUFx2_ASAP7_75t_L g4279 ( 
.A(n_3070),
.Y(n_4279)
);

AOI21xp5_ASAP7_75t_L g4280 ( 
.A1(n_3243),
.A2(n_3198),
.B(n_3197),
.Y(n_4280)
);

INVx1_ASAP7_75t_L g4281 ( 
.A(n_2746),
.Y(n_4281)
);

AOI21xp5_ASAP7_75t_L g4282 ( 
.A1(n_3243),
.A2(n_3198),
.B(n_3197),
.Y(n_4282)
);

AOI21xp5_ASAP7_75t_L g4283 ( 
.A1(n_3243),
.A2(n_3198),
.B(n_3197),
.Y(n_4283)
);

AND2x4_ASAP7_75t_L g4284 ( 
.A(n_2764),
.B(n_2813),
.Y(n_4284)
);

NAND2xp5_ASAP7_75t_L g4285 ( 
.A(n_3295),
.B(n_3073),
.Y(n_4285)
);

AOI22x1_ASAP7_75t_L g4286 ( 
.A1(n_2841),
.A2(n_3216),
.B1(n_3145),
.B2(n_3153),
.Y(n_4286)
);

NAND2xp5_ASAP7_75t_L g4287 ( 
.A(n_3073),
.B(n_3459),
.Y(n_4287)
);

BUFx6f_ASAP7_75t_L g4288 ( 
.A(n_2718),
.Y(n_4288)
);

NAND2xp5_ASAP7_75t_L g4289 ( 
.A(n_3459),
.B(n_3461),
.Y(n_4289)
);

AO32x1_ASAP7_75t_L g4290 ( 
.A1(n_3385),
.A2(n_3396),
.A3(n_3388),
.B1(n_2940),
.B2(n_2954),
.Y(n_4290)
);

NAND2xp5_ASAP7_75t_SL g4291 ( 
.A(n_3374),
.B(n_2965),
.Y(n_4291)
);

AOI21xp5_ASAP7_75t_L g4292 ( 
.A1(n_3243),
.A2(n_3198),
.B(n_3197),
.Y(n_4292)
);

OAI221xp5_ASAP7_75t_L g4293 ( 
.A1(n_2841),
.A2(n_3469),
.B1(n_3303),
.B2(n_3145),
.C(n_3191),
.Y(n_4293)
);

NOR2xp33_ASAP7_75t_L g4294 ( 
.A(n_2813),
.B(n_2823),
.Y(n_4294)
);

NOR2xp33_ASAP7_75t_L g4295 ( 
.A(n_2823),
.B(n_2869),
.Y(n_4295)
);

NAND2xp5_ASAP7_75t_L g4296 ( 
.A(n_3461),
.B(n_3443),
.Y(n_4296)
);

AOI21xp5_ASAP7_75t_L g4297 ( 
.A1(n_3243),
.A2(n_3198),
.B(n_3197),
.Y(n_4297)
);

BUFx6f_ASAP7_75t_L g4298 ( 
.A(n_2718),
.Y(n_4298)
);

OAI22xp5_ASAP7_75t_L g4299 ( 
.A1(n_2662),
.A2(n_2677),
.B1(n_2676),
.B2(n_3163),
.Y(n_4299)
);

NOR3xp33_ASAP7_75t_L g4300 ( 
.A(n_3469),
.B(n_2915),
.C(n_2859),
.Y(n_4300)
);

AOI21x1_ASAP7_75t_L g4301 ( 
.A1(n_3192),
.A2(n_3231),
.B(n_3369),
.Y(n_4301)
);

NOR2xp33_ASAP7_75t_L g4302 ( 
.A(n_2823),
.B(n_2869),
.Y(n_4302)
);

INVxp67_ASAP7_75t_L g4303 ( 
.A(n_3397),
.Y(n_4303)
);

OA22x2_ASAP7_75t_L g4304 ( 
.A1(n_3047),
.A2(n_3065),
.B1(n_3078),
.B2(n_2981),
.Y(n_4304)
);

BUFx2_ASAP7_75t_L g4305 ( 
.A(n_3317),
.Y(n_4305)
);

INVx1_ASAP7_75t_SL g4306 ( 
.A(n_3423),
.Y(n_4306)
);

NAND2xp5_ASAP7_75t_L g4307 ( 
.A(n_3443),
.B(n_3445),
.Y(n_4307)
);

NAND2xp5_ASAP7_75t_SL g4308 ( 
.A(n_3374),
.B(n_2965),
.Y(n_4308)
);

INVx1_ASAP7_75t_L g4309 ( 
.A(n_3224),
.Y(n_4309)
);

O2A1O1Ixp33_ASAP7_75t_L g4310 ( 
.A1(n_3220),
.A2(n_3248),
.B(n_3261),
.C(n_3251),
.Y(n_4310)
);

NOR2xp33_ASAP7_75t_L g4311 ( 
.A(n_2823),
.B(n_2869),
.Y(n_4311)
);

AOI21xp5_ASAP7_75t_L g4312 ( 
.A1(n_3197),
.A2(n_3241),
.B(n_3198),
.Y(n_4312)
);

OAI21xp5_ASAP7_75t_L g4313 ( 
.A1(n_3445),
.A2(n_3450),
.B(n_3447),
.Y(n_4313)
);

BUFx12f_ASAP7_75t_L g4314 ( 
.A(n_2854),
.Y(n_4314)
);

NAND2xp5_ASAP7_75t_L g4315 ( 
.A(n_3445),
.B(n_3447),
.Y(n_4315)
);

BUFx6f_ASAP7_75t_L g4316 ( 
.A(n_2718),
.Y(n_4316)
);

NAND2xp5_ASAP7_75t_SL g4317 ( 
.A(n_3374),
.B(n_2965),
.Y(n_4317)
);

NOR2xp33_ASAP7_75t_L g4318 ( 
.A(n_2823),
.B(n_2869),
.Y(n_4318)
);

INVx4_ASAP7_75t_L g4319 ( 
.A(n_2684),
.Y(n_4319)
);

OAI21xp33_ASAP7_75t_L g4320 ( 
.A1(n_2841),
.A2(n_3463),
.B(n_3450),
.Y(n_4320)
);

NAND2xp5_ASAP7_75t_SL g4321 ( 
.A(n_3374),
.B(n_2965),
.Y(n_4321)
);

AOI22xp5_ASAP7_75t_L g4322 ( 
.A1(n_3175),
.A2(n_2986),
.B1(n_2854),
.B2(n_2901),
.Y(n_4322)
);

NOR2xp33_ASAP7_75t_L g4323 ( 
.A(n_2869),
.B(n_2901),
.Y(n_4323)
);

BUFx3_ASAP7_75t_L g4324 ( 
.A(n_2756),
.Y(n_4324)
);

NAND2xp5_ASAP7_75t_SL g4325 ( 
.A(n_2965),
.B(n_3469),
.Y(n_4325)
);

AOI221xp5_ASAP7_75t_L g4326 ( 
.A1(n_3467),
.A2(n_2676),
.B1(n_2662),
.B2(n_2677),
.C(n_2981),
.Y(n_4326)
);

NAND2xp5_ASAP7_75t_L g4327 ( 
.A(n_3397),
.B(n_3408),
.Y(n_4327)
);

NAND3xp33_ASAP7_75t_L g4328 ( 
.A(n_2964),
.B(n_3436),
.C(n_3309),
.Y(n_4328)
);

NAND2xp5_ASAP7_75t_SL g4329 ( 
.A(n_2965),
.B(n_3469),
.Y(n_4329)
);

AOI22xp5_ASAP7_75t_L g4330 ( 
.A1(n_2986),
.A2(n_2901),
.B1(n_2905),
.B2(n_2869),
.Y(n_4330)
);

AND2x2_ASAP7_75t_L g4331 ( 
.A(n_2965),
.B(n_2662),
.Y(n_4331)
);

NAND2xp5_ASAP7_75t_L g4332 ( 
.A(n_3408),
.B(n_3234),
.Y(n_4332)
);

AOI21xp5_ASAP7_75t_L g4333 ( 
.A1(n_3197),
.A2(n_3241),
.B(n_2914),
.Y(n_4333)
);

NAND2xp5_ASAP7_75t_L g4334 ( 
.A(n_3240),
.B(n_3254),
.Y(n_4334)
);

NAND3xp33_ASAP7_75t_SL g4335 ( 
.A(n_3113),
.B(n_3153),
.C(n_3145),
.Y(n_4335)
);

AOI21xp33_ASAP7_75t_L g4336 ( 
.A1(n_2964),
.A2(n_3436),
.B(n_3309),
.Y(n_4336)
);

AOI21xp5_ASAP7_75t_L g4337 ( 
.A1(n_3241),
.A2(n_2914),
.B(n_2904),
.Y(n_4337)
);

INVx1_ASAP7_75t_L g4338 ( 
.A(n_3224),
.Y(n_4338)
);

INVx3_ASAP7_75t_L g4339 ( 
.A(n_2718),
.Y(n_4339)
);

AOI221xp5_ASAP7_75t_L g4340 ( 
.A1(n_2662),
.A2(n_2677),
.B1(n_2676),
.B2(n_2981),
.C(n_3224),
.Y(n_4340)
);

INVx3_ASAP7_75t_SL g4341 ( 
.A(n_3216),
.Y(n_4341)
);

BUFx12f_ASAP7_75t_L g4342 ( 
.A(n_2986),
.Y(n_4342)
);

AOI21xp5_ASAP7_75t_L g4343 ( 
.A1(n_3241),
.A2(n_2914),
.B(n_2904),
.Y(n_4343)
);

NOR2xp33_ASAP7_75t_L g4344 ( 
.A(n_2869),
.B(n_2901),
.Y(n_4344)
);

NAND2xp5_ASAP7_75t_L g4345 ( 
.A(n_3240),
.B(n_3254),
.Y(n_4345)
);

O2A1O1Ixp5_ASAP7_75t_L g4346 ( 
.A1(n_2672),
.A2(n_2788),
.B(n_2792),
.C(n_2840),
.Y(n_4346)
);

OAI21xp33_ASAP7_75t_L g4347 ( 
.A1(n_2790),
.A2(n_3248),
.B(n_3220),
.Y(n_4347)
);

NAND2xp5_ASAP7_75t_L g4348 ( 
.A(n_3240),
.B(n_3254),
.Y(n_4348)
);

AND2x2_ASAP7_75t_L g4349 ( 
.A(n_2676),
.B(n_2677),
.Y(n_4349)
);

NOR2xp33_ASAP7_75t_L g4350 ( 
.A(n_2869),
.B(n_2901),
.Y(n_4350)
);

NAND2xp5_ASAP7_75t_L g4351 ( 
.A(n_3254),
.B(n_3268),
.Y(n_4351)
);

OA22x2_ASAP7_75t_L g4352 ( 
.A1(n_3047),
.A2(n_3065),
.B1(n_3078),
.B2(n_2981),
.Y(n_4352)
);

NAND2xp5_ASAP7_75t_L g4353 ( 
.A(n_3268),
.B(n_3274),
.Y(n_4353)
);

NAND2xp5_ASAP7_75t_SL g4354 ( 
.A(n_3120),
.B(n_3148),
.Y(n_4354)
);

AO21x1_ASAP7_75t_L g4355 ( 
.A1(n_3220),
.A2(n_3251),
.B(n_3248),
.Y(n_4355)
);

INVx3_ASAP7_75t_L g4356 ( 
.A(n_2718),
.Y(n_4356)
);

AOI22xp33_ASAP7_75t_L g4357 ( 
.A1(n_2869),
.A2(n_2905),
.B1(n_2917),
.B2(n_2901),
.Y(n_4357)
);

AOI21xp5_ASAP7_75t_L g4358 ( 
.A1(n_3241),
.A2(n_2914),
.B(n_2904),
.Y(n_4358)
);

BUFx2_ASAP7_75t_L g4359 ( 
.A(n_3317),
.Y(n_4359)
);

AND2x2_ASAP7_75t_L g4360 ( 
.A(n_2790),
.B(n_2901),
.Y(n_4360)
);

NOR2xp33_ASAP7_75t_L g4361 ( 
.A(n_2901),
.B(n_2905),
.Y(n_4361)
);

AND2x2_ASAP7_75t_L g4362 ( 
.A(n_2790),
.B(n_2901),
.Y(n_4362)
);

NAND2xp5_ASAP7_75t_L g4363 ( 
.A(n_3268),
.B(n_3274),
.Y(n_4363)
);

AOI21xp5_ASAP7_75t_L g4364 ( 
.A1(n_3241),
.A2(n_2940),
.B(n_2904),
.Y(n_4364)
);

AOI21xp5_ASAP7_75t_L g4365 ( 
.A1(n_3241),
.A2(n_2954),
.B(n_2940),
.Y(n_4365)
);

NOR2xp67_ASAP7_75t_L g4366 ( 
.A(n_2698),
.B(n_2729),
.Y(n_4366)
);

OAI21xp5_ASAP7_75t_L g4367 ( 
.A1(n_2940),
.A2(n_2957),
.B(n_2954),
.Y(n_4367)
);

NAND2xp5_ASAP7_75t_SL g4368 ( 
.A(n_3120),
.B(n_3148),
.Y(n_4368)
);

HB1xp67_ASAP7_75t_L g4369 ( 
.A(n_3423),
.Y(n_4369)
);

OAI21xp5_ASAP7_75t_L g4370 ( 
.A1(n_2954),
.A2(n_2969),
.B(n_2957),
.Y(n_4370)
);

INVx2_ASAP7_75t_SL g4371 ( 
.A(n_4218),
.Y(n_4371)
);

OAI21x1_ASAP7_75t_L g4372 ( 
.A1(n_4005),
.A2(n_4057),
.B(n_4017),
.Y(n_4372)
);

AOI21x1_ASAP7_75t_L g4373 ( 
.A1(n_3716),
.A2(n_3231),
.B(n_3192),
.Y(n_4373)
);

INVxp67_ASAP7_75t_L g4374 ( 
.A(n_3525),
.Y(n_4374)
);

O2A1O1Ixp5_ASAP7_75t_L g4375 ( 
.A1(n_3725),
.A2(n_2788),
.B(n_2672),
.C(n_3161),
.Y(n_4375)
);

A2O1A1Ixp33_ASAP7_75t_L g4376 ( 
.A1(n_4326),
.A2(n_4340),
.B(n_3687),
.C(n_3756),
.Y(n_4376)
);

NAND2xp5_ASAP7_75t_L g4377 ( 
.A(n_3558),
.B(n_2936),
.Y(n_4377)
);

OAI22xp5_ASAP7_75t_L g4378 ( 
.A1(n_3756),
.A2(n_2911),
.B1(n_2981),
.B2(n_3164),
.Y(n_4378)
);

AOI221xp5_ASAP7_75t_SL g4379 ( 
.A1(n_3566),
.A2(n_3454),
.B1(n_3317),
.B2(n_2917),
.C(n_2979),
.Y(n_4379)
);

OAI21xp5_ASAP7_75t_L g4380 ( 
.A1(n_3665),
.A2(n_2969),
.B(n_2957),
.Y(n_4380)
);

BUFx12f_ASAP7_75t_L g4381 ( 
.A(n_3491),
.Y(n_4381)
);

OAI21xp5_ASAP7_75t_L g4382 ( 
.A1(n_3665),
.A2(n_2969),
.B(n_2957),
.Y(n_4382)
);

NAND2xp5_ASAP7_75t_L g4383 ( 
.A(n_3558),
.B(n_2936),
.Y(n_4383)
);

INVx2_ASAP7_75t_L g4384 ( 
.A(n_3690),
.Y(n_4384)
);

AND2x2_ASAP7_75t_L g4385 ( 
.A(n_4349),
.B(n_2905),
.Y(n_4385)
);

A2O1A1Ixp33_ASAP7_75t_L g4386 ( 
.A1(n_4326),
.A2(n_3164),
.B(n_3169),
.C(n_3097),
.Y(n_4386)
);

OAI22xp33_ASAP7_75t_L g4387 ( 
.A1(n_3762),
.A2(n_2986),
.B1(n_2751),
.B2(n_2881),
.Y(n_4387)
);

BUFx6f_ASAP7_75t_L g4388 ( 
.A(n_4218),
.Y(n_4388)
);

AOI21xp5_ASAP7_75t_L g4389 ( 
.A1(n_3482),
.A2(n_3105),
.B(n_3102),
.Y(n_4389)
);

NAND2xp5_ASAP7_75t_L g4390 ( 
.A(n_3990),
.B(n_2936),
.Y(n_4390)
);

AOI21xp5_ASAP7_75t_L g4391 ( 
.A1(n_3482),
.A2(n_3105),
.B(n_3102),
.Y(n_4391)
);

HB1xp67_ASAP7_75t_L g4392 ( 
.A(n_4268),
.Y(n_4392)
);

AOI21xp33_ASAP7_75t_L g4393 ( 
.A1(n_3605),
.A2(n_3309),
.B(n_2964),
.Y(n_4393)
);

AOI21xp5_ASAP7_75t_L g4394 ( 
.A1(n_3624),
.A2(n_3105),
.B(n_3102),
.Y(n_4394)
);

AND2x2_ASAP7_75t_L g4395 ( 
.A(n_4349),
.B(n_2905),
.Y(n_4395)
);

A2O1A1Ixp33_ASAP7_75t_L g4396 ( 
.A1(n_4340),
.A2(n_3169),
.B(n_3097),
.C(n_3105),
.Y(n_4396)
);

NAND2xp5_ASAP7_75t_L g4397 ( 
.A(n_4035),
.B(n_3990),
.Y(n_4397)
);

NAND2xp5_ASAP7_75t_L g4398 ( 
.A(n_4035),
.B(n_3274),
.Y(n_4398)
);

OAI21x1_ASAP7_75t_L g4399 ( 
.A1(n_4005),
.A2(n_3267),
.B(n_3290),
.Y(n_4399)
);

OAI22xp5_ASAP7_75t_L g4400 ( 
.A1(n_3577),
.A2(n_3454),
.B1(n_3317),
.B2(n_3013),
.Y(n_4400)
);

OAI21xp5_ASAP7_75t_L g4401 ( 
.A1(n_3577),
.A2(n_2988),
.B(n_2969),
.Y(n_4401)
);

AO32x2_ASAP7_75t_L g4402 ( 
.A1(n_4271),
.A2(n_3396),
.A3(n_3388),
.B1(n_3385),
.B2(n_2729),
.Y(n_4402)
);

AOI21xp5_ASAP7_75t_L g4403 ( 
.A1(n_3624),
.A2(n_3105),
.B(n_3102),
.Y(n_4403)
);

NOR2xp67_ASAP7_75t_L g4404 ( 
.A(n_4337),
.B(n_2698),
.Y(n_4404)
);

OAI21x1_ASAP7_75t_L g4405 ( 
.A1(n_4017),
.A2(n_3267),
.B(n_3290),
.Y(n_4405)
);

OAI21x1_ASAP7_75t_SL g4406 ( 
.A1(n_4028),
.A2(n_2729),
.B(n_2698),
.Y(n_4406)
);

OAI22xp5_ASAP7_75t_L g4407 ( 
.A1(n_3737),
.A2(n_3454),
.B1(n_3013),
.B2(n_2751),
.Y(n_4407)
);

AOI22xp5_ASAP7_75t_L g4408 ( 
.A1(n_3605),
.A2(n_3353),
.B1(n_3013),
.B2(n_3018),
.Y(n_4408)
);

NAND2xp5_ASAP7_75t_L g4409 ( 
.A(n_3571),
.B(n_3290),
.Y(n_4409)
);

AND2x2_ASAP7_75t_L g4410 ( 
.A(n_3873),
.B(n_2905),
.Y(n_4410)
);

OAI21x1_ASAP7_75t_L g4411 ( 
.A1(n_4057),
.A2(n_3267),
.B(n_3290),
.Y(n_4411)
);

INVx1_ASAP7_75t_L g4412 ( 
.A(n_4309),
.Y(n_4412)
);

NAND2xp5_ASAP7_75t_L g4413 ( 
.A(n_3571),
.B(n_3297),
.Y(n_4413)
);

OAI21xp5_ASAP7_75t_L g4414 ( 
.A1(n_3585),
.A2(n_3002),
.B(n_2988),
.Y(n_4414)
);

AND2x2_ASAP7_75t_L g4415 ( 
.A(n_3873),
.B(n_2905),
.Y(n_4415)
);

A2O1A1Ixp33_ASAP7_75t_L g4416 ( 
.A1(n_3687),
.A2(n_3169),
.B(n_3097),
.C(n_3105),
.Y(n_4416)
);

INVx1_ASAP7_75t_L g4417 ( 
.A(n_4309),
.Y(n_4417)
);

AOI21xp5_ASAP7_75t_L g4418 ( 
.A1(n_3741),
.A2(n_3105),
.B(n_3102),
.Y(n_4418)
);

INVxp67_ASAP7_75t_SL g4419 ( 
.A(n_3698),
.Y(n_4419)
);

NAND2xp5_ASAP7_75t_L g4420 ( 
.A(n_3595),
.B(n_3297),
.Y(n_4420)
);

NAND2xp5_ASAP7_75t_SL g4421 ( 
.A(n_3740),
.B(n_2905),
.Y(n_4421)
);

AND2x4_ASAP7_75t_SL g4422 ( 
.A(n_3844),
.B(n_3366),
.Y(n_4422)
);

OAI21x1_ASAP7_75t_L g4423 ( 
.A1(n_4149),
.A2(n_3267),
.B(n_3297),
.Y(n_4423)
);

NAND2xp5_ASAP7_75t_SL g4424 ( 
.A(n_3740),
.B(n_2905),
.Y(n_4424)
);

CKINVDCx6p67_ASAP7_75t_R g4425 ( 
.A(n_4135),
.Y(n_4425)
);

NAND2xp5_ASAP7_75t_L g4426 ( 
.A(n_3595),
.B(n_3297),
.Y(n_4426)
);

AND2x4_ASAP7_75t_L g4427 ( 
.A(n_3873),
.B(n_2917),
.Y(n_4427)
);

INVx1_ASAP7_75t_L g4428 ( 
.A(n_4338),
.Y(n_4428)
);

NAND2xp5_ASAP7_75t_L g4429 ( 
.A(n_3814),
.B(n_3302),
.Y(n_4429)
);

OAI21x1_ASAP7_75t_L g4430 ( 
.A1(n_4149),
.A2(n_3306),
.B(n_3302),
.Y(n_4430)
);

AO31x2_ASAP7_75t_L g4431 ( 
.A1(n_3780),
.A2(n_3962),
.A3(n_4355),
.B(n_3570),
.Y(n_4431)
);

INVx1_ASAP7_75t_SL g4432 ( 
.A(n_3711),
.Y(n_4432)
);

OAI21xp33_ASAP7_75t_L g4433 ( 
.A1(n_3730),
.A2(n_3261),
.B(n_3251),
.Y(n_4433)
);

AOI21xp5_ASAP7_75t_L g4434 ( 
.A1(n_3741),
.A2(n_3102),
.B(n_3278),
.Y(n_4434)
);

NAND2xp5_ASAP7_75t_L g4435 ( 
.A(n_3814),
.B(n_3302),
.Y(n_4435)
);

AOI21xp33_ASAP7_75t_L g4436 ( 
.A1(n_3734),
.A2(n_3309),
.B(n_2964),
.Y(n_4436)
);

AO31x2_ASAP7_75t_L g4437 ( 
.A1(n_3780),
.A2(n_3312),
.A3(n_3313),
.B(n_3306),
.Y(n_4437)
);

INVx1_ASAP7_75t_L g4438 ( 
.A(n_4338),
.Y(n_4438)
);

NAND2xp5_ASAP7_75t_L g4439 ( 
.A(n_3829),
.B(n_3835),
.Y(n_4439)
);

OAI22xp5_ASAP7_75t_L g4440 ( 
.A1(n_3566),
.A2(n_3013),
.B1(n_2751),
.B2(n_2881),
.Y(n_4440)
);

INVx3_ASAP7_75t_L g4441 ( 
.A(n_4218),
.Y(n_4441)
);

OAI21x1_ASAP7_75t_L g4442 ( 
.A1(n_4174),
.A2(n_3312),
.B(n_3306),
.Y(n_4442)
);

AOI21xp5_ASAP7_75t_L g4443 ( 
.A1(n_3599),
.A2(n_3102),
.B(n_3278),
.Y(n_4443)
);

AOI21xp5_ASAP7_75t_L g4444 ( 
.A1(n_3599),
.A2(n_3370),
.B(n_3315),
.Y(n_4444)
);

AOI21xp5_ASAP7_75t_L g4445 ( 
.A1(n_3824),
.A2(n_3370),
.B(n_3315),
.Y(n_4445)
);

AOI211x1_ASAP7_75t_L g4446 ( 
.A1(n_3924),
.A2(n_3263),
.B(n_3289),
.C(n_3261),
.Y(n_4446)
);

NAND2xp33_ASAP7_75t_L g4447 ( 
.A(n_3807),
.B(n_2980),
.Y(n_4447)
);

OAI21x1_ASAP7_75t_L g4448 ( 
.A1(n_4174),
.A2(n_3312),
.B(n_3306),
.Y(n_4448)
);

AOI21xp5_ASAP7_75t_L g4449 ( 
.A1(n_3824),
.A2(n_3002),
.B(n_2988),
.Y(n_4449)
);

NAND2xp5_ASAP7_75t_L g4450 ( 
.A(n_3829),
.B(n_3306),
.Y(n_4450)
);

CKINVDCx5p33_ASAP7_75t_R g4451 ( 
.A(n_3501),
.Y(n_4451)
);

OAI21xp5_ASAP7_75t_L g4452 ( 
.A1(n_3585),
.A2(n_3002),
.B(n_2988),
.Y(n_4452)
);

AOI21xp5_ASAP7_75t_L g4453 ( 
.A1(n_3827),
.A2(n_3007),
.B(n_3002),
.Y(n_4453)
);

OAI21xp5_ASAP7_75t_L g4454 ( 
.A1(n_3725),
.A2(n_3040),
.B(n_3007),
.Y(n_4454)
);

OAI21x1_ASAP7_75t_L g4455 ( 
.A1(n_3830),
.A2(n_4187),
.B(n_4186),
.Y(n_4455)
);

AND2x2_ASAP7_75t_L g4456 ( 
.A(n_3873),
.B(n_2917),
.Y(n_4456)
);

INVx1_ASAP7_75t_L g4457 ( 
.A(n_3847),
.Y(n_4457)
);

NAND2x1_ASAP7_75t_L g4458 ( 
.A(n_3586),
.B(n_3108),
.Y(n_4458)
);

NAND2xp5_ASAP7_75t_L g4459 ( 
.A(n_3835),
.B(n_3313),
.Y(n_4459)
);

OA21x2_ASAP7_75t_L g4460 ( 
.A1(n_4042),
.A2(n_3244),
.B(n_3233),
.Y(n_4460)
);

NAND2xp5_ASAP7_75t_L g4461 ( 
.A(n_3842),
.B(n_3316),
.Y(n_4461)
);

INVx4_ASAP7_75t_L g4462 ( 
.A(n_4094),
.Y(n_4462)
);

AOI211x1_ASAP7_75t_L g4463 ( 
.A1(n_3924),
.A2(n_3289),
.B(n_3291),
.C(n_3263),
.Y(n_4463)
);

BUFx3_ASAP7_75t_L g4464 ( 
.A(n_4240),
.Y(n_4464)
);

INVx1_ASAP7_75t_SL g4465 ( 
.A(n_3711),
.Y(n_4465)
);

NAND2xp5_ASAP7_75t_L g4466 ( 
.A(n_3842),
.B(n_3316),
.Y(n_4466)
);

NAND2xp5_ASAP7_75t_L g4467 ( 
.A(n_3845),
.B(n_3316),
.Y(n_4467)
);

NAND2xp5_ASAP7_75t_SL g4468 ( 
.A(n_3762),
.B(n_2917),
.Y(n_4468)
);

NAND2xp33_ASAP7_75t_SL g4469 ( 
.A(n_4222),
.B(n_3353),
.Y(n_4469)
);

AOI21xp5_ASAP7_75t_L g4470 ( 
.A1(n_3827),
.A2(n_3040),
.B(n_3007),
.Y(n_4470)
);

NAND2x1p5_ASAP7_75t_L g4471 ( 
.A(n_4267),
.B(n_2794),
.Y(n_4471)
);

OAI21xp5_ASAP7_75t_L g4472 ( 
.A1(n_3770),
.A2(n_3040),
.B(n_3007),
.Y(n_4472)
);

CKINVDCx5p33_ASAP7_75t_R g4473 ( 
.A(n_3883),
.Y(n_4473)
);

AOI31xp67_ASAP7_75t_L g4474 ( 
.A1(n_4063),
.A2(n_2695),
.A3(n_2703),
.B(n_2702),
.Y(n_4474)
);

NAND2xp5_ASAP7_75t_L g4475 ( 
.A(n_3845),
.B(n_3322),
.Y(n_4475)
);

AOI21xp5_ASAP7_75t_L g4476 ( 
.A1(n_3736),
.A2(n_3052),
.B(n_3040),
.Y(n_4476)
);

INVx5_ASAP7_75t_L g4477 ( 
.A(n_3703),
.Y(n_4477)
);

OAI21xp5_ASAP7_75t_L g4478 ( 
.A1(n_3770),
.A2(n_3089),
.B(n_3052),
.Y(n_4478)
);

INVx1_ASAP7_75t_L g4479 ( 
.A(n_3847),
.Y(n_4479)
);

OR2x2_ASAP7_75t_L g4480 ( 
.A(n_4268),
.B(n_2917),
.Y(n_4480)
);

INVx5_ASAP7_75t_L g4481 ( 
.A(n_3703),
.Y(n_4481)
);

OAI21x1_ASAP7_75t_L g4482 ( 
.A1(n_4196),
.A2(n_4203),
.B(n_4201),
.Y(n_4482)
);

INVx3_ASAP7_75t_L g4483 ( 
.A(n_4218),
.Y(n_4483)
);

NAND2xp5_ASAP7_75t_L g4484 ( 
.A(n_3848),
.B(n_3339),
.Y(n_4484)
);

BUFx2_ASAP7_75t_L g4485 ( 
.A(n_3847),
.Y(n_4485)
);

OAI21x1_ASAP7_75t_L g4486 ( 
.A1(n_4203),
.A2(n_4229),
.B(n_4224),
.Y(n_4486)
);

AOI21x1_ASAP7_75t_L g4487 ( 
.A1(n_3716),
.A2(n_3231),
.B(n_3366),
.Y(n_4487)
);

OAI21x1_ASAP7_75t_L g4488 ( 
.A1(n_4224),
.A2(n_3349),
.B(n_3347),
.Y(n_4488)
);

A2O1A1Ixp33_ASAP7_75t_L g4489 ( 
.A1(n_3745),
.A2(n_3169),
.B(n_3097),
.C(n_3286),
.Y(n_4489)
);

NAND2x1_ASAP7_75t_L g4490 ( 
.A(n_3586),
.B(n_3108),
.Y(n_4490)
);

AOI21xp5_ASAP7_75t_L g4491 ( 
.A1(n_3736),
.A2(n_3089),
.B(n_3052),
.Y(n_4491)
);

NAND2xp5_ASAP7_75t_L g4492 ( 
.A(n_3848),
.B(n_3347),
.Y(n_4492)
);

OAI21xp33_ASAP7_75t_L g4493 ( 
.A1(n_3600),
.A2(n_3289),
.B(n_3263),
.Y(n_4493)
);

AOI21xp5_ASAP7_75t_L g4494 ( 
.A1(n_3748),
.A2(n_3089),
.B(n_3052),
.Y(n_4494)
);

AND2x4_ASAP7_75t_L g4495 ( 
.A(n_3873),
.B(n_2917),
.Y(n_4495)
);

BUFx6f_ASAP7_75t_L g4496 ( 
.A(n_4218),
.Y(n_4496)
);

INVx1_ASAP7_75t_L g4497 ( 
.A(n_3847),
.Y(n_4497)
);

OAI21x1_ASAP7_75t_L g4498 ( 
.A1(n_4229),
.A2(n_3349),
.B(n_3347),
.Y(n_4498)
);

AOI21xp5_ASAP7_75t_L g4499 ( 
.A1(n_3748),
.A2(n_3091),
.B(n_3089),
.Y(n_4499)
);

AOI21xp5_ASAP7_75t_L g4500 ( 
.A1(n_3752),
.A2(n_3132),
.B(n_3091),
.Y(n_4500)
);

AOI21x1_ASAP7_75t_L g4501 ( 
.A1(n_3724),
.A2(n_3366),
.B(n_3293),
.Y(n_4501)
);

AOI21xp5_ASAP7_75t_L g4502 ( 
.A1(n_3752),
.A2(n_3132),
.B(n_3091),
.Y(n_4502)
);

NAND2xp5_ASAP7_75t_L g4503 ( 
.A(n_3859),
.B(n_3347),
.Y(n_4503)
);

NAND2xp5_ASAP7_75t_L g4504 ( 
.A(n_3859),
.B(n_3349),
.Y(n_4504)
);

AOI21xp5_ASAP7_75t_L g4505 ( 
.A1(n_3755),
.A2(n_3132),
.B(n_3091),
.Y(n_4505)
);

AOI21xp5_ASAP7_75t_L g4506 ( 
.A1(n_3755),
.A2(n_3139),
.B(n_3132),
.Y(n_4506)
);

AOI22xp5_ASAP7_75t_L g4507 ( 
.A1(n_3623),
.A2(n_3353),
.B1(n_3018),
.B2(n_2842),
.Y(n_4507)
);

INVx1_ASAP7_75t_L g4508 ( 
.A(n_3847),
.Y(n_4508)
);

INVx3_ASAP7_75t_L g4509 ( 
.A(n_4218),
.Y(n_4509)
);

AOI22xp5_ASAP7_75t_L g4510 ( 
.A1(n_3627),
.A2(n_3353),
.B1(n_3018),
.B2(n_2842),
.Y(n_4510)
);

OAI21xp5_ASAP7_75t_L g4511 ( 
.A1(n_3745),
.A2(n_3142),
.B(n_3139),
.Y(n_4511)
);

INVx1_ASAP7_75t_L g4512 ( 
.A(n_3847),
.Y(n_4512)
);

NOR2xp33_ASAP7_75t_L g4513 ( 
.A(n_3850),
.B(n_2917),
.Y(n_4513)
);

INVx5_ASAP7_75t_L g4514 ( 
.A(n_3703),
.Y(n_4514)
);

CKINVDCx5p33_ASAP7_75t_R g4515 ( 
.A(n_3753),
.Y(n_4515)
);

INVx1_ASAP7_75t_L g4516 ( 
.A(n_3847),
.Y(n_4516)
);

CKINVDCx5p33_ASAP7_75t_R g4517 ( 
.A(n_3818),
.Y(n_4517)
);

AOI21xp5_ASAP7_75t_L g4518 ( 
.A1(n_4337),
.A2(n_3142),
.B(n_3139),
.Y(n_4518)
);

AOI21xp5_ASAP7_75t_L g4519 ( 
.A1(n_4343),
.A2(n_3142),
.B(n_3139),
.Y(n_4519)
);

BUFx2_ASAP7_75t_L g4520 ( 
.A(n_3749),
.Y(n_4520)
);

BUFx3_ASAP7_75t_L g4521 ( 
.A(n_4240),
.Y(n_4521)
);

OAI21xp5_ASAP7_75t_L g4522 ( 
.A1(n_3746),
.A2(n_3181),
.B(n_3142),
.Y(n_4522)
);

NAND2x1p5_ASAP7_75t_L g4523 ( 
.A(n_4267),
.B(n_2794),
.Y(n_4523)
);

BUFx12f_ASAP7_75t_L g4524 ( 
.A(n_3615),
.Y(n_4524)
);

AOI21xp5_ASAP7_75t_L g4525 ( 
.A1(n_4358),
.A2(n_3201),
.B(n_3181),
.Y(n_4525)
);

AOI21xp5_ASAP7_75t_L g4526 ( 
.A1(n_4358),
.A2(n_3201),
.B(n_3181),
.Y(n_4526)
);

OR2x6_ASAP7_75t_L g4527 ( 
.A(n_3479),
.B(n_2672),
.Y(n_4527)
);

AOI22xp33_ASAP7_75t_L g4528 ( 
.A1(n_3757),
.A2(n_2951),
.B1(n_2979),
.B2(n_2917),
.Y(n_4528)
);

NAND2xp5_ASAP7_75t_L g4529 ( 
.A(n_3863),
.B(n_3349),
.Y(n_4529)
);

NOR2xp67_ASAP7_75t_L g4530 ( 
.A(n_4343),
.B(n_4364),
.Y(n_4530)
);

INVx3_ASAP7_75t_L g4531 ( 
.A(n_4218),
.Y(n_4531)
);

INVx2_ASAP7_75t_L g4532 ( 
.A(n_3690),
.Y(n_4532)
);

BUFx2_ASAP7_75t_L g4533 ( 
.A(n_3749),
.Y(n_4533)
);

BUFx12f_ASAP7_75t_L g4534 ( 
.A(n_4027),
.Y(n_4534)
);

OAI21xp5_ASAP7_75t_L g4535 ( 
.A1(n_3764),
.A2(n_3201),
.B(n_3181),
.Y(n_4535)
);

NOR2xp33_ASAP7_75t_L g4536 ( 
.A(n_3850),
.B(n_3757),
.Y(n_4536)
);

AOI21xp5_ASAP7_75t_L g4537 ( 
.A1(n_4364),
.A2(n_3201),
.B(n_3161),
.Y(n_4537)
);

INVx1_ASAP7_75t_L g4538 ( 
.A(n_3690),
.Y(n_4538)
);

INVx1_ASAP7_75t_L g4539 ( 
.A(n_3784),
.Y(n_4539)
);

OR2x2_ASAP7_75t_L g4540 ( 
.A(n_4268),
.B(n_2917),
.Y(n_4540)
);

AOI21xp33_ASAP7_75t_L g4541 ( 
.A1(n_3779),
.A2(n_3309),
.B(n_2964),
.Y(n_4541)
);

AND2x2_ASAP7_75t_L g4542 ( 
.A(n_3873),
.B(n_2951),
.Y(n_4542)
);

NAND2xp5_ASAP7_75t_L g4543 ( 
.A(n_4106),
.B(n_4117),
.Y(n_4543)
);

INVx1_ASAP7_75t_L g4544 ( 
.A(n_3784),
.Y(n_4544)
);

NOR2xp33_ASAP7_75t_SL g4545 ( 
.A(n_3610),
.B(n_2964),
.Y(n_4545)
);

O2A1O1Ixp5_ASAP7_75t_L g4546 ( 
.A1(n_3776),
.A2(n_2788),
.B(n_3161),
.C(n_2855),
.Y(n_4546)
);

AOI21xp5_ASAP7_75t_L g4547 ( 
.A1(n_4365),
.A2(n_3161),
.B(n_3148),
.Y(n_4547)
);

AOI22xp33_ASAP7_75t_L g4548 ( 
.A1(n_3729),
.A2(n_3852),
.B1(n_3858),
.B2(n_3826),
.Y(n_4548)
);

AOI21x1_ASAP7_75t_L g4549 ( 
.A1(n_3724),
.A2(n_3366),
.B(n_3293),
.Y(n_4549)
);

INVx1_ASAP7_75t_L g4550 ( 
.A(n_3784),
.Y(n_4550)
);

INVx2_ASAP7_75t_L g4551 ( 
.A(n_3790),
.Y(n_4551)
);

NAND2xp5_ASAP7_75t_SL g4552 ( 
.A(n_3836),
.B(n_2951),
.Y(n_4552)
);

INVx1_ASAP7_75t_L g4553 ( 
.A(n_3790),
.Y(n_4553)
);

AOI22xp5_ASAP7_75t_L g4554 ( 
.A1(n_3729),
.A2(n_3813),
.B1(n_3836),
.B2(n_3771),
.Y(n_4554)
);

AND2x6_ASAP7_75t_SL g4555 ( 
.A(n_4211),
.B(n_3366),
.Y(n_4555)
);

HB1xp67_ASAP7_75t_L g4556 ( 
.A(n_4268),
.Y(n_4556)
);

OA21x2_ASAP7_75t_L g4557 ( 
.A1(n_4042),
.A2(n_3252),
.B(n_3247),
.Y(n_4557)
);

OR2x2_ASAP7_75t_L g4558 ( 
.A(n_4268),
.B(n_2951),
.Y(n_4558)
);

AOI21xp5_ASAP7_75t_L g4559 ( 
.A1(n_4365),
.A2(n_3161),
.B(n_3148),
.Y(n_4559)
);

INVx3_ASAP7_75t_L g4560 ( 
.A(n_4226),
.Y(n_4560)
);

NAND3xp33_ASAP7_75t_L g4561 ( 
.A(n_3807),
.B(n_2979),
.C(n_2951),
.Y(n_4561)
);

NAND2x1_ASAP7_75t_L g4562 ( 
.A(n_3586),
.B(n_3108),
.Y(n_4562)
);

HB1xp67_ASAP7_75t_L g4563 ( 
.A(n_3525),
.Y(n_4563)
);

OAI21xp5_ASAP7_75t_L g4564 ( 
.A1(n_3767),
.A2(n_3145),
.B(n_3113),
.Y(n_4564)
);

AOI21xp5_ASAP7_75t_L g4565 ( 
.A1(n_3560),
.A2(n_3733),
.B(n_4044),
.Y(n_4565)
);

NAND2xp5_ASAP7_75t_SL g4566 ( 
.A(n_3759),
.B(n_2951),
.Y(n_4566)
);

OR2x2_ASAP7_75t_L g4567 ( 
.A(n_3930),
.B(n_2951),
.Y(n_4567)
);

AOI21xp33_ASAP7_75t_L g4568 ( 
.A1(n_3779),
.A2(n_3309),
.B(n_2964),
.Y(n_4568)
);

OAI21xp5_ASAP7_75t_L g4569 ( 
.A1(n_3767),
.A2(n_3153),
.B(n_3113),
.Y(n_4569)
);

NAND2x1_ASAP7_75t_L g4570 ( 
.A(n_3586),
.B(n_3108),
.Y(n_4570)
);

NOR2xp33_ASAP7_75t_L g4571 ( 
.A(n_3935),
.B(n_2951),
.Y(n_4571)
);

OAI21x1_ASAP7_75t_L g4572 ( 
.A1(n_4262),
.A2(n_3378),
.B(n_3372),
.Y(n_4572)
);

AOI21xp5_ASAP7_75t_L g4573 ( 
.A1(n_3560),
.A2(n_3161),
.B(n_3148),
.Y(n_4573)
);

OAI21x1_ASAP7_75t_L g4574 ( 
.A1(n_4262),
.A2(n_3378),
.B(n_3372),
.Y(n_4574)
);

A2O1A1Ixp33_ASAP7_75t_L g4575 ( 
.A1(n_3560),
.A2(n_3287),
.B(n_3286),
.C(n_3211),
.Y(n_4575)
);

NAND3x1_ASAP7_75t_L g4576 ( 
.A(n_4111),
.B(n_3402),
.C(n_3399),
.Y(n_4576)
);

NAND2xp5_ASAP7_75t_SL g4577 ( 
.A(n_3759),
.B(n_2951),
.Y(n_4577)
);

CKINVDCx20_ASAP7_75t_R g4578 ( 
.A(n_3529),
.Y(n_4578)
);

OA22x2_ASAP7_75t_L g4579 ( 
.A1(n_4263),
.A2(n_3366),
.B1(n_3065),
.B2(n_3078),
.Y(n_4579)
);

AO31x2_ASAP7_75t_L g4580 ( 
.A1(n_3570),
.A2(n_3386),
.A3(n_3387),
.B(n_3378),
.Y(n_4580)
);

OR2x2_ASAP7_75t_L g4581 ( 
.A(n_3930),
.B(n_2951),
.Y(n_4581)
);

INVxp67_ASAP7_75t_SL g4582 ( 
.A(n_3698),
.Y(n_4582)
);

OAI21x1_ASAP7_75t_L g4583 ( 
.A1(n_3892),
.A2(n_3387),
.B(n_3386),
.Y(n_4583)
);

NOR2xp67_ASAP7_75t_L g4584 ( 
.A(n_4333),
.B(n_2729),
.Y(n_4584)
);

OAI21x1_ASAP7_75t_L g4585 ( 
.A1(n_3892),
.A2(n_3959),
.B(n_3914),
.Y(n_4585)
);

OAI21x1_ASAP7_75t_L g4586 ( 
.A1(n_3914),
.A2(n_3387),
.B(n_3386),
.Y(n_4586)
);

AND2x2_ASAP7_75t_L g4587 ( 
.A(n_3900),
.B(n_2979),
.Y(n_4587)
);

OAI21x1_ASAP7_75t_L g4588 ( 
.A1(n_3914),
.A2(n_3403),
.B(n_3391),
.Y(n_4588)
);

AND2x2_ASAP7_75t_L g4589 ( 
.A(n_3900),
.B(n_2979),
.Y(n_4589)
);

BUFx3_ASAP7_75t_L g4590 ( 
.A(n_4240),
.Y(n_4590)
);

AOI22xp33_ASAP7_75t_L g4591 ( 
.A1(n_3779),
.A2(n_2979),
.B1(n_3353),
.B2(n_3309),
.Y(n_4591)
);

AOI21xp5_ASAP7_75t_L g4592 ( 
.A1(n_3560),
.A2(n_3148),
.B(n_3120),
.Y(n_4592)
);

OAI21x1_ASAP7_75t_SL g4593 ( 
.A1(n_4028),
.A2(n_2759),
.B(n_2740),
.Y(n_4593)
);

OAI21x1_ASAP7_75t_L g4594 ( 
.A1(n_3959),
.A2(n_3403),
.B(n_3391),
.Y(n_4594)
);

OAI21x1_ASAP7_75t_L g4595 ( 
.A1(n_3959),
.A2(n_3403),
.B(n_3391),
.Y(n_4595)
);

INVx2_ASAP7_75t_L g4596 ( 
.A(n_3790),
.Y(n_4596)
);

OAI21x1_ASAP7_75t_L g4597 ( 
.A1(n_4280),
.A2(n_3420),
.B(n_3403),
.Y(n_4597)
);

OA21x2_ASAP7_75t_L g4598 ( 
.A1(n_4051),
.A2(n_3252),
.B(n_3247),
.Y(n_4598)
);

OAI21x1_ASAP7_75t_L g4599 ( 
.A1(n_4280),
.A2(n_3420),
.B(n_3403),
.Y(n_4599)
);

AND2x2_ASAP7_75t_L g4600 ( 
.A(n_3900),
.B(n_2979),
.Y(n_4600)
);

A2O1A1Ixp33_ASAP7_75t_L g4601 ( 
.A1(n_3733),
.A2(n_3287),
.B(n_3286),
.C(n_3211),
.Y(n_4601)
);

INVx2_ASAP7_75t_L g4602 ( 
.A(n_3817),
.Y(n_4602)
);

OAI21x1_ASAP7_75t_L g4603 ( 
.A1(n_4282),
.A2(n_4292),
.B(n_4283),
.Y(n_4603)
);

INVx4_ASAP7_75t_L g4604 ( 
.A(n_4094),
.Y(n_4604)
);

AOI21xp5_ASAP7_75t_L g4605 ( 
.A1(n_3733),
.A2(n_3148),
.B(n_3120),
.Y(n_4605)
);

OAI21xp5_ASAP7_75t_L g4606 ( 
.A1(n_3866),
.A2(n_3782),
.B(n_3743),
.Y(n_4606)
);

OAI21xp5_ASAP7_75t_L g4607 ( 
.A1(n_3866),
.A2(n_3153),
.B(n_3113),
.Y(n_4607)
);

AOI22xp5_ASAP7_75t_L g4608 ( 
.A1(n_3771),
.A2(n_3353),
.B1(n_3018),
.B2(n_2842),
.Y(n_4608)
);

OAI21xp5_ASAP7_75t_L g4609 ( 
.A1(n_3782),
.A2(n_3191),
.B(n_3113),
.Y(n_4609)
);

HB1xp67_ASAP7_75t_L g4610 ( 
.A(n_3667),
.Y(n_4610)
);

AOI21xp5_ASAP7_75t_L g4611 ( 
.A1(n_3733),
.A2(n_3148),
.B(n_3120),
.Y(n_4611)
);

OAI21x1_ASAP7_75t_L g4612 ( 
.A1(n_4283),
.A2(n_3422),
.B(n_3420),
.Y(n_4612)
);

OAI22xp5_ASAP7_75t_L g4613 ( 
.A1(n_4304),
.A2(n_2751),
.B1(n_2881),
.B2(n_2684),
.Y(n_4613)
);

INVx2_ASAP7_75t_L g4614 ( 
.A(n_3817),
.Y(n_4614)
);

BUFx2_ASAP7_75t_L g4615 ( 
.A(n_3749),
.Y(n_4615)
);

AOI21xp5_ASAP7_75t_L g4616 ( 
.A1(n_4044),
.A2(n_3148),
.B(n_3120),
.Y(n_4616)
);

INVx1_ASAP7_75t_L g4617 ( 
.A(n_3817),
.Y(n_4617)
);

INVx2_ASAP7_75t_L g4618 ( 
.A(n_3837),
.Y(n_4618)
);

BUFx6f_ASAP7_75t_L g4619 ( 
.A(n_4226),
.Y(n_4619)
);

OAI22xp5_ASAP7_75t_L g4620 ( 
.A1(n_4304),
.A2(n_2751),
.B1(n_2881),
.B2(n_2684),
.Y(n_4620)
);

AOI22xp5_ASAP7_75t_L g4621 ( 
.A1(n_4103),
.A2(n_3353),
.B1(n_3018),
.B2(n_2842),
.Y(n_4621)
);

INVx1_ASAP7_75t_L g4622 ( 
.A(n_3837),
.Y(n_4622)
);

OAI21xp5_ASAP7_75t_L g4623 ( 
.A1(n_3743),
.A2(n_3191),
.B(n_3385),
.Y(n_4623)
);

NAND2xp5_ASAP7_75t_L g4624 ( 
.A(n_4128),
.B(n_2979),
.Y(n_4624)
);

INVx1_ASAP7_75t_L g4625 ( 
.A(n_3837),
.Y(n_4625)
);

AOI21xp5_ASAP7_75t_L g4626 ( 
.A1(n_4053),
.A2(n_3148),
.B(n_3120),
.Y(n_4626)
);

INVx1_ASAP7_75t_L g4627 ( 
.A(n_3862),
.Y(n_4627)
);

O2A1O1Ixp5_ASAP7_75t_L g4628 ( 
.A1(n_3796),
.A2(n_2855),
.B(n_2840),
.C(n_3249),
.Y(n_4628)
);

AOI21xp5_ASAP7_75t_L g4629 ( 
.A1(n_4053),
.A2(n_3120),
.B(n_3367),
.Y(n_4629)
);

NAND2xp5_ASAP7_75t_L g4630 ( 
.A(n_4102),
.B(n_2979),
.Y(n_4630)
);

INVx2_ASAP7_75t_SL g4631 ( 
.A(n_4226),
.Y(n_4631)
);

NAND2xp5_ASAP7_75t_L g4632 ( 
.A(n_4102),
.B(n_2979),
.Y(n_4632)
);

INVx1_ASAP7_75t_SL g4633 ( 
.A(n_3722),
.Y(n_4633)
);

AOI21xp5_ASAP7_75t_L g4634 ( 
.A1(n_4099),
.A2(n_3120),
.B(n_3367),
.Y(n_4634)
);

NAND2xp5_ASAP7_75t_L g4635 ( 
.A(n_3906),
.B(n_3910),
.Y(n_4635)
);

INVx2_ASAP7_75t_SL g4636 ( 
.A(n_4226),
.Y(n_4636)
);

HB1xp67_ASAP7_75t_L g4637 ( 
.A(n_3667),
.Y(n_4637)
);

INVx2_ASAP7_75t_L g4638 ( 
.A(n_3862),
.Y(n_4638)
);

INVx2_ASAP7_75t_SL g4639 ( 
.A(n_4226),
.Y(n_4639)
);

NAND2xp5_ASAP7_75t_L g4640 ( 
.A(n_3906),
.B(n_3388),
.Y(n_4640)
);

AOI21xp5_ASAP7_75t_L g4641 ( 
.A1(n_4099),
.A2(n_3120),
.B(n_3367),
.Y(n_4641)
);

AND2x4_ASAP7_75t_L g4642 ( 
.A(n_3900),
.B(n_3366),
.Y(n_4642)
);

AOI21x1_ASAP7_75t_L g4643 ( 
.A1(n_3498),
.A2(n_3366),
.B(n_3293),
.Y(n_4643)
);

INVx1_ASAP7_75t_L g4644 ( 
.A(n_3862),
.Y(n_4644)
);

AOI21xp5_ASAP7_75t_L g4645 ( 
.A1(n_4195),
.A2(n_3367),
.B(n_3211),
.Y(n_4645)
);

INVx1_ASAP7_75t_L g4646 ( 
.A(n_3867),
.Y(n_4646)
);

O2A1O1Ixp5_ASAP7_75t_L g4647 ( 
.A1(n_3796),
.A2(n_2855),
.B(n_2840),
.C(n_3249),
.Y(n_4647)
);

OAI21x1_ASAP7_75t_L g4648 ( 
.A1(n_4292),
.A2(n_4297),
.B(n_3607),
.Y(n_4648)
);

OAI21xp5_ASAP7_75t_L g4649 ( 
.A1(n_3761),
.A2(n_3191),
.B(n_3396),
.Y(n_4649)
);

AOI21xp5_ASAP7_75t_L g4650 ( 
.A1(n_4195),
.A2(n_3367),
.B(n_3211),
.Y(n_4650)
);

OAI21x1_ASAP7_75t_L g4651 ( 
.A1(n_3607),
.A2(n_2855),
.B(n_2840),
.Y(n_4651)
);

NOR2xp33_ASAP7_75t_L g4652 ( 
.A(n_3935),
.B(n_3423),
.Y(n_4652)
);

OAI21xp5_ASAP7_75t_L g4653 ( 
.A1(n_3661),
.A2(n_3191),
.B(n_3396),
.Y(n_4653)
);

OAI21xp33_ASAP7_75t_L g4654 ( 
.A1(n_3779),
.A2(n_3318),
.B(n_3291),
.Y(n_4654)
);

AOI21xp5_ASAP7_75t_L g4655 ( 
.A1(n_4250),
.A2(n_3367),
.B(n_3211),
.Y(n_4655)
);

AOI21xp33_ASAP7_75t_L g4656 ( 
.A1(n_3697),
.A2(n_3436),
.B(n_3395),
.Y(n_4656)
);

AOI21xp5_ASAP7_75t_L g4657 ( 
.A1(n_4250),
.A2(n_3213),
.B(n_3183),
.Y(n_4657)
);

OAI21x1_ASAP7_75t_L g4658 ( 
.A1(n_4255),
.A2(n_2855),
.B(n_2840),
.Y(n_4658)
);

NAND2xp5_ASAP7_75t_SL g4659 ( 
.A(n_3697),
.B(n_3436),
.Y(n_4659)
);

A2O1A1Ixp33_ASAP7_75t_L g4660 ( 
.A1(n_4172),
.A2(n_3287),
.B(n_3286),
.C(n_3213),
.Y(n_4660)
);

AOI21xp5_ASAP7_75t_SL g4661 ( 
.A1(n_3601),
.A2(n_3246),
.B(n_3191),
.Y(n_4661)
);

OA22x2_ASAP7_75t_L g4662 ( 
.A1(n_4263),
.A2(n_3065),
.B1(n_3078),
.B2(n_3047),
.Y(n_4662)
);

NAND2xp5_ASAP7_75t_L g4663 ( 
.A(n_3910),
.B(n_3253),
.Y(n_4663)
);

AOI21xp5_ASAP7_75t_L g4664 ( 
.A1(n_4255),
.A2(n_3213),
.B(n_3183),
.Y(n_4664)
);

NAND2xp5_ASAP7_75t_L g4665 ( 
.A(n_4015),
.B(n_3253),
.Y(n_4665)
);

OAI21xp5_ASAP7_75t_L g4666 ( 
.A1(n_3661),
.A2(n_2831),
.B(n_2824),
.Y(n_4666)
);

AND3x4_ASAP7_75t_L g4667 ( 
.A(n_4111),
.B(n_3065),
.C(n_3047),
.Y(n_4667)
);

A2O1A1Ixp33_ASAP7_75t_L g4668 ( 
.A1(n_4320),
.A2(n_3287),
.B(n_3286),
.C(n_3213),
.Y(n_4668)
);

OAI21x1_ASAP7_75t_L g4669 ( 
.A1(n_4312),
.A2(n_2855),
.B(n_2840),
.Y(n_4669)
);

NAND2xp5_ASAP7_75t_L g4670 ( 
.A(n_4015),
.B(n_3256),
.Y(n_4670)
);

OA21x2_ASAP7_75t_L g4671 ( 
.A1(n_4051),
.A2(n_3262),
.B(n_3256),
.Y(n_4671)
);

BUFx2_ASAP7_75t_L g4672 ( 
.A(n_3749),
.Y(n_4672)
);

NAND2xp5_ASAP7_75t_L g4673 ( 
.A(n_4056),
.B(n_3262),
.Y(n_4673)
);

NAND2xp5_ASAP7_75t_L g4674 ( 
.A(n_4056),
.B(n_3262),
.Y(n_4674)
);

BUFx6f_ASAP7_75t_L g4675 ( 
.A(n_4226),
.Y(n_4675)
);

AND2x2_ASAP7_75t_L g4676 ( 
.A(n_3900),
.B(n_4284),
.Y(n_4676)
);

NAND2x1p5_ASAP7_75t_L g4677 ( 
.A(n_4286),
.B(n_2794),
.Y(n_4677)
);

NAND2x1p5_ASAP7_75t_L g4678 ( 
.A(n_4286),
.B(n_4319),
.Y(n_4678)
);

AND2x2_ASAP7_75t_L g4679 ( 
.A(n_3900),
.B(n_2703),
.Y(n_4679)
);

O2A1O1Ixp5_ASAP7_75t_L g4680 ( 
.A1(n_3800),
.A2(n_3255),
.B(n_3249),
.C(n_2889),
.Y(n_4680)
);

INVxp67_ASAP7_75t_SL g4681 ( 
.A(n_4278),
.Y(n_4681)
);

BUFx2_ASAP7_75t_L g4682 ( 
.A(n_3749),
.Y(n_4682)
);

AOI21xp5_ASAP7_75t_L g4683 ( 
.A1(n_3893),
.A2(n_3213),
.B(n_3183),
.Y(n_4683)
);

OAI22xp5_ASAP7_75t_SL g4684 ( 
.A1(n_4103),
.A2(n_3047),
.B1(n_3078),
.B2(n_3065),
.Y(n_4684)
);

OAI21xp33_ASAP7_75t_L g4685 ( 
.A1(n_3783),
.A2(n_3318),
.B(n_3291),
.Y(n_4685)
);

NAND2xp5_ASAP7_75t_L g4686 ( 
.A(n_3806),
.B(n_3270),
.Y(n_4686)
);

OAI22xp5_ASAP7_75t_L g4687 ( 
.A1(n_4304),
.A2(n_2751),
.B1(n_2881),
.B2(n_2684),
.Y(n_4687)
);

AOI21xp5_ASAP7_75t_L g4688 ( 
.A1(n_3893),
.A2(n_3805),
.B(n_3795),
.Y(n_4688)
);

O2A1O1Ixp5_ASAP7_75t_L g4689 ( 
.A1(n_3791),
.A2(n_3255),
.B(n_3249),
.C(n_2889),
.Y(n_4689)
);

INVxp67_ASAP7_75t_SL g4690 ( 
.A(n_4278),
.Y(n_4690)
);

NAND2xp5_ASAP7_75t_L g4691 ( 
.A(n_3806),
.B(n_3270),
.Y(n_4691)
);

NAND2xp5_ASAP7_75t_L g4692 ( 
.A(n_3915),
.B(n_3270),
.Y(n_4692)
);

NAND2xp5_ASAP7_75t_SL g4693 ( 
.A(n_3619),
.B(n_3436),
.Y(n_4693)
);

OAI21x1_ASAP7_75t_SL g4694 ( 
.A1(n_4032),
.A2(n_2759),
.B(n_2740),
.Y(n_4694)
);

HB1xp67_ASAP7_75t_L g4695 ( 
.A(n_4238),
.Y(n_4695)
);

NAND2xp5_ASAP7_75t_L g4696 ( 
.A(n_3915),
.B(n_3280),
.Y(n_4696)
);

NAND2xp5_ASAP7_75t_L g4697 ( 
.A(n_3927),
.B(n_3280),
.Y(n_4697)
);

BUFx5_ASAP7_75t_L g4698 ( 
.A(n_3598),
.Y(n_4698)
);

OAI21x1_ASAP7_75t_SL g4699 ( 
.A1(n_4032),
.A2(n_2759),
.B(n_2740),
.Y(n_4699)
);

NAND2xp5_ASAP7_75t_L g4700 ( 
.A(n_3927),
.B(n_3280),
.Y(n_4700)
);

NAND2xp5_ASAP7_75t_L g4701 ( 
.A(n_3895),
.B(n_3283),
.Y(n_4701)
);

INVx1_ASAP7_75t_L g4702 ( 
.A(n_3867),
.Y(n_4702)
);

NAND2xp5_ASAP7_75t_L g4703 ( 
.A(n_3895),
.B(n_3283),
.Y(n_4703)
);

AOI21x1_ASAP7_75t_SL g4704 ( 
.A1(n_3544),
.A2(n_3255),
.B(n_3249),
.Y(n_4704)
);

INVx3_ASAP7_75t_L g4705 ( 
.A(n_4226),
.Y(n_4705)
);

OAI22xp5_ASAP7_75t_L g4706 ( 
.A1(n_4304),
.A2(n_4352),
.B1(n_3786),
.B2(n_4085),
.Y(n_4706)
);

BUFx3_ASAP7_75t_L g4707 ( 
.A(n_4240),
.Y(n_4707)
);

NAND2xp5_ASAP7_75t_SL g4708 ( 
.A(n_3619),
.B(n_3436),
.Y(n_4708)
);

NAND2x1p5_ASAP7_75t_L g4709 ( 
.A(n_4319),
.B(n_2794),
.Y(n_4709)
);

INVx2_ASAP7_75t_L g4710 ( 
.A(n_3867),
.Y(n_4710)
);

OAI21xp33_ASAP7_75t_SL g4711 ( 
.A1(n_4352),
.A2(n_2759),
.B(n_2824),
.Y(n_4711)
);

NOR2xp33_ASAP7_75t_L g4712 ( 
.A(n_3926),
.B(n_3922),
.Y(n_4712)
);

AOI22xp5_ASAP7_75t_L g4713 ( 
.A1(n_3822),
.A2(n_3018),
.B1(n_2842),
.B2(n_2847),
.Y(n_4713)
);

OAI21x1_ASAP7_75t_L g4714 ( 
.A1(n_4346),
.A2(n_2726),
.B(n_2725),
.Y(n_4714)
);

AOI21xp5_ASAP7_75t_L g4715 ( 
.A1(n_3795),
.A2(n_3218),
.B(n_3183),
.Y(n_4715)
);

NAND2xp5_ASAP7_75t_L g4716 ( 
.A(n_3838),
.B(n_3283),
.Y(n_4716)
);

OAI21x1_ASAP7_75t_L g4717 ( 
.A1(n_4346),
.A2(n_2736),
.B(n_2726),
.Y(n_4717)
);

BUFx6f_ASAP7_75t_L g4718 ( 
.A(n_4233),
.Y(n_4718)
);

AOI211x1_ASAP7_75t_L g4719 ( 
.A1(n_3868),
.A2(n_3321),
.B(n_3325),
.C(n_3318),
.Y(n_4719)
);

BUFx3_ASAP7_75t_L g4720 ( 
.A(n_3801),
.Y(n_4720)
);

AOI21x1_ASAP7_75t_L g4721 ( 
.A1(n_3884),
.A2(n_4301),
.B(n_4264),
.Y(n_4721)
);

NAND2xp5_ASAP7_75t_L g4722 ( 
.A(n_4033),
.B(n_3285),
.Y(n_4722)
);

NOR2xp33_ASAP7_75t_L g4723 ( 
.A(n_3926),
.B(n_3423),
.Y(n_4723)
);

AOI21xp5_ASAP7_75t_L g4724 ( 
.A1(n_3805),
.A2(n_3218),
.B(n_3183),
.Y(n_4724)
);

NAND2xp5_ASAP7_75t_L g4725 ( 
.A(n_4033),
.B(n_3285),
.Y(n_4725)
);

OAI21xp5_ASAP7_75t_L g4726 ( 
.A1(n_3812),
.A2(n_2831),
.B(n_2824),
.Y(n_4726)
);

NAND2x1p5_ASAP7_75t_L g4727 ( 
.A(n_4319),
.B(n_2794),
.Y(n_4727)
);

OAI21xp5_ASAP7_75t_L g4728 ( 
.A1(n_3868),
.A2(n_2831),
.B(n_2824),
.Y(n_4728)
);

BUFx3_ASAP7_75t_L g4729 ( 
.A(n_3801),
.Y(n_4729)
);

AOI21xp5_ASAP7_75t_L g4730 ( 
.A1(n_3808),
.A2(n_3222),
.B(n_3218),
.Y(n_4730)
);

NOR2xp33_ASAP7_75t_L g4731 ( 
.A(n_3922),
.B(n_3423),
.Y(n_4731)
);

AOI21xp5_ASAP7_75t_SL g4732 ( 
.A1(n_3555),
.A2(n_3246),
.B(n_3442),
.Y(n_4732)
);

NAND2xp5_ASAP7_75t_L g4733 ( 
.A(n_3875),
.B(n_3285),
.Y(n_4733)
);

OAI21x1_ASAP7_75t_L g4734 ( 
.A1(n_3978),
.A2(n_2743),
.B(n_2736),
.Y(n_4734)
);

OAI22xp5_ASAP7_75t_L g4735 ( 
.A1(n_4352),
.A2(n_2684),
.B1(n_2881),
.B2(n_2751),
.Y(n_4735)
);

INVxp67_ASAP7_75t_SL g4736 ( 
.A(n_3870),
.Y(n_4736)
);

OAI21x1_ASAP7_75t_L g4737 ( 
.A1(n_3978),
.A2(n_2750),
.B(n_2743),
.Y(n_4737)
);

NAND2x1_ASAP7_75t_L g4738 ( 
.A(n_3586),
.B(n_3108),
.Y(n_4738)
);

NAND2xp5_ASAP7_75t_L g4739 ( 
.A(n_3875),
.B(n_3298),
.Y(n_4739)
);

INVx3_ASAP7_75t_L g4740 ( 
.A(n_4233),
.Y(n_4740)
);

BUFx4f_ASAP7_75t_L g4741 ( 
.A(n_4152),
.Y(n_4741)
);

AO22x2_ASAP7_75t_L g4742 ( 
.A1(n_4194),
.A2(n_3065),
.B1(n_3078),
.B2(n_3047),
.Y(n_4742)
);

AND2x4_ASAP7_75t_L g4743 ( 
.A(n_3479),
.B(n_2798),
.Y(n_4743)
);

NOR2xp33_ASAP7_75t_L g4744 ( 
.A(n_3849),
.B(n_3423),
.Y(n_4744)
);

NAND2xp5_ASAP7_75t_L g4745 ( 
.A(n_3903),
.B(n_3298),
.Y(n_4745)
);

INVxp67_ASAP7_75t_L g4746 ( 
.A(n_4199),
.Y(n_4746)
);

AOI21xp5_ASAP7_75t_L g4747 ( 
.A1(n_3808),
.A2(n_3222),
.B(n_3218),
.Y(n_4747)
);

AOI21xp5_ASAP7_75t_L g4748 ( 
.A1(n_3816),
.A2(n_3222),
.B(n_3218),
.Y(n_4748)
);

NAND2xp5_ASAP7_75t_L g4749 ( 
.A(n_3903),
.B(n_3298),
.Y(n_4749)
);

NAND2xp5_ASAP7_75t_L g4750 ( 
.A(n_3912),
.B(n_3300),
.Y(n_4750)
);

NAND2xp5_ASAP7_75t_L g4751 ( 
.A(n_3912),
.B(n_4006),
.Y(n_4751)
);

NAND2xp5_ASAP7_75t_L g4752 ( 
.A(n_4006),
.B(n_3300),
.Y(n_4752)
);

AOI21xp5_ASAP7_75t_L g4753 ( 
.A1(n_3816),
.A2(n_3489),
.B(n_3916),
.Y(n_4753)
);

INVxp67_ASAP7_75t_SL g4754 ( 
.A(n_3870),
.Y(n_4754)
);

AOI22xp5_ASAP7_75t_L g4755 ( 
.A1(n_3822),
.A2(n_3833),
.B1(n_3846),
.B2(n_3840),
.Y(n_4755)
);

BUFx2_ASAP7_75t_L g4756 ( 
.A(n_3749),
.Y(n_4756)
);

INVx2_ASAP7_75t_L g4757 ( 
.A(n_3869),
.Y(n_4757)
);

INVx1_ASAP7_75t_L g4758 ( 
.A(n_3869),
.Y(n_4758)
);

AND2x2_ASAP7_75t_SL g4759 ( 
.A(n_3939),
.B(n_2859),
.Y(n_4759)
);

NAND2xp5_ASAP7_75t_L g4760 ( 
.A(n_4008),
.B(n_3300),
.Y(n_4760)
);

OAI21x1_ASAP7_75t_L g4761 ( 
.A1(n_4264),
.A2(n_2761),
.B(n_2750),
.Y(n_4761)
);

INVx2_ASAP7_75t_L g4762 ( 
.A(n_3869),
.Y(n_4762)
);

BUFx2_ASAP7_75t_L g4763 ( 
.A(n_3749),
.Y(n_4763)
);

BUFx3_ASAP7_75t_L g4764 ( 
.A(n_3801),
.Y(n_4764)
);

NAND2xp5_ASAP7_75t_L g4765 ( 
.A(n_4008),
.B(n_3301),
.Y(n_4765)
);

BUFx3_ASAP7_75t_L g4766 ( 
.A(n_3991),
.Y(n_4766)
);

OA21x2_ASAP7_75t_L g4767 ( 
.A1(n_4202),
.A2(n_3305),
.B(n_3301),
.Y(n_4767)
);

AND3x4_ASAP7_75t_L g4768 ( 
.A(n_4161),
.B(n_3078),
.C(n_3047),
.Y(n_4768)
);

BUFx3_ASAP7_75t_L g4769 ( 
.A(n_3991),
.Y(n_4769)
);

AOI21xp5_ASAP7_75t_L g4770 ( 
.A1(n_3489),
.A2(n_3237),
.B(n_3222),
.Y(n_4770)
);

OA21x2_ASAP7_75t_L g4771 ( 
.A1(n_4202),
.A2(n_3865),
.B(n_3552),
.Y(n_4771)
);

INVx1_ASAP7_75t_L g4772 ( 
.A(n_3877),
.Y(n_4772)
);

NAND2xp5_ASAP7_75t_L g4773 ( 
.A(n_4029),
.B(n_3301),
.Y(n_4773)
);

CKINVDCx8_ASAP7_75t_R g4774 ( 
.A(n_4007),
.Y(n_4774)
);

BUFx4f_ASAP7_75t_L g4775 ( 
.A(n_4152),
.Y(n_4775)
);

OA22x2_ASAP7_75t_L g4776 ( 
.A1(n_4322),
.A2(n_3404),
.B1(n_3428),
.B2(n_3427),
.Y(n_4776)
);

AND2x4_ASAP7_75t_L g4777 ( 
.A(n_3479),
.B(n_2798),
.Y(n_4777)
);

INVx1_ASAP7_75t_SL g4778 ( 
.A(n_3722),
.Y(n_4778)
);

AOI21xp5_ASAP7_75t_L g4779 ( 
.A1(n_3916),
.A2(n_3237),
.B(n_3222),
.Y(n_4779)
);

BUFx6f_ASAP7_75t_L g4780 ( 
.A(n_4233),
.Y(n_4780)
);

INVx1_ASAP7_75t_L g4781 ( 
.A(n_3877),
.Y(n_4781)
);

INVx1_ASAP7_75t_L g4782 ( 
.A(n_3877),
.Y(n_4782)
);

AOI21xp5_ASAP7_75t_L g4783 ( 
.A1(n_3928),
.A2(n_3237),
.B(n_2805),
.Y(n_4783)
);

NAND2xp5_ASAP7_75t_L g4784 ( 
.A(n_4029),
.B(n_3305),
.Y(n_4784)
);

OAI21x1_ASAP7_75t_L g4785 ( 
.A1(n_4100),
.A2(n_3483),
.B(n_4156),
.Y(n_4785)
);

NAND2xp5_ASAP7_75t_L g4786 ( 
.A(n_4060),
.B(n_3305),
.Y(n_4786)
);

AOI21x1_ASAP7_75t_SL g4787 ( 
.A1(n_3544),
.A2(n_3255),
.B(n_3249),
.Y(n_4787)
);

INVx1_ASAP7_75t_L g4788 ( 
.A(n_3880),
.Y(n_4788)
);

AO21x1_ASAP7_75t_L g4789 ( 
.A1(n_4259),
.A2(n_3319),
.B(n_3308),
.Y(n_4789)
);

INVxp67_ASAP7_75t_SL g4790 ( 
.A(n_3871),
.Y(n_4790)
);

INVxp67_ASAP7_75t_SL g4791 ( 
.A(n_3871),
.Y(n_4791)
);

NAND2xp5_ASAP7_75t_L g4792 ( 
.A(n_4060),
.B(n_3308),
.Y(n_4792)
);

OAI21xp5_ASAP7_75t_L g4793 ( 
.A1(n_3638),
.A2(n_3428),
.B(n_3427),
.Y(n_4793)
);

NAND2xp5_ASAP7_75t_L g4794 ( 
.A(n_4074),
.B(n_3308),
.Y(n_4794)
);

NOR2xp33_ASAP7_75t_L g4795 ( 
.A(n_3578),
.B(n_3423),
.Y(n_4795)
);

NAND2xp5_ASAP7_75t_L g4796 ( 
.A(n_4074),
.B(n_3319),
.Y(n_4796)
);

NAND2xp5_ASAP7_75t_L g4797 ( 
.A(n_4077),
.B(n_3319),
.Y(n_4797)
);

INVx4_ASAP7_75t_L g4798 ( 
.A(n_4094),
.Y(n_4798)
);

OAI21xp5_ASAP7_75t_L g4799 ( 
.A1(n_3638),
.A2(n_3428),
.B(n_3427),
.Y(n_4799)
);

OAI21xp5_ASAP7_75t_L g4800 ( 
.A1(n_3646),
.A2(n_3428),
.B(n_3427),
.Y(n_4800)
);

AOI21xp5_ASAP7_75t_SL g4801 ( 
.A1(n_3810),
.A2(n_3246),
.B(n_3442),
.Y(n_4801)
);

NAND2xp5_ASAP7_75t_L g4802 ( 
.A(n_4077),
.B(n_3324),
.Y(n_4802)
);

NAND2xp5_ASAP7_75t_L g4803 ( 
.A(n_4089),
.B(n_3324),
.Y(n_4803)
);

NAND2xp5_ASAP7_75t_L g4804 ( 
.A(n_4089),
.B(n_3324),
.Y(n_4804)
);

NOR2xp33_ASAP7_75t_L g4805 ( 
.A(n_4086),
.B(n_3423),
.Y(n_4805)
);

CKINVDCx20_ASAP7_75t_R g4806 ( 
.A(n_3920),
.Y(n_4806)
);

AOI21xp5_ASAP7_75t_L g4807 ( 
.A1(n_3928),
.A2(n_3237),
.B(n_2805),
.Y(n_4807)
);

INVx1_ASAP7_75t_L g4808 ( 
.A(n_3880),
.Y(n_4808)
);

NOR2xp67_ASAP7_75t_L g4809 ( 
.A(n_4293),
.B(n_3452),
.Y(n_4809)
);

INVx1_ASAP7_75t_L g4810 ( 
.A(n_3880),
.Y(n_4810)
);

HB1xp67_ASAP7_75t_L g4811 ( 
.A(n_4238),
.Y(n_4811)
);

NAND2xp5_ASAP7_75t_L g4812 ( 
.A(n_3941),
.B(n_3332),
.Y(n_4812)
);

OAI22xp5_ASAP7_75t_L g4813 ( 
.A1(n_3594),
.A2(n_2903),
.B1(n_2948),
.B2(n_2921),
.Y(n_4813)
);

A2O1A1Ixp33_ASAP7_75t_L g4814 ( 
.A1(n_4320),
.A2(n_3622),
.B(n_4347),
.C(n_4160),
.Y(n_4814)
);

INVx2_ASAP7_75t_SL g4815 ( 
.A(n_4233),
.Y(n_4815)
);

OAI21xp5_ASAP7_75t_L g4816 ( 
.A1(n_3646),
.A2(n_3592),
.B(n_3510),
.Y(n_4816)
);

NOR2x1_ASAP7_75t_L g4817 ( 
.A(n_4217),
.B(n_3112),
.Y(n_4817)
);

AOI21x1_ASAP7_75t_L g4818 ( 
.A1(n_3884),
.A2(n_3325),
.B(n_3321),
.Y(n_4818)
);

INVx1_ASAP7_75t_L g4819 ( 
.A(n_3907),
.Y(n_4819)
);

AO21x1_ASAP7_75t_L g4820 ( 
.A1(n_4259),
.A2(n_3340),
.B(n_3332),
.Y(n_4820)
);

NOR2x1_ASAP7_75t_L g4821 ( 
.A(n_4217),
.B(n_3112),
.Y(n_4821)
);

INVxp67_ASAP7_75t_L g4822 ( 
.A(n_4199),
.Y(n_4822)
);

OAI22xp5_ASAP7_75t_L g4823 ( 
.A1(n_3594),
.A2(n_2903),
.B1(n_2948),
.B2(n_2921),
.Y(n_4823)
);

OAI21x1_ASAP7_75t_L g4824 ( 
.A1(n_4170),
.A2(n_4183),
.B(n_4171),
.Y(n_4824)
);

NAND2x1p5_ASAP7_75t_L g4825 ( 
.A(n_4319),
.B(n_2798),
.Y(n_4825)
);

NAND2xp5_ASAP7_75t_L g4826 ( 
.A(n_3941),
.B(n_3332),
.Y(n_4826)
);

AOI21xp5_ASAP7_75t_L g4827 ( 
.A1(n_3929),
.A2(n_3947),
.B(n_3940),
.Y(n_4827)
);

OAI22xp5_ASAP7_75t_L g4828 ( 
.A1(n_3478),
.A2(n_2903),
.B1(n_2948),
.B2(n_2921),
.Y(n_4828)
);

AOI21xp5_ASAP7_75t_L g4829 ( 
.A1(n_3929),
.A2(n_3947),
.B(n_3940),
.Y(n_4829)
);

OAI21xp5_ASAP7_75t_L g4830 ( 
.A1(n_3592),
.A2(n_3455),
.B(n_3452),
.Y(n_4830)
);

INVx2_ASAP7_75t_L g4831 ( 
.A(n_3907),
.Y(n_4831)
);

OAI21x1_ASAP7_75t_L g4832 ( 
.A1(n_4171),
.A2(n_4183),
.B(n_3874),
.Y(n_4832)
);

AOI21xp5_ASAP7_75t_SL g4833 ( 
.A1(n_3810),
.A2(n_3246),
.B(n_3442),
.Y(n_4833)
);

A2O1A1Ixp33_ASAP7_75t_L g4834 ( 
.A1(n_3622),
.A2(n_3287),
.B(n_3237),
.C(n_2798),
.Y(n_4834)
);

NAND2xp5_ASAP7_75t_L g4835 ( 
.A(n_3951),
.B(n_3340),
.Y(n_4835)
);

NAND2xp5_ASAP7_75t_L g4836 ( 
.A(n_3951),
.B(n_3340),
.Y(n_4836)
);

AOI21xp5_ASAP7_75t_L g4837 ( 
.A1(n_3952),
.A2(n_2805),
.B(n_2798),
.Y(n_4837)
);

INVx1_ASAP7_75t_L g4838 ( 
.A(n_3907),
.Y(n_4838)
);

NAND2xp5_ASAP7_75t_L g4839 ( 
.A(n_3969),
.B(n_3343),
.Y(n_4839)
);

NOR2xp67_ASAP7_75t_SL g4840 ( 
.A(n_4314),
.B(n_2903),
.Y(n_4840)
);

NAND2xp5_ASAP7_75t_L g4841 ( 
.A(n_3969),
.B(n_3343),
.Y(n_4841)
);

NOR2x1_ASAP7_75t_SL g4842 ( 
.A(n_3931),
.B(n_2718),
.Y(n_4842)
);

AOI21xp33_ASAP7_75t_L g4843 ( 
.A1(n_3854),
.A2(n_3436),
.B(n_3395),
.Y(n_4843)
);

INVx2_ASAP7_75t_SL g4844 ( 
.A(n_4241),
.Y(n_4844)
);

NAND2xp5_ASAP7_75t_L g4845 ( 
.A(n_3954),
.B(n_3343),
.Y(n_4845)
);

AOI21xp5_ASAP7_75t_L g4846 ( 
.A1(n_3952),
.A2(n_3766),
.B(n_3765),
.Y(n_4846)
);

NAND2xp5_ASAP7_75t_L g4847 ( 
.A(n_3954),
.B(n_3346),
.Y(n_4847)
);

NOR2xp67_ASAP7_75t_SL g4848 ( 
.A(n_4314),
.B(n_2903),
.Y(n_4848)
);

OAI22xp5_ASAP7_75t_L g4849 ( 
.A1(n_3548),
.A2(n_2903),
.B1(n_2948),
.B2(n_2921),
.Y(n_4849)
);

BUFx2_ASAP7_75t_L g4850 ( 
.A(n_3985),
.Y(n_4850)
);

A2O1A1Ixp33_ASAP7_75t_L g4851 ( 
.A1(n_4347),
.A2(n_2812),
.B(n_2822),
.C(n_2805),
.Y(n_4851)
);

O2A1O1Ixp33_ASAP7_75t_L g4852 ( 
.A1(n_3843),
.A2(n_3321),
.B(n_3327),
.C(n_3325),
.Y(n_4852)
);

NAND2xp5_ASAP7_75t_L g4853 ( 
.A(n_4062),
.B(n_3346),
.Y(n_4853)
);

INVx3_ASAP7_75t_L g4854 ( 
.A(n_4241),
.Y(n_4854)
);

AND2x2_ASAP7_75t_L g4855 ( 
.A(n_3703),
.B(n_2799),
.Y(n_4855)
);

NAND2xp5_ASAP7_75t_L g4856 ( 
.A(n_4062),
.B(n_3346),
.Y(n_4856)
);

BUFx3_ASAP7_75t_L g4857 ( 
.A(n_3991),
.Y(n_4857)
);

INVx1_ASAP7_75t_L g4858 ( 
.A(n_3918),
.Y(n_4858)
);

INVx2_ASAP7_75t_SL g4859 ( 
.A(n_4241),
.Y(n_4859)
);

NAND2xp5_ASAP7_75t_L g4860 ( 
.A(n_4065),
.B(n_3352),
.Y(n_4860)
);

NAND2xp5_ASAP7_75t_L g4861 ( 
.A(n_4065),
.B(n_4139),
.Y(n_4861)
);

INVx1_ASAP7_75t_L g4862 ( 
.A(n_3918),
.Y(n_4862)
);

A2O1A1Ixp33_ASAP7_75t_L g4863 ( 
.A1(n_4118),
.A2(n_2812),
.B(n_2822),
.C(n_2903),
.Y(n_4863)
);

HB1xp67_ASAP7_75t_L g4864 ( 
.A(n_4247),
.Y(n_4864)
);

AOI21xp5_ASAP7_75t_L g4865 ( 
.A1(n_3766),
.A2(n_2822),
.B(n_2812),
.Y(n_4865)
);

INVx2_ASAP7_75t_L g4866 ( 
.A(n_3918),
.Y(n_4866)
);

AND2x4_ASAP7_75t_L g4867 ( 
.A(n_3479),
.B(n_2822),
.Y(n_4867)
);

NAND2xp5_ASAP7_75t_L g4868 ( 
.A(n_4139),
.B(n_3352),
.Y(n_4868)
);

NAND2xp5_ASAP7_75t_L g4869 ( 
.A(n_4143),
.B(n_4215),
.Y(n_4869)
);

INVx2_ASAP7_75t_L g4870 ( 
.A(n_3934),
.Y(n_4870)
);

NAND2xp5_ASAP7_75t_L g4871 ( 
.A(n_4143),
.B(n_4215),
.Y(n_4871)
);

NAND2xp5_ASAP7_75t_L g4872 ( 
.A(n_4221),
.B(n_3352),
.Y(n_4872)
);

NAND2xp5_ASAP7_75t_L g4873 ( 
.A(n_4221),
.B(n_3355),
.Y(n_4873)
);

AOI21xp5_ASAP7_75t_L g4874 ( 
.A1(n_3492),
.A2(n_3246),
.B(n_3249),
.Y(n_4874)
);

INVx1_ASAP7_75t_L g4875 ( 
.A(n_3934),
.Y(n_4875)
);

OAI21xp5_ASAP7_75t_L g4876 ( 
.A1(n_3510),
.A2(n_3455),
.B(n_3452),
.Y(n_4876)
);

OAI21x1_ASAP7_75t_L g4877 ( 
.A1(n_3887),
.A2(n_3891),
.B(n_3888),
.Y(n_4877)
);

AND2x2_ASAP7_75t_L g4878 ( 
.A(n_3703),
.B(n_2802),
.Y(n_4878)
);

CKINVDCx5p33_ASAP7_75t_R g4879 ( 
.A(n_3617),
.Y(n_4879)
);

AND2x4_ASAP7_75t_L g4880 ( 
.A(n_3479),
.B(n_2921),
.Y(n_4880)
);

AOI21x1_ASAP7_75t_L g4881 ( 
.A1(n_3498),
.A2(n_3328),
.B(n_3327),
.Y(n_4881)
);

NAND2xp5_ASAP7_75t_SL g4882 ( 
.A(n_3636),
.B(n_3423),
.Y(n_4882)
);

AOI21xp5_ASAP7_75t_L g4883 ( 
.A1(n_3492),
.A2(n_3246),
.B(n_3255),
.Y(n_4883)
);

NAND2xp5_ASAP7_75t_SL g4884 ( 
.A(n_3854),
.B(n_3423),
.Y(n_4884)
);

INVx1_ASAP7_75t_L g4885 ( 
.A(n_3934),
.Y(n_4885)
);

INVx5_ASAP7_75t_L g4886 ( 
.A(n_3703),
.Y(n_4886)
);

AND2x2_ASAP7_75t_L g4887 ( 
.A(n_4274),
.B(n_2802),
.Y(n_4887)
);

INVx2_ASAP7_75t_L g4888 ( 
.A(n_3937),
.Y(n_4888)
);

INVx3_ASAP7_75t_L g4889 ( 
.A(n_4248),
.Y(n_4889)
);

NAND2xp5_ASAP7_75t_L g4890 ( 
.A(n_4072),
.B(n_3885),
.Y(n_4890)
);

OAI21x1_ASAP7_75t_SL g4891 ( 
.A1(n_4046),
.A2(n_3328),
.B(n_3327),
.Y(n_4891)
);

INVx2_ASAP7_75t_L g4892 ( 
.A(n_3937),
.Y(n_4892)
);

AOI22xp5_ASAP7_75t_L g4893 ( 
.A1(n_3833),
.A2(n_3018),
.B1(n_2842),
.B2(n_2847),
.Y(n_4893)
);

AO31x2_ASAP7_75t_L g4894 ( 
.A1(n_4271),
.A2(n_2830),
.A3(n_2827),
.B(n_2829),
.Y(n_4894)
);

OAI22xp5_ASAP7_75t_L g4895 ( 
.A1(n_3939),
.A2(n_2921),
.B1(n_2961),
.B2(n_2948),
.Y(n_4895)
);

OAI21x1_ASAP7_75t_L g4896 ( 
.A1(n_4031),
.A2(n_2829),
.B(n_2830),
.Y(n_4896)
);

OA22x2_ASAP7_75t_L g4897 ( 
.A1(n_4322),
.A2(n_3404),
.B1(n_3455),
.B2(n_3452),
.Y(n_4897)
);

INVx1_ASAP7_75t_L g4898 ( 
.A(n_3937),
.Y(n_4898)
);

O2A1O1Ixp5_ASAP7_75t_L g4899 ( 
.A1(n_4054),
.A2(n_3255),
.B(n_2889),
.C(n_2916),
.Y(n_4899)
);

A2O1A1Ixp33_ASAP7_75t_L g4900 ( 
.A1(n_4116),
.A2(n_2948),
.B(n_2961),
.C(n_2921),
.Y(n_4900)
);

NOR3xp33_ASAP7_75t_L g4901 ( 
.A(n_3550),
.B(n_3455),
.C(n_3402),
.Y(n_4901)
);

NAND2xp5_ASAP7_75t_SL g4902 ( 
.A(n_3851),
.B(n_3426),
.Y(n_4902)
);

OA22x2_ASAP7_75t_L g4903 ( 
.A1(n_3621),
.A2(n_4059),
.B1(n_4084),
.B2(n_3580),
.Y(n_4903)
);

AND2x2_ASAP7_75t_L g4904 ( 
.A(n_4274),
.B(n_2830),
.Y(n_4904)
);

AOI21xp5_ASAP7_75t_L g4905 ( 
.A1(n_4013),
.A2(n_3246),
.B(n_3255),
.Y(n_4905)
);

AND2x2_ASAP7_75t_L g4906 ( 
.A(n_4274),
.B(n_2830),
.Y(n_4906)
);

OAI21x1_ASAP7_75t_L g4907 ( 
.A1(n_4031),
.A2(n_4251),
.B(n_4242),
.Y(n_4907)
);

OAI21x1_ASAP7_75t_L g4908 ( 
.A1(n_4031),
.A2(n_2838),
.B(n_2832),
.Y(n_4908)
);

AOI21xp33_ASAP7_75t_L g4909 ( 
.A1(n_3851),
.A2(n_3395),
.B(n_3390),
.Y(n_4909)
);

AOI21x1_ASAP7_75t_L g4910 ( 
.A1(n_3534),
.A2(n_3329),
.B(n_3328),
.Y(n_4910)
);

NAND2xp5_ASAP7_75t_SL g4911 ( 
.A(n_3635),
.B(n_3426),
.Y(n_4911)
);

OAI21x1_ASAP7_75t_L g4912 ( 
.A1(n_4031),
.A2(n_2838),
.B(n_2832),
.Y(n_4912)
);

NAND2xp5_ASAP7_75t_L g4913 ( 
.A(n_3885),
.B(n_3362),
.Y(n_4913)
);

NAND2xp5_ASAP7_75t_L g4914 ( 
.A(n_3894),
.B(n_3362),
.Y(n_4914)
);

AOI21xp5_ASAP7_75t_L g4915 ( 
.A1(n_4013),
.A2(n_2948),
.B(n_2921),
.Y(n_4915)
);

A2O1A1Ixp33_ASAP7_75t_L g4916 ( 
.A1(n_3477),
.A2(n_2948),
.B(n_2961),
.C(n_2921),
.Y(n_4916)
);

OAI21xp5_ASAP7_75t_L g4917 ( 
.A1(n_3481),
.A2(n_3602),
.B(n_3504),
.Y(n_4917)
);

OAI21x1_ASAP7_75t_SL g4918 ( 
.A1(n_4046),
.A2(n_3331),
.B(n_3329),
.Y(n_4918)
);

INVx2_ASAP7_75t_SL g4919 ( 
.A(n_4248),
.Y(n_4919)
);

OAI21x1_ASAP7_75t_L g4920 ( 
.A1(n_4242),
.A2(n_2838),
.B(n_2832),
.Y(n_4920)
);

AOI21xp5_ASAP7_75t_L g4921 ( 
.A1(n_4024),
.A2(n_2961),
.B(n_2948),
.Y(n_4921)
);

NAND3xp33_ASAP7_75t_SL g4922 ( 
.A(n_3488),
.B(n_3331),
.C(n_3329),
.Y(n_4922)
);

OAI21x1_ASAP7_75t_L g4923 ( 
.A1(n_4242),
.A2(n_2843),
.B(n_2838),
.Y(n_4923)
);

OAI21xp33_ASAP7_75t_L g4924 ( 
.A1(n_3839),
.A2(n_3334),
.B(n_3331),
.Y(n_4924)
);

OAI21x1_ASAP7_75t_L g4925 ( 
.A1(n_4242),
.A2(n_4251),
.B(n_3547),
.Y(n_4925)
);

OAI21x1_ASAP7_75t_L g4926 ( 
.A1(n_4251),
.A2(n_2843),
.B(n_2838),
.Y(n_4926)
);

AOI21xp33_ASAP7_75t_L g4927 ( 
.A1(n_3602),
.A2(n_3834),
.B(n_3825),
.Y(n_4927)
);

NAND2xp5_ASAP7_75t_L g4928 ( 
.A(n_3894),
.B(n_3365),
.Y(n_4928)
);

A2O1A1Ixp33_ASAP7_75t_L g4929 ( 
.A1(n_3477),
.A2(n_2982),
.B(n_3044),
.C(n_2961),
.Y(n_4929)
);

INVx1_ASAP7_75t_L g4930 ( 
.A(n_3945),
.Y(n_4930)
);

OAI21x1_ASAP7_75t_L g4931 ( 
.A1(n_4251),
.A2(n_2846),
.B(n_2843),
.Y(n_4931)
);

OAI21xp33_ASAP7_75t_L g4932 ( 
.A1(n_3840),
.A2(n_3335),
.B(n_3334),
.Y(n_4932)
);

CKINVDCx5p33_ASAP7_75t_R g4933 ( 
.A(n_3617),
.Y(n_4933)
);

INVx1_ASAP7_75t_L g4934 ( 
.A(n_4036),
.Y(n_4934)
);

INVx1_ASAP7_75t_L g4935 ( 
.A(n_4036),
.Y(n_4935)
);

OAI21x1_ASAP7_75t_L g4936 ( 
.A1(n_4098),
.A2(n_2850),
.B(n_2846),
.Y(n_4936)
);

AOI21xp5_ASAP7_75t_L g4937 ( 
.A1(n_4024),
.A2(n_2982),
.B(n_2961),
.Y(n_4937)
);

OAI21x1_ASAP7_75t_L g4938 ( 
.A1(n_4098),
.A2(n_2852),
.B(n_2850),
.Y(n_4938)
);

NAND2xp5_ASAP7_75t_L g4939 ( 
.A(n_3896),
.B(n_3365),
.Y(n_4939)
);

AOI22xp5_ASAP7_75t_L g4940 ( 
.A1(n_3846),
.A2(n_2847),
.B1(n_2836),
.B2(n_2842),
.Y(n_4940)
);

NAND2xp5_ASAP7_75t_SL g4941 ( 
.A(n_3635),
.B(n_3426),
.Y(n_4941)
);

A2O1A1Ixp33_ASAP7_75t_L g4942 ( 
.A1(n_3621),
.A2(n_2982),
.B(n_3044),
.C(n_2961),
.Y(n_4942)
);

AOI22xp5_ASAP7_75t_L g4943 ( 
.A1(n_3490),
.A2(n_2836),
.B1(n_2862),
.B2(n_2847),
.Y(n_4943)
);

NAND2xp5_ASAP7_75t_L g4944 ( 
.A(n_3896),
.B(n_3365),
.Y(n_4944)
);

NOR2xp33_ASAP7_75t_L g4945 ( 
.A(n_3948),
.B(n_3426),
.Y(n_4945)
);

NAND2xp5_ASAP7_75t_L g4946 ( 
.A(n_3897),
.B(n_3368),
.Y(n_4946)
);

BUFx3_ASAP7_75t_L g4947 ( 
.A(n_4248),
.Y(n_4947)
);

INVx3_ASAP7_75t_L g4948 ( 
.A(n_4248),
.Y(n_4948)
);

OAI21xp5_ASAP7_75t_L g4949 ( 
.A1(n_3481),
.A2(n_3335),
.B(n_3334),
.Y(n_4949)
);

AOI21xp5_ASAP7_75t_L g4950 ( 
.A1(n_4198),
.A2(n_2982),
.B(n_2961),
.Y(n_4950)
);

NAND2xp5_ASAP7_75t_L g4951 ( 
.A(n_3897),
.B(n_3878),
.Y(n_4951)
);

CKINVDCx5p33_ASAP7_75t_R g4952 ( 
.A(n_3696),
.Y(n_4952)
);

NAND2xp5_ASAP7_75t_SL g4953 ( 
.A(n_3828),
.B(n_3426),
.Y(n_4953)
);

NAND2x1p5_ASAP7_75t_L g4954 ( 
.A(n_3744),
.B(n_2961),
.Y(n_4954)
);

NAND2xp5_ASAP7_75t_L g4955 ( 
.A(n_3886),
.B(n_3368),
.Y(n_4955)
);

NAND2xp5_ASAP7_75t_SL g4956 ( 
.A(n_3828),
.B(n_3426),
.Y(n_4956)
);

OA22x2_ASAP7_75t_L g4957 ( 
.A1(n_3580),
.A2(n_3404),
.B1(n_3395),
.B2(n_3390),
.Y(n_4957)
);

NAND2xp5_ASAP7_75t_L g4958 ( 
.A(n_3878),
.B(n_3368),
.Y(n_4958)
);

AOI21x1_ASAP7_75t_SL g4959 ( 
.A1(n_3629),
.A2(n_3273),
.B(n_3269),
.Y(n_4959)
);

NAND2xp5_ASAP7_75t_L g4960 ( 
.A(n_3889),
.B(n_4068),
.Y(n_4960)
);

BUFx2_ASAP7_75t_L g4961 ( 
.A(n_3985),
.Y(n_4961)
);

NOR2xp33_ASAP7_75t_L g4962 ( 
.A(n_3948),
.B(n_3426),
.Y(n_4962)
);

INVx2_ASAP7_75t_SL g4963 ( 
.A(n_4288),
.Y(n_4963)
);

OAI22xp5_ASAP7_75t_L g4964 ( 
.A1(n_3939),
.A2(n_2961),
.B1(n_3044),
.B2(n_2982),
.Y(n_4964)
);

OAI22xp5_ASAP7_75t_L g4965 ( 
.A1(n_3872),
.A2(n_2961),
.B1(n_3044),
.B2(n_2982),
.Y(n_4965)
);

OAI22x1_ASAP7_75t_L g4966 ( 
.A1(n_4080),
.A2(n_3495),
.B1(n_3554),
.B2(n_4113),
.Y(n_4966)
);

OAI21xp5_ASAP7_75t_L g4967 ( 
.A1(n_3504),
.A2(n_3342),
.B(n_3335),
.Y(n_4967)
);

OAI21xp5_ASAP7_75t_L g4968 ( 
.A1(n_3487),
.A2(n_3350),
.B(n_3342),
.Y(n_4968)
);

O2A1O1Ixp5_ASAP7_75t_L g4969 ( 
.A1(n_4001),
.A2(n_2889),
.B(n_2916),
.C(n_2908),
.Y(n_4969)
);

AOI21xp5_ASAP7_75t_L g4970 ( 
.A1(n_4293),
.A2(n_3044),
.B(n_2982),
.Y(n_4970)
);

INVx5_ASAP7_75t_L g4971 ( 
.A(n_4288),
.Y(n_4971)
);

AOI21xp5_ASAP7_75t_L g4972 ( 
.A1(n_3516),
.A2(n_3044),
.B(n_2982),
.Y(n_4972)
);

NAND2xp5_ASAP7_75t_L g4973 ( 
.A(n_3886),
.B(n_3373),
.Y(n_4973)
);

OAI21xp5_ASAP7_75t_L g4974 ( 
.A1(n_3487),
.A2(n_3350),
.B(n_3342),
.Y(n_4974)
);

AO31x2_ASAP7_75t_L g4975 ( 
.A1(n_4277),
.A2(n_2858),
.A3(n_2883),
.B(n_2863),
.Y(n_4975)
);

AO31x2_ASAP7_75t_L g4976 ( 
.A1(n_4277),
.A2(n_2858),
.A3(n_2883),
.B(n_2863),
.Y(n_4976)
);

BUFx4_ASAP7_75t_SL g4977 ( 
.A(n_4083),
.Y(n_4977)
);

AND2x2_ASAP7_75t_L g4978 ( 
.A(n_4331),
.B(n_3988),
.Y(n_4978)
);

NAND2xp5_ASAP7_75t_L g4979 ( 
.A(n_3889),
.B(n_3373),
.Y(n_4979)
);

NAND2xp5_ASAP7_75t_L g4980 ( 
.A(n_4020),
.B(n_3373),
.Y(n_4980)
);

AOI21x1_ASAP7_75t_L g4981 ( 
.A1(n_3534),
.A2(n_3351),
.B(n_3350),
.Y(n_4981)
);

INVx1_ASAP7_75t_SL g4982 ( 
.A(n_3754),
.Y(n_4982)
);

NAND2xp5_ASAP7_75t_L g4983 ( 
.A(n_4068),
.B(n_3377),
.Y(n_4983)
);

OAI21xp5_ASAP7_75t_L g4984 ( 
.A1(n_3484),
.A2(n_3361),
.B(n_3351),
.Y(n_4984)
);

INVx1_ASAP7_75t_L g4985 ( 
.A(n_4037),
.Y(n_4985)
);

NAND2xp5_ASAP7_75t_L g4986 ( 
.A(n_4020),
.B(n_3377),
.Y(n_4986)
);

AOI21xp5_ASAP7_75t_L g4987 ( 
.A1(n_3516),
.A2(n_3044),
.B(n_2982),
.Y(n_4987)
);

INVx1_ASAP7_75t_L g4988 ( 
.A(n_4090),
.Y(n_4988)
);

NAND2xp5_ASAP7_75t_L g4989 ( 
.A(n_4034),
.B(n_3377),
.Y(n_4989)
);

BUFx3_ASAP7_75t_L g4990 ( 
.A(n_4288),
.Y(n_4990)
);

INVx2_ASAP7_75t_SL g4991 ( 
.A(n_4288),
.Y(n_4991)
);

NAND2xp5_ASAP7_75t_L g4992 ( 
.A(n_4034),
.B(n_3379),
.Y(n_4992)
);

NAND3xp33_ASAP7_75t_SL g4993 ( 
.A(n_3488),
.B(n_3533),
.C(n_3515),
.Y(n_4993)
);

NAND2xp5_ASAP7_75t_L g4994 ( 
.A(n_3739),
.B(n_3379),
.Y(n_4994)
);

OA22x2_ASAP7_75t_L g4995 ( 
.A1(n_3659),
.A2(n_3404),
.B1(n_3395),
.B2(n_3390),
.Y(n_4995)
);

OAI21x1_ASAP7_75t_L g4996 ( 
.A1(n_4205),
.A2(n_2887),
.B(n_2883),
.Y(n_4996)
);

OAI21x1_ASAP7_75t_L g4997 ( 
.A1(n_4205),
.A2(n_2887),
.B(n_2883),
.Y(n_4997)
);

NAND2xp5_ASAP7_75t_L g4998 ( 
.A(n_3739),
.B(n_3379),
.Y(n_4998)
);

OAI21xp5_ASAP7_75t_L g4999 ( 
.A1(n_3484),
.A2(n_3376),
.B(n_3361),
.Y(n_4999)
);

AOI221xp5_ASAP7_75t_SL g5000 ( 
.A1(n_4261),
.A2(n_3410),
.B1(n_3413),
.B2(n_3393),
.C(n_3382),
.Y(n_5000)
);

OAI21xp5_ASAP7_75t_L g5001 ( 
.A1(n_3637),
.A2(n_3394),
.B(n_3376),
.Y(n_5001)
);

NAND2xp33_ASAP7_75t_L g5002 ( 
.A(n_3495),
.B(n_2980),
.Y(n_5002)
);

INVx1_ASAP7_75t_L g5003 ( 
.A(n_4140),
.Y(n_5003)
);

NAND2x1p5_ASAP7_75t_L g5004 ( 
.A(n_3744),
.B(n_2982),
.Y(n_5004)
);

OAI21xp5_ASAP7_75t_L g5005 ( 
.A1(n_3637),
.A2(n_3394),
.B(n_3376),
.Y(n_5005)
);

OAI21xp5_ASAP7_75t_L g5006 ( 
.A1(n_3645),
.A2(n_3405),
.B(n_3394),
.Y(n_5006)
);

INVx1_ASAP7_75t_L g5007 ( 
.A(n_4140),
.Y(n_5007)
);

INVx1_ASAP7_75t_L g5008 ( 
.A(n_4148),
.Y(n_5008)
);

AOI21xp5_ASAP7_75t_L g5009 ( 
.A1(n_3518),
.A2(n_3044),
.B(n_2982),
.Y(n_5009)
);

OAI21x1_ASAP7_75t_L g5010 ( 
.A1(n_3768),
.A2(n_2893),
.B(n_2887),
.Y(n_5010)
);

NAND2xp5_ASAP7_75t_SL g5011 ( 
.A(n_3499),
.B(n_3426),
.Y(n_5011)
);

NOR2xp33_ASAP7_75t_L g5012 ( 
.A(n_3642),
.B(n_3649),
.Y(n_5012)
);

NAND2xp5_ASAP7_75t_L g5013 ( 
.A(n_3787),
.B(n_3382),
.Y(n_5013)
);

OAI21xp5_ASAP7_75t_L g5014 ( 
.A1(n_3645),
.A2(n_3414),
.B(n_3405),
.Y(n_5014)
);

AND2x4_ASAP7_75t_L g5015 ( 
.A(n_3479),
.B(n_3579),
.Y(n_5015)
);

AOI221xp5_ASAP7_75t_L g5016 ( 
.A1(n_3865),
.A2(n_3382),
.B1(n_3413),
.B2(n_3410),
.C(n_3393),
.Y(n_5016)
);

A2O1A1Ixp33_ASAP7_75t_L g5017 ( 
.A1(n_3650),
.A2(n_3080),
.B(n_3092),
.C(n_3044),
.Y(n_5017)
);

INVx1_ASAP7_75t_L g5018 ( 
.A(n_4165),
.Y(n_5018)
);

A2O1A1Ixp33_ASAP7_75t_L g5019 ( 
.A1(n_3650),
.A2(n_3080),
.B(n_3092),
.C(n_3044),
.Y(n_5019)
);

OAI22xp5_ASAP7_75t_L g5020 ( 
.A1(n_3882),
.A2(n_3044),
.B1(n_3092),
.B2(n_3080),
.Y(n_5020)
);

NAND2xp5_ASAP7_75t_L g5021 ( 
.A(n_3787),
.B(n_3393),
.Y(n_5021)
);

NOR2xp33_ASAP7_75t_L g5022 ( 
.A(n_3655),
.B(n_3426),
.Y(n_5022)
);

AND2x2_ASAP7_75t_L g5023 ( 
.A(n_4331),
.B(n_3988),
.Y(n_5023)
);

NAND2xp5_ASAP7_75t_L g5024 ( 
.A(n_3798),
.B(n_3410),
.Y(n_5024)
);

BUFx3_ASAP7_75t_L g5025 ( 
.A(n_4288),
.Y(n_5025)
);

OAI21x1_ASAP7_75t_L g5026 ( 
.A1(n_3793),
.A2(n_2920),
.B(n_2900),
.Y(n_5026)
);

OAI21xp5_ASAP7_75t_L g5027 ( 
.A1(n_3706),
.A2(n_3414),
.B(n_3405),
.Y(n_5027)
);

OAI21x1_ASAP7_75t_L g5028 ( 
.A1(n_3793),
.A2(n_3556),
.B(n_3604),
.Y(n_5028)
);

AOI21xp5_ASAP7_75t_L g5029 ( 
.A1(n_3518),
.A2(n_3092),
.B(n_3080),
.Y(n_5029)
);

NAND2xp5_ASAP7_75t_L g5030 ( 
.A(n_3798),
.B(n_3832),
.Y(n_5030)
);

INVx1_ASAP7_75t_L g5031 ( 
.A(n_4165),
.Y(n_5031)
);

NAND2xp5_ASAP7_75t_L g5032 ( 
.A(n_3832),
.B(n_3413),
.Y(n_5032)
);

OAI21xp5_ASAP7_75t_L g5033 ( 
.A1(n_3706),
.A2(n_3429),
.B(n_3414),
.Y(n_5033)
);

AOI22xp5_ASAP7_75t_L g5034 ( 
.A1(n_3506),
.A2(n_2836),
.B1(n_2862),
.B2(n_2847),
.Y(n_5034)
);

NOR2xp33_ASAP7_75t_L g5035 ( 
.A(n_3537),
.B(n_3426),
.Y(n_5035)
);

AOI21xp5_ASAP7_75t_L g5036 ( 
.A1(n_3856),
.A2(n_3092),
.B(n_3080),
.Y(n_5036)
);

AO21x1_ASAP7_75t_L g5037 ( 
.A1(n_4261),
.A2(n_3431),
.B(n_3418),
.Y(n_5037)
);

AOI211x1_ASAP7_75t_L g5038 ( 
.A1(n_4038),
.A2(n_3429),
.B(n_3439),
.C(n_3438),
.Y(n_5038)
);

NOR2xp67_ASAP7_75t_L g5039 ( 
.A(n_3993),
.B(n_3080),
.Y(n_5039)
);

NOR2xp67_ASAP7_75t_SL g5040 ( 
.A(n_4314),
.B(n_3080),
.Y(n_5040)
);

INVx3_ASAP7_75t_L g5041 ( 
.A(n_4288),
.Y(n_5041)
);

CKINVDCx5p33_ASAP7_75t_R g5042 ( 
.A(n_3513),
.Y(n_5042)
);

NAND2xp5_ASAP7_75t_L g5043 ( 
.A(n_4045),
.B(n_3418),
.Y(n_5043)
);

BUFx8_ASAP7_75t_L g5044 ( 
.A(n_4342),
.Y(n_5044)
);

CKINVDCx5p33_ASAP7_75t_R g5045 ( 
.A(n_3513),
.Y(n_5045)
);

AOI22xp5_ASAP7_75t_L g5046 ( 
.A1(n_3562),
.A2(n_2836),
.B1(n_2862),
.B2(n_2847),
.Y(n_5046)
);

A2O1A1Ixp33_ASAP7_75t_L g5047 ( 
.A1(n_4164),
.A2(n_3092),
.B(n_3080),
.C(n_3345),
.Y(n_5047)
);

NAND2x1p5_ASAP7_75t_L g5048 ( 
.A(n_3744),
.B(n_3080),
.Y(n_5048)
);

OAI21xp5_ASAP7_75t_L g5049 ( 
.A1(n_3604),
.A2(n_3480),
.B(n_3568),
.Y(n_5049)
);

AOI21xp5_ASAP7_75t_L g5050 ( 
.A1(n_3856),
.A2(n_3092),
.B(n_3080),
.Y(n_5050)
);

OAI21x1_ASAP7_75t_L g5051 ( 
.A1(n_3898),
.A2(n_2926),
.B(n_2920),
.Y(n_5051)
);

OAI21x1_ASAP7_75t_L g5052 ( 
.A1(n_3898),
.A2(n_2926),
.B(n_2920),
.Y(n_5052)
);

INVx1_ASAP7_75t_L g5053 ( 
.A(n_4182),
.Y(n_5053)
);

OAI21x1_ASAP7_75t_L g5054 ( 
.A1(n_3898),
.A2(n_2930),
.B(n_2926),
.Y(n_5054)
);

NAND2xp5_ASAP7_75t_L g5055 ( 
.A(n_4045),
.B(n_3418),
.Y(n_5055)
);

OAI21x1_ASAP7_75t_L g5056 ( 
.A1(n_3898),
.A2(n_2930),
.B(n_2926),
.Y(n_5056)
);

NAND2xp5_ASAP7_75t_L g5057 ( 
.A(n_3543),
.B(n_3431),
.Y(n_5057)
);

INVxp67_ASAP7_75t_L g5058 ( 
.A(n_4199),
.Y(n_5058)
);

INVx5_ASAP7_75t_L g5059 ( 
.A(n_4298),
.Y(n_5059)
);

INVx2_ASAP7_75t_SL g5060 ( 
.A(n_4298),
.Y(n_5060)
);

OAI21xp5_ASAP7_75t_L g5061 ( 
.A1(n_3568),
.A2(n_3663),
.B(n_3658),
.Y(n_5061)
);

OAI21xp5_ASAP7_75t_L g5062 ( 
.A1(n_3658),
.A2(n_3438),
.B(n_3429),
.Y(n_5062)
);

NAND2xp5_ASAP7_75t_L g5063 ( 
.A(n_3763),
.B(n_3432),
.Y(n_5063)
);

AOI21x1_ASAP7_75t_SL g5064 ( 
.A1(n_3629),
.A2(n_3273),
.B(n_3269),
.Y(n_5064)
);

A2O1A1Ixp33_ASAP7_75t_L g5065 ( 
.A1(n_4164),
.A2(n_3092),
.B(n_3080),
.C(n_3345),
.Y(n_5065)
);

OAI21xp5_ASAP7_75t_L g5066 ( 
.A1(n_3663),
.A2(n_3710),
.B(n_3825),
.Y(n_5066)
);

NAND2x1p5_ASAP7_75t_L g5067 ( 
.A(n_3744),
.B(n_3944),
.Y(n_5067)
);

O2A1O1Ixp5_ASAP7_75t_L g5068 ( 
.A1(n_4039),
.A2(n_2908),
.B(n_2916),
.C(n_2889),
.Y(n_5068)
);

AOI21xp5_ASAP7_75t_L g5069 ( 
.A1(n_4213),
.A2(n_3092),
.B(n_3345),
.Y(n_5069)
);

BUFx3_ASAP7_75t_L g5070 ( 
.A(n_4298),
.Y(n_5070)
);

NAND2xp5_ASAP7_75t_L g5071 ( 
.A(n_4132),
.B(n_4313),
.Y(n_5071)
);

NAND2xp5_ASAP7_75t_L g5072 ( 
.A(n_4313),
.B(n_3432),
.Y(n_5072)
);

CKINVDCx5p33_ASAP7_75t_R g5073 ( 
.A(n_3513),
.Y(n_5073)
);

NAND2xp5_ASAP7_75t_L g5074 ( 
.A(n_3804),
.B(n_3437),
.Y(n_5074)
);

NAND2xp5_ASAP7_75t_L g5075 ( 
.A(n_3804),
.B(n_3965),
.Y(n_5075)
);

INVxp67_ASAP7_75t_L g5076 ( 
.A(n_3781),
.Y(n_5076)
);

NOR2x1_ASAP7_75t_SL g5077 ( 
.A(n_3931),
.B(n_3092),
.Y(n_5077)
);

OAI21x1_ASAP7_75t_L g5078 ( 
.A1(n_3709),
.A2(n_3967),
.B(n_4047),
.Y(n_5078)
);

BUFx3_ASAP7_75t_L g5079 ( 
.A(n_4298),
.Y(n_5079)
);

BUFx12f_ASAP7_75t_L g5080 ( 
.A(n_4027),
.Y(n_5080)
);

CKINVDCx11_ASAP7_75t_R g5081 ( 
.A(n_4135),
.Y(n_5081)
);

OAI21x1_ASAP7_75t_L g5082 ( 
.A1(n_3967),
.A2(n_4052),
.B(n_4047),
.Y(n_5082)
);

NAND2xp5_ASAP7_75t_L g5083 ( 
.A(n_3965),
.B(n_3437),
.Y(n_5083)
);

NAND2xp5_ASAP7_75t_L g5084 ( 
.A(n_4003),
.B(n_4315),
.Y(n_5084)
);

NAND2xp5_ASAP7_75t_L g5085 ( 
.A(n_4003),
.B(n_3437),
.Y(n_5085)
);

INVxp67_ASAP7_75t_L g5086 ( 
.A(n_3475),
.Y(n_5086)
);

AOI21x1_ASAP7_75t_L g5087 ( 
.A1(n_4119),
.A2(n_4120),
.B(n_3997),
.Y(n_5087)
);

OAI22xp5_ASAP7_75t_L g5088 ( 
.A1(n_3972),
.A2(n_3165),
.B1(n_2876),
.B2(n_3005),
.Y(n_5088)
);

AND2x4_ASAP7_75t_L g5089 ( 
.A(n_3479),
.B(n_3112),
.Y(n_5089)
);

AND2x4_ASAP7_75t_L g5090 ( 
.A(n_3579),
.B(n_3112),
.Y(n_5090)
);

BUFx5_ASAP7_75t_L g5091 ( 
.A(n_3598),
.Y(n_5091)
);

INVxp67_ASAP7_75t_SL g5092 ( 
.A(n_4214),
.Y(n_5092)
);

OAI21x1_ASAP7_75t_L g5093 ( 
.A1(n_4052),
.A2(n_2958),
.B(n_2949),
.Y(n_5093)
);

BUFx3_ASAP7_75t_L g5094 ( 
.A(n_4298),
.Y(n_5094)
);

NAND2x1p5_ASAP7_75t_L g5095 ( 
.A(n_3944),
.B(n_3112),
.Y(n_5095)
);

AOI21x1_ASAP7_75t_L g5096 ( 
.A1(n_3983),
.A2(n_3439),
.B(n_3438),
.Y(n_5096)
);

AOI21xp5_ASAP7_75t_L g5097 ( 
.A1(n_4219),
.A2(n_3375),
.B(n_3345),
.Y(n_5097)
);

AOI21xp5_ASAP7_75t_L g5098 ( 
.A1(n_4223),
.A2(n_3375),
.B(n_3345),
.Y(n_5098)
);

AND2x6_ASAP7_75t_L g5099 ( 
.A(n_3497),
.B(n_3375),
.Y(n_5099)
);

OAI21x1_ASAP7_75t_L g5100 ( 
.A1(n_4075),
.A2(n_2967),
.B(n_2958),
.Y(n_5100)
);

AOI21xp5_ASAP7_75t_L g5101 ( 
.A1(n_4232),
.A2(n_3380),
.B(n_3375),
.Y(n_5101)
);

OAI21x1_ASAP7_75t_SL g5102 ( 
.A1(n_4079),
.A2(n_3439),
.B(n_2915),
.Y(n_5102)
);

AOI21xp5_ASAP7_75t_L g5103 ( 
.A1(n_4237),
.A2(n_3380),
.B(n_3375),
.Y(n_5103)
);

NAND2x1p5_ASAP7_75t_L g5104 ( 
.A(n_3944),
.B(n_3129),
.Y(n_5104)
);

AOI21xp5_ASAP7_75t_L g5105 ( 
.A1(n_4252),
.A2(n_3380),
.B(n_3167),
.Y(n_5105)
);

INVx1_ASAP7_75t_SL g5106 ( 
.A(n_3754),
.Y(n_5106)
);

INVx1_ASAP7_75t_SL g5107 ( 
.A(n_4306),
.Y(n_5107)
);

AOI22xp33_ASAP7_75t_L g5108 ( 
.A1(n_4146),
.A2(n_2980),
.B1(n_2836),
.B2(n_2862),
.Y(n_5108)
);

AOI21xp5_ASAP7_75t_L g5109 ( 
.A1(n_4276),
.A2(n_3380),
.B(n_3167),
.Y(n_5109)
);

CKINVDCx9p33_ASAP7_75t_R g5110 ( 
.A(n_3960),
.Y(n_5110)
);

OAI22xp5_ASAP7_75t_L g5111 ( 
.A1(n_3974),
.A2(n_3165),
.B1(n_2876),
.B2(n_3005),
.Y(n_5111)
);

OAI21x1_ASAP7_75t_L g5112 ( 
.A1(n_4091),
.A2(n_3710),
.B(n_4104),
.Y(n_5112)
);

NAND3xp33_ASAP7_75t_L g5113 ( 
.A(n_3597),
.B(n_3440),
.C(n_3330),
.Y(n_5113)
);

OAI21x1_ASAP7_75t_L g5114 ( 
.A1(n_4114),
.A2(n_4012),
.B(n_3993),
.Y(n_5114)
);

OAI21x1_ASAP7_75t_L g5115 ( 
.A1(n_4114),
.A2(n_3006),
.B(n_3004),
.Y(n_5115)
);

BUFx3_ASAP7_75t_L g5116 ( 
.A(n_4298),
.Y(n_5116)
);

OAI21xp5_ASAP7_75t_L g5117 ( 
.A1(n_3834),
.A2(n_3536),
.B(n_3549),
.Y(n_5117)
);

INVx4_ASAP7_75t_L g5118 ( 
.A(n_4094),
.Y(n_5118)
);

NAND2xp5_ASAP7_75t_L g5119 ( 
.A(n_4038),
.B(n_3006),
.Y(n_5119)
);

INVxp67_ASAP7_75t_SL g5120 ( 
.A(n_4214),
.Y(n_5120)
);

AOI21xp5_ASAP7_75t_L g5121 ( 
.A1(n_4291),
.A2(n_3380),
.B(n_3167),
.Y(n_5121)
);

OAI22xp5_ASAP7_75t_L g5122 ( 
.A1(n_3572),
.A2(n_3165),
.B1(n_2876),
.B2(n_3005),
.Y(n_5122)
);

OAI21xp5_ASAP7_75t_L g5123 ( 
.A1(n_3536),
.A2(n_3363),
.B(n_3357),
.Y(n_5123)
);

A2O1A1Ixp33_ASAP7_75t_L g5124 ( 
.A1(n_4244),
.A2(n_3005),
.B(n_3017),
.C(n_2992),
.Y(n_5124)
);

BUFx3_ASAP7_75t_L g5125 ( 
.A(n_4316),
.Y(n_5125)
);

NOR2xp33_ASAP7_75t_L g5126 ( 
.A(n_3574),
.B(n_3433),
.Y(n_5126)
);

INVx6_ASAP7_75t_L g5127 ( 
.A(n_3844),
.Y(n_5127)
);

AO31x2_ASAP7_75t_L g5128 ( 
.A1(n_4123),
.A2(n_4101),
.A3(n_4247),
.B(n_4299),
.Y(n_5128)
);

INVx2_ASAP7_75t_SL g5129 ( 
.A(n_4316),
.Y(n_5129)
);

NAND2xp5_ASAP7_75t_SL g5130 ( 
.A(n_3499),
.B(n_3433),
.Y(n_5130)
);

AOI22xp5_ASAP7_75t_L g5131 ( 
.A1(n_3976),
.A2(n_3550),
.B1(n_3546),
.B2(n_3542),
.Y(n_5131)
);

OAI21x1_ASAP7_75t_L g5132 ( 
.A1(n_4012),
.A2(n_3022),
.B(n_3020),
.Y(n_5132)
);

AOI21xp5_ASAP7_75t_L g5133 ( 
.A1(n_4308),
.A2(n_3167),
.B(n_3390),
.Y(n_5133)
);

BUFx2_ASAP7_75t_L g5134 ( 
.A(n_3985),
.Y(n_5134)
);

NOR2x1_ASAP7_75t_SL g5135 ( 
.A(n_3626),
.B(n_3390),
.Y(n_5135)
);

OA21x2_ASAP7_75t_L g5136 ( 
.A1(n_3905),
.A2(n_3046),
.B(n_3024),
.Y(n_5136)
);

OAI21x1_ASAP7_75t_SL g5137 ( 
.A1(n_3860),
.A2(n_2915),
.B(n_2859),
.Y(n_5137)
);

OAI21xp5_ASAP7_75t_L g5138 ( 
.A1(n_3549),
.A2(n_3363),
.B(n_3357),
.Y(n_5138)
);

NOR2xp33_ASAP7_75t_L g5139 ( 
.A(n_3640),
.B(n_3433),
.Y(n_5139)
);

AOI21xp5_ASAP7_75t_L g5140 ( 
.A1(n_4317),
.A2(n_3167),
.B(n_3390),
.Y(n_5140)
);

OA21x2_ASAP7_75t_L g5141 ( 
.A1(n_3905),
.A2(n_3057),
.B(n_3046),
.Y(n_5141)
);

BUFx6f_ASAP7_75t_L g5142 ( 
.A(n_4316),
.Y(n_5142)
);

INVx5_ASAP7_75t_L g5143 ( 
.A(n_4316),
.Y(n_5143)
);

NAND3xp33_ASAP7_75t_SL g5144 ( 
.A(n_5131),
.B(n_3659),
.C(n_3528),
.Y(n_5144)
);

AOI21xp5_ASAP7_75t_L g5145 ( 
.A1(n_4732),
.A2(n_3802),
.B(n_4290),
.Y(n_5145)
);

OAI22xp5_ASAP7_75t_L g5146 ( 
.A1(n_4376),
.A2(n_4554),
.B1(n_4548),
.B2(n_5131),
.Y(n_5146)
);

NOR2x1_ASAP7_75t_R g5147 ( 
.A(n_4381),
.B(n_4342),
.Y(n_5147)
);

OA21x2_ASAP7_75t_L g5148 ( 
.A1(n_4372),
.A2(n_4266),
.B(n_3966),
.Y(n_5148)
);

HB1xp67_ASAP7_75t_L g5149 ( 
.A(n_4695),
.Y(n_5149)
);

OAI21x1_ASAP7_75t_L g5150 ( 
.A1(n_4721),
.A2(n_4113),
.B(n_3760),
.Y(n_5150)
);

AOI21xp5_ASAP7_75t_L g5151 ( 
.A1(n_4816),
.A2(n_3802),
.B(n_4321),
.Y(n_5151)
);

AOI21x1_ASAP7_75t_L g5152 ( 
.A1(n_4721),
.A2(n_4549),
.B(n_4501),
.Y(n_5152)
);

OAI21x1_ASAP7_75t_L g5153 ( 
.A1(n_4721),
.A2(n_3760),
.B(n_3731),
.Y(n_5153)
);

OAI21xp5_ASAP7_75t_SL g5154 ( 
.A1(n_4554),
.A2(n_3958),
.B(n_3809),
.Y(n_5154)
);

O2A1O1Ixp33_ASAP7_75t_L g5155 ( 
.A1(n_4993),
.A2(n_3925),
.B(n_3819),
.C(n_3932),
.Y(n_5155)
);

OAI21xp5_ASAP7_75t_L g5156 ( 
.A1(n_4917),
.A2(n_3712),
.B(n_3634),
.Y(n_5156)
);

OAI22xp5_ASAP7_75t_L g5157 ( 
.A1(n_4376),
.A2(n_3913),
.B1(n_3831),
.B2(n_3572),
.Y(n_5157)
);

AOI21xp5_ASAP7_75t_L g5158 ( 
.A1(n_4816),
.A2(n_3610),
.B(n_4244),
.Y(n_5158)
);

CKINVDCx5p33_ASAP7_75t_R g5159 ( 
.A(n_4451),
.Y(n_5159)
);

NOR4xp25_ASAP7_75t_L g5160 ( 
.A(n_4993),
.B(n_4917),
.C(n_5117),
.D(n_4927),
.Y(n_5160)
);

NAND2xp5_ASAP7_75t_L g5161 ( 
.A(n_4681),
.B(n_4225),
.Y(n_5161)
);

AOI21xp5_ASAP7_75t_L g5162 ( 
.A1(n_5061),
.A2(n_3820),
.B(n_4142),
.Y(n_5162)
);

O2A1O1Ixp5_ASAP7_75t_L g5163 ( 
.A1(n_5117),
.A2(n_3625),
.B(n_3668),
.C(n_4121),
.Y(n_5163)
);

AOI21x1_ASAP7_75t_L g5164 ( 
.A1(n_4549),
.A2(n_3502),
.B(n_4368),
.Y(n_5164)
);

AOI21xp5_ASAP7_75t_L g5165 ( 
.A1(n_5061),
.A2(n_5065),
.B(n_5047),
.Y(n_5165)
);

A2O1A1Ixp33_ASAP7_75t_L g5166 ( 
.A1(n_4536),
.A2(n_4146),
.B(n_3977),
.C(n_3982),
.Y(n_5166)
);

INVx2_ASAP7_75t_L g5167 ( 
.A(n_4384),
.Y(n_5167)
);

OAI21x1_ASAP7_75t_L g5168 ( 
.A1(n_4950),
.A2(n_3760),
.B(n_3731),
.Y(n_5168)
);

INVx3_ASAP7_75t_SL g5169 ( 
.A(n_4952),
.Y(n_5169)
);

A2O1A1Ixp33_ASAP7_75t_L g5170 ( 
.A1(n_4536),
.A2(n_3977),
.B(n_3982),
.C(n_4161),
.Y(n_5170)
);

NAND2x1p5_ASAP7_75t_L g5171 ( 
.A(n_4840),
.B(n_4848),
.Y(n_5171)
);

AOI21xp5_ASAP7_75t_L g5172 ( 
.A1(n_5047),
.A2(n_3820),
.B(n_3973),
.Y(n_5172)
);

OAI21xp33_ASAP7_75t_L g5173 ( 
.A1(n_4548),
.A2(n_3785),
.B(n_4023),
.Y(n_5173)
);

NAND2xp5_ASAP7_75t_L g5174 ( 
.A(n_4681),
.B(n_4225),
.Y(n_5174)
);

NAND2xp5_ASAP7_75t_L g5175 ( 
.A(n_4690),
.B(n_4234),
.Y(n_5175)
);

INVx1_ASAP7_75t_L g5176 ( 
.A(n_4412),
.Y(n_5176)
);

AOI221xp5_ASAP7_75t_L g5177 ( 
.A1(n_4606),
.A2(n_4023),
.B1(n_4004),
.B2(n_4101),
.C(n_3955),
.Y(n_5177)
);

AOI21xp5_ASAP7_75t_SL g5178 ( 
.A1(n_4814),
.A2(n_3943),
.B(n_3936),
.Y(n_5178)
);

NAND2x1p5_ASAP7_75t_L g5179 ( 
.A(n_4840),
.B(n_4257),
.Y(n_5179)
);

CKINVDCx11_ASAP7_75t_R g5180 ( 
.A(n_4806),
.Y(n_5180)
);

AND2x2_ASAP7_75t_L g5181 ( 
.A(n_4978),
.B(n_4305),
.Y(n_5181)
);

OR2x2_ASAP7_75t_L g5182 ( 
.A(n_4567),
.B(n_3519),
.Y(n_5182)
);

AOI21xp5_ASAP7_75t_L g5183 ( 
.A1(n_5065),
.A2(n_3981),
.B(n_3973),
.Y(n_5183)
);

CKINVDCx5p33_ASAP7_75t_R g5184 ( 
.A(n_4381),
.Y(n_5184)
);

INVx2_ASAP7_75t_L g5185 ( 
.A(n_4384),
.Y(n_5185)
);

OAI22x1_ASAP7_75t_L g5186 ( 
.A1(n_4667),
.A2(n_4080),
.B1(n_4330),
.B2(n_3554),
.Y(n_5186)
);

CKINVDCx16_ASAP7_75t_R g5187 ( 
.A(n_4381),
.Y(n_5187)
);

NAND3xp33_ASAP7_75t_L g5188 ( 
.A(n_4606),
.B(n_3573),
.C(n_3565),
.Y(n_5188)
);

INVx3_ASAP7_75t_L g5189 ( 
.A(n_5142),
.Y(n_5189)
);

OAI22xp33_ASAP7_75t_L g5190 ( 
.A1(n_4903),
.A2(n_3949),
.B1(n_3981),
.B2(n_3541),
.Y(n_5190)
);

AND2x4_ASAP7_75t_L g5191 ( 
.A(n_5015),
.B(n_3579),
.Y(n_5191)
);

OAI21xp5_ASAP7_75t_L g5192 ( 
.A1(n_5049),
.A2(n_3713),
.B(n_3590),
.Y(n_5192)
);

INVx2_ASAP7_75t_SL g5193 ( 
.A(n_5127),
.Y(n_5193)
);

NAND2x1p5_ASAP7_75t_L g5194 ( 
.A(n_4848),
.B(n_4257),
.Y(n_5194)
);

O2A1O1Ixp5_ASAP7_75t_L g5195 ( 
.A1(n_4693),
.A2(n_4354),
.B(n_4230),
.C(n_4243),
.Y(n_5195)
);

OAI221xp5_ASAP7_75t_L g5196 ( 
.A1(n_5049),
.A2(n_3541),
.B1(n_3949),
.B2(n_3677),
.C(n_4016),
.Y(n_5196)
);

INVx1_ASAP7_75t_L g5197 ( 
.A(n_4412),
.Y(n_5197)
);

A2O1A1Ixp33_ASAP7_75t_L g5198 ( 
.A1(n_4814),
.A2(n_4254),
.B(n_4109),
.C(n_3961),
.Y(n_5198)
);

INVx3_ASAP7_75t_SL g5199 ( 
.A(n_5042),
.Y(n_5199)
);

OR2x6_ASAP7_75t_L g5200 ( 
.A(n_4592),
.B(n_3956),
.Y(n_5200)
);

AOI22xp5_ASAP7_75t_L g5201 ( 
.A1(n_4378),
.A2(n_3955),
.B1(n_4112),
.B2(n_3546),
.Y(n_5201)
);

AOI22xp5_ASAP7_75t_L g5202 ( 
.A1(n_4378),
.A2(n_4112),
.B1(n_3583),
.B2(n_4019),
.Y(n_5202)
);

AOI21xp5_ASAP7_75t_L g5203 ( 
.A1(n_4693),
.A2(n_4370),
.B(n_4367),
.Y(n_5203)
);

OAI21x1_ASAP7_75t_L g5204 ( 
.A1(n_4950),
.A2(n_3760),
.B(n_3731),
.Y(n_5204)
);

AOI21xp5_ASAP7_75t_L g5205 ( 
.A1(n_4708),
.A2(n_4900),
.B(n_4942),
.Y(n_5205)
);

INVx1_ASAP7_75t_L g5206 ( 
.A(n_4417),
.Y(n_5206)
);

INVxp67_ASAP7_75t_L g5207 ( 
.A(n_5030),
.Y(n_5207)
);

NAND2xp5_ASAP7_75t_L g5208 ( 
.A(n_4690),
.B(n_4951),
.Y(n_5208)
);

INVx4_ASAP7_75t_L g5209 ( 
.A(n_4425),
.Y(n_5209)
);

AOI21xp5_ASAP7_75t_L g5210 ( 
.A1(n_4708),
.A2(n_4370),
.B(n_4367),
.Y(n_5210)
);

INVx2_ASAP7_75t_L g5211 ( 
.A(n_4384),
.Y(n_5211)
);

BUFx8_ASAP7_75t_L g5212 ( 
.A(n_4534),
.Y(n_5212)
);

NAND2xp5_ASAP7_75t_L g5213 ( 
.A(n_4951),
.B(n_4234),
.Y(n_5213)
);

OAI21xp5_ASAP7_75t_L g5214 ( 
.A1(n_4927),
.A2(n_4903),
.B(n_4755),
.Y(n_5214)
);

OA21x2_ASAP7_75t_L g5215 ( 
.A1(n_4372),
.A2(n_4105),
.B(n_4178),
.Y(n_5215)
);

OAI22xp5_ASAP7_75t_L g5216 ( 
.A1(n_4755),
.A2(n_3831),
.B1(n_3913),
.B2(n_3572),
.Y(n_5216)
);

A2O1A1Ixp33_ASAP7_75t_L g5217 ( 
.A1(n_4654),
.A2(n_4254),
.B(n_3502),
.C(n_3901),
.Y(n_5217)
);

OAI21xp5_ASAP7_75t_L g5218 ( 
.A1(n_4903),
.A2(n_4922),
.B(n_4960),
.Y(n_5218)
);

INVxp67_ASAP7_75t_SL g5219 ( 
.A(n_4665),
.Y(n_5219)
);

AOI21xp5_ASAP7_75t_L g5220 ( 
.A1(n_4753),
.A2(n_4290),
.B(n_4249),
.Y(n_5220)
);

AND3x2_ASAP7_75t_L g5221 ( 
.A(n_4801),
.B(n_3582),
.C(n_3551),
.Y(n_5221)
);

INVx4_ASAP7_75t_L g5222 ( 
.A(n_4425),
.Y(n_5222)
);

INVx2_ASAP7_75t_SL g5223 ( 
.A(n_5127),
.Y(n_5223)
);

OAI21x1_ASAP7_75t_L g5224 ( 
.A1(n_4585),
.A2(n_3731),
.B(n_3675),
.Y(n_5224)
);

NAND2xp5_ASAP7_75t_L g5225 ( 
.A(n_4736),
.B(n_4272),
.Y(n_5225)
);

INVx2_ASAP7_75t_L g5226 ( 
.A(n_4532),
.Y(n_5226)
);

OAI21x1_ASAP7_75t_L g5227 ( 
.A1(n_4585),
.A2(n_3675),
.B(n_3672),
.Y(n_5227)
);

AND2x6_ASAP7_75t_L g5228 ( 
.A(n_4464),
.B(n_3497),
.Y(n_5228)
);

INVx1_ASAP7_75t_L g5229 ( 
.A(n_4417),
.Y(n_5229)
);

INVx1_ASAP7_75t_L g5230 ( 
.A(n_4428),
.Y(n_5230)
);

O2A1O1Ixp33_ASAP7_75t_SL g5231 ( 
.A1(n_4806),
.A2(n_3987),
.B(n_3958),
.C(n_3971),
.Y(n_5231)
);

AOI22xp5_ASAP7_75t_L g5232 ( 
.A1(n_4903),
.A2(n_3583),
.B1(n_3949),
.B2(n_4107),
.Y(n_5232)
);

OAI21x1_ASAP7_75t_L g5233 ( 
.A1(n_4585),
.A2(n_3682),
.B(n_3678),
.Y(n_5233)
);

AOI21xp5_ASAP7_75t_L g5234 ( 
.A1(n_4753),
.A2(n_4290),
.B(n_4010),
.Y(n_5234)
);

HB1xp67_ASAP7_75t_L g5235 ( 
.A(n_4695),
.Y(n_5235)
);

BUFx2_ASAP7_75t_L g5236 ( 
.A(n_4711),
.Y(n_5236)
);

CKINVDCx5p33_ASAP7_75t_R g5237 ( 
.A(n_4473),
.Y(n_5237)
);

O2A1O1Ixp33_ASAP7_75t_L g5238 ( 
.A1(n_4960),
.A2(n_3573),
.B(n_3565),
.C(n_3643),
.Y(n_5238)
);

NOR2xp33_ASAP7_75t_L g5239 ( 
.A(n_4879),
.B(n_3987),
.Y(n_5239)
);

NAND2xp5_ASAP7_75t_L g5240 ( 
.A(n_4736),
.B(n_4754),
.Y(n_5240)
);

NOR2xp33_ASAP7_75t_L g5241 ( 
.A(n_4933),
.B(n_3511),
.Y(n_5241)
);

INVx3_ASAP7_75t_L g5242 ( 
.A(n_4388),
.Y(n_5242)
);

OAI21x1_ASAP7_75t_L g5243 ( 
.A1(n_4372),
.A2(n_3682),
.B(n_3678),
.Y(n_5243)
);

INVx1_ASAP7_75t_L g5244 ( 
.A(n_4428),
.Y(n_5244)
);

AOI21xp5_ASAP7_75t_L g5245 ( 
.A1(n_4972),
.A2(n_4290),
.B(n_4227),
.Y(n_5245)
);

AND2x2_ASAP7_75t_L g5246 ( 
.A(n_4978),
.B(n_4359),
.Y(n_5246)
);

AOI22xp5_ASAP7_75t_L g5247 ( 
.A1(n_4712),
.A2(n_3584),
.B1(n_3542),
.B2(n_3589),
.Y(n_5247)
);

O2A1O1Ixp5_ASAP7_75t_SL g5248 ( 
.A1(n_4902),
.A2(n_3890),
.B(n_3520),
.C(n_3938),
.Y(n_5248)
);

AOI21xp5_ASAP7_75t_L g5249 ( 
.A1(n_4972),
.A2(n_4290),
.B(n_3699),
.Y(n_5249)
);

NAND2xp5_ASAP7_75t_L g5250 ( 
.A(n_4754),
.B(n_4272),
.Y(n_5250)
);

INVx3_ASAP7_75t_SL g5251 ( 
.A(n_5045),
.Y(n_5251)
);

O2A1O1Ixp33_ASAP7_75t_SL g5252 ( 
.A1(n_4882),
.A2(n_3902),
.B(n_3953),
.C(n_3917),
.Y(n_5252)
);

INVxp67_ASAP7_75t_L g5253 ( 
.A(n_5030),
.Y(n_5253)
);

AOI21xp5_ASAP7_75t_L g5254 ( 
.A1(n_4987),
.A2(n_4290),
.B(n_3699),
.Y(n_5254)
);

OAI22xp33_ASAP7_75t_L g5255 ( 
.A1(n_4621),
.A2(n_4330),
.B1(n_3582),
.B2(n_3551),
.Y(n_5255)
);

BUFx10_ASAP7_75t_L g5256 ( 
.A(n_5073),
.Y(n_5256)
);

BUFx2_ASAP7_75t_L g5257 ( 
.A(n_4711),
.Y(n_5257)
);

AOI22xp5_ASAP7_75t_L g5258 ( 
.A1(n_4712),
.A2(n_3575),
.B1(n_3553),
.B2(n_3853),
.Y(n_5258)
);

OAI21x1_ASAP7_75t_L g5259 ( 
.A1(n_4487),
.A2(n_3688),
.B(n_3684),
.Y(n_5259)
);

AOI21xp5_ASAP7_75t_L g5260 ( 
.A1(n_4987),
.A2(n_3699),
.B(n_4048),
.Y(n_5260)
);

NOR2xp33_ASAP7_75t_L g5261 ( 
.A(n_4578),
.B(n_3695),
.Y(n_5261)
);

AND3x2_ASAP7_75t_L g5262 ( 
.A(n_4833),
.B(n_3879),
.C(n_3719),
.Y(n_5262)
);

AOI21x1_ASAP7_75t_L g5263 ( 
.A1(n_4501),
.A2(n_4373),
.B(n_4487),
.Y(n_5263)
);

INVx4_ASAP7_75t_SL g5264 ( 
.A(n_5099),
.Y(n_5264)
);

NAND2xp5_ASAP7_75t_L g5265 ( 
.A(n_4790),
.B(n_4281),
.Y(n_5265)
);

NAND2xp5_ASAP7_75t_L g5266 ( 
.A(n_4790),
.B(n_4281),
.Y(n_5266)
);

OAI21xp5_ASAP7_75t_L g5267 ( 
.A1(n_4922),
.A2(n_3713),
.B(n_3509),
.Y(n_5267)
);

INVx1_ASAP7_75t_L g5268 ( 
.A(n_4438),
.Y(n_5268)
);

INVx1_ASAP7_75t_L g5269 ( 
.A(n_4438),
.Y(n_5269)
);

O2A1O1Ixp33_ASAP7_75t_SL g5270 ( 
.A1(n_4882),
.A2(n_3938),
.B(n_3520),
.C(n_3890),
.Y(n_5270)
);

OAI21xp5_ASAP7_75t_L g5271 ( 
.A1(n_5066),
.A2(n_3509),
.B(n_3508),
.Y(n_5271)
);

NAND2xp5_ASAP7_75t_SL g5272 ( 
.A(n_4377),
.B(n_4133),
.Y(n_5272)
);

NAND2xp5_ASAP7_75t_L g5273 ( 
.A(n_4791),
.B(n_4246),
.Y(n_5273)
);

NAND2xp5_ASAP7_75t_L g5274 ( 
.A(n_4791),
.B(n_4246),
.Y(n_5274)
);

INVx2_ASAP7_75t_L g5275 ( 
.A(n_4532),
.Y(n_5275)
);

AOI21xp5_ASAP7_75t_L g5276 ( 
.A1(n_5009),
.A2(n_3699),
.B(n_4064),
.Y(n_5276)
);

NAND2xp5_ASAP7_75t_L g5277 ( 
.A(n_4751),
.B(n_4861),
.Y(n_5277)
);

AOI21xp5_ASAP7_75t_L g5278 ( 
.A1(n_5009),
.A2(n_3699),
.B(n_4093),
.Y(n_5278)
);

BUFx3_ASAP7_75t_L g5279 ( 
.A(n_4425),
.Y(n_5279)
);

INVx1_ASAP7_75t_L g5280 ( 
.A(n_4538),
.Y(n_5280)
);

AOI21xp5_ASAP7_75t_SL g5281 ( 
.A1(n_4900),
.A2(n_4025),
.B(n_4000),
.Y(n_5281)
);

OAI221xp5_ASAP7_75t_L g5282 ( 
.A1(n_4901),
.A2(n_3631),
.B1(n_4105),
.B2(n_3671),
.C(n_3708),
.Y(n_5282)
);

O2A1O1Ixp33_ASAP7_75t_L g5283 ( 
.A1(n_5066),
.A2(n_3643),
.B(n_3700),
.C(n_3662),
.Y(n_5283)
);

AOI21xp5_ASAP7_75t_L g5284 ( 
.A1(n_5029),
.A2(n_3699),
.B(n_4231),
.Y(n_5284)
);

INVx1_ASAP7_75t_L g5285 ( 
.A(n_4538),
.Y(n_5285)
);

BUFx3_ASAP7_75t_L g5286 ( 
.A(n_4534),
.Y(n_5286)
);

OAI21x1_ASAP7_75t_SL g5287 ( 
.A1(n_4789),
.A2(n_4310),
.B(n_4124),
.Y(n_5287)
);

AOI21xp5_ASAP7_75t_L g5288 ( 
.A1(n_5029),
.A2(n_4453),
.B(n_4449),
.Y(n_5288)
);

OAI21x1_ASAP7_75t_L g5289 ( 
.A1(n_4373),
.A2(n_3688),
.B(n_3684),
.Y(n_5289)
);

AOI21xp5_ASAP7_75t_L g5290 ( 
.A1(n_4449),
.A2(n_4335),
.B(n_4231),
.Y(n_5290)
);

INVx4_ASAP7_75t_L g5291 ( 
.A(n_4462),
.Y(n_5291)
);

INVx1_ASAP7_75t_L g5292 ( 
.A(n_4539),
.Y(n_5292)
);

NOR2xp33_ASAP7_75t_L g5293 ( 
.A(n_4578),
.B(n_4066),
.Y(n_5293)
);

O2A1O1Ixp33_ASAP7_75t_SL g5294 ( 
.A1(n_5124),
.A2(n_4076),
.B(n_3742),
.C(n_4141),
.Y(n_5294)
);

OAI21x1_ASAP7_75t_L g5295 ( 
.A1(n_4373),
.A2(n_3689),
.B(n_3587),
.Y(n_5295)
);

NAND2xp5_ASAP7_75t_L g5296 ( 
.A(n_4751),
.B(n_4178),
.Y(n_5296)
);

NAND2xp5_ASAP7_75t_SL g5297 ( 
.A(n_4377),
.B(n_4078),
.Y(n_5297)
);

OA21x2_ASAP7_75t_L g5298 ( 
.A1(n_4648),
.A2(n_4004),
.B(n_3689),
.Y(n_5298)
);

INVx1_ASAP7_75t_L g5299 ( 
.A(n_4539),
.Y(n_5299)
);

AOI21xp5_ASAP7_75t_L g5300 ( 
.A1(n_4453),
.A2(n_4335),
.B(n_4329),
.Y(n_5300)
);

NAND2xp5_ASAP7_75t_L g5301 ( 
.A(n_4861),
.B(n_3532),
.Y(n_5301)
);

INVx1_ASAP7_75t_L g5302 ( 
.A(n_4544),
.Y(n_5302)
);

CKINVDCx20_ASAP7_75t_R g5303 ( 
.A(n_5081),
.Y(n_5303)
);

INVx3_ASAP7_75t_L g5304 ( 
.A(n_4388),
.Y(n_5304)
);

AND2x2_ASAP7_75t_L g5305 ( 
.A(n_4978),
.B(n_4253),
.Y(n_5305)
);

AOI21x1_ASAP7_75t_L g5306 ( 
.A1(n_4501),
.A2(n_4366),
.B(n_4073),
.Y(n_5306)
);

AO21x2_ASAP7_75t_L g5307 ( 
.A1(n_4476),
.A2(n_4366),
.B(n_4073),
.Y(n_5307)
);

AND2x4_ASAP7_75t_L g5308 ( 
.A(n_5015),
.B(n_3579),
.Y(n_5308)
);

OAI21x1_ASAP7_75t_L g5309 ( 
.A1(n_4455),
.A2(n_5082),
.B(n_5078),
.Y(n_5309)
);

O2A1O1Ixp33_ASAP7_75t_L g5310 ( 
.A1(n_4541),
.A2(n_3662),
.B(n_3653),
.C(n_3508),
.Y(n_5310)
);

NAND2xp5_ASAP7_75t_SL g5311 ( 
.A(n_4383),
.B(n_4390),
.Y(n_5311)
);

NAND2xp5_ASAP7_75t_L g5312 ( 
.A(n_4439),
.B(n_4543),
.Y(n_5312)
);

AND2x4_ASAP7_75t_L g5313 ( 
.A(n_5015),
.B(n_3579),
.Y(n_5313)
);

OAI21x1_ASAP7_75t_L g5314 ( 
.A1(n_4455),
.A2(n_5082),
.B(n_5078),
.Y(n_5314)
);

AOI21xp5_ASAP7_75t_L g5315 ( 
.A1(n_4942),
.A2(n_4328),
.B(n_3540),
.Y(n_5315)
);

OAI22xp5_ASAP7_75t_L g5316 ( 
.A1(n_4396),
.A2(n_3831),
.B1(n_3913),
.B2(n_3591),
.Y(n_5316)
);

BUFx2_ASAP7_75t_L g5317 ( 
.A(n_4947),
.Y(n_5317)
);

BUFx10_ASAP7_75t_L g5318 ( 
.A(n_4422),
.Y(n_5318)
);

NOR2xp33_ASAP7_75t_L g5319 ( 
.A(n_4524),
.B(n_4135),
.Y(n_5319)
);

OAI21x1_ASAP7_75t_L g5320 ( 
.A1(n_4455),
.A2(n_3587),
.B(n_3647),
.Y(n_5320)
);

A2O1A1Ixp33_ASAP7_75t_L g5321 ( 
.A1(n_4654),
.A2(n_4180),
.B(n_3591),
.C(n_4328),
.Y(n_5321)
);

INVx1_ASAP7_75t_L g5322 ( 
.A(n_4544),
.Y(n_5322)
);

INVx4_ASAP7_75t_L g5323 ( 
.A(n_4462),
.Y(n_5323)
);

BUFx3_ASAP7_75t_L g5324 ( 
.A(n_4534),
.Y(n_5324)
);

AOI21xp5_ASAP7_75t_L g5325 ( 
.A1(n_4470),
.A2(n_3540),
.B(n_3532),
.Y(n_5325)
);

A2O1A1Ixp33_ASAP7_75t_L g5326 ( 
.A1(n_4396),
.A2(n_3591),
.B(n_4122),
.C(n_4058),
.Y(n_5326)
);

NAND3xp33_ASAP7_75t_SL g5327 ( 
.A(n_4901),
.B(n_3683),
.C(n_3681),
.Y(n_5327)
);

AOI21xp5_ASAP7_75t_L g5328 ( 
.A1(n_4470),
.A2(n_4325),
.B(n_4134),
.Y(n_5328)
);

AOI22xp33_ASAP7_75t_L g5329 ( 
.A1(n_4447),
.A2(n_4097),
.B1(n_4081),
.B2(n_3612),
.Y(n_5329)
);

A2O1A1Ixp33_ASAP7_75t_L g5330 ( 
.A1(n_4386),
.A2(n_4122),
.B(n_3714),
.C(n_3579),
.Y(n_5330)
);

AOI21xp5_ASAP7_75t_L g5331 ( 
.A1(n_4915),
.A2(n_4145),
.B(n_4129),
.Y(n_5331)
);

A2O1A1Ixp33_ASAP7_75t_L g5332 ( 
.A1(n_4386),
.A2(n_3579),
.B(n_3639),
.C(n_3612),
.Y(n_5332)
);

AO31x2_ASAP7_75t_L g5333 ( 
.A1(n_4820),
.A2(n_4270),
.A3(n_4273),
.B(n_4245),
.Y(n_5333)
);

INVx5_ASAP7_75t_L g5334 ( 
.A(n_4971),
.Y(n_5334)
);

BUFx3_ASAP7_75t_L g5335 ( 
.A(n_5080),
.Y(n_5335)
);

NAND2xp5_ASAP7_75t_L g5336 ( 
.A(n_4439),
.B(n_4543),
.Y(n_5336)
);

CKINVDCx20_ASAP7_75t_R g5337 ( 
.A(n_5081),
.Y(n_5337)
);

OAI21x1_ASAP7_75t_L g5338 ( 
.A1(n_5082),
.A2(n_3587),
.B(n_3647),
.Y(n_5338)
);

INVx2_ASAP7_75t_L g5339 ( 
.A(n_4532),
.Y(n_5339)
);

INVx2_ASAP7_75t_L g5340 ( 
.A(n_4551),
.Y(n_5340)
);

AOI21xp5_ASAP7_75t_L g5341 ( 
.A1(n_4518),
.A2(n_4166),
.B(n_3596),
.Y(n_5341)
);

OAI21xp5_ASAP7_75t_L g5342 ( 
.A1(n_4968),
.A2(n_4147),
.B(n_3596),
.Y(n_5342)
);

AO31x2_ASAP7_75t_L g5343 ( 
.A1(n_5037),
.A2(n_4295),
.A3(n_4302),
.B(n_4294),
.Y(n_5343)
);

AOI21xp5_ASAP7_75t_L g5344 ( 
.A1(n_4915),
.A2(n_4336),
.B(n_4216),
.Y(n_5344)
);

INVx1_ASAP7_75t_L g5345 ( 
.A(n_4550),
.Y(n_5345)
);

AOI21xp5_ASAP7_75t_L g5346 ( 
.A1(n_4518),
.A2(n_4336),
.B(n_3630),
.Y(n_5346)
);

INVx1_ASAP7_75t_L g5347 ( 
.A(n_4550),
.Y(n_5347)
);

INVx5_ASAP7_75t_L g5348 ( 
.A(n_4971),
.Y(n_5348)
);

OAI21xp5_ASAP7_75t_L g5349 ( 
.A1(n_4968),
.A2(n_4147),
.B(n_3563),
.Y(n_5349)
);

AOI21xp5_ASAP7_75t_L g5350 ( 
.A1(n_4519),
.A2(n_3630),
.B(n_3626),
.Y(n_5350)
);

HB1xp67_ASAP7_75t_L g5351 ( 
.A(n_4811),
.Y(n_5351)
);

INVx2_ASAP7_75t_L g5352 ( 
.A(n_4551),
.Y(n_5352)
);

INVx1_ASAP7_75t_SL g5353 ( 
.A(n_4432),
.Y(n_5353)
);

AOI221xp5_ASAP7_75t_SL g5354 ( 
.A1(n_4706),
.A2(n_3957),
.B1(n_3686),
.B2(n_3841),
.C(n_3633),
.Y(n_5354)
);

OAI21x1_ASAP7_75t_L g5355 ( 
.A1(n_5078),
.A2(n_3647),
.B(n_3701),
.Y(n_5355)
);

INVx1_ASAP7_75t_L g5356 ( 
.A(n_4553),
.Y(n_5356)
);

INVx3_ASAP7_75t_L g5357 ( 
.A(n_5142),
.Y(n_5357)
);

OAI21xp5_ASAP7_75t_L g5358 ( 
.A1(n_4974),
.A2(n_4552),
.B(n_4401),
.Y(n_5358)
);

INVx3_ASAP7_75t_L g5359 ( 
.A(n_5142),
.Y(n_5359)
);

AOI22xp5_ASAP7_75t_L g5360 ( 
.A1(n_5012),
.A2(n_4552),
.B1(n_4685),
.B2(n_4932),
.Y(n_5360)
);

A2O1A1Ixp33_ASAP7_75t_L g5361 ( 
.A1(n_4541),
.A2(n_3612),
.B(n_3670),
.C(n_3639),
.Y(n_5361)
);

CKINVDCx5p33_ASAP7_75t_R g5362 ( 
.A(n_4515),
.Y(n_5362)
);

OAI21x1_ASAP7_75t_L g5363 ( 
.A1(n_4648),
.A2(n_3647),
.B(n_3701),
.Y(n_5363)
);

INVx1_ASAP7_75t_L g5364 ( 
.A(n_4553),
.Y(n_5364)
);

OAI21x1_ASAP7_75t_L g5365 ( 
.A1(n_4648),
.A2(n_3701),
.B(n_4115),
.Y(n_5365)
);

AND2x4_ASAP7_75t_L g5366 ( 
.A(n_5015),
.B(n_3612),
.Y(n_5366)
);

OAI21x1_ASAP7_75t_L g5367 ( 
.A1(n_4603),
.A2(n_3701),
.B(n_4126),
.Y(n_5367)
);

AO31x2_ASAP7_75t_L g5368 ( 
.A1(n_5037),
.A2(n_4318),
.A3(n_4323),
.B(n_4311),
.Y(n_5368)
);

OAI22x1_ASAP7_75t_L g5369 ( 
.A1(n_4667),
.A2(n_3702),
.B1(n_3723),
.B2(n_3519),
.Y(n_5369)
);

AOI21xp5_ASAP7_75t_L g5370 ( 
.A1(n_4921),
.A2(n_4193),
.B(n_4152),
.Y(n_5370)
);

AND2x4_ASAP7_75t_L g5371 ( 
.A(n_5015),
.B(n_3612),
.Y(n_5371)
);

OAI21xp5_ASAP7_75t_L g5372 ( 
.A1(n_4974),
.A2(n_3563),
.B(n_3660),
.Y(n_5372)
);

OR2x2_ASAP7_75t_L g5373 ( 
.A(n_4567),
.B(n_3702),
.Y(n_5373)
);

AOI22xp5_ASAP7_75t_SL g5374 ( 
.A1(n_4706),
.A2(n_4957),
.B1(n_4662),
.B2(n_4579),
.Y(n_5374)
);

CKINVDCx16_ASAP7_75t_R g5375 ( 
.A(n_5080),
.Y(n_5375)
);

AOI21xp5_ASAP7_75t_L g5376 ( 
.A1(n_4937),
.A2(n_4193),
.B(n_4152),
.Y(n_5376)
);

INVx2_ASAP7_75t_L g5377 ( 
.A(n_4551),
.Y(n_5377)
);

BUFx2_ASAP7_75t_L g5378 ( 
.A(n_4947),
.Y(n_5378)
);

OAI21xp33_ASAP7_75t_L g5379 ( 
.A1(n_4685),
.A2(n_3980),
.B(n_3975),
.Y(n_5379)
);

BUFx2_ASAP7_75t_L g5380 ( 
.A(n_4947),
.Y(n_5380)
);

AOI21xp5_ASAP7_75t_L g5381 ( 
.A1(n_4937),
.A2(n_4193),
.B(n_4152),
.Y(n_5381)
);

AOI21xp5_ASAP7_75t_L g5382 ( 
.A1(n_4970),
.A2(n_4193),
.B(n_3630),
.Y(n_5382)
);

INVx1_ASAP7_75t_L g5383 ( 
.A(n_4617),
.Y(n_5383)
);

INVx1_ASAP7_75t_L g5384 ( 
.A(n_4617),
.Y(n_5384)
);

OR2x6_ASAP7_75t_L g5385 ( 
.A(n_4592),
.B(n_3612),
.Y(n_5385)
);

AO22x1_ASAP7_75t_L g5386 ( 
.A1(n_5044),
.A2(n_4300),
.B1(n_3598),
.B2(n_3676),
.Y(n_5386)
);

OR2x2_ASAP7_75t_L g5387 ( 
.A(n_4567),
.B(n_3723),
.Y(n_5387)
);

NAND2xp5_ASAP7_75t_L g5388 ( 
.A(n_4383),
.B(n_4275),
.Y(n_5388)
);

NOR2xp67_ASAP7_75t_L g5389 ( 
.A(n_4561),
.B(n_3612),
.Y(n_5389)
);

OAI21x1_ASAP7_75t_L g5390 ( 
.A1(n_4482),
.A2(n_4151),
.B(n_4130),
.Y(n_5390)
);

AND2x2_ASAP7_75t_L g5391 ( 
.A(n_5023),
.B(n_4253),
.Y(n_5391)
);

A2O1A1Ixp33_ASAP7_75t_L g5392 ( 
.A1(n_4568),
.A2(n_3639),
.B(n_3685),
.C(n_3670),
.Y(n_5392)
);

INVx1_ASAP7_75t_L g5393 ( 
.A(n_4622),
.Y(n_5393)
);

INVx2_ASAP7_75t_L g5394 ( 
.A(n_4596),
.Y(n_5394)
);

NAND3xp33_ASAP7_75t_SL g5395 ( 
.A(n_4774),
.B(n_3633),
.C(n_3632),
.Y(n_5395)
);

AO31x2_ASAP7_75t_L g5396 ( 
.A1(n_5037),
.A2(n_4350),
.A3(n_4361),
.B(n_4344),
.Y(n_5396)
);

AOI21xp5_ASAP7_75t_L g5397 ( 
.A1(n_4519),
.A2(n_3630),
.B(n_3626),
.Y(n_5397)
);

INVx1_ASAP7_75t_L g5398 ( 
.A(n_4622),
.Y(n_5398)
);

INVx1_ASAP7_75t_L g5399 ( 
.A(n_4625),
.Y(n_5399)
);

OA21x2_ASAP7_75t_L g5400 ( 
.A1(n_5028),
.A2(n_4151),
.B(n_4130),
.Y(n_5400)
);

OAI21xp5_ASAP7_75t_L g5401 ( 
.A1(n_4401),
.A2(n_3660),
.B(n_3485),
.Y(n_5401)
);

NOR4xp25_ASAP7_75t_L g5402 ( 
.A(n_4433),
.B(n_3632),
.C(n_3957),
.D(n_3975),
.Y(n_5402)
);

OAI21xp5_ASAP7_75t_L g5403 ( 
.A1(n_4561),
.A2(n_3485),
.B(n_3474),
.Y(n_5403)
);

INVx1_ASAP7_75t_L g5404 ( 
.A(n_4625),
.Y(n_5404)
);

A2O1A1Ixp33_ASAP7_75t_L g5405 ( 
.A1(n_4568),
.A2(n_3639),
.B(n_3685),
.C(n_3670),
.Y(n_5405)
);

OAI21xp5_ASAP7_75t_L g5406 ( 
.A1(n_5012),
.A2(n_3493),
.B(n_3474),
.Y(n_5406)
);

OAI21xp5_ASAP7_75t_L g5407 ( 
.A1(n_5124),
.A2(n_4659),
.B(n_4390),
.Y(n_5407)
);

INVx1_ASAP7_75t_L g5408 ( 
.A(n_4627),
.Y(n_5408)
);

OAI22xp5_ASAP7_75t_L g5409 ( 
.A1(n_4591),
.A2(n_3980),
.B1(n_3994),
.B2(n_3984),
.Y(n_5409)
);

INVx1_ASAP7_75t_L g5410 ( 
.A(n_4627),
.Y(n_5410)
);

NOR2xp67_ASAP7_75t_L g5411 ( 
.A(n_4525),
.B(n_3639),
.Y(n_5411)
);

NOR2xp33_ASAP7_75t_L g5412 ( 
.A(n_4524),
.B(n_4027),
.Y(n_5412)
);

O2A1O1Ixp33_ASAP7_75t_SL g5413 ( 
.A1(n_4660),
.A2(n_4834),
.B(n_4489),
.C(n_4977),
.Y(n_5413)
);

INVx2_ASAP7_75t_L g5414 ( 
.A(n_4596),
.Y(n_5414)
);

OAI21xp5_ASAP7_75t_L g5415 ( 
.A1(n_5006),
.A2(n_5014),
.B(n_4967),
.Y(n_5415)
);

A2O1A1Ixp33_ASAP7_75t_L g5416 ( 
.A1(n_4932),
.A2(n_3639),
.B(n_3685),
.C(n_3670),
.Y(n_5416)
);

AOI21xp5_ASAP7_75t_L g5417 ( 
.A1(n_4525),
.A2(n_3630),
.B(n_3626),
.Y(n_5417)
);

AND2x2_ASAP7_75t_L g5418 ( 
.A(n_5023),
.B(n_4253),
.Y(n_5418)
);

OAI21xp5_ASAP7_75t_L g5419 ( 
.A1(n_5006),
.A2(n_3505),
.B(n_3493),
.Y(n_5419)
);

INVx2_ASAP7_75t_L g5420 ( 
.A(n_4596),
.Y(n_5420)
);

OAI22xp5_ASAP7_75t_L g5421 ( 
.A1(n_4591),
.A2(n_3984),
.B1(n_3995),
.B2(n_3994),
.Y(n_5421)
);

AOI21xp5_ASAP7_75t_L g5422 ( 
.A1(n_4526),
.A2(n_4661),
.B(n_4565),
.Y(n_5422)
);

NOR2xp67_ASAP7_75t_L g5423 ( 
.A(n_4526),
.B(n_3639),
.Y(n_5423)
);

BUFx10_ASAP7_75t_L g5424 ( 
.A(n_4422),
.Y(n_5424)
);

NAND2xp5_ASAP7_75t_SL g5425 ( 
.A(n_4397),
.B(n_4621),
.Y(n_5425)
);

NOR2xp67_ASAP7_75t_L g5426 ( 
.A(n_4613),
.B(n_3670),
.Y(n_5426)
);

BUFx3_ASAP7_75t_L g5427 ( 
.A(n_5080),
.Y(n_5427)
);

AOI22xp5_ASAP7_75t_L g5428 ( 
.A1(n_4513),
.A2(n_4447),
.B1(n_4684),
.B2(n_4468),
.Y(n_5428)
);

INVx1_ASAP7_75t_L g5429 ( 
.A(n_4644),
.Y(n_5429)
);

INVx2_ASAP7_75t_L g5430 ( 
.A(n_4602),
.Y(n_5430)
);

A2O1A1Ixp33_ASAP7_75t_L g5431 ( 
.A1(n_4660),
.A2(n_3670),
.B(n_3693),
.C(n_3685),
.Y(n_5431)
);

BUFx12f_ASAP7_75t_L g5432 ( 
.A(n_4524),
.Y(n_5432)
);

NAND2xp5_ASAP7_75t_L g5433 ( 
.A(n_4397),
.B(n_4275),
.Y(n_5433)
);

OAI21xp5_ASAP7_75t_L g5434 ( 
.A1(n_5014),
.A2(n_3512),
.B(n_3505),
.Y(n_5434)
);

OAI21x1_ASAP7_75t_L g5435 ( 
.A1(n_4486),
.A2(n_3721),
.B(n_3618),
.Y(n_5435)
);

AOI21xp5_ASAP7_75t_L g5436 ( 
.A1(n_4827),
.A2(n_3630),
.B(n_3626),
.Y(n_5436)
);

A2O1A1Ixp33_ASAP7_75t_L g5437 ( 
.A1(n_4809),
.A2(n_3670),
.B(n_3693),
.C(n_3685),
.Y(n_5437)
);

AOI211xp5_ASAP7_75t_L g5438 ( 
.A1(n_4393),
.A2(n_3693),
.B(n_3685),
.C(n_3995),
.Y(n_5438)
);

NOR2xp33_ASAP7_75t_SL g5439 ( 
.A(n_4774),
.B(n_4342),
.Y(n_5439)
);

INVx1_ASAP7_75t_L g5440 ( 
.A(n_4644),
.Y(n_5440)
);

OR2x2_ASAP7_75t_L g5441 ( 
.A(n_4581),
.B(n_4159),
.Y(n_5441)
);

NAND2xp5_ASAP7_75t_SL g5442 ( 
.A(n_4774),
.B(n_4809),
.Y(n_5442)
);

NAND2xp5_ASAP7_75t_SL g5443 ( 
.A(n_4684),
.B(n_3676),
.Y(n_5443)
);

A2O1A1Ixp33_ASAP7_75t_L g5444 ( 
.A1(n_4680),
.A2(n_3685),
.B(n_3693),
.C(n_3535),
.Y(n_5444)
);

AND2x4_ASAP7_75t_L g5445 ( 
.A(n_4642),
.B(n_3693),
.Y(n_5445)
);

AOI21xp5_ASAP7_75t_L g5446 ( 
.A1(n_4827),
.A2(n_3626),
.B(n_3693),
.Y(n_5446)
);

OR2x2_ASAP7_75t_L g5447 ( 
.A(n_4581),
.B(n_4159),
.Y(n_5447)
);

OAI21x1_ASAP7_75t_L g5448 ( 
.A1(n_4486),
.A2(n_3933),
.B(n_3792),
.Y(n_5448)
);

INVx1_ASAP7_75t_L g5449 ( 
.A(n_4646),
.Y(n_5449)
);

AOI21xp5_ASAP7_75t_L g5450 ( 
.A1(n_4565),
.A2(n_3517),
.B(n_3512),
.Y(n_5450)
);

HB1xp67_ASAP7_75t_L g5451 ( 
.A(n_4811),
.Y(n_5451)
);

OR2x2_ASAP7_75t_L g5452 ( 
.A(n_4480),
.B(n_4168),
.Y(n_5452)
);

NAND2xp5_ASAP7_75t_L g5453 ( 
.A(n_5071),
.B(n_4092),
.Y(n_5453)
);

NOR2xp33_ASAP7_75t_L g5454 ( 
.A(n_4517),
.B(n_4110),
.Y(n_5454)
);

INVx1_ASAP7_75t_L g5455 ( 
.A(n_4646),
.Y(n_5455)
);

NAND3x1_ASAP7_75t_L g5456 ( 
.A(n_4817),
.B(n_4300),
.C(n_4002),
.Y(n_5456)
);

INVxp67_ASAP7_75t_SL g5457 ( 
.A(n_4665),
.Y(n_5457)
);

INVx1_ASAP7_75t_L g5458 ( 
.A(n_4702),
.Y(n_5458)
);

CKINVDCx5p33_ASAP7_75t_R g5459 ( 
.A(n_4977),
.Y(n_5459)
);

AOI21xp5_ASAP7_75t_L g5460 ( 
.A1(n_4829),
.A2(n_3693),
.B(n_3517),
.Y(n_5460)
);

AOI221x1_ASAP7_75t_L g5461 ( 
.A1(n_4966),
.A2(n_3651),
.B1(n_3656),
.B2(n_3654),
.C(n_3679),
.Y(n_5461)
);

AOI21xp5_ASAP7_75t_L g5462 ( 
.A1(n_4829),
.A2(n_4306),
.B(n_3507),
.Y(n_5462)
);

AOI21x1_ASAP7_75t_L g5463 ( 
.A1(n_4818),
.A2(n_3654),
.B(n_3651),
.Y(n_5463)
);

BUFx2_ASAP7_75t_L g5464 ( 
.A(n_4990),
.Y(n_5464)
);

NAND2xp5_ASAP7_75t_L g5465 ( 
.A(n_5071),
.B(n_4287),
.Y(n_5465)
);

OAI21xp5_ASAP7_75t_L g5466 ( 
.A1(n_4967),
.A2(n_3523),
.B(n_3522),
.Y(n_5466)
);

NAND2x1p5_ASAP7_75t_L g5467 ( 
.A(n_5040),
.B(n_4316),
.Y(n_5467)
);

AOI21xp5_ASAP7_75t_SL g5468 ( 
.A1(n_4834),
.A2(n_3503),
.B(n_3497),
.Y(n_5468)
);

NOR2xp33_ASAP7_75t_L g5469 ( 
.A(n_4635),
.B(n_4110),
.Y(n_5469)
);

AOI22xp5_ASAP7_75t_L g5470 ( 
.A1(n_4513),
.A2(n_3564),
.B1(n_3535),
.B2(n_3996),
.Y(n_5470)
);

INVx2_ASAP7_75t_L g5471 ( 
.A(n_4602),
.Y(n_5471)
);

NOR2xp33_ASAP7_75t_L g5472 ( 
.A(n_4635),
.B(n_4110),
.Y(n_5472)
);

INVxp67_ASAP7_75t_SL g5473 ( 
.A(n_4670),
.Y(n_5473)
);

NAND2xp5_ASAP7_75t_L g5474 ( 
.A(n_4869),
.B(n_4287),
.Y(n_5474)
);

BUFx2_ASAP7_75t_L g5475 ( 
.A(n_4990),
.Y(n_5475)
);

AOI21xp5_ASAP7_75t_L g5476 ( 
.A1(n_4830),
.A2(n_4966),
.B(n_4537),
.Y(n_5476)
);

AOI221x1_ASAP7_75t_L g5477 ( 
.A1(n_4966),
.A2(n_3656),
.B1(n_3679),
.B2(n_3593),
.C(n_3569),
.Y(n_5477)
);

NAND2xp5_ASAP7_75t_L g5478 ( 
.A(n_4869),
.B(n_3857),
.Y(n_5478)
);

OAI21x1_ASAP7_75t_L g5479 ( 
.A1(n_5112),
.A2(n_3933),
.B(n_3792),
.Y(n_5479)
);

AOI21xp5_ASAP7_75t_L g5480 ( 
.A1(n_4830),
.A2(n_3564),
.B(n_4144),
.Y(n_5480)
);

INVx1_ASAP7_75t_L g5481 ( 
.A(n_4702),
.Y(n_5481)
);

AOI21xp5_ASAP7_75t_L g5482 ( 
.A1(n_4537),
.A2(n_3564),
.B(n_4144),
.Y(n_5482)
);

AND2x2_ASAP7_75t_L g5483 ( 
.A(n_5023),
.B(n_4360),
.Y(n_5483)
);

AOI21xp5_ASAP7_75t_L g5484 ( 
.A1(n_4793),
.A2(n_4153),
.B(n_4150),
.Y(n_5484)
);

NAND2xp5_ASAP7_75t_L g5485 ( 
.A(n_4871),
.B(n_3857),
.Y(n_5485)
);

AOI21xp5_ASAP7_75t_SL g5486 ( 
.A1(n_4851),
.A2(n_3530),
.B(n_3503),
.Y(n_5486)
);

A2O1A1Ixp33_ASAP7_75t_L g5487 ( 
.A1(n_4680),
.A2(n_3535),
.B(n_4169),
.C(n_3507),
.Y(n_5487)
);

INVx1_ASAP7_75t_L g5488 ( 
.A(n_4758),
.Y(n_5488)
);

NOR2xp33_ASAP7_75t_SL g5489 ( 
.A(n_4545),
.B(n_3503),
.Y(n_5489)
);

NAND2xp5_ASAP7_75t_L g5490 ( 
.A(n_4871),
.B(n_4420),
.Y(n_5490)
);

OAI21x1_ASAP7_75t_L g5491 ( 
.A1(n_5112),
.A2(n_3933),
.B(n_3792),
.Y(n_5491)
);

AOI22xp33_ASAP7_75t_L g5492 ( 
.A1(n_4393),
.A2(n_3738),
.B1(n_3950),
.B2(n_3919),
.Y(n_5492)
);

AND2x2_ASAP7_75t_L g5493 ( 
.A(n_4742),
.B(n_4360),
.Y(n_5493)
);

AOI21xp5_ASAP7_75t_L g5494 ( 
.A1(n_4616),
.A2(n_4626),
.B(n_5114),
.Y(n_5494)
);

NAND3xp33_ASAP7_75t_L g5495 ( 
.A(n_4446),
.B(n_3692),
.C(n_3680),
.Y(n_5495)
);

OAI21x1_ASAP7_75t_SL g5496 ( 
.A1(n_4949),
.A2(n_4181),
.B(n_4177),
.Y(n_5496)
);

NOR2xp33_ASAP7_75t_SL g5497 ( 
.A(n_4545),
.B(n_3530),
.Y(n_5497)
);

O2A1O1Ixp33_ASAP7_75t_SL g5498 ( 
.A1(n_4489),
.A2(n_3531),
.B(n_3628),
.C(n_3996),
.Y(n_5498)
);

INVx2_ASAP7_75t_SL g5499 ( 
.A(n_5127),
.Y(n_5499)
);

AOI21xp5_ASAP7_75t_L g5500 ( 
.A1(n_4616),
.A2(n_4626),
.B(n_5114),
.Y(n_5500)
);

INVx2_ASAP7_75t_L g5501 ( 
.A(n_4602),
.Y(n_5501)
);

OA21x2_ASAP7_75t_L g5502 ( 
.A1(n_5028),
.A2(n_4189),
.B(n_4357),
.Y(n_5502)
);

NAND2x1_ASAP7_75t_L g5503 ( 
.A(n_4406),
.B(n_3718),
.Y(n_5503)
);

AOI21xp5_ASAP7_75t_L g5504 ( 
.A1(n_5114),
.A2(n_3557),
.B(n_3494),
.Y(n_5504)
);

CKINVDCx20_ASAP7_75t_R g5505 ( 
.A(n_5110),
.Y(n_5505)
);

NOR2xp67_ASAP7_75t_L g5506 ( 
.A(n_4620),
.B(n_4687),
.Y(n_5506)
);

NOR2xp33_ASAP7_75t_L g5507 ( 
.A(n_5076),
.B(n_4131),
.Y(n_5507)
);

BUFx2_ASAP7_75t_R g5508 ( 
.A(n_4464),
.Y(n_5508)
);

AOI21x1_ASAP7_75t_L g5509 ( 
.A1(n_4818),
.A2(n_4369),
.B(n_4327),
.Y(n_5509)
);

NAND3xp33_ASAP7_75t_L g5510 ( 
.A(n_4446),
.B(n_3692),
.C(n_3680),
.Y(n_5510)
);

NAND2xp5_ASAP7_75t_L g5511 ( 
.A(n_4420),
.B(n_3861),
.Y(n_5511)
);

BUFx3_ASAP7_75t_L g5512 ( 
.A(n_5044),
.Y(n_5512)
);

OAI21xp5_ASAP7_75t_L g5513 ( 
.A1(n_4440),
.A2(n_4924),
.B(n_4876),
.Y(n_5513)
);

A2O1A1Ixp33_ASAP7_75t_L g5514 ( 
.A1(n_4689),
.A2(n_4169),
.B(n_3557),
.C(n_3657),
.Y(n_5514)
);

CKINVDCx20_ASAP7_75t_R g5515 ( 
.A(n_5110),
.Y(n_5515)
);

INVx3_ASAP7_75t_L g5516 ( 
.A(n_4388),
.Y(n_5516)
);

NAND2xp33_ASAP7_75t_L g5517 ( 
.A(n_4493),
.B(n_2980),
.Y(n_5517)
);

AOI21xp5_ASAP7_75t_L g5518 ( 
.A1(n_4476),
.A2(n_3657),
.B(n_3494),
.Y(n_5518)
);

INVx1_ASAP7_75t_L g5519 ( 
.A(n_4758),
.Y(n_5519)
);

OAI21x1_ASAP7_75t_L g5520 ( 
.A1(n_4785),
.A2(n_4155),
.B(n_4137),
.Y(n_5520)
);

OAI21x1_ASAP7_75t_L g5521 ( 
.A1(n_5036),
.A2(n_4155),
.B(n_4137),
.Y(n_5521)
);

NOR2xp33_ASAP7_75t_L g5522 ( 
.A(n_5076),
.B(n_4131),
.Y(n_5522)
);

INVx1_ASAP7_75t_L g5523 ( 
.A(n_4772),
.Y(n_5523)
);

NOR2x1_ASAP7_75t_SL g5524 ( 
.A(n_4620),
.B(n_4235),
.Y(n_5524)
);

A2O1A1Ixp33_ASAP7_75t_L g5525 ( 
.A1(n_4689),
.A2(n_4169),
.B(n_3774),
.C(n_3720),
.Y(n_5525)
);

HB1xp67_ASAP7_75t_L g5526 ( 
.A(n_4563),
.Y(n_5526)
);

NAND2xp5_ASAP7_75t_L g5527 ( 
.A(n_4426),
.B(n_3861),
.Y(n_5527)
);

AOI221xp5_ASAP7_75t_L g5528 ( 
.A1(n_4924),
.A2(n_3773),
.B1(n_3789),
.B2(n_3788),
.C(n_3778),
.Y(n_5528)
);

NAND2xp5_ASAP7_75t_L g5529 ( 
.A(n_4426),
.B(n_4200),
.Y(n_5529)
);

OAI21xp5_ASAP7_75t_L g5530 ( 
.A1(n_4440),
.A2(n_3523),
.B(n_3522),
.Y(n_5530)
);

OAI22x1_ASAP7_75t_L g5531 ( 
.A1(n_4667),
.A2(n_4279),
.B1(n_4188),
.B2(n_3738),
.Y(n_5531)
);

AOI21x1_ASAP7_75t_L g5532 ( 
.A1(n_4818),
.A2(n_4327),
.B(n_3717),
.Y(n_5532)
);

O2A1O1Ixp5_ASAP7_75t_SL g5533 ( 
.A1(n_4902),
.A2(n_4303),
.B(n_4228),
.C(n_3402),
.Y(n_5533)
);

OAI21xp5_ASAP7_75t_SL g5534 ( 
.A1(n_4608),
.A2(n_2836),
.B(n_2847),
.Y(n_5534)
);

INVx1_ASAP7_75t_L g5535 ( 
.A(n_4772),
.Y(n_5535)
);

AOI22xp33_ASAP7_75t_L g5536 ( 
.A1(n_4407),
.A2(n_3738),
.B1(n_3950),
.B2(n_3919),
.Y(n_5536)
);

OR2x6_ASAP7_75t_L g5537 ( 
.A(n_4605),
.B(n_4235),
.Y(n_5537)
);

OAI22xp5_ASAP7_75t_L g5538 ( 
.A1(n_5113),
.A2(n_4009),
.B1(n_4021),
.B2(n_4002),
.Y(n_5538)
);

AND2x2_ASAP7_75t_L g5539 ( 
.A(n_4742),
.B(n_4362),
.Y(n_5539)
);

BUFx3_ASAP7_75t_L g5540 ( 
.A(n_5044),
.Y(n_5540)
);

A2O1A1Ixp33_ASAP7_75t_L g5541 ( 
.A1(n_4688),
.A2(n_3728),
.B(n_3727),
.C(n_3620),
.Y(n_5541)
);

OAI21x1_ASAP7_75t_L g5542 ( 
.A1(n_5050),
.A2(n_4256),
.B(n_4239),
.Y(n_5542)
);

OAI21x1_ASAP7_75t_L g5543 ( 
.A1(n_5050),
.A2(n_4256),
.B(n_4239),
.Y(n_5543)
);

OAI21x1_ASAP7_75t_SL g5544 ( 
.A1(n_4949),
.A2(n_4176),
.B(n_4175),
.Y(n_5544)
);

INVx4_ASAP7_75t_L g5545 ( 
.A(n_4462),
.Y(n_5545)
);

NAND2xp5_ASAP7_75t_L g5546 ( 
.A(n_4890),
.B(n_4200),
.Y(n_5546)
);

INVx2_ASAP7_75t_L g5547 ( 
.A(n_4614),
.Y(n_5547)
);

NAND2xp5_ASAP7_75t_L g5548 ( 
.A(n_4890),
.B(n_4212),
.Y(n_5548)
);

OA21x2_ASAP7_75t_L g5549 ( 
.A1(n_4824),
.A2(n_4491),
.B(n_4846),
.Y(n_5549)
);

AO31x2_ASAP7_75t_L g5550 ( 
.A1(n_4842),
.A2(n_3908),
.A3(n_3921),
.B(n_3899),
.Y(n_5550)
);

NAND2xp33_ASAP7_75t_R g5551 ( 
.A(n_4850),
.B(n_3676),
.Y(n_5551)
);

INVx8_ASAP7_75t_L g5552 ( 
.A(n_5099),
.Y(n_5552)
);

INVx1_ASAP7_75t_L g5553 ( 
.A(n_4781),
.Y(n_5553)
);

AOI21xp5_ASAP7_75t_L g5554 ( 
.A1(n_4547),
.A2(n_4153),
.B(n_4150),
.Y(n_5554)
);

HB1xp67_ASAP7_75t_L g5555 ( 
.A(n_4563),
.Y(n_5555)
);

BUFx6f_ASAP7_75t_L g5556 ( 
.A(n_4388),
.Y(n_5556)
);

O2A1O1Ixp33_ASAP7_75t_SL g5557 ( 
.A1(n_4421),
.A2(n_4009),
.B(n_4022),
.C(n_4021),
.Y(n_5557)
);

A2O1A1Ixp33_ASAP7_75t_L g5558 ( 
.A1(n_4851),
.A2(n_3728),
.B(n_3727),
.C(n_3620),
.Y(n_5558)
);

O2A1O1Ixp5_ASAP7_75t_L g5559 ( 
.A1(n_4884),
.A2(n_4941),
.B(n_4911),
.C(n_4577),
.Y(n_5559)
);

OAI21x1_ASAP7_75t_L g5560 ( 
.A1(n_4444),
.A2(n_4256),
.B(n_4239),
.Y(n_5560)
);

AOI21xp5_ASAP7_75t_L g5561 ( 
.A1(n_4547),
.A2(n_4162),
.B(n_4158),
.Y(n_5561)
);

NOR2xp33_ASAP7_75t_L g5562 ( 
.A(n_4805),
.B(n_4131),
.Y(n_5562)
);

AOI21xp5_ASAP7_75t_L g5563 ( 
.A1(n_4559),
.A2(n_4162),
.B(n_4158),
.Y(n_5563)
);

AND2x2_ASAP7_75t_L g5564 ( 
.A(n_4742),
.B(n_4362),
.Y(n_5564)
);

BUFx10_ASAP7_75t_L g5565 ( 
.A(n_4422),
.Y(n_5565)
);

NOR2xp67_ASAP7_75t_L g5566 ( 
.A(n_4687),
.B(n_4269),
.Y(n_5566)
);

A2O1A1Ixp33_ASAP7_75t_L g5567 ( 
.A1(n_4605),
.A2(n_4611),
.B(n_4929),
.C(n_4916),
.Y(n_5567)
);

INVx1_ASAP7_75t_L g5568 ( 
.A(n_4781),
.Y(n_5568)
);

AOI22xp33_ASAP7_75t_L g5569 ( 
.A1(n_4407),
.A2(n_3738),
.B1(n_3950),
.B2(n_3919),
.Y(n_5569)
);

NAND2xp5_ASAP7_75t_L g5570 ( 
.A(n_4812),
.B(n_4212),
.Y(n_5570)
);

NAND2xp5_ASAP7_75t_L g5571 ( 
.A(n_4812),
.B(n_4188),
.Y(n_5571)
);

O2A1O1Ixp33_ASAP7_75t_SL g5572 ( 
.A1(n_4421),
.A2(n_4022),
.B(n_4030),
.C(n_4026),
.Y(n_5572)
);

O2A1O1Ixp33_ASAP7_75t_L g5573 ( 
.A1(n_4566),
.A2(n_4026),
.B(n_4041),
.C(n_4030),
.Y(n_5573)
);

O2A1O1Ixp33_ASAP7_75t_SL g5574 ( 
.A1(n_4424),
.A2(n_4041),
.B(n_4061),
.C(n_4043),
.Y(n_5574)
);

AND2x2_ASAP7_75t_L g5575 ( 
.A(n_4742),
.B(n_4235),
.Y(n_5575)
);

NAND2xp5_ASAP7_75t_L g5576 ( 
.A(n_4826),
.B(n_4279),
.Y(n_5576)
);

NAND2xp5_ASAP7_75t_L g5577 ( 
.A(n_4826),
.B(n_4835),
.Y(n_5577)
);

NOR2xp33_ASAP7_75t_L g5578 ( 
.A(n_4805),
.B(n_4138),
.Y(n_5578)
);

BUFx6f_ASAP7_75t_L g5579 ( 
.A(n_4388),
.Y(n_5579)
);

OAI22x1_ASAP7_75t_L g5580 ( 
.A1(n_4667),
.A2(n_3950),
.B1(n_4049),
.B2(n_3919),
.Y(n_5580)
);

INVx1_ASAP7_75t_L g5581 ( 
.A(n_4782),
.Y(n_5581)
);

AOI21xp5_ASAP7_75t_SL g5582 ( 
.A1(n_5017),
.A2(n_3620),
.B(n_3530),
.Y(n_5582)
);

BUFx2_ASAP7_75t_L g5583 ( 
.A(n_4990),
.Y(n_5583)
);

A2O1A1Ixp33_ASAP7_75t_L g5584 ( 
.A1(n_4611),
.A2(n_3727),
.B(n_3728),
.C(n_3704),
.Y(n_5584)
);

INVx2_ASAP7_75t_L g5585 ( 
.A(n_4614),
.Y(n_5585)
);

NOR2x1_ASAP7_75t_SL g5586 ( 
.A(n_4735),
.B(n_4235),
.Y(n_5586)
);

A2O1A1Ixp33_ASAP7_75t_L g5587 ( 
.A1(n_4916),
.A2(n_3727),
.B(n_3728),
.C(n_3704),
.Y(n_5587)
);

CKINVDCx5p33_ASAP7_75t_R g5588 ( 
.A(n_5044),
.Y(n_5588)
);

AOI21xp5_ASAP7_75t_L g5589 ( 
.A1(n_4793),
.A2(n_4173),
.B(n_4167),
.Y(n_5589)
);

NOR2xp67_ASAP7_75t_L g5590 ( 
.A(n_4735),
.B(n_4269),
.Y(n_5590)
);

OAI21xp5_ASAP7_75t_L g5591 ( 
.A1(n_4876),
.A2(n_3526),
.B(n_3664),
.Y(n_5591)
);

AOI21xp5_ASAP7_75t_L g5592 ( 
.A1(n_4799),
.A2(n_4173),
.B(n_4167),
.Y(n_5592)
);

AO31x2_ASAP7_75t_L g5593 ( 
.A1(n_4842),
.A2(n_3923),
.A3(n_3946),
.B(n_3921),
.Y(n_5593)
);

AOI21xp5_ASAP7_75t_L g5594 ( 
.A1(n_4799),
.A2(n_3735),
.B(n_3732),
.Y(n_5594)
);

INVx1_ASAP7_75t_SL g5595 ( 
.A(n_4432),
.Y(n_5595)
);

AOI221x1_ASAP7_75t_L g5596 ( 
.A1(n_4493),
.A2(n_3963),
.B1(n_3964),
.B2(n_3946),
.C(n_3923),
.Y(n_5596)
);

AND2x4_ASAP7_75t_L g5597 ( 
.A(n_4642),
.B(n_4235),
.Y(n_5597)
);

BUFx6f_ASAP7_75t_L g5598 ( 
.A(n_4388),
.Y(n_5598)
);

INVx1_ASAP7_75t_L g5599 ( 
.A(n_4782),
.Y(n_5599)
);

AOI21xp5_ASAP7_75t_L g5600 ( 
.A1(n_4800),
.A2(n_3735),
.B(n_3732),
.Y(n_5600)
);

INVx1_ASAP7_75t_L g5601 ( 
.A(n_4788),
.Y(n_5601)
);

INVx2_ASAP7_75t_SL g5602 ( 
.A(n_5127),
.Y(n_5602)
);

OAI21xp5_ASAP7_75t_L g5603 ( 
.A1(n_4813),
.A2(n_3526),
.B(n_3664),
.Y(n_5603)
);

INVx3_ASAP7_75t_L g5604 ( 
.A(n_5142),
.Y(n_5604)
);

AND2x2_ASAP7_75t_L g5605 ( 
.A(n_4742),
.B(n_4235),
.Y(n_5605)
);

INVx3_ASAP7_75t_SL g5606 ( 
.A(n_5127),
.Y(n_5606)
);

BUFx12f_ASAP7_75t_L g5607 ( 
.A(n_5044),
.Y(n_5607)
);

BUFx2_ASAP7_75t_L g5608 ( 
.A(n_5025),
.Y(n_5608)
);

NAND2xp5_ASAP7_75t_SL g5609 ( 
.A(n_4379),
.B(n_3676),
.Y(n_5609)
);

NAND2xp5_ASAP7_75t_SL g5610 ( 
.A(n_4379),
.B(n_4049),
.Y(n_5610)
);

INVxp67_ASAP7_75t_L g5611 ( 
.A(n_5063),
.Y(n_5611)
);

AND2x2_ASAP7_75t_L g5612 ( 
.A(n_4742),
.B(n_4049),
.Y(n_5612)
);

OAI21x1_ASAP7_75t_L g5613 ( 
.A1(n_4925),
.A2(n_4356),
.B(n_4339),
.Y(n_5613)
);

NAND2x1p5_ASAP7_75t_L g5614 ( 
.A(n_5040),
.B(n_4817),
.Y(n_5614)
);

INVx2_ASAP7_75t_L g5615 ( 
.A(n_4614),
.Y(n_5615)
);

OAI21x1_ASAP7_75t_L g5616 ( 
.A1(n_4925),
.A2(n_4356),
.B(n_3751),
.Y(n_5616)
);

INVx3_ASAP7_75t_SL g5617 ( 
.A(n_5127),
.Y(n_5617)
);

BUFx3_ASAP7_75t_L g5618 ( 
.A(n_5025),
.Y(n_5618)
);

OAI22xp5_ASAP7_75t_L g5619 ( 
.A1(n_5113),
.A2(n_4061),
.B1(n_4067),
.B2(n_4043),
.Y(n_5619)
);

INVxp67_ASAP7_75t_SL g5620 ( 
.A(n_4670),
.Y(n_5620)
);

OAI21x1_ASAP7_75t_L g5621 ( 
.A1(n_4925),
.A2(n_4356),
.B(n_3751),
.Y(n_5621)
);

O2A1O1Ixp33_ASAP7_75t_SL g5622 ( 
.A1(n_4424),
.A2(n_4067),
.B(n_4070),
.C(n_4069),
.Y(n_5622)
);

AOI21xp5_ASAP7_75t_L g5623 ( 
.A1(n_4800),
.A2(n_3769),
.B(n_3747),
.Y(n_5623)
);

AOI21xp5_ASAP7_75t_L g5624 ( 
.A1(n_4929),
.A2(n_3769),
.B(n_3747),
.Y(n_5624)
);

AND2x2_ASAP7_75t_L g5625 ( 
.A(n_4385),
.B(n_4049),
.Y(n_5625)
);

NAND3xp33_ASAP7_75t_SL g5626 ( 
.A(n_4768),
.B(n_4070),
.C(n_4069),
.Y(n_5626)
);

AOI21xp5_ASAP7_75t_L g5627 ( 
.A1(n_5017),
.A2(n_3775),
.B(n_3772),
.Y(n_5627)
);

NAND2xp5_ASAP7_75t_L g5628 ( 
.A(n_4836),
.B(n_4839),
.Y(n_5628)
);

CKINVDCx20_ASAP7_75t_R g5629 ( 
.A(n_4720),
.Y(n_5629)
);

INVx1_ASAP7_75t_L g5630 ( 
.A(n_4788),
.Y(n_5630)
);

OAI21xp5_ASAP7_75t_L g5631 ( 
.A1(n_4813),
.A2(n_4823),
.B(n_4577),
.Y(n_5631)
);

OAI21x1_ASAP7_75t_L g5632 ( 
.A1(n_4445),
.A2(n_3775),
.B(n_3772),
.Y(n_5632)
);

HB1xp67_ASAP7_75t_L g5633 ( 
.A(n_4610),
.Y(n_5633)
);

INVx2_ASAP7_75t_L g5634 ( 
.A(n_4618),
.Y(n_5634)
);

AOI21xp5_ASAP7_75t_L g5635 ( 
.A1(n_5019),
.A2(n_3794),
.B(n_3777),
.Y(n_5635)
);

OAI22xp5_ASAP7_75t_L g5636 ( 
.A1(n_4468),
.A2(n_4087),
.B1(n_4095),
.B2(n_4082),
.Y(n_5636)
);

AO21x2_ASAP7_75t_L g5637 ( 
.A1(n_4419),
.A2(n_3794),
.B(n_3777),
.Y(n_5637)
);

NAND2xp5_ASAP7_75t_L g5638 ( 
.A(n_4839),
.B(n_4841),
.Y(n_5638)
);

A2O1A1Ixp33_ASAP7_75t_L g5639 ( 
.A1(n_4846),
.A2(n_3727),
.B(n_3728),
.C(n_3704),
.Y(n_5639)
);

O2A1O1Ixp33_ASAP7_75t_L g5640 ( 
.A1(n_4566),
.A2(n_4087),
.B(n_4095),
.C(n_4082),
.Y(n_5640)
);

AOI21xp5_ASAP7_75t_L g5641 ( 
.A1(n_5019),
.A2(n_4307),
.B(n_4289),
.Y(n_5641)
);

NAND2xp33_ASAP7_75t_SL g5642 ( 
.A(n_4768),
.B(n_3003),
.Y(n_5642)
);

INVx3_ASAP7_75t_L g5643 ( 
.A(n_5142),
.Y(n_5643)
);

OAI21x1_ASAP7_75t_L g5644 ( 
.A1(n_4445),
.A2(n_4332),
.B(n_3707),
.Y(n_5644)
);

AOI21xp5_ASAP7_75t_SL g5645 ( 
.A1(n_4575),
.A2(n_4108),
.B(n_3911),
.Y(n_5645)
);

BUFx8_ASAP7_75t_L g5646 ( 
.A(n_4850),
.Y(n_5646)
);

OAI21xp5_ASAP7_75t_L g5647 ( 
.A1(n_4823),
.A2(n_4828),
.B(n_4400),
.Y(n_5647)
);

NAND2xp5_ASAP7_75t_L g5648 ( 
.A(n_5084),
.B(n_3486),
.Y(n_5648)
);

BUFx2_ASAP7_75t_L g5649 ( 
.A(n_5025),
.Y(n_5649)
);

OAI21xp5_ASAP7_75t_L g5650 ( 
.A1(n_4828),
.A2(n_3669),
.B(n_3694),
.Y(n_5650)
);

AOI21xp5_ASAP7_75t_L g5651 ( 
.A1(n_4559),
.A2(n_4307),
.B(n_4316),
.Y(n_5651)
);

O2A1O1Ixp33_ASAP7_75t_SL g5652 ( 
.A1(n_4575),
.A2(n_4303),
.B(n_3496),
.C(n_3674),
.Y(n_5652)
);

INVx1_ASAP7_75t_L g5653 ( 
.A(n_4808),
.Y(n_5653)
);

CKINVDCx5p33_ASAP7_75t_R g5654 ( 
.A(n_4465),
.Y(n_5654)
);

AOI21xp5_ASAP7_75t_L g5655 ( 
.A1(n_4494),
.A2(n_4220),
.B(n_4332),
.Y(n_5655)
);

AOI221x1_ASAP7_75t_L g5656 ( 
.A1(n_5122),
.A2(n_4454),
.B1(n_4511),
.B2(n_4666),
.C(n_4414),
.Y(n_5656)
);

INVx1_ASAP7_75t_L g5657 ( 
.A(n_4808),
.Y(n_5657)
);

OAI21x1_ASAP7_75t_L g5658 ( 
.A1(n_4832),
.A2(n_3707),
.B(n_3694),
.Y(n_5658)
);

OAI21x1_ASAP7_75t_L g5659 ( 
.A1(n_4832),
.A2(n_3669),
.B(n_4175),
.Y(n_5659)
);

NAND2xp5_ASAP7_75t_L g5660 ( 
.A(n_5084),
.B(n_3521),
.Y(n_5660)
);

AOI21xp5_ASAP7_75t_L g5661 ( 
.A1(n_4494),
.A2(n_4220),
.B(n_4289),
.Y(n_5661)
);

BUFx8_ASAP7_75t_L g5662 ( 
.A(n_4850),
.Y(n_5662)
);

AOI21xp5_ASAP7_75t_L g5663 ( 
.A1(n_4499),
.A2(n_4220),
.B(n_4197),
.Y(n_5663)
);

NAND3xp33_ASAP7_75t_L g5664 ( 
.A(n_4463),
.B(n_4571),
.C(n_4652),
.Y(n_5664)
);

NOR2xp33_ASAP7_75t_L g5665 ( 
.A(n_4624),
.B(n_4138),
.Y(n_5665)
);

AOI22xp33_ASAP7_75t_L g5666 ( 
.A1(n_4400),
.A2(n_4050),
.B1(n_3718),
.B2(n_3876),
.Y(n_5666)
);

INVx1_ASAP7_75t_L g5667 ( 
.A(n_4810),
.Y(n_5667)
);

AND2x2_ASAP7_75t_L g5668 ( 
.A(n_4385),
.B(n_4050),
.Y(n_5668)
);

NAND3x1_ASAP7_75t_L g5669 ( 
.A(n_4821),
.B(n_3674),
.C(n_4176),
.Y(n_5669)
);

AOI22xp5_ASAP7_75t_L g5670 ( 
.A1(n_4571),
.A2(n_3718),
.B1(n_3876),
.B2(n_3815),
.Y(n_5670)
);

INVx1_ASAP7_75t_L g5671 ( 
.A(n_4810),
.Y(n_5671)
);

INVx1_ASAP7_75t_L g5672 ( 
.A(n_4819),
.Y(n_5672)
);

INVx1_ASAP7_75t_L g5673 ( 
.A(n_4819),
.Y(n_5673)
);

OAI22xp5_ASAP7_75t_L g5674 ( 
.A1(n_4957),
.A2(n_3823),
.B1(n_3811),
.B2(n_4157),
.Y(n_5674)
);

OAI21x1_ASAP7_75t_L g5675 ( 
.A1(n_4832),
.A2(n_4345),
.B(n_4334),
.Y(n_5675)
);

OAI21x1_ASAP7_75t_L g5676 ( 
.A1(n_4678),
.A2(n_4345),
.B(n_4334),
.Y(n_5676)
);

AOI21xp5_ASAP7_75t_L g5677 ( 
.A1(n_4443),
.A2(n_4296),
.B(n_4197),
.Y(n_5677)
);

NAND2xp33_ASAP7_75t_SL g5678 ( 
.A(n_4768),
.B(n_3003),
.Y(n_5678)
);

INVx2_ASAP7_75t_L g5679 ( 
.A(n_4618),
.Y(n_5679)
);

INVx1_ASAP7_75t_L g5680 ( 
.A(n_4838),
.Y(n_5680)
);

AOI22xp5_ASAP7_75t_L g5681 ( 
.A1(n_4713),
.A2(n_3718),
.B1(n_3876),
.B2(n_2980),
.Y(n_5681)
);

O2A1O1Ixp5_ASAP7_75t_L g5682 ( 
.A1(n_4884),
.A2(n_4941),
.B(n_4911),
.C(n_5087),
.Y(n_5682)
);

CKINVDCx11_ASAP7_75t_R g5683 ( 
.A(n_4555),
.Y(n_5683)
);

OR2x6_ASAP7_75t_L g5684 ( 
.A(n_5039),
.B(n_3718),
.Y(n_5684)
);

BUFx6f_ASAP7_75t_L g5685 ( 
.A(n_4388),
.Y(n_5685)
);

AOI21xp5_ASAP7_75t_L g5686 ( 
.A1(n_4443),
.A2(n_4296),
.B(n_4204),
.Y(n_5686)
);

NAND2xp5_ASAP7_75t_L g5687 ( 
.A(n_5057),
.B(n_3521),
.Y(n_5687)
);

OAI21x1_ASAP7_75t_L g5688 ( 
.A1(n_4678),
.A2(n_4351),
.B(n_4348),
.Y(n_5688)
);

BUFx2_ASAP7_75t_R g5689 ( 
.A(n_4464),
.Y(n_5689)
);

O2A1O1Ixp33_ASAP7_75t_SL g5690 ( 
.A1(n_4601),
.A2(n_3496),
.B(n_3970),
.C(n_3968),
.Y(n_5690)
);

OR2x2_ASAP7_75t_L g5691 ( 
.A(n_4480),
.B(n_3864),
.Y(n_5691)
);

NAND2xp5_ASAP7_75t_L g5692 ( 
.A(n_5057),
.B(n_3539),
.Y(n_5692)
);

INVx1_ASAP7_75t_L g5693 ( 
.A(n_4838),
.Y(n_5693)
);

AO22x2_ASAP7_75t_L g5694 ( 
.A1(n_4768),
.A2(n_4050),
.B1(n_3979),
.B2(n_3986),
.Y(n_5694)
);

AOI21xp5_ASAP7_75t_L g5695 ( 
.A1(n_4511),
.A2(n_4204),
.B(n_4192),
.Y(n_5695)
);

A2O1A1Ixp33_ASAP7_75t_L g5696 ( 
.A1(n_4899),
.A2(n_4108),
.B(n_4127),
.C(n_3911),
.Y(n_5696)
);

BUFx2_ASAP7_75t_L g5697 ( 
.A(n_5070),
.Y(n_5697)
);

AOI21xp5_ASAP7_75t_L g5698 ( 
.A1(n_4645),
.A2(n_4208),
.B(n_4192),
.Y(n_5698)
);

HB1xp67_ASAP7_75t_L g5699 ( 
.A(n_4610),
.Y(n_5699)
);

AOI21xp5_ASAP7_75t_L g5700 ( 
.A1(n_4645),
.A2(n_4209),
.B(n_4208),
.Y(n_5700)
);

INVx1_ASAP7_75t_SL g5701 ( 
.A(n_4465),
.Y(n_5701)
);

AOI21xp5_ASAP7_75t_L g5702 ( 
.A1(n_4650),
.A2(n_4210),
.B(n_4209),
.Y(n_5702)
);

INVx2_ASAP7_75t_L g5703 ( 
.A(n_4618),
.Y(n_5703)
);

INVxp67_ASAP7_75t_L g5704 ( 
.A(n_5063),
.Y(n_5704)
);

OAI22xp5_ASAP7_75t_L g5705 ( 
.A1(n_4957),
.A2(n_4157),
.B1(n_4096),
.B2(n_3608),
.Y(n_5705)
);

INVx4_ASAP7_75t_SL g5706 ( 
.A(n_5099),
.Y(n_5706)
);

BUFx2_ASAP7_75t_L g5707 ( 
.A(n_5070),
.Y(n_5707)
);

NOR2xp33_ASAP7_75t_L g5708 ( 
.A(n_4624),
.B(n_4138),
.Y(n_5708)
);

INVx1_ASAP7_75t_L g5709 ( 
.A(n_4858),
.Y(n_5709)
);

NOR2xp67_ASAP7_75t_L g5710 ( 
.A(n_4971),
.B(n_5059),
.Y(n_5710)
);

NAND3xp33_ASAP7_75t_L g5711 ( 
.A(n_4463),
.B(n_3608),
.C(n_3476),
.Y(n_5711)
);

AOI21xp5_ASAP7_75t_L g5712 ( 
.A1(n_4650),
.A2(n_4210),
.B(n_4348),
.Y(n_5712)
);

AOI21xp5_ASAP7_75t_L g5713 ( 
.A1(n_4499),
.A2(n_4353),
.B(n_4351),
.Y(n_5713)
);

AOI21xp5_ASAP7_75t_L g5714 ( 
.A1(n_4500),
.A2(n_4363),
.B(n_4353),
.Y(n_5714)
);

OAI22xp33_ASAP7_75t_L g5715 ( 
.A1(n_4408),
.A2(n_3750),
.B1(n_3758),
.B2(n_3715),
.Y(n_5715)
);

AOI21xp5_ASAP7_75t_L g5716 ( 
.A1(n_4500),
.A2(n_4363),
.B(n_4191),
.Y(n_5716)
);

INVx1_ASAP7_75t_L g5717 ( 
.A(n_4858),
.Y(n_5717)
);

OA21x2_ASAP7_75t_L g5718 ( 
.A1(n_4502),
.A2(n_3992),
.B(n_3989),
.Y(n_5718)
);

AOI21xp5_ASAP7_75t_L g5719 ( 
.A1(n_4502),
.A2(n_4191),
.B(n_4228),
.Y(n_5719)
);

AOI221xp5_ASAP7_75t_L g5720 ( 
.A1(n_4719),
.A2(n_3998),
.B1(n_3999),
.B2(n_3527),
.C(n_4011),
.Y(n_5720)
);

AO21x2_ASAP7_75t_L g5721 ( 
.A1(n_4419),
.A2(n_4582),
.B(n_4530),
.Y(n_5721)
);

OAI22xp5_ASAP7_75t_L g5722 ( 
.A1(n_4957),
.A2(n_4096),
.B1(n_4285),
.B2(n_3476),
.Y(n_5722)
);

BUFx6f_ASAP7_75t_L g5723 ( 
.A(n_4388),
.Y(n_5723)
);

OR2x2_ASAP7_75t_L g5724 ( 
.A(n_4480),
.B(n_4055),
.Y(n_5724)
);

A2O1A1Ixp33_ASAP7_75t_L g5725 ( 
.A1(n_4899),
.A2(n_4108),
.B(n_4127),
.C(n_3911),
.Y(n_5725)
);

AOI21xp5_ASAP7_75t_L g5726 ( 
.A1(n_4505),
.A2(n_3167),
.B(n_3390),
.Y(n_5726)
);

INVx2_ASAP7_75t_SL g5727 ( 
.A(n_4637),
.Y(n_5727)
);

AND2x2_ASAP7_75t_L g5728 ( 
.A(n_4385),
.B(n_4050),
.Y(n_5728)
);

NOR2xp33_ASAP7_75t_L g5729 ( 
.A(n_4630),
.B(n_4154),
.Y(n_5729)
);

INVx1_ASAP7_75t_L g5730 ( 
.A(n_4862),
.Y(n_5730)
);

A2O1A1Ixp33_ASAP7_75t_L g5731 ( 
.A1(n_4608),
.A2(n_4179),
.B(n_4236),
.C(n_4127),
.Y(n_5731)
);

OAI21x1_ASAP7_75t_L g5732 ( 
.A1(n_4678),
.A2(n_4071),
.B(n_4014),
.Y(n_5732)
);

AOI21xp5_ASAP7_75t_L g5733 ( 
.A1(n_4505),
.A2(n_3167),
.B(n_3390),
.Y(n_5733)
);

BUFx2_ASAP7_75t_L g5734 ( 
.A(n_5070),
.Y(n_5734)
);

INVx3_ASAP7_75t_L g5735 ( 
.A(n_5142),
.Y(n_5735)
);

AO21x1_ASAP7_75t_L g5736 ( 
.A1(n_4582),
.A2(n_4088),
.B(n_4071),
.Y(n_5736)
);

NAND2xp33_ASAP7_75t_L g5737 ( 
.A(n_4469),
.B(n_2980),
.Y(n_5737)
);

NOR4xp25_ASAP7_75t_L g5738 ( 
.A(n_4852),
.B(n_4088),
.C(n_4163),
.D(n_4136),
.Y(n_5738)
);

INVx1_ASAP7_75t_L g5739 ( 
.A(n_4862),
.Y(n_5739)
);

AOI21xp5_ASAP7_75t_L g5740 ( 
.A1(n_4506),
.A2(n_3167),
.B(n_3390),
.Y(n_5740)
);

INVx5_ASAP7_75t_SL g5741 ( 
.A(n_4527),
.Y(n_5741)
);

AOI21xp5_ASAP7_75t_L g5742 ( 
.A1(n_4629),
.A2(n_4641),
.B(n_4634),
.Y(n_5742)
);

AOI21xp5_ASAP7_75t_L g5743 ( 
.A1(n_4634),
.A2(n_4641),
.B(n_5039),
.Y(n_5743)
);

NAND2xp5_ASAP7_75t_L g5744 ( 
.A(n_4633),
.B(n_3545),
.Y(n_5744)
);

BUFx3_ASAP7_75t_L g5745 ( 
.A(n_5079),
.Y(n_5745)
);

INVx1_ASAP7_75t_L g5746 ( 
.A(n_4875),
.Y(n_5746)
);

INVx1_ASAP7_75t_L g5747 ( 
.A(n_4875),
.Y(n_5747)
);

INVx2_ASAP7_75t_L g5748 ( 
.A(n_4638),
.Y(n_5748)
);

AOI21xp33_ASAP7_75t_L g5749 ( 
.A1(n_4852),
.A2(n_4185),
.B(n_4184),
.Y(n_5749)
);

AOI22xp5_ASAP7_75t_L g5750 ( 
.A1(n_4713),
.A2(n_3876),
.B1(n_2980),
.B2(n_2862),
.Y(n_5750)
);

A2O1A1Ixp33_ASAP7_75t_L g5751 ( 
.A1(n_4408),
.A2(n_4236),
.B(n_4324),
.C(n_4179),
.Y(n_5751)
);

OAI21xp5_ASAP7_75t_L g5752 ( 
.A1(n_4770),
.A2(n_3363),
.B(n_3357),
.Y(n_5752)
);

BUFx2_ASAP7_75t_L g5753 ( 
.A(n_5079),
.Y(n_5753)
);

AOI22xp5_ASAP7_75t_L g5754 ( 
.A1(n_4893),
.A2(n_3876),
.B1(n_2980),
.B2(n_2862),
.Y(n_5754)
);

NAND2xp5_ASAP7_75t_L g5755 ( 
.A(n_4633),
.B(n_3611),
.Y(n_5755)
);

NOR2x1_ASAP7_75t_L g5756 ( 
.A(n_4404),
.B(n_4584),
.Y(n_5756)
);

A2O1A1Ixp33_ASAP7_75t_L g5757 ( 
.A1(n_4668),
.A2(n_4236),
.B(n_4324),
.C(n_4179),
.Y(n_5757)
);

OR2x2_ASAP7_75t_L g5758 ( 
.A(n_4540),
.B(n_4285),
.Y(n_5758)
);

A2O1A1Ixp33_ASAP7_75t_L g5759 ( 
.A1(n_4668),
.A2(n_4324),
.B(n_2862),
.C(n_2885),
.Y(n_5759)
);

INVx5_ASAP7_75t_L g5760 ( 
.A(n_4971),
.Y(n_5760)
);

AND2x4_ASAP7_75t_L g5761 ( 
.A(n_4642),
.B(n_3715),
.Y(n_5761)
);

A2O1A1Ixp33_ASAP7_75t_L g5762 ( 
.A1(n_5002),
.A2(n_2885),
.B(n_2913),
.C(n_2836),
.Y(n_5762)
);

AO22x2_ASAP7_75t_L g5763 ( 
.A1(n_5122),
.A2(n_4185),
.B1(n_4190),
.B2(n_4184),
.Y(n_5763)
);

BUFx6f_ASAP7_75t_L g5764 ( 
.A(n_4496),
.Y(n_5764)
);

NAND2xp5_ASAP7_75t_L g5765 ( 
.A(n_4778),
.B(n_3611),
.Y(n_5765)
);

AOI21xp5_ASAP7_75t_L g5766 ( 
.A1(n_5002),
.A2(n_3167),
.B(n_3395),
.Y(n_5766)
);

NAND2xp5_ASAP7_75t_SL g5767 ( 
.A(n_4759),
.B(n_3527),
.Y(n_5767)
);

INVx3_ASAP7_75t_L g5768 ( 
.A(n_5142),
.Y(n_5768)
);

AOI21xp5_ASAP7_75t_L g5769 ( 
.A1(n_4380),
.A2(n_4382),
.B(n_4434),
.Y(n_5769)
);

CKINVDCx11_ASAP7_75t_R g5770 ( 
.A(n_4555),
.Y(n_5770)
);

AOI221x1_ASAP7_75t_L g5771 ( 
.A1(n_4454),
.A2(n_4207),
.B1(n_4206),
.B2(n_3691),
.C(n_3705),
.Y(n_5771)
);

AOI21xp5_ASAP7_75t_L g5772 ( 
.A1(n_4382),
.A2(n_3395),
.B(n_3715),
.Y(n_5772)
);

OAI21xp5_ASAP7_75t_L g5773 ( 
.A1(n_4472),
.A2(n_3363),
.B(n_3357),
.Y(n_5773)
);

NOR2xp33_ASAP7_75t_L g5774 ( 
.A(n_4630),
.B(n_4154),
.Y(n_5774)
);

AOI21xp5_ASAP7_75t_L g5775 ( 
.A1(n_4434),
.A2(n_4452),
.B(n_4414),
.Y(n_5775)
);

CKINVDCx5p33_ASAP7_75t_R g5776 ( 
.A(n_4778),
.Y(n_5776)
);

AOI21xp5_ASAP7_75t_L g5777 ( 
.A1(n_4452),
.A2(n_4837),
.B(n_4389),
.Y(n_5777)
);

O2A1O1Ixp33_ASAP7_75t_L g5778 ( 
.A1(n_4863),
.A2(n_4341),
.B(n_3402),
.C(n_3415),
.Y(n_5778)
);

O2A1O1Ixp33_ASAP7_75t_L g5779 ( 
.A1(n_4843),
.A2(n_4341),
.B(n_3415),
.C(n_3399),
.Y(n_5779)
);

AOI22xp5_ASAP7_75t_L g5780 ( 
.A1(n_4893),
.A2(n_2980),
.B1(n_2913),
.B2(n_2922),
.Y(n_5780)
);

OAI22xp5_ASAP7_75t_L g5781 ( 
.A1(n_4528),
.A2(n_4258),
.B1(n_4265),
.B2(n_4260),
.Y(n_5781)
);

AOI21xp5_ASAP7_75t_L g5782 ( 
.A1(n_4837),
.A2(n_4391),
.B(n_4389),
.Y(n_5782)
);

NOR2xp33_ASAP7_75t_SL g5783 ( 
.A(n_4462),
.B(n_2859),
.Y(n_5783)
);

AOI21xp5_ASAP7_75t_L g5784 ( 
.A1(n_4391),
.A2(n_3395),
.B(n_3715),
.Y(n_5784)
);

A2O1A1Ixp33_ASAP7_75t_L g5785 ( 
.A1(n_4940),
.A2(n_2913),
.B(n_2922),
.C(n_2885),
.Y(n_5785)
);

INVx2_ASAP7_75t_L g5786 ( 
.A(n_4638),
.Y(n_5786)
);

NAND2xp5_ASAP7_75t_L g5787 ( 
.A(n_4982),
.B(n_3614),
.Y(n_5787)
);

INVx1_ASAP7_75t_L g5788 ( 
.A(n_4885),
.Y(n_5788)
);

BUFx2_ASAP7_75t_L g5789 ( 
.A(n_5079),
.Y(n_5789)
);

AOI21xp5_ASAP7_75t_L g5790 ( 
.A1(n_4573),
.A2(n_3442),
.B(n_2915),
.Y(n_5790)
);

AOI21xp5_ASAP7_75t_L g5791 ( 
.A1(n_4573),
.A2(n_3442),
.B(n_2915),
.Y(n_5791)
);

A2O1A1Ixp33_ASAP7_75t_L g5792 ( 
.A1(n_4940),
.A2(n_2913),
.B(n_2922),
.C(n_2885),
.Y(n_5792)
);

INVx1_ASAP7_75t_L g5793 ( 
.A(n_4885),
.Y(n_5793)
);

O2A1O1Ixp33_ASAP7_75t_SL g5794 ( 
.A1(n_4601),
.A2(n_4207),
.B(n_4154),
.C(n_4258),
.Y(n_5794)
);

AOI21xp5_ASAP7_75t_L g5795 ( 
.A1(n_4387),
.A2(n_2915),
.B(n_2859),
.Y(n_5795)
);

NOR2xp33_ASAP7_75t_L g5796 ( 
.A(n_4632),
.B(n_2885),
.Y(n_5796)
);

A2O1A1Ixp33_ASAP7_75t_L g5797 ( 
.A1(n_4666),
.A2(n_4653),
.B(n_4656),
.C(n_4478),
.Y(n_5797)
);

AOI21xp5_ASAP7_75t_L g5798 ( 
.A1(n_4387),
.A2(n_2915),
.B(n_2859),
.Y(n_5798)
);

OA21x2_ASAP7_75t_L g5799 ( 
.A1(n_4628),
.A2(n_3673),
.B(n_3614),
.Y(n_5799)
);

NAND2xp5_ASAP7_75t_SL g5800 ( 
.A(n_4759),
.B(n_3433),
.Y(n_5800)
);

BUFx3_ASAP7_75t_L g5801 ( 
.A(n_5094),
.Y(n_5801)
);

INVx2_ASAP7_75t_SL g5802 ( 
.A(n_4637),
.Y(n_5802)
);

BUFx2_ASAP7_75t_L g5803 ( 
.A(n_5094),
.Y(n_5803)
);

AOI21xp5_ASAP7_75t_L g5804 ( 
.A1(n_4649),
.A2(n_2927),
.B(n_2859),
.Y(n_5804)
);

INVx2_ASAP7_75t_SL g5805 ( 
.A(n_5094),
.Y(n_5805)
);

AO31x2_ASAP7_75t_L g5806 ( 
.A1(n_5077),
.A2(n_3691),
.A3(n_3705),
.B(n_3673),
.Y(n_5806)
);

NAND2xp33_ASAP7_75t_SL g5807 ( 
.A(n_4961),
.B(n_3003),
.Y(n_5807)
);

AOI21xp5_ASAP7_75t_L g5808 ( 
.A1(n_4649),
.A2(n_2943),
.B(n_2927),
.Y(n_5808)
);

AOI21xp5_ASAP7_75t_L g5809 ( 
.A1(n_4623),
.A2(n_2943),
.B(n_2927),
.Y(n_5809)
);

NAND2xp5_ASAP7_75t_L g5810 ( 
.A(n_4982),
.B(n_3799),
.Y(n_5810)
);

BUFx10_ASAP7_75t_L g5811 ( 
.A(n_5099),
.Y(n_5811)
);

OAI21x1_ASAP7_75t_L g5812 ( 
.A1(n_4399),
.A2(n_4411),
.B(n_4405),
.Y(n_5812)
);

O2A1O1Ixp33_ASAP7_75t_SL g5813 ( 
.A1(n_5011),
.A2(n_4265),
.B(n_4260),
.C(n_4007),
.Y(n_5813)
);

INVx1_ASAP7_75t_L g5814 ( 
.A(n_4898),
.Y(n_5814)
);

O2A1O1Ixp33_ASAP7_75t_L g5815 ( 
.A1(n_4843),
.A2(n_4341),
.B(n_3415),
.C(n_3399),
.Y(n_5815)
);

A2O1A1Ixp33_ASAP7_75t_L g5816 ( 
.A1(n_4653),
.A2(n_2913),
.B(n_2922),
.C(n_2885),
.Y(n_5816)
);

AO31x2_ASAP7_75t_L g5817 ( 
.A1(n_5077),
.A2(n_3514),
.A3(n_3538),
.B(n_3500),
.Y(n_5817)
);

AOI21xp5_ASAP7_75t_L g5818 ( 
.A1(n_4623),
.A2(n_2943),
.B(n_2927),
.Y(n_5818)
);

OAI21x1_ASAP7_75t_SL g5819 ( 
.A1(n_5135),
.A2(n_3219),
.B(n_3203),
.Y(n_5819)
);

A2O1A1Ixp33_ASAP7_75t_L g5820 ( 
.A1(n_4656),
.A2(n_2913),
.B(n_2922),
.C(n_2885),
.Y(n_5820)
);

NOR2x1_ASAP7_75t_R g5821 ( 
.A(n_4720),
.B(n_2876),
.Y(n_5821)
);

OA21x2_ASAP7_75t_L g5822 ( 
.A1(n_4628),
.A2(n_3514),
.B(n_3500),
.Y(n_5822)
);

OAI21xp5_ASAP7_75t_L g5823 ( 
.A1(n_4472),
.A2(n_3363),
.B(n_3357),
.Y(n_5823)
);

INVx2_ASAP7_75t_SL g5824 ( 
.A(n_5116),
.Y(n_5824)
);

INVx1_ASAP7_75t_L g5825 ( 
.A(n_4898),
.Y(n_5825)
);

AOI21xp5_ASAP7_75t_L g5826 ( 
.A1(n_4865),
.A2(n_3750),
.B(n_3715),
.Y(n_5826)
);

AOI21xp5_ASAP7_75t_L g5827 ( 
.A1(n_4865),
.A2(n_3758),
.B(n_3750),
.Y(n_5827)
);

NOR2xp33_ASAP7_75t_SL g5828 ( 
.A(n_4462),
.B(n_2927),
.Y(n_5828)
);

OAI21x1_ASAP7_75t_L g5829 ( 
.A1(n_4399),
.A2(n_3538),
.B(n_3514),
.Y(n_5829)
);

O2A1O1Ixp33_ASAP7_75t_L g5830 ( 
.A1(n_4478),
.A2(n_3415),
.B(n_3399),
.C(n_3363),
.Y(n_5830)
);

INVx2_ASAP7_75t_L g5831 ( 
.A(n_4638),
.Y(n_5831)
);

INVxp67_ASAP7_75t_L g5832 ( 
.A(n_5043),
.Y(n_5832)
);

INVx1_ASAP7_75t_L g5833 ( 
.A(n_4930),
.Y(n_5833)
);

BUFx12f_ASAP7_75t_L g5834 ( 
.A(n_4604),
.Y(n_5834)
);

OAI22xp5_ASAP7_75t_L g5835 ( 
.A1(n_4528),
.A2(n_4040),
.B1(n_4011),
.B2(n_3999),
.Y(n_5835)
);

INVx1_ASAP7_75t_L g5836 ( 
.A(n_4930),
.Y(n_5836)
);

INVx5_ASAP7_75t_L g5837 ( 
.A(n_4971),
.Y(n_5837)
);

NAND2xp5_ASAP7_75t_L g5838 ( 
.A(n_5106),
.B(n_3799),
.Y(n_5838)
);

BUFx6f_ASAP7_75t_L g5839 ( 
.A(n_4496),
.Y(n_5839)
);

NAND2xp5_ASAP7_75t_L g5840 ( 
.A(n_5106),
.B(n_3726),
.Y(n_5840)
);

AOI21x1_ASAP7_75t_L g5841 ( 
.A1(n_4910),
.A2(n_3219),
.B(n_3538),
.Y(n_5841)
);

OAI21x1_ASAP7_75t_L g5842 ( 
.A1(n_4399),
.A2(n_3561),
.B(n_3559),
.Y(n_5842)
);

AOI21x1_ASAP7_75t_L g5843 ( 
.A1(n_4910),
.A2(n_3219),
.B(n_3559),
.Y(n_5843)
);

CKINVDCx5p33_ASAP7_75t_R g5844 ( 
.A(n_5075),
.Y(n_5844)
);

AOI21xp5_ASAP7_75t_L g5845 ( 
.A1(n_4874),
.A2(n_2943),
.B(n_2927),
.Y(n_5845)
);

INVx3_ASAP7_75t_L g5846 ( 
.A(n_5142),
.Y(n_5846)
);

CKINVDCx5p33_ASAP7_75t_R g5847 ( 
.A(n_5075),
.Y(n_5847)
);

O2A1O1Ixp33_ASAP7_75t_L g5848 ( 
.A1(n_4918),
.A2(n_3399),
.B(n_2908),
.C(n_2916),
.Y(n_5848)
);

NOR2xp67_ASAP7_75t_L g5849 ( 
.A(n_4971),
.B(n_3559),
.Y(n_5849)
);

INVx3_ASAP7_75t_L g5850 ( 
.A(n_4496),
.Y(n_5850)
);

AND2x4_ASAP7_75t_L g5851 ( 
.A(n_4642),
.B(n_3750),
.Y(n_5851)
);

INVx2_ASAP7_75t_L g5852 ( 
.A(n_4710),
.Y(n_5852)
);

NOR2xp67_ASAP7_75t_SL g5853 ( 
.A(n_4521),
.B(n_3003),
.Y(n_5853)
);

AND2x2_ASAP7_75t_L g5854 ( 
.A(n_4395),
.B(n_3998),
.Y(n_5854)
);

AO32x2_ASAP7_75t_L g5855 ( 
.A1(n_4371),
.A2(n_3726),
.A3(n_3797),
.B1(n_3524),
.B2(n_4040),
.Y(n_5855)
);

BUFx6f_ASAP7_75t_SL g5856 ( 
.A(n_4604),
.Y(n_5856)
);

AOI21xp33_ASAP7_75t_L g5857 ( 
.A1(n_4652),
.A2(n_3603),
.B(n_3567),
.Y(n_5857)
);

O2A1O1Ixp33_ASAP7_75t_SL g5858 ( 
.A1(n_5011),
.A2(n_4018),
.B(n_3576),
.C(n_3581),
.Y(n_5858)
);

OAI21x1_ASAP7_75t_L g5859 ( 
.A1(n_4405),
.A2(n_3576),
.B(n_3561),
.Y(n_5859)
);

O2A1O1Ixp33_ASAP7_75t_L g5860 ( 
.A1(n_4891),
.A2(n_2908),
.B(n_2916),
.C(n_2889),
.Y(n_5860)
);

INVx1_ASAP7_75t_L g5861 ( 
.A(n_4934),
.Y(n_5861)
);

NOR2xp33_ASAP7_75t_L g5862 ( 
.A(n_4632),
.B(n_2913),
.Y(n_5862)
);

OAI22xp5_ASAP7_75t_L g5863 ( 
.A1(n_5108),
.A2(n_3758),
.B1(n_3821),
.B2(n_3803),
.Y(n_5863)
);

AOI21xp5_ASAP7_75t_L g5864 ( 
.A1(n_4874),
.A2(n_2943),
.B(n_2927),
.Y(n_5864)
);

OAI22xp5_ASAP7_75t_L g5865 ( 
.A1(n_5108),
.A2(n_3758),
.B1(n_3821),
.B2(n_3803),
.Y(n_5865)
);

NAND2xp5_ASAP7_75t_L g5866 ( 
.A(n_4701),
.B(n_3797),
.Y(n_5866)
);

INVx1_ASAP7_75t_L g5867 ( 
.A(n_4934),
.Y(n_5867)
);

INVx1_ASAP7_75t_L g5868 ( 
.A(n_4935),
.Y(n_5868)
);

INVxp67_ASAP7_75t_SL g5869 ( 
.A(n_4673),
.Y(n_5869)
);

O2A1O1Ixp33_ASAP7_75t_L g5870 ( 
.A1(n_4891),
.A2(n_2908),
.B(n_2916),
.C(n_2889),
.Y(n_5870)
);

NAND2xp5_ASAP7_75t_L g5871 ( 
.A(n_4701),
.B(n_3581),
.Y(n_5871)
);

INVx1_ASAP7_75t_L g5872 ( 
.A(n_4935),
.Y(n_5872)
);

NAND2xp5_ASAP7_75t_L g5873 ( 
.A(n_4703),
.B(n_3606),
.Y(n_5873)
);

NOR2xp67_ASAP7_75t_L g5874 ( 
.A(n_4971),
.B(n_3606),
.Y(n_5874)
);

NOR2xp33_ASAP7_75t_L g5875 ( 
.A(n_4744),
.B(n_2922),
.Y(n_5875)
);

BUFx12f_ASAP7_75t_L g5876 ( 
.A(n_4604),
.Y(n_5876)
);

AOI21xp5_ASAP7_75t_SL g5877 ( 
.A1(n_4416),
.A2(n_3005),
.B(n_2992),
.Y(n_5877)
);

NOR2xp33_ASAP7_75t_L g5878 ( 
.A(n_4744),
.B(n_2922),
.Y(n_5878)
);

INVx3_ASAP7_75t_L g5879 ( 
.A(n_4496),
.Y(n_5879)
);

OAI21xp5_ASAP7_75t_L g5880 ( 
.A1(n_4522),
.A2(n_3273),
.B(n_3269),
.Y(n_5880)
);

OAI21xp5_ASAP7_75t_L g5881 ( 
.A1(n_4522),
.A2(n_3273),
.B(n_3269),
.Y(n_5881)
);

A2O1A1Ixp33_ASAP7_75t_L g5882 ( 
.A1(n_4564),
.A2(n_2945),
.B(n_2970),
.C(n_2938),
.Y(n_5882)
);

AO32x2_ASAP7_75t_L g5883 ( 
.A1(n_4371),
.A2(n_3524),
.A3(n_3588),
.B1(n_3613),
.B2(n_3648),
.Y(n_5883)
);

A2O1A1Ixp33_ASAP7_75t_L g5884 ( 
.A1(n_4564),
.A2(n_2945),
.B(n_2970),
.C(n_2938),
.Y(n_5884)
);

CKINVDCx11_ASAP7_75t_R g5885 ( 
.A(n_4720),
.Y(n_5885)
);

A2O1A1Ixp33_ASAP7_75t_L g5886 ( 
.A1(n_4569),
.A2(n_4728),
.B(n_4647),
.C(n_4945),
.Y(n_5886)
);

INVx5_ASAP7_75t_L g5887 ( 
.A(n_4971),
.Y(n_5887)
);

NAND2xp5_ASAP7_75t_L g5888 ( 
.A(n_4703),
.B(n_3609),
.Y(n_5888)
);

A2O1A1Ixp33_ASAP7_75t_L g5889 ( 
.A1(n_4569),
.A2(n_2945),
.B(n_2970),
.C(n_2938),
.Y(n_5889)
);

OR2x6_ASAP7_75t_L g5890 ( 
.A(n_4579),
.B(n_3758),
.Y(n_5890)
);

INVx3_ASAP7_75t_L g5891 ( 
.A(n_4496),
.Y(n_5891)
);

HB1xp67_ASAP7_75t_L g5892 ( 
.A(n_4887),
.Y(n_5892)
);

OAI21xp5_ASAP7_75t_SL g5893 ( 
.A1(n_4507),
.A2(n_2945),
.B(n_2938),
.Y(n_5893)
);

AND2x2_ASAP7_75t_L g5894 ( 
.A(n_4395),
.B(n_3588),
.Y(n_5894)
);

AOI21xp5_ASAP7_75t_L g5895 ( 
.A1(n_4883),
.A2(n_2975),
.B(n_2943),
.Y(n_5895)
);

NOR2xp67_ASAP7_75t_L g5896 ( 
.A(n_5059),
.B(n_3641),
.Y(n_5896)
);

BUFx4f_ASAP7_75t_L g5897 ( 
.A(n_4759),
.Y(n_5897)
);

INVx2_ASAP7_75t_L g5898 ( 
.A(n_4710),
.Y(n_5898)
);

AOI21xp5_ASAP7_75t_L g5899 ( 
.A1(n_4883),
.A2(n_2975),
.B(n_2943),
.Y(n_5899)
);

NAND2xp5_ASAP7_75t_L g5900 ( 
.A(n_4955),
.B(n_3641),
.Y(n_5900)
);

HB1xp67_ASAP7_75t_L g5901 ( 
.A(n_4887),
.Y(n_5901)
);

OR2x6_ASAP7_75t_L g5902 ( 
.A(n_4579),
.B(n_3758),
.Y(n_5902)
);

BUFx8_ASAP7_75t_L g5903 ( 
.A(n_4961),
.Y(n_5903)
);

NOR2xp33_ASAP7_75t_L g5904 ( 
.A(n_4795),
.B(n_2938),
.Y(n_5904)
);

NAND2xp5_ASAP7_75t_L g5905 ( 
.A(n_4958),
.B(n_3644),
.Y(n_5905)
);

AND2x2_ASAP7_75t_L g5906 ( 
.A(n_4395),
.B(n_3644),
.Y(n_5906)
);

AOI21xp5_ASAP7_75t_L g5907 ( 
.A1(n_4416),
.A2(n_3067),
.B(n_2975),
.Y(n_5907)
);

NAND2x1p5_ASAP7_75t_L g5908 ( 
.A(n_5059),
.B(n_5143),
.Y(n_5908)
);

AO21x1_ASAP7_75t_L g5909 ( 
.A1(n_4958),
.A2(n_4979),
.B(n_4973),
.Y(n_5909)
);

A2O1A1Ixp33_ASAP7_75t_L g5910 ( 
.A1(n_4728),
.A2(n_2945),
.B(n_2970),
.C(n_2938),
.Y(n_5910)
);

OAI22xp33_ASAP7_75t_L g5911 ( 
.A1(n_4943),
.A2(n_3821),
.B1(n_3855),
.B2(n_3803),
.Y(n_5911)
);

AOI21x1_ASAP7_75t_L g5912 ( 
.A1(n_4981),
.A2(n_3652),
.B(n_3648),
.Y(n_5912)
);

HB1xp67_ASAP7_75t_L g5913 ( 
.A(n_4887),
.Y(n_5913)
);

OR2x6_ASAP7_75t_L g5914 ( 
.A(n_4579),
.B(n_3803),
.Y(n_5914)
);

BUFx12f_ASAP7_75t_L g5915 ( 
.A(n_4604),
.Y(n_5915)
);

NAND2xp5_ASAP7_75t_L g5916 ( 
.A(n_4973),
.B(n_4979),
.Y(n_5916)
);

AOI221xp5_ASAP7_75t_SL g5917 ( 
.A1(n_4746),
.A2(n_3616),
.B1(n_3666),
.B2(n_3942),
.C(n_3909),
.Y(n_5917)
);

NAND2xp5_ASAP7_75t_L g5918 ( 
.A(n_4980),
.B(n_3616),
.Y(n_5918)
);

AOI21xp5_ASAP7_75t_L g5919 ( 
.A1(n_4783),
.A2(n_4807),
.B(n_4647),
.Y(n_5919)
);

INVx2_ASAP7_75t_L g5920 ( 
.A(n_4710),
.Y(n_5920)
);

AO21x2_ASAP7_75t_L g5921 ( 
.A1(n_4807),
.A2(n_2878),
.B(n_2875),
.Y(n_5921)
);

BUFx6f_ASAP7_75t_L g5922 ( 
.A(n_4496),
.Y(n_5922)
);

INVx4_ASAP7_75t_L g5923 ( 
.A(n_4604),
.Y(n_5923)
);

BUFx2_ASAP7_75t_L g5924 ( 
.A(n_5116),
.Y(n_5924)
);

INVx2_ASAP7_75t_L g5925 ( 
.A(n_4757),
.Y(n_5925)
);

A2O1A1Ixp33_ASAP7_75t_L g5926 ( 
.A1(n_4945),
.A2(n_2945),
.B(n_2970),
.C(n_2938),
.Y(n_5926)
);

OAI22xp5_ASAP7_75t_L g5927 ( 
.A1(n_4995),
.A2(n_3821),
.B1(n_3855),
.B2(n_3803),
.Y(n_5927)
);

AND2x4_ASAP7_75t_L g5928 ( 
.A(n_4642),
.B(n_3803),
.Y(n_5928)
);

OAI21x1_ASAP7_75t_L g5929 ( 
.A1(n_4411),
.A2(n_2916),
.B(n_2908),
.Y(n_5929)
);

OAI21x1_ASAP7_75t_L g5930 ( 
.A1(n_4423),
.A2(n_2932),
.B(n_2908),
.Y(n_5930)
);

AOI221x1_ASAP7_75t_L g5931 ( 
.A1(n_4535),
.A2(n_3026),
.B1(n_3054),
.B2(n_3058),
.C(n_3079),
.Y(n_5931)
);

AND2x2_ASAP7_75t_L g5932 ( 
.A(n_4662),
.B(n_3666),
.Y(n_5932)
);

OA21x2_ASAP7_75t_L g5933 ( 
.A1(n_4423),
.A2(n_3057),
.B(n_3046),
.Y(n_5933)
);

INVx1_ASAP7_75t_L g5934 ( 
.A(n_4985),
.Y(n_5934)
);

NOR2xp33_ASAP7_75t_L g5935 ( 
.A(n_4795),
.B(n_2945),
.Y(n_5935)
);

O2A1O1Ixp5_ASAP7_75t_L g5936 ( 
.A1(n_5087),
.A2(n_2973),
.B(n_2974),
.C(n_2970),
.Y(n_5936)
);

OAI21xp5_ASAP7_75t_L g5937 ( 
.A1(n_4535),
.A2(n_3273),
.B(n_3269),
.Y(n_5937)
);

NAND2x1_ASAP7_75t_L g5938 ( 
.A(n_4406),
.B(n_3598),
.Y(n_5938)
);

AOI21xp5_ASAP7_75t_L g5939 ( 
.A1(n_5069),
.A2(n_4418),
.B(n_4895),
.Y(n_5939)
);

BUFx8_ASAP7_75t_L g5940 ( 
.A(n_5134),
.Y(n_5940)
);

INVx1_ASAP7_75t_L g5941 ( 
.A(n_4985),
.Y(n_5941)
);

OAI21xp5_ASAP7_75t_L g5942 ( 
.A1(n_4984),
.A2(n_3273),
.B(n_3269),
.Y(n_5942)
);

OA21x2_ASAP7_75t_L g5943 ( 
.A1(n_4423),
.A2(n_5000),
.B(n_4442),
.Y(n_5943)
);

BUFx3_ASAP7_75t_L g5944 ( 
.A(n_5116),
.Y(n_5944)
);

NAND2xp5_ASAP7_75t_L g5945 ( 
.A(n_4980),
.B(n_3821),
.Y(n_5945)
);

NAND2xp5_ASAP7_75t_L g5946 ( 
.A(n_4983),
.B(n_3855),
.Y(n_5946)
);

INVx1_ASAP7_75t_L g5947 ( 
.A(n_4988),
.Y(n_5947)
);

INVx2_ASAP7_75t_L g5948 ( 
.A(n_4757),
.Y(n_5948)
);

NAND2xp5_ASAP7_75t_L g5949 ( 
.A(n_4983),
.B(n_3855),
.Y(n_5949)
);

OAI221xp5_ASAP7_75t_L g5950 ( 
.A1(n_4607),
.A2(n_4943),
.B1(n_5046),
.B2(n_5034),
.C(n_4510),
.Y(n_5950)
);

BUFx10_ASAP7_75t_L g5951 ( 
.A(n_5099),
.Y(n_5951)
);

NAND2x1p5_ASAP7_75t_L g5952 ( 
.A(n_5059),
.B(n_3855),
.Y(n_5952)
);

AOI22xp5_ASAP7_75t_L g5953 ( 
.A1(n_4731),
.A2(n_2980),
.B1(n_2970),
.B2(n_2974),
.Y(n_5953)
);

NOR2x1_ASAP7_75t_SL g5954 ( 
.A(n_4881),
.B(n_3881),
.Y(n_5954)
);

NAND2xp5_ASAP7_75t_L g5955 ( 
.A(n_4986),
.B(n_3881),
.Y(n_5955)
);

INVx2_ASAP7_75t_SL g5956 ( 
.A(n_5125),
.Y(n_5956)
);

AOI21xp5_ASAP7_75t_L g5957 ( 
.A1(n_4895),
.A2(n_3904),
.B(n_3881),
.Y(n_5957)
);

OAI22xp5_ASAP7_75t_L g5958 ( 
.A1(n_4995),
.A2(n_3904),
.B1(n_3909),
.B2(n_3881),
.Y(n_5958)
);

CKINVDCx20_ASAP7_75t_R g5959 ( 
.A(n_4729),
.Y(n_5959)
);

A2O1A1Ixp33_ASAP7_75t_L g5960 ( 
.A1(n_4962),
.A2(n_2974),
.B(n_3009),
.C(n_2973),
.Y(n_5960)
);

NAND3xp33_ASAP7_75t_L g5961 ( 
.A(n_4962),
.B(n_5000),
.C(n_5016),
.Y(n_5961)
);

BUFx3_ASAP7_75t_L g5962 ( 
.A(n_5125),
.Y(n_5962)
);

OAI22xp33_ASAP7_75t_L g5963 ( 
.A1(n_5034),
.A2(n_3904),
.B1(n_3909),
.B2(n_3881),
.Y(n_5963)
);

OAI21x1_ASAP7_75t_L g5964 ( 
.A1(n_4877),
.A2(n_2966),
.B(n_2932),
.Y(n_5964)
);

AO32x2_ASAP7_75t_L g5965 ( 
.A1(n_4371),
.A2(n_4018),
.A3(n_2975),
.B1(n_3072),
.B2(n_3067),
.Y(n_5965)
);

OAI22xp5_ASAP7_75t_L g5966 ( 
.A1(n_4995),
.A2(n_3909),
.B1(n_3942),
.B2(n_3904),
.Y(n_5966)
);

AOI22xp33_ASAP7_75t_L g5967 ( 
.A1(n_4759),
.A2(n_3909),
.B1(n_3942),
.B2(n_3904),
.Y(n_5967)
);

AOI21xp5_ASAP7_75t_L g5968 ( 
.A1(n_4964),
.A2(n_3909),
.B(n_3904),
.Y(n_5968)
);

OAI21x1_ASAP7_75t_L g5969 ( 
.A1(n_4877),
.A2(n_2966),
.B(n_2932),
.Y(n_5969)
);

AND2x4_ASAP7_75t_L g5970 ( 
.A(n_4676),
.B(n_3904),
.Y(n_5970)
);

INVx1_ASAP7_75t_L g5971 ( 
.A(n_4988),
.Y(n_5971)
);

A2O1A1Ixp33_ASAP7_75t_L g5972 ( 
.A1(n_4969),
.A2(n_2974),
.B(n_3009),
.C(n_2973),
.Y(n_5972)
);

OAI21x1_ASAP7_75t_L g5973 ( 
.A1(n_4877),
.A2(n_2966),
.B(n_2932),
.Y(n_5973)
);

NAND2xp5_ASAP7_75t_L g5974 ( 
.A(n_4986),
.B(n_3942),
.Y(n_5974)
);

AOI22xp33_ASAP7_75t_L g5975 ( 
.A1(n_5134),
.A2(n_4125),
.B1(n_3942),
.B2(n_3598),
.Y(n_5975)
);

OAI21x1_ASAP7_75t_L g5976 ( 
.A1(n_4657),
.A2(n_2966),
.B(n_2932),
.Y(n_5976)
);

AO31x2_ASAP7_75t_L g5977 ( 
.A1(n_4485),
.A2(n_3060),
.A3(n_3066),
.B(n_3057),
.Y(n_5977)
);

AOI21x1_ASAP7_75t_L g5978 ( 
.A1(n_4981),
.A2(n_3203),
.B(n_3186),
.Y(n_5978)
);

INVx1_ASAP7_75t_L g5979 ( 
.A(n_5003),
.Y(n_5979)
);

NAND2x1p5_ASAP7_75t_L g5980 ( 
.A(n_5059),
.B(n_3942),
.Y(n_5980)
);

NAND2xp5_ASAP7_75t_L g5981 ( 
.A(n_4989),
.B(n_4125),
.Y(n_5981)
);

OAI22xp5_ASAP7_75t_L g5982 ( 
.A1(n_4995),
.A2(n_4125),
.B1(n_3165),
.B2(n_2876),
.Y(n_5982)
);

AOI21xp5_ASAP7_75t_L g5983 ( 
.A1(n_5062),
.A2(n_3067),
.B(n_2975),
.Y(n_5983)
);

OAI21x1_ASAP7_75t_L g5984 ( 
.A1(n_4657),
.A2(n_2966),
.B(n_2932),
.Y(n_5984)
);

OA21x2_ASAP7_75t_L g5985 ( 
.A1(n_4430),
.A2(n_3066),
.B(n_3060),
.Y(n_5985)
);

CKINVDCx5p33_ASAP7_75t_R g5986 ( 
.A(n_4729),
.Y(n_5986)
);

AOI21xp5_ASAP7_75t_L g5987 ( 
.A1(n_5062),
.A2(n_3067),
.B(n_2975),
.Y(n_5987)
);

AOI21x1_ASAP7_75t_L g5988 ( 
.A1(n_4881),
.A2(n_3203),
.B(n_3186),
.Y(n_5988)
);

NAND2xp5_ASAP7_75t_SL g5989 ( 
.A(n_4507),
.B(n_3433),
.Y(n_5989)
);

O2A1O1Ixp5_ASAP7_75t_SL g5990 ( 
.A1(n_4864),
.A2(n_2966),
.B(n_2977),
.C(n_2932),
.Y(n_5990)
);

AO31x2_ASAP7_75t_L g5991 ( 
.A1(n_4485),
.A2(n_3066),
.A3(n_3084),
.B(n_3060),
.Y(n_5991)
);

AOI221xp5_ASAP7_75t_L g5992 ( 
.A1(n_4719),
.A2(n_3440),
.B1(n_3330),
.B2(n_4125),
.C(n_3014),
.Y(n_5992)
);

OAI21x1_ASAP7_75t_L g5993 ( 
.A1(n_4664),
.A2(n_2977),
.B(n_2966),
.Y(n_5993)
);

NOR2xp33_ASAP7_75t_L g5994 ( 
.A(n_5022),
.B(n_2973),
.Y(n_5994)
);

OAI21x1_ASAP7_75t_L g5995 ( 
.A1(n_4664),
.A2(n_2995),
.B(n_2977),
.Y(n_5995)
);

INVx1_ASAP7_75t_L g5996 ( 
.A(n_5003),
.Y(n_5996)
);

OAI22xp5_ASAP7_75t_L g5997 ( 
.A1(n_4520),
.A2(n_4125),
.B1(n_3165),
.B2(n_2876),
.Y(n_5997)
);

CKINVDCx5p33_ASAP7_75t_R g5998 ( 
.A(n_4729),
.Y(n_5998)
);

OAI21xp5_ASAP7_75t_L g5999 ( 
.A1(n_4984),
.A2(n_3273),
.B(n_3269),
.Y(n_5999)
);

OAI21xp5_ASAP7_75t_L g6000 ( 
.A1(n_4999),
.A2(n_3336),
.B(n_3326),
.Y(n_6000)
);

INVx2_ASAP7_75t_L g6001 ( 
.A(n_4757),
.Y(n_6001)
);

BUFx3_ASAP7_75t_L g6002 ( 
.A(n_5125),
.Y(n_6002)
);

BUFx3_ASAP7_75t_L g6003 ( 
.A(n_4764),
.Y(n_6003)
);

AOI21xp5_ASAP7_75t_L g6004 ( 
.A1(n_4999),
.A2(n_3067),
.B(n_2975),
.Y(n_6004)
);

OAI21x1_ASAP7_75t_L g6005 ( 
.A1(n_4655),
.A2(n_2995),
.B(n_2977),
.Y(n_6005)
);

CKINVDCx11_ASAP7_75t_R g6006 ( 
.A(n_4764),
.Y(n_6006)
);

AOI21xp5_ASAP7_75t_L g6007 ( 
.A1(n_4716),
.A2(n_3072),
.B(n_3067),
.Y(n_6007)
);

INVx5_ASAP7_75t_L g6008 ( 
.A(n_5059),
.Y(n_6008)
);

AOI21xp5_ASAP7_75t_L g6009 ( 
.A1(n_4716),
.A2(n_3072),
.B(n_3067),
.Y(n_6009)
);

AOI22xp5_ASAP7_75t_L g6010 ( 
.A1(n_4731),
.A2(n_2980),
.B1(n_2973),
.B2(n_2974),
.Y(n_6010)
);

A2O1A1Ixp33_ASAP7_75t_L g6011 ( 
.A1(n_4969),
.A2(n_2974),
.B(n_3009),
.C(n_3014),
.Y(n_6011)
);

NOR2xp33_ASAP7_75t_L g6012 ( 
.A(n_5022),
.B(n_2973),
.Y(n_6012)
);

AO31x2_ASAP7_75t_L g6013 ( 
.A1(n_5105),
.A2(n_5121),
.A3(n_5109),
.B(n_4533),
.Y(n_6013)
);

BUFx2_ASAP7_75t_L g6014 ( 
.A(n_5134),
.Y(n_6014)
);

AOI21xp5_ASAP7_75t_L g6015 ( 
.A1(n_5001),
.A2(n_3072),
.B(n_4125),
.Y(n_6015)
);

INVx3_ASAP7_75t_L g6016 ( 
.A(n_4496),
.Y(n_6016)
);

AOI22xp5_ASAP7_75t_L g6017 ( 
.A1(n_5046),
.A2(n_2974),
.B1(n_3014),
.B2(n_2973),
.Y(n_6017)
);

AND2x2_ASAP7_75t_L g6018 ( 
.A(n_4662),
.B(n_3844),
.Y(n_6018)
);

AO22x2_ASAP7_75t_L g6019 ( 
.A1(n_4822),
.A2(n_3172),
.B1(n_2977),
.B2(n_3166),
.Y(n_6019)
);

AOI22xp5_ASAP7_75t_L g6020 ( 
.A1(n_4723),
.A2(n_3014),
.B1(n_3009),
.B2(n_3598),
.Y(n_6020)
);

NAND2xp5_ASAP7_75t_L g6021 ( 
.A(n_4989),
.B(n_3598),
.Y(n_6021)
);

BUFx4f_ASAP7_75t_L g6022 ( 
.A(n_4954),
.Y(n_6022)
);

O2A1O1Ixp33_ASAP7_75t_SL g6023 ( 
.A1(n_5130),
.A2(n_3131),
.B(n_2995),
.C(n_3026),
.Y(n_6023)
);

OAI22xp33_ASAP7_75t_L g6024 ( 
.A1(n_4510),
.A2(n_3165),
.B1(n_2876),
.B2(n_3075),
.Y(n_6024)
);

INVx1_ASAP7_75t_L g6025 ( 
.A(n_5007),
.Y(n_6025)
);

INVx4_ASAP7_75t_SL g6026 ( 
.A(n_5099),
.Y(n_6026)
);

INVx1_ASAP7_75t_L g6027 ( 
.A(n_5007),
.Y(n_6027)
);

AOI21xp5_ASAP7_75t_L g6028 ( 
.A1(n_4394),
.A2(n_3411),
.B(n_3407),
.Y(n_6028)
);

OA21x2_ASAP7_75t_L g6029 ( 
.A1(n_4430),
.A2(n_3066),
.B(n_3060),
.Y(n_6029)
);

NAND2xp5_ASAP7_75t_L g6030 ( 
.A(n_5208),
.B(n_4864),
.Y(n_6030)
);

INVx2_ASAP7_75t_L g6031 ( 
.A(n_5883),
.Y(n_6031)
);

AOI22xp33_ASAP7_75t_L g6032 ( 
.A1(n_5146),
.A2(n_4662),
.B1(n_4436),
.B2(n_4723),
.Y(n_6032)
);

INVx4_ASAP7_75t_L g6033 ( 
.A(n_5607),
.Y(n_6033)
);

AO31x2_ASAP7_75t_L g6034 ( 
.A1(n_5909),
.A2(n_4533),
.A3(n_4615),
.B(n_4520),
.Y(n_6034)
);

OAI21xp5_ASAP7_75t_L g6035 ( 
.A1(n_5160),
.A2(n_4576),
.B(n_4403),
.Y(n_6035)
);

INVx3_ASAP7_75t_L g6036 ( 
.A(n_5890),
.Y(n_6036)
);

INVx1_ASAP7_75t_L g6037 ( 
.A(n_5280),
.Y(n_6037)
);

BUFx6f_ASAP7_75t_L g6038 ( 
.A(n_5334),
.Y(n_6038)
);

BUFx8_ASAP7_75t_L g6039 ( 
.A(n_5856),
.Y(n_6039)
);

BUFx6f_ASAP7_75t_L g6040 ( 
.A(n_5334),
.Y(n_6040)
);

INVx2_ASAP7_75t_L g6041 ( 
.A(n_5883),
.Y(n_6041)
);

BUFx6f_ASAP7_75t_L g6042 ( 
.A(n_5334),
.Y(n_6042)
);

AOI22xp33_ASAP7_75t_L g6043 ( 
.A1(n_5146),
.A2(n_4436),
.B1(n_4909),
.B2(n_4739),
.Y(n_6043)
);

INVx1_ASAP7_75t_L g6044 ( 
.A(n_5280),
.Y(n_6044)
);

OAI21x1_ASAP7_75t_L g6045 ( 
.A1(n_5309),
.A2(n_4643),
.B(n_4442),
.Y(n_6045)
);

O2A1O1Ixp33_ASAP7_75t_SL g6046 ( 
.A1(n_5218),
.A2(n_5130),
.B(n_4953),
.C(n_4956),
.Y(n_6046)
);

OA21x2_ASAP7_75t_L g6047 ( 
.A1(n_5220),
.A2(n_4479),
.B(n_4457),
.Y(n_6047)
);

OAI21x1_ASAP7_75t_L g6048 ( 
.A1(n_5309),
.A2(n_4643),
.B(n_4442),
.Y(n_6048)
);

NOR2xp33_ASAP7_75t_SL g6049 ( 
.A(n_5508),
.B(n_4798),
.Y(n_6049)
);

INVx2_ASAP7_75t_L g6050 ( 
.A(n_5883),
.Y(n_6050)
);

BUFx3_ASAP7_75t_L g6051 ( 
.A(n_5646),
.Y(n_6051)
);

HB1xp67_ASAP7_75t_L g6052 ( 
.A(n_5550),
.Y(n_6052)
);

AOI22xp5_ASAP7_75t_L g6053 ( 
.A1(n_5154),
.A2(n_5126),
.B1(n_5035),
.B2(n_4965),
.Y(n_6053)
);

AOI222xp33_ASAP7_75t_L g6054 ( 
.A1(n_5214),
.A2(n_4739),
.B1(n_4733),
.B2(n_5033),
.C1(n_5027),
.C2(n_5005),
.Y(n_6054)
);

OAI22xp33_ASAP7_75t_L g6055 ( 
.A1(n_5247),
.A2(n_5360),
.B1(n_5201),
.B2(n_5202),
.Y(n_6055)
);

OAI21x1_ASAP7_75t_L g6056 ( 
.A1(n_5314),
.A2(n_4448),
.B(n_4576),
.Y(n_6056)
);

OAI21x1_ASAP7_75t_L g6057 ( 
.A1(n_5152),
.A2(n_4448),
.B(n_4576),
.Y(n_6057)
);

OAI21x1_ASAP7_75t_SL g6058 ( 
.A1(n_5156),
.A2(n_5135),
.B(n_5137),
.Y(n_6058)
);

INVx1_ASAP7_75t_L g6059 ( 
.A(n_5285),
.Y(n_6059)
);

OAI21x1_ASAP7_75t_L g6060 ( 
.A1(n_5152),
.A2(n_4737),
.B(n_4734),
.Y(n_6060)
);

AND2x4_ASAP7_75t_L g6061 ( 
.A(n_5710),
.B(n_4477),
.Y(n_6061)
);

BUFx12f_ASAP7_75t_L g6062 ( 
.A(n_5184),
.Y(n_6062)
);

OAI21x1_ASAP7_75t_L g6063 ( 
.A1(n_5263),
.A2(n_4737),
.B(n_4734),
.Y(n_6063)
);

OAI21x1_ASAP7_75t_L g6064 ( 
.A1(n_5263),
.A2(n_4737),
.B(n_4734),
.Y(n_6064)
);

AND2x4_ASAP7_75t_L g6065 ( 
.A(n_5710),
.B(n_4477),
.Y(n_6065)
);

NAND3xp33_ASAP7_75t_L g6066 ( 
.A(n_5160),
.B(n_5016),
.C(n_4771),
.Y(n_6066)
);

INVx1_ASAP7_75t_L g6067 ( 
.A(n_5285),
.Y(n_6067)
);

NAND2x1p5_ASAP7_75t_L g6068 ( 
.A(n_5334),
.B(n_4477),
.Y(n_6068)
);

OAI21x1_ASAP7_75t_L g6069 ( 
.A1(n_5812),
.A2(n_4907),
.B(n_4717),
.Y(n_6069)
);

NAND2xp5_ASAP7_75t_L g6070 ( 
.A(n_5208),
.B(n_4392),
.Y(n_6070)
);

BUFx3_ASAP7_75t_L g6071 ( 
.A(n_5646),
.Y(n_6071)
);

NAND2xp5_ASAP7_75t_L g6072 ( 
.A(n_5219),
.B(n_4392),
.Y(n_6072)
);

NAND2x1p5_ASAP7_75t_L g6073 ( 
.A(n_5334),
.B(n_4477),
.Y(n_6073)
);

INVxp67_ASAP7_75t_SL g6074 ( 
.A(n_5736),
.Y(n_6074)
);

INVx1_ASAP7_75t_L g6075 ( 
.A(n_5292),
.Y(n_6075)
);

BUFx6f_ASAP7_75t_L g6076 ( 
.A(n_5334),
.Y(n_6076)
);

OAI21x1_ASAP7_75t_L g6077 ( 
.A1(n_5812),
.A2(n_4907),
.B(n_4717),
.Y(n_6077)
);

AOI22xp33_ASAP7_75t_L g6078 ( 
.A1(n_5214),
.A2(n_4909),
.B1(n_4733),
.B2(n_4965),
.Y(n_6078)
);

INVx8_ASAP7_75t_L g6079 ( 
.A(n_5607),
.Y(n_6079)
);

OAI21x1_ASAP7_75t_L g6080 ( 
.A1(n_5150),
.A2(n_4907),
.B(n_4717),
.Y(n_6080)
);

NAND2xp5_ASAP7_75t_L g6081 ( 
.A(n_5457),
.B(n_5473),
.Y(n_6081)
);

NOR2xp33_ASAP7_75t_L g6082 ( 
.A(n_5277),
.B(n_4822),
.Y(n_6082)
);

OAI22xp5_ASAP7_75t_L g6083 ( 
.A1(n_5247),
.A2(n_4533),
.B1(n_4615),
.B2(n_4520),
.Y(n_6083)
);

OAI22xp5_ASAP7_75t_SL g6084 ( 
.A1(n_5505),
.A2(n_5058),
.B1(n_4672),
.B2(n_4682),
.Y(n_6084)
);

A2O1A1Ixp33_ASAP7_75t_L g6085 ( 
.A1(n_5155),
.A2(n_5068),
.B(n_4394),
.C(n_4403),
.Y(n_6085)
);

OAI21x1_ASAP7_75t_L g6086 ( 
.A1(n_5150),
.A2(n_4714),
.B(n_4881),
.Y(n_6086)
);

BUFx2_ASAP7_75t_L g6087 ( 
.A(n_5890),
.Y(n_6087)
);

NOR2xp33_ASAP7_75t_L g6088 ( 
.A(n_5277),
.B(n_5058),
.Y(n_6088)
);

BUFx12f_ASAP7_75t_L g6089 ( 
.A(n_5212),
.Y(n_6089)
);

AOI221xp5_ASAP7_75t_L g6090 ( 
.A1(n_5218),
.A2(n_4682),
.B1(n_4756),
.B2(n_4672),
.C(n_4615),
.Y(n_6090)
);

BUFx3_ASAP7_75t_L g6091 ( 
.A(n_5646),
.Y(n_6091)
);

INVx1_ASAP7_75t_SL g6092 ( 
.A(n_5353),
.Y(n_6092)
);

OAI21x1_ASAP7_75t_L g6093 ( 
.A1(n_5243),
.A2(n_4714),
.B(n_4523),
.Y(n_6093)
);

A2O1A1Ixp33_ASAP7_75t_L g6094 ( 
.A1(n_5156),
.A2(n_5068),
.B(n_4607),
.C(n_4609),
.Y(n_6094)
);

OAI21xp5_ASAP7_75t_L g6095 ( 
.A1(n_5158),
.A2(n_5140),
.B(n_5133),
.Y(n_6095)
);

AOI21x1_ASAP7_75t_L g6096 ( 
.A1(n_5220),
.A2(n_4556),
.B(n_5121),
.Y(n_6096)
);

OAI21x1_ASAP7_75t_L g6097 ( 
.A1(n_5243),
.A2(n_4714),
.B(n_4523),
.Y(n_6097)
);

OA21x2_ASAP7_75t_L g6098 ( 
.A1(n_5249),
.A2(n_4479),
.B(n_4457),
.Y(n_6098)
);

INVx1_ASAP7_75t_L g6099 ( 
.A(n_5292),
.Y(n_6099)
);

INVx2_ASAP7_75t_L g6100 ( 
.A(n_5883),
.Y(n_6100)
);

BUFx6f_ASAP7_75t_L g6101 ( 
.A(n_5348),
.Y(n_6101)
);

INVx1_ASAP7_75t_L g6102 ( 
.A(n_5299),
.Y(n_6102)
);

INVx4_ASAP7_75t_L g6103 ( 
.A(n_5607),
.Y(n_6103)
);

BUFx8_ASAP7_75t_L g6104 ( 
.A(n_5856),
.Y(n_6104)
);

INVx1_ASAP7_75t_SL g6105 ( 
.A(n_5353),
.Y(n_6105)
);

OA21x2_ASAP7_75t_L g6106 ( 
.A1(n_5249),
.A2(n_4508),
.B(n_4497),
.Y(n_6106)
);

OAI22xp5_ASAP7_75t_L g6107 ( 
.A1(n_5360),
.A2(n_4682),
.B1(n_4756),
.B2(n_4672),
.Y(n_6107)
);

AO21x2_ASAP7_75t_L g6108 ( 
.A1(n_5234),
.A2(n_4918),
.B(n_4891),
.Y(n_6108)
);

NOR2xp33_ASAP7_75t_R g6109 ( 
.A(n_5187),
.B(n_5515),
.Y(n_6109)
);

OA21x2_ASAP7_75t_L g6110 ( 
.A1(n_5254),
.A2(n_5500),
.B(n_5494),
.Y(n_6110)
);

INVx3_ASAP7_75t_L g6111 ( 
.A(n_5890),
.Y(n_6111)
);

INVx4_ASAP7_75t_L g6112 ( 
.A(n_5221),
.Y(n_6112)
);

INVx2_ASAP7_75t_L g6113 ( 
.A(n_5883),
.Y(n_6113)
);

NAND2xp33_ASAP7_75t_SL g6114 ( 
.A(n_5303),
.B(n_4763),
.Y(n_6114)
);

HB1xp67_ASAP7_75t_L g6115 ( 
.A(n_5550),
.Y(n_6115)
);

INVx1_ASAP7_75t_L g6116 ( 
.A(n_5299),
.Y(n_6116)
);

OAI21xp5_ASAP7_75t_L g6117 ( 
.A1(n_5188),
.A2(n_5140),
.B(n_5133),
.Y(n_6117)
);

OAI21x1_ASAP7_75t_L g6118 ( 
.A1(n_5295),
.A2(n_4523),
.B(n_4471),
.Y(n_6118)
);

OAI21x1_ASAP7_75t_L g6119 ( 
.A1(n_5295),
.A2(n_4523),
.B(n_4471),
.Y(n_6119)
);

NAND4xp25_ASAP7_75t_L g6120 ( 
.A(n_5271),
.B(n_5415),
.C(n_5188),
.D(n_5177),
.Y(n_6120)
);

NAND2xp5_ASAP7_75t_L g6121 ( 
.A(n_5620),
.B(n_4556),
.Y(n_6121)
);

OAI22xp5_ASAP7_75t_L g6122 ( 
.A1(n_5201),
.A2(n_4763),
.B1(n_4897),
.B2(n_4776),
.Y(n_6122)
);

AOI22xp33_ASAP7_75t_L g6123 ( 
.A1(n_5144),
.A2(n_5173),
.B1(n_5177),
.B2(n_5271),
.Y(n_6123)
);

OAI21x1_ASAP7_75t_L g6124 ( 
.A1(n_5227),
.A2(n_4677),
.B(n_4471),
.Y(n_6124)
);

INVx1_ASAP7_75t_L g6125 ( 
.A(n_5302),
.Y(n_6125)
);

CKINVDCx11_ASAP7_75t_R g6126 ( 
.A(n_5169),
.Y(n_6126)
);

INVx1_ASAP7_75t_L g6127 ( 
.A(n_5302),
.Y(n_6127)
);

INVx4_ASAP7_75t_SL g6128 ( 
.A(n_5228),
.Y(n_6128)
);

OAI21x1_ASAP7_75t_L g6129 ( 
.A1(n_5227),
.A2(n_4677),
.B(n_4471),
.Y(n_6129)
);

AOI21xp5_ASAP7_75t_L g6130 ( 
.A1(n_5782),
.A2(n_4546),
.B(n_4905),
.Y(n_6130)
);

CKINVDCx20_ASAP7_75t_R g6131 ( 
.A(n_5180),
.Y(n_6131)
);

INVx1_ASAP7_75t_L g6132 ( 
.A(n_5322),
.Y(n_6132)
);

AOI21xp5_ASAP7_75t_L g6133 ( 
.A1(n_5782),
.A2(n_5777),
.B(n_5165),
.Y(n_6133)
);

NAND2x1p5_ASAP7_75t_L g6134 ( 
.A(n_5348),
.B(n_4477),
.Y(n_6134)
);

OA21x2_ASAP7_75t_L g6135 ( 
.A1(n_5254),
.A2(n_4512),
.B(n_4508),
.Y(n_6135)
);

BUFx3_ASAP7_75t_L g6136 ( 
.A(n_5646),
.Y(n_6136)
);

BUFx4f_ASAP7_75t_L g6137 ( 
.A(n_5432),
.Y(n_6137)
);

AOI22xp33_ASAP7_75t_L g6138 ( 
.A1(n_5173),
.A2(n_5118),
.B1(n_4798),
.B2(n_5123),
.Y(n_6138)
);

INVx2_ASAP7_75t_L g6139 ( 
.A(n_5883),
.Y(n_6139)
);

CKINVDCx5p33_ASAP7_75t_R g6140 ( 
.A(n_5459),
.Y(n_6140)
);

BUFx3_ASAP7_75t_L g6141 ( 
.A(n_5662),
.Y(n_6141)
);

AOI22xp33_ASAP7_75t_L g6142 ( 
.A1(n_5372),
.A2(n_5118),
.B1(n_4798),
.B2(n_5123),
.Y(n_6142)
);

INVx1_ASAP7_75t_L g6143 ( 
.A(n_5322),
.Y(n_6143)
);

AND2x2_ASAP7_75t_L g6144 ( 
.A(n_5890),
.B(n_4402),
.Y(n_6144)
);

INVx6_ASAP7_75t_L g6145 ( 
.A(n_5811),
.Y(n_6145)
);

OAI21xp5_ASAP7_75t_L g6146 ( 
.A1(n_5415),
.A2(n_5098),
.B(n_5097),
.Y(n_6146)
);

OAI21x1_ASAP7_75t_L g6147 ( 
.A1(n_5233),
.A2(n_5259),
.B(n_5743),
.Y(n_6147)
);

OAI22xp5_ASAP7_75t_L g6148 ( 
.A1(n_5202),
.A2(n_4776),
.B1(n_4897),
.B2(n_5035),
.Y(n_6148)
);

INVx1_ASAP7_75t_SL g6149 ( 
.A(n_5595),
.Y(n_6149)
);

OAI21xp5_ASAP7_75t_L g6150 ( 
.A1(n_5178),
.A2(n_5098),
.B(n_5097),
.Y(n_6150)
);

AOI222xp33_ASAP7_75t_L g6151 ( 
.A1(n_5372),
.A2(n_5033),
.B1(n_5027),
.B2(n_5005),
.C1(n_5001),
.C2(n_4853),
.Y(n_6151)
);

AND2x4_ASAP7_75t_L g6152 ( 
.A(n_5348),
.B(n_4477),
.Y(n_6152)
);

INVx1_ASAP7_75t_L g6153 ( 
.A(n_5345),
.Y(n_6153)
);

OAI21x1_ASAP7_75t_L g6154 ( 
.A1(n_5259),
.A2(n_4677),
.B(n_4761),
.Y(n_6154)
);

OAI21x1_ASAP7_75t_L g6155 ( 
.A1(n_5743),
.A2(n_5289),
.B(n_5479),
.Y(n_6155)
);

AOI21xp5_ASAP7_75t_L g6156 ( 
.A1(n_5777),
.A2(n_4546),
.B(n_4905),
.Y(n_6156)
);

INVx1_ASAP7_75t_L g6157 ( 
.A(n_5345),
.Y(n_6157)
);

OAI21xp5_ASAP7_75t_L g6158 ( 
.A1(n_5178),
.A2(n_5103),
.B(n_5101),
.Y(n_6158)
);

AOI22xp33_ASAP7_75t_L g6159 ( 
.A1(n_5327),
.A2(n_5118),
.B1(n_4798),
.B2(n_4469),
.Y(n_6159)
);

NOR2xp33_ASAP7_75t_L g6160 ( 
.A(n_5311),
.B(n_4953),
.Y(n_6160)
);

INVx1_ASAP7_75t_SL g6161 ( 
.A(n_5595),
.Y(n_6161)
);

INVx2_ASAP7_75t_L g6162 ( 
.A(n_5977),
.Y(n_6162)
);

INVx1_ASAP7_75t_L g6163 ( 
.A(n_5347),
.Y(n_6163)
);

AND2x4_ASAP7_75t_L g6164 ( 
.A(n_5348),
.B(n_4477),
.Y(n_6164)
);

AND2x2_ASAP7_75t_L g6165 ( 
.A(n_5890),
.B(n_4402),
.Y(n_6165)
);

NOR2xp67_ASAP7_75t_L g6166 ( 
.A(n_5927),
.B(n_4477),
.Y(n_6166)
);

AOI22x1_ASAP7_75t_L g6167 ( 
.A1(n_5186),
.A2(n_4609),
.B1(n_4593),
.B2(n_4406),
.Y(n_6167)
);

BUFx4f_ASAP7_75t_SL g6168 ( 
.A(n_5432),
.Y(n_6168)
);

OA21x2_ASAP7_75t_L g6169 ( 
.A1(n_5494),
.A2(n_4516),
.B(n_4512),
.Y(n_6169)
);

AO31x2_ASAP7_75t_L g6170 ( 
.A1(n_5639),
.A2(n_4516),
.A3(n_4779),
.B(n_5101),
.Y(n_6170)
);

INVx1_ASAP7_75t_L g6171 ( 
.A(n_5347),
.Y(n_6171)
);

INVx2_ASAP7_75t_L g6172 ( 
.A(n_5977),
.Y(n_6172)
);

AOI21x1_ASAP7_75t_L g6173 ( 
.A1(n_5234),
.A2(n_5096),
.B(n_4956),
.Y(n_6173)
);

AO21x2_ASAP7_75t_L g6174 ( 
.A1(n_5288),
.A2(n_4694),
.B(n_4593),
.Y(n_6174)
);

INVx2_ASAP7_75t_L g6175 ( 
.A(n_5977),
.Y(n_6175)
);

NOR2xp33_ASAP7_75t_SL g6176 ( 
.A(n_5508),
.B(n_4798),
.Y(n_6176)
);

INVx1_ASAP7_75t_L g6177 ( 
.A(n_5356),
.Y(n_6177)
);

BUFx2_ASAP7_75t_L g6178 ( 
.A(n_5902),
.Y(n_6178)
);

INVx1_ASAP7_75t_L g6179 ( 
.A(n_5356),
.Y(n_6179)
);

INVx1_ASAP7_75t_SL g6180 ( 
.A(n_5701),
.Y(n_6180)
);

INVx2_ASAP7_75t_SL g6181 ( 
.A(n_5348),
.Y(n_6181)
);

BUFx4f_ASAP7_75t_L g6182 ( 
.A(n_5432),
.Y(n_6182)
);

NAND2x1p5_ASAP7_75t_L g6183 ( 
.A(n_5348),
.B(n_4481),
.Y(n_6183)
);

INVx2_ASAP7_75t_L g6184 ( 
.A(n_5977),
.Y(n_6184)
);

OAI22xp5_ASAP7_75t_L g6185 ( 
.A1(n_5232),
.A2(n_4897),
.B1(n_4776),
.B2(n_5126),
.Y(n_6185)
);

INVx1_ASAP7_75t_L g6186 ( 
.A(n_5364),
.Y(n_6186)
);

AND2x2_ASAP7_75t_L g6187 ( 
.A(n_5902),
.B(n_4402),
.Y(n_6187)
);

OAI21x1_ASAP7_75t_L g6188 ( 
.A1(n_5491),
.A2(n_4787),
.B(n_4704),
.Y(n_6188)
);

CKINVDCx6p67_ASAP7_75t_R g6189 ( 
.A(n_5187),
.Y(n_6189)
);

AOI22xp33_ASAP7_75t_L g6190 ( 
.A1(n_5358),
.A2(n_5118),
.B1(n_5088),
.B2(n_5111),
.Y(n_6190)
);

OAI21x1_ASAP7_75t_L g6191 ( 
.A1(n_5224),
.A2(n_4787),
.B(n_4704),
.Y(n_6191)
);

INVx1_ASAP7_75t_L g6192 ( 
.A(n_5364),
.Y(n_6192)
);

AND2x4_ASAP7_75t_L g6193 ( 
.A(n_5760),
.B(n_4481),
.Y(n_6193)
);

OAI21x1_ASAP7_75t_L g6194 ( 
.A1(n_5224),
.A2(n_5153),
.B(n_5168),
.Y(n_6194)
);

NOR2xp33_ASAP7_75t_L g6195 ( 
.A(n_5272),
.B(n_5086),
.Y(n_6195)
);

AOI21xp5_ASAP7_75t_L g6196 ( 
.A1(n_6028),
.A2(n_5775),
.B(n_5769),
.Y(n_6196)
);

AOI21x1_ASAP7_75t_L g6197 ( 
.A1(n_5509),
.A2(n_5096),
.B(n_4779),
.Y(n_6197)
);

INVx4_ASAP7_75t_SL g6198 ( 
.A(n_5228),
.Y(n_6198)
);

INVx1_ASAP7_75t_L g6199 ( 
.A(n_5383),
.Y(n_6199)
);

O2A1O1Ixp33_ASAP7_75t_L g6200 ( 
.A1(n_5154),
.A2(n_4992),
.B(n_4847),
.C(n_4853),
.Y(n_6200)
);

INVx2_ASAP7_75t_L g6201 ( 
.A(n_5977),
.Y(n_6201)
);

AOI21xp5_ASAP7_75t_L g6202 ( 
.A1(n_6028),
.A2(n_4683),
.B(n_4715),
.Y(n_6202)
);

OAI21x1_ASAP7_75t_L g6203 ( 
.A1(n_5153),
.A2(n_5064),
.B(n_4959),
.Y(n_6203)
);

BUFx2_ASAP7_75t_R g6204 ( 
.A(n_5169),
.Y(n_6204)
);

NAND2xp5_ASAP7_75t_L g6205 ( 
.A(n_5869),
.B(n_4374),
.Y(n_6205)
);

AOI22xp33_ASAP7_75t_L g6206 ( 
.A1(n_5358),
.A2(n_5118),
.B1(n_5088),
.B2(n_5111),
.Y(n_6206)
);

AO31x2_ASAP7_75t_L g6207 ( 
.A1(n_5541),
.A2(n_5103),
.A3(n_4992),
.B(n_4762),
.Y(n_6207)
);

OAI21x1_ASAP7_75t_L g6208 ( 
.A1(n_5168),
.A2(n_5064),
.B(n_4959),
.Y(n_6208)
);

INVx2_ASAP7_75t_L g6209 ( 
.A(n_5977),
.Y(n_6209)
);

OAI21x1_ASAP7_75t_L g6210 ( 
.A1(n_5204),
.A2(n_4655),
.B(n_4583),
.Y(n_6210)
);

INVx1_ASAP7_75t_SL g6211 ( 
.A(n_5701),
.Y(n_6211)
);

AOI21xp5_ASAP7_75t_L g6212 ( 
.A1(n_5775),
.A2(n_4683),
.B(n_4715),
.Y(n_6212)
);

NOR2xp33_ASAP7_75t_L g6213 ( 
.A(n_5301),
.B(n_5086),
.Y(n_6213)
);

AO31x2_ASAP7_75t_L g6214 ( 
.A1(n_5558),
.A2(n_4831),
.A3(n_4866),
.B(n_4762),
.Y(n_6214)
);

NOR2xp33_ASAP7_75t_L g6215 ( 
.A(n_5301),
.B(n_5139),
.Y(n_6215)
);

INVx2_ASAP7_75t_L g6216 ( 
.A(n_5991),
.Y(n_6216)
);

INVx2_ASAP7_75t_L g6217 ( 
.A(n_5991),
.Y(n_6217)
);

A2O1A1Ixp33_ASAP7_75t_L g6218 ( 
.A1(n_5283),
.A2(n_5138),
.B(n_4724),
.C(n_4747),
.Y(n_6218)
);

OAI22xp33_ASAP7_75t_L g6219 ( 
.A1(n_5232),
.A2(n_4897),
.B1(n_4776),
.B2(n_4725),
.Y(n_6219)
);

AND2x2_ASAP7_75t_L g6220 ( 
.A(n_5902),
.B(n_4402),
.Y(n_6220)
);

NAND2xp5_ASAP7_75t_L g6221 ( 
.A(n_5916),
.B(n_4374),
.Y(n_6221)
);

INVx2_ASAP7_75t_L g6222 ( 
.A(n_5991),
.Y(n_6222)
);

INVx1_ASAP7_75t_L g6223 ( 
.A(n_5383),
.Y(n_6223)
);

AO21x2_ASAP7_75t_L g6224 ( 
.A1(n_5919),
.A2(n_4694),
.B(n_4593),
.Y(n_6224)
);

OA21x2_ASAP7_75t_L g6225 ( 
.A1(n_5284),
.A2(n_4599),
.B(n_4597),
.Y(n_6225)
);

INVx1_ASAP7_75t_L g6226 ( 
.A(n_5384),
.Y(n_6226)
);

BUFx3_ASAP7_75t_L g6227 ( 
.A(n_5662),
.Y(n_6227)
);

NAND2xp5_ASAP7_75t_SL g6228 ( 
.A(n_5354),
.B(n_4481),
.Y(n_6228)
);

INVx1_ASAP7_75t_L g6229 ( 
.A(n_5384),
.Y(n_6229)
);

A2O1A1Ixp33_ASAP7_75t_L g6230 ( 
.A1(n_5163),
.A2(n_5138),
.B(n_4724),
.C(n_4747),
.Y(n_6230)
);

AOI22xp33_ASAP7_75t_L g6231 ( 
.A1(n_5192),
.A2(n_4771),
.B1(n_5139),
.B2(n_4495),
.Y(n_6231)
);

BUFx3_ASAP7_75t_L g6232 ( 
.A(n_5662),
.Y(n_6232)
);

NAND2x1p5_ASAP7_75t_L g6233 ( 
.A(n_5760),
.B(n_4481),
.Y(n_6233)
);

INVx1_ASAP7_75t_SL g6234 ( 
.A(n_5317),
.Y(n_6234)
);

INVx2_ASAP7_75t_SL g6235 ( 
.A(n_5760),
.Y(n_6235)
);

INVx2_ASAP7_75t_SL g6236 ( 
.A(n_5760),
.Y(n_6236)
);

AO21x2_ASAP7_75t_L g6237 ( 
.A1(n_5919),
.A2(n_4699),
.B(n_4694),
.Y(n_6237)
);

AOI21xp5_ASAP7_75t_L g6238 ( 
.A1(n_5769),
.A2(n_5422),
.B(n_5784),
.Y(n_6238)
);

OAI21xp5_ASAP7_75t_L g6239 ( 
.A1(n_5267),
.A2(n_4748),
.B(n_4730),
.Y(n_6239)
);

BUFx3_ASAP7_75t_L g6240 ( 
.A(n_5662),
.Y(n_6240)
);

OAI21x1_ASAP7_75t_L g6241 ( 
.A1(n_5290),
.A2(n_4588),
.B(n_4586),
.Y(n_6241)
);

CKINVDCx20_ASAP7_75t_R g6242 ( 
.A(n_5337),
.Y(n_6242)
);

NAND2xp5_ASAP7_75t_L g6243 ( 
.A(n_5916),
.B(n_4431),
.Y(n_6243)
);

OAI21x1_ASAP7_75t_L g6244 ( 
.A1(n_5290),
.A2(n_4594),
.B(n_4588),
.Y(n_6244)
);

INVx3_ASAP7_75t_L g6245 ( 
.A(n_5902),
.Y(n_6245)
);

OR2x2_ASAP7_75t_L g6246 ( 
.A(n_5236),
.B(n_4975),
.Y(n_6246)
);

OAI21x1_ASAP7_75t_L g6247 ( 
.A1(n_5990),
.A2(n_4595),
.B(n_4594),
.Y(n_6247)
);

OAI21x1_ASAP7_75t_L g6248 ( 
.A1(n_5990),
.A2(n_4595),
.B(n_4594),
.Y(n_6248)
);

OAI21xp5_ASAP7_75t_L g6249 ( 
.A1(n_5267),
.A2(n_4748),
.B(n_4730),
.Y(n_6249)
);

BUFx2_ASAP7_75t_L g6250 ( 
.A(n_5902),
.Y(n_6250)
);

INVx2_ASAP7_75t_L g6251 ( 
.A(n_5991),
.Y(n_6251)
);

INVx1_ASAP7_75t_L g6252 ( 
.A(n_5393),
.Y(n_6252)
);

OAI211xp5_ASAP7_75t_L g6253 ( 
.A1(n_5354),
.A2(n_4771),
.B(n_4726),
.C(n_5096),
.Y(n_6253)
);

NAND2xp5_ASAP7_75t_L g6254 ( 
.A(n_5213),
.B(n_4431),
.Y(n_6254)
);

OAI22xp5_ASAP7_75t_L g6255 ( 
.A1(n_5258),
.A2(n_4726),
.B1(n_4558),
.B2(n_4540),
.Y(n_6255)
);

OAI22xp5_ASAP7_75t_L g6256 ( 
.A1(n_5258),
.A2(n_4558),
.B1(n_4847),
.B2(n_4845),
.Y(n_6256)
);

AO21x2_ASAP7_75t_L g6257 ( 
.A1(n_5349),
.A2(n_4699),
.B(n_5102),
.Y(n_6257)
);

INVx2_ASAP7_75t_L g6258 ( 
.A(n_5991),
.Y(n_6258)
);

INVx1_ASAP7_75t_L g6259 ( 
.A(n_5393),
.Y(n_6259)
);

NOR2xp67_ASAP7_75t_SL g6260 ( 
.A(n_5281),
.B(n_4764),
.Y(n_6260)
);

INVx2_ASAP7_75t_L g6261 ( 
.A(n_5991),
.Y(n_6261)
);

OAI21x1_ASAP7_75t_L g6262 ( 
.A1(n_5742),
.A2(n_4599),
.B(n_4597),
.Y(n_6262)
);

AO31x2_ASAP7_75t_L g6263 ( 
.A1(n_5587),
.A2(n_4866),
.A3(n_4870),
.B(n_4831),
.Y(n_6263)
);

INVx1_ASAP7_75t_L g6264 ( 
.A(n_5398),
.Y(n_6264)
);

OA21x2_ASAP7_75t_L g6265 ( 
.A1(n_5284),
.A2(n_4612),
.B(n_4574),
.Y(n_6265)
);

BUFx6f_ASAP7_75t_L g6266 ( 
.A(n_5760),
.Y(n_6266)
);

INVx1_ASAP7_75t_L g6267 ( 
.A(n_5398),
.Y(n_6267)
);

BUFx3_ASAP7_75t_L g6268 ( 
.A(n_5903),
.Y(n_6268)
);

INVx4_ASAP7_75t_L g6269 ( 
.A(n_5262),
.Y(n_6269)
);

HB1xp67_ASAP7_75t_L g6270 ( 
.A(n_5550),
.Y(n_6270)
);

INVx1_ASAP7_75t_L g6271 ( 
.A(n_5399),
.Y(n_6271)
);

INVx4_ASAP7_75t_SL g6272 ( 
.A(n_5228),
.Y(n_6272)
);

OAI21x1_ASAP7_75t_L g6273 ( 
.A1(n_5245),
.A2(n_5390),
.B(n_5365),
.Y(n_6273)
);

OAI21x1_ASAP7_75t_L g6274 ( 
.A1(n_5245),
.A2(n_4574),
.B(n_4572),
.Y(n_6274)
);

INVx1_ASAP7_75t_L g6275 ( 
.A(n_5399),
.Y(n_6275)
);

AO21x2_ASAP7_75t_L g6276 ( 
.A1(n_5349),
.A2(n_4699),
.B(n_5102),
.Y(n_6276)
);

BUFx6f_ASAP7_75t_L g6277 ( 
.A(n_5760),
.Y(n_6277)
);

AND2x2_ASAP7_75t_L g6278 ( 
.A(n_5914),
.B(n_4402),
.Y(n_6278)
);

INVx1_ASAP7_75t_L g6279 ( 
.A(n_5404),
.Y(n_6279)
);

OAI21xp5_ASAP7_75t_L g6280 ( 
.A1(n_5166),
.A2(n_4474),
.B(n_4845),
.Y(n_6280)
);

AO21x2_ASAP7_75t_L g6281 ( 
.A1(n_5342),
.A2(n_5102),
.B(n_4674),
.Y(n_6281)
);

INVx1_ASAP7_75t_L g6282 ( 
.A(n_5404),
.Y(n_6282)
);

OAI21x1_ASAP7_75t_L g6283 ( 
.A1(n_5367),
.A2(n_5306),
.B(n_5504),
.Y(n_6283)
);

INVx2_ASAP7_75t_L g6284 ( 
.A(n_5718),
.Y(n_6284)
);

NOR2xp33_ASAP7_75t_SL g6285 ( 
.A(n_5689),
.B(n_5020),
.Y(n_6285)
);

OAI21xp5_ASAP7_75t_L g6286 ( 
.A1(n_5192),
.A2(n_4474),
.B(n_4856),
.Y(n_6286)
);

OAI21x1_ASAP7_75t_L g6287 ( 
.A1(n_5306),
.A2(n_5504),
.B(n_5320),
.Y(n_6287)
);

AOI22xp5_ASAP7_75t_L g6288 ( 
.A1(n_5190),
.A2(n_5020),
.B1(n_4849),
.B2(n_5099),
.Y(n_6288)
);

OA21x2_ASAP7_75t_L g6289 ( 
.A1(n_5260),
.A2(n_5278),
.B(n_5276),
.Y(n_6289)
);

NAND2xp5_ASAP7_75t_SL g6290 ( 
.A(n_5897),
.B(n_4481),
.Y(n_6290)
);

INVx1_ASAP7_75t_L g6291 ( 
.A(n_5408),
.Y(n_6291)
);

AOI221x1_ASAP7_75t_L g6292 ( 
.A1(n_5157),
.A2(n_4750),
.B1(n_4752),
.B2(n_4749),
.C(n_4745),
.Y(n_6292)
);

BUFx2_ASAP7_75t_L g6293 ( 
.A(n_5914),
.Y(n_6293)
);

INVx2_ASAP7_75t_L g6294 ( 
.A(n_5718),
.Y(n_6294)
);

OAI22xp5_ASAP7_75t_L g6295 ( 
.A1(n_5157),
.A2(n_4558),
.B1(n_4860),
.B2(n_4856),
.Y(n_6295)
);

AO21x2_ASAP7_75t_L g6296 ( 
.A1(n_5342),
.A2(n_4674),
.B(n_4673),
.Y(n_6296)
);

AOI21xp5_ASAP7_75t_L g6297 ( 
.A1(n_5784),
.A2(n_4849),
.B(n_4771),
.Y(n_6297)
);

AND2x2_ASAP7_75t_L g6298 ( 
.A(n_5914),
.B(n_4402),
.Y(n_6298)
);

OR2x2_ASAP7_75t_L g6299 ( 
.A(n_5236),
.B(n_4975),
.Y(n_6299)
);

OAI22xp33_ASAP7_75t_L g6300 ( 
.A1(n_5428),
.A2(n_4725),
.B1(n_4722),
.B2(n_4860),
.Y(n_6300)
);

HB1xp67_ASAP7_75t_L g6301 ( 
.A(n_5550),
.Y(n_6301)
);

INVx1_ASAP7_75t_L g6302 ( 
.A(n_5408),
.Y(n_6302)
);

A2O1A1Ixp33_ASAP7_75t_L g6303 ( 
.A1(n_5162),
.A2(n_4375),
.B(n_4722),
.C(n_4481),
.Y(n_6303)
);

INVx1_ASAP7_75t_L g6304 ( 
.A(n_5410),
.Y(n_6304)
);

INVx2_ASAP7_75t_L g6305 ( 
.A(n_5718),
.Y(n_6305)
);

OAI22xp5_ASAP7_75t_L g6306 ( 
.A1(n_5584),
.A2(n_5038),
.B1(n_4749),
.B2(n_4750),
.Y(n_6306)
);

AO32x2_ASAP7_75t_L g6307 ( 
.A1(n_5927),
.A2(n_4639),
.A3(n_4815),
.B1(n_4636),
.B2(n_4631),
.Y(n_6307)
);

NOR2xp33_ASAP7_75t_SL g6308 ( 
.A(n_5689),
.B(n_5059),
.Y(n_6308)
);

INVx1_ASAP7_75t_L g6309 ( 
.A(n_5410),
.Y(n_6309)
);

INVx2_ASAP7_75t_L g6310 ( 
.A(n_5718),
.Y(n_6310)
);

OAI21x1_ASAP7_75t_L g6311 ( 
.A1(n_5520),
.A2(n_5912),
.B(n_5338),
.Y(n_6311)
);

AO32x2_ASAP7_75t_L g6312 ( 
.A1(n_5958),
.A2(n_4639),
.A3(n_4815),
.B1(n_4636),
.B2(n_4631),
.Y(n_6312)
);

AOI21xp5_ASAP7_75t_L g6313 ( 
.A1(n_5733),
.A2(n_4771),
.B(n_4527),
.Y(n_6313)
);

INVx2_ASAP7_75t_L g6314 ( 
.A(n_5822),
.Y(n_6314)
);

INVx2_ASAP7_75t_L g6315 ( 
.A(n_5822),
.Y(n_6315)
);

INVx2_ASAP7_75t_L g6316 ( 
.A(n_5822),
.Y(n_6316)
);

INVx2_ASAP7_75t_SL g6317 ( 
.A(n_5837),
.Y(n_6317)
);

A2O1A1Ixp33_ASAP7_75t_L g6318 ( 
.A1(n_5145),
.A2(n_4375),
.B(n_4514),
.C(n_4481),
.Y(n_6318)
);

INVx8_ASAP7_75t_L g6319 ( 
.A(n_5834),
.Y(n_6319)
);

INVx3_ASAP7_75t_L g6320 ( 
.A(n_5914),
.Y(n_6320)
);

INVx1_ASAP7_75t_L g6321 ( 
.A(n_5429),
.Y(n_6321)
);

AO21x2_ASAP7_75t_L g6322 ( 
.A1(n_5287),
.A2(n_4938),
.B(n_4936),
.Y(n_6322)
);

INVx1_ASAP7_75t_L g6323 ( 
.A(n_5429),
.Y(n_6323)
);

AO21x2_ASAP7_75t_L g6324 ( 
.A1(n_5287),
.A2(n_4938),
.B(n_4936),
.Y(n_6324)
);

NAND2xp5_ASAP7_75t_L g6325 ( 
.A(n_5213),
.B(n_4431),
.Y(n_6325)
);

AO31x2_ASAP7_75t_L g6326 ( 
.A1(n_5656),
.A2(n_4888),
.A3(n_4892),
.B(n_4870),
.Y(n_6326)
);

OA21x2_ASAP7_75t_L g6327 ( 
.A1(n_5260),
.A2(n_4997),
.B(n_4996),
.Y(n_6327)
);

BUFx6f_ASAP7_75t_L g6328 ( 
.A(n_5837),
.Y(n_6328)
);

OAI21x1_ASAP7_75t_L g6329 ( 
.A1(n_5344),
.A2(n_4498),
.B(n_4488),
.Y(n_6329)
);

NAND2xp5_ASAP7_75t_L g6330 ( 
.A(n_5240),
.B(n_4431),
.Y(n_6330)
);

AOI21x1_ASAP7_75t_L g6331 ( 
.A1(n_5509),
.A2(n_4557),
.B(n_4460),
.Y(n_6331)
);

NAND2xp5_ASAP7_75t_L g6332 ( 
.A(n_5240),
.B(n_4431),
.Y(n_6332)
);

OR2x2_ASAP7_75t_L g6333 ( 
.A(n_5257),
.B(n_5914),
.Y(n_6333)
);

CKINVDCx16_ASAP7_75t_R g6334 ( 
.A(n_5551),
.Y(n_6334)
);

CKINVDCx5p33_ASAP7_75t_R g6335 ( 
.A(n_5159),
.Y(n_6335)
);

NAND2xp5_ASAP7_75t_L g6336 ( 
.A(n_5611),
.B(n_4431),
.Y(n_6336)
);

INVx1_ASAP7_75t_L g6337 ( 
.A(n_5440),
.Y(n_6337)
);

INVx1_ASAP7_75t_SL g6338 ( 
.A(n_5317),
.Y(n_6338)
);

OAI21x1_ASAP7_75t_SL g6339 ( 
.A1(n_5172),
.A2(n_5137),
.B(n_4752),
.Y(n_6339)
);

OR2x6_ASAP7_75t_L g6340 ( 
.A(n_5582),
.B(n_4527),
.Y(n_6340)
);

BUFx3_ASAP7_75t_L g6341 ( 
.A(n_5903),
.Y(n_6341)
);

OAI22xp5_ASAP7_75t_L g6342 ( 
.A1(n_5198),
.A2(n_5038),
.B1(n_4760),
.B2(n_4765),
.Y(n_6342)
);

AOI22xp33_ASAP7_75t_L g6343 ( 
.A1(n_5282),
.A2(n_5216),
.B1(n_5379),
.B2(n_5626),
.Y(n_6343)
);

BUFx6f_ASAP7_75t_L g6344 ( 
.A(n_5837),
.Y(n_6344)
);

AND2x2_ASAP7_75t_L g6345 ( 
.A(n_5855),
.B(n_4402),
.Y(n_6345)
);

INVx2_ASAP7_75t_SL g6346 ( 
.A(n_5837),
.Y(n_6346)
);

OAI21xp5_ASAP7_75t_L g6347 ( 
.A1(n_5961),
.A2(n_4474),
.B(n_4745),
.Y(n_6347)
);

AOI22xp33_ASAP7_75t_L g6348 ( 
.A1(n_5282),
.A2(n_4495),
.B1(n_4427),
.B2(n_4521),
.Y(n_6348)
);

OAI21x1_ASAP7_75t_L g6349 ( 
.A1(n_5435),
.A2(n_5448),
.B(n_5462),
.Y(n_6349)
);

INVx1_ASAP7_75t_L g6350 ( 
.A(n_5440),
.Y(n_6350)
);

NOR2xp33_ASAP7_75t_L g6351 ( 
.A(n_5469),
.B(n_4904),
.Y(n_6351)
);

INVx2_ASAP7_75t_L g6352 ( 
.A(n_5822),
.Y(n_6352)
);

AOI21x1_ASAP7_75t_L g6353 ( 
.A1(n_5532),
.A2(n_4557),
.B(n_4460),
.Y(n_6353)
);

AND2x2_ASAP7_75t_L g6354 ( 
.A(n_5855),
.B(n_4402),
.Y(n_6354)
);

BUFx2_ASAP7_75t_L g6355 ( 
.A(n_5694),
.Y(n_6355)
);

OAI21x1_ASAP7_75t_L g6356 ( 
.A1(n_5462),
.A2(n_5939),
.B(n_5436),
.Y(n_6356)
);

NAND2xp5_ASAP7_75t_L g6357 ( 
.A(n_5704),
.B(n_4431),
.Y(n_6357)
);

NOR2xp33_ASAP7_75t_L g6358 ( 
.A(n_5472),
.B(n_4904),
.Y(n_6358)
);

CKINVDCx5p33_ASAP7_75t_R g6359 ( 
.A(n_5237),
.Y(n_6359)
);

INVx2_ASAP7_75t_L g6360 ( 
.A(n_5817),
.Y(n_6360)
);

INVx2_ASAP7_75t_L g6361 ( 
.A(n_5817),
.Y(n_6361)
);

INVx1_ASAP7_75t_L g6362 ( 
.A(n_5449),
.Y(n_6362)
);

INVx2_ASAP7_75t_L g6363 ( 
.A(n_5817),
.Y(n_6363)
);

INVx1_ASAP7_75t_L g6364 ( 
.A(n_5449),
.Y(n_6364)
);

AO21x1_ASAP7_75t_L g6365 ( 
.A1(n_5216),
.A2(n_4765),
.B(n_4760),
.Y(n_6365)
);

INVx1_ASAP7_75t_L g6366 ( 
.A(n_5455),
.Y(n_6366)
);

INVx2_ASAP7_75t_L g6367 ( 
.A(n_5817),
.Y(n_6367)
);

CKINVDCx5p33_ASAP7_75t_R g6368 ( 
.A(n_5362),
.Y(n_6368)
);

OR2x2_ASAP7_75t_L g6369 ( 
.A(n_5257),
.B(n_4975),
.Y(n_6369)
);

O2A1O1Ixp33_ASAP7_75t_SL g6370 ( 
.A1(n_5217),
.A2(n_4490),
.B(n_4562),
.C(n_4458),
.Y(n_6370)
);

NAND3xp33_ASAP7_75t_L g6371 ( 
.A(n_5961),
.B(n_4784),
.C(n_4773),
.Y(n_6371)
);

INVx1_ASAP7_75t_L g6372 ( 
.A(n_5455),
.Y(n_6372)
);

OAI21x1_ASAP7_75t_L g6373 ( 
.A1(n_5436),
.A2(n_5363),
.B(n_5732),
.Y(n_6373)
);

OAI21xp5_ASAP7_75t_L g6374 ( 
.A1(n_5170),
.A2(n_4784),
.B(n_4773),
.Y(n_6374)
);

AOI22xp33_ASAP7_75t_L g6375 ( 
.A1(n_5379),
.A2(n_4495),
.B1(n_4427),
.B2(n_4521),
.Y(n_6375)
);

AND2x4_ASAP7_75t_L g6376 ( 
.A(n_5837),
.B(n_4481),
.Y(n_6376)
);

INVx3_ASAP7_75t_L g6377 ( 
.A(n_5597),
.Y(n_6377)
);

INVx3_ASAP7_75t_L g6378 ( 
.A(n_5597),
.Y(n_6378)
);

INVx2_ASAP7_75t_L g6379 ( 
.A(n_5817),
.Y(n_6379)
);

AND2x2_ASAP7_75t_L g6380 ( 
.A(n_5855),
.B(n_5128),
.Y(n_6380)
);

OA21x2_ASAP7_75t_L g6381 ( 
.A1(n_5276),
.A2(n_4938),
.B(n_4936),
.Y(n_6381)
);

BUFx6f_ASAP7_75t_L g6382 ( 
.A(n_5837),
.Y(n_6382)
);

INVx1_ASAP7_75t_L g6383 ( 
.A(n_5458),
.Y(n_6383)
);

INVx2_ASAP7_75t_L g6384 ( 
.A(n_5817),
.Y(n_6384)
);

OAI21x1_ASAP7_75t_L g6385 ( 
.A1(n_5355),
.A2(n_5988),
.B(n_5908),
.Y(n_6385)
);

INVx2_ASAP7_75t_L g6386 ( 
.A(n_5550),
.Y(n_6386)
);

AND2x2_ASAP7_75t_L g6387 ( 
.A(n_5855),
.B(n_5128),
.Y(n_6387)
);

BUFx8_ASAP7_75t_L g6388 ( 
.A(n_5856),
.Y(n_6388)
);

HB1xp67_ASAP7_75t_L g6389 ( 
.A(n_5550),
.Y(n_6389)
);

INVx1_ASAP7_75t_L g6390 ( 
.A(n_5458),
.Y(n_6390)
);

HB1xp67_ASAP7_75t_L g6391 ( 
.A(n_5593),
.Y(n_6391)
);

HB1xp67_ASAP7_75t_L g6392 ( 
.A(n_5593),
.Y(n_6392)
);

AOI21xp5_ASAP7_75t_L g6393 ( 
.A1(n_5726),
.A2(n_4527),
.B(n_5136),
.Y(n_6393)
);

BUFx3_ASAP7_75t_L g6394 ( 
.A(n_5903),
.Y(n_6394)
);

NAND2xp5_ASAP7_75t_L g6395 ( 
.A(n_5161),
.B(n_4431),
.Y(n_6395)
);

NOR2x1_ASAP7_75t_SL g6396 ( 
.A(n_5537),
.B(n_5059),
.Y(n_6396)
);

NAND2x1p5_ASAP7_75t_L g6397 ( 
.A(n_5887),
.B(n_4514),
.Y(n_6397)
);

AOI22xp33_ASAP7_75t_L g6398 ( 
.A1(n_5196),
.A2(n_4495),
.B1(n_4427),
.B2(n_4590),
.Y(n_6398)
);

AND2x2_ASAP7_75t_L g6399 ( 
.A(n_5855),
.B(n_5128),
.Y(n_6399)
);

INVx1_ASAP7_75t_SL g6400 ( 
.A(n_5378),
.Y(n_6400)
);

INVx1_ASAP7_75t_L g6401 ( 
.A(n_5481),
.Y(n_6401)
);

OAI22xp5_ASAP7_75t_L g6402 ( 
.A1(n_5428),
.A2(n_4792),
.B1(n_4794),
.B2(n_4786),
.Y(n_6402)
);

AOI22xp33_ASAP7_75t_L g6403 ( 
.A1(n_5196),
.A2(n_4495),
.B1(n_4427),
.B2(n_4590),
.Y(n_6403)
);

AOI22xp33_ASAP7_75t_L g6404 ( 
.A1(n_5425),
.A2(n_4427),
.B1(n_4707),
.B2(n_4590),
.Y(n_6404)
);

OR2x2_ASAP7_75t_L g6405 ( 
.A(n_6013),
.B(n_4975),
.Y(n_6405)
);

INVx2_ASAP7_75t_L g6406 ( 
.A(n_5593),
.Y(n_6406)
);

INVx3_ASAP7_75t_L g6407 ( 
.A(n_5597),
.Y(n_6407)
);

AOI21x1_ASAP7_75t_L g6408 ( 
.A1(n_5532),
.A2(n_4557),
.B(n_4460),
.Y(n_6408)
);

INVx2_ASAP7_75t_SL g6409 ( 
.A(n_5887),
.Y(n_6409)
);

BUFx2_ASAP7_75t_L g6410 ( 
.A(n_5694),
.Y(n_6410)
);

INVx6_ASAP7_75t_L g6411 ( 
.A(n_5811),
.Y(n_6411)
);

INVx1_ASAP7_75t_L g6412 ( 
.A(n_5481),
.Y(n_6412)
);

NAND2xp5_ASAP7_75t_L g6413 ( 
.A(n_5161),
.B(n_5092),
.Y(n_6413)
);

INVx1_ASAP7_75t_L g6414 ( 
.A(n_5488),
.Y(n_6414)
);

INVx2_ASAP7_75t_L g6415 ( 
.A(n_5593),
.Y(n_6415)
);

HB1xp67_ASAP7_75t_L g6416 ( 
.A(n_5593),
.Y(n_6416)
);

AOI221xp5_ASAP7_75t_L g6417 ( 
.A1(n_5402),
.A2(n_4794),
.B1(n_4796),
.B2(n_4792),
.C(n_4786),
.Y(n_6417)
);

AOI21x1_ASAP7_75t_L g6418 ( 
.A1(n_5841),
.A2(n_4557),
.B(n_4460),
.Y(n_6418)
);

BUFx6f_ASAP7_75t_L g6419 ( 
.A(n_5887),
.Y(n_6419)
);

AOI22xp5_ASAP7_75t_L g6420 ( 
.A1(n_5517),
.A2(n_5099),
.B1(n_3009),
.B2(n_3014),
.Y(n_6420)
);

INVx1_ASAP7_75t_L g6421 ( 
.A(n_5488),
.Y(n_6421)
);

BUFx3_ASAP7_75t_L g6422 ( 
.A(n_5903),
.Y(n_6422)
);

AND2x4_ASAP7_75t_L g6423 ( 
.A(n_5887),
.B(n_4514),
.Y(n_6423)
);

AOI22xp5_ASAP7_75t_L g6424 ( 
.A1(n_5316),
.A2(n_5099),
.B1(n_3009),
.B2(n_3014),
.Y(n_6424)
);

OAI21xp5_ASAP7_75t_L g6425 ( 
.A1(n_5476),
.A2(n_4797),
.B(n_4796),
.Y(n_6425)
);

AND2x4_ASAP7_75t_L g6426 ( 
.A(n_5887),
.B(n_4514),
.Y(n_6426)
);

BUFx2_ASAP7_75t_R g6427 ( 
.A(n_5169),
.Y(n_6427)
);

OAI22xp5_ASAP7_75t_L g6428 ( 
.A1(n_5321),
.A2(n_4802),
.B1(n_4803),
.B2(n_4797),
.Y(n_6428)
);

INVx1_ASAP7_75t_L g6429 ( 
.A(n_5519),
.Y(n_6429)
);

INVx1_ASAP7_75t_L g6430 ( 
.A(n_5519),
.Y(n_6430)
);

OAI21x1_ASAP7_75t_SL g6431 ( 
.A1(n_5205),
.A2(n_5137),
.B(n_4803),
.Y(n_6431)
);

OAI21x1_ASAP7_75t_SL g6432 ( 
.A1(n_5183),
.A2(n_4804),
.B(n_4802),
.Y(n_6432)
);

INVx1_ASAP7_75t_L g6433 ( 
.A(n_5523),
.Y(n_6433)
);

A2O1A1Ixp33_ASAP7_75t_L g6434 ( 
.A1(n_5145),
.A2(n_4886),
.B(n_4514),
.C(n_4804),
.Y(n_6434)
);

INVx3_ASAP7_75t_L g6435 ( 
.A(n_5597),
.Y(n_6435)
);

A2O1A1Ixp33_ASAP7_75t_L g6436 ( 
.A1(n_5374),
.A2(n_5759),
.B(n_5534),
.C(n_5238),
.Y(n_6436)
);

INVx4_ASAP7_75t_L g6437 ( 
.A(n_5834),
.Y(n_6437)
);

INVx1_ASAP7_75t_L g6438 ( 
.A(n_5523),
.Y(n_6438)
);

NAND2xp5_ASAP7_75t_L g6439 ( 
.A(n_5174),
.B(n_5092),
.Y(n_6439)
);

INVx2_ASAP7_75t_L g6440 ( 
.A(n_5593),
.Y(n_6440)
);

OAI21x1_ASAP7_75t_L g6441 ( 
.A1(n_5521),
.A2(n_4658),
.B(n_4669),
.Y(n_6441)
);

O2A1O1Ixp33_ASAP7_75t_SL g6442 ( 
.A1(n_5330),
.A2(n_4490),
.B(n_4562),
.C(n_4458),
.Y(n_6442)
);

INVx1_ASAP7_75t_L g6443 ( 
.A(n_5535),
.Y(n_6443)
);

OAI22xp5_ASAP7_75t_L g6444 ( 
.A1(n_5374),
.A2(n_5694),
.B1(n_5296),
.B2(n_5664),
.Y(n_6444)
);

INVx2_ASAP7_75t_L g6445 ( 
.A(n_5855),
.Y(n_6445)
);

INVx4_ASAP7_75t_SL g6446 ( 
.A(n_5228),
.Y(n_6446)
);

NOR2x1_ASAP7_75t_SL g6447 ( 
.A(n_5537),
.B(n_5143),
.Y(n_6447)
);

OAI21xp5_ASAP7_75t_L g6448 ( 
.A1(n_5252),
.A2(n_5072),
.B(n_4398),
.Y(n_6448)
);

OAI22xp5_ASAP7_75t_L g6449 ( 
.A1(n_5694),
.A2(n_5072),
.B1(n_5055),
.B2(n_5043),
.Y(n_6449)
);

INVx1_ASAP7_75t_L g6450 ( 
.A(n_5535),
.Y(n_6450)
);

A2O1A1Ixp33_ASAP7_75t_L g6451 ( 
.A1(n_5534),
.A2(n_4886),
.B(n_4514),
.C(n_4904),
.Y(n_6451)
);

BUFx4_ASAP7_75t_SL g6452 ( 
.A(n_5286),
.Y(n_6452)
);

AOI221xp5_ASAP7_75t_L g6453 ( 
.A1(n_5402),
.A2(n_4906),
.B1(n_4696),
.B2(n_4700),
.C(n_4697),
.Y(n_6453)
);

AOI22xp33_ASAP7_75t_L g6454 ( 
.A1(n_5296),
.A2(n_4707),
.B1(n_4906),
.B2(n_4775),
.Y(n_6454)
);

INVx1_ASAP7_75t_L g6455 ( 
.A(n_5553),
.Y(n_6455)
);

AND3x2_ASAP7_75t_L g6456 ( 
.A(n_5439),
.B(n_4906),
.C(n_5120),
.Y(n_6456)
);

CKINVDCx11_ASAP7_75t_R g6457 ( 
.A(n_5199),
.Y(n_6457)
);

NAND2x1p5_ASAP7_75t_L g6458 ( 
.A(n_5887),
.B(n_4514),
.Y(n_6458)
);

AOI21x1_ASAP7_75t_L g6459 ( 
.A1(n_5841),
.A2(n_4557),
.B(n_4460),
.Y(n_6459)
);

NAND3xp33_ASAP7_75t_L g6460 ( 
.A(n_5656),
.B(n_4696),
.C(n_4692),
.Y(n_6460)
);

INVx2_ASAP7_75t_SL g6461 ( 
.A(n_6008),
.Y(n_6461)
);

INVx2_ASAP7_75t_L g6462 ( 
.A(n_5985),
.Y(n_6462)
);

OAI221xp5_ASAP7_75t_L g6463 ( 
.A1(n_5407),
.A2(n_4857),
.B1(n_4769),
.B2(n_4766),
.C(n_4398),
.Y(n_6463)
);

AOI22x1_ASAP7_75t_L g6464 ( 
.A1(n_5186),
.A2(n_5004),
.B1(n_5048),
.B2(n_4954),
.Y(n_6464)
);

INVx1_ASAP7_75t_L g6465 ( 
.A(n_5553),
.Y(n_6465)
);

NAND2xp5_ASAP7_75t_L g6466 ( 
.A(n_5174),
.B(n_5120),
.Y(n_6466)
);

AND2x2_ASAP7_75t_L g6467 ( 
.A(n_5694),
.B(n_5128),
.Y(n_6467)
);

INVx1_ASAP7_75t_L g6468 ( 
.A(n_5568),
.Y(n_6468)
);

CKINVDCx20_ASAP7_75t_R g6469 ( 
.A(n_5885),
.Y(n_6469)
);

NOR2xp33_ASAP7_75t_L g6470 ( 
.A(n_5312),
.B(n_4676),
.Y(n_6470)
);

INVx1_ASAP7_75t_L g6471 ( 
.A(n_5568),
.Y(n_6471)
);

BUFx3_ASAP7_75t_L g6472 ( 
.A(n_5940),
.Y(n_6472)
);

AOI21xp5_ASAP7_75t_L g6473 ( 
.A1(n_5726),
.A2(n_4527),
.B(n_5136),
.Y(n_6473)
);

NAND2x1p5_ASAP7_75t_L g6474 ( 
.A(n_6008),
.B(n_4514),
.Y(n_6474)
);

OA21x2_ASAP7_75t_L g6475 ( 
.A1(n_5461),
.A2(n_5132),
.B(n_5010),
.Y(n_6475)
);

INVx2_ASAP7_75t_SL g6476 ( 
.A(n_6008),
.Y(n_6476)
);

OAI22xp5_ASAP7_75t_L g6477 ( 
.A1(n_5664),
.A2(n_5055),
.B1(n_4686),
.B2(n_4691),
.Y(n_6477)
);

OAI22xp5_ASAP7_75t_L g6478 ( 
.A1(n_5316),
.A2(n_4686),
.B1(n_4691),
.B2(n_4692),
.Y(n_6478)
);

INVx2_ASAP7_75t_L g6479 ( 
.A(n_5985),
.Y(n_6479)
);

INVx1_ASAP7_75t_L g6480 ( 
.A(n_5581),
.Y(n_6480)
);

OAI22xp33_ASAP7_75t_L g6481 ( 
.A1(n_5950),
.A2(n_4707),
.B1(n_4738),
.B2(n_4570),
.Y(n_6481)
);

OAI21x1_ASAP7_75t_L g6482 ( 
.A1(n_5542),
.A2(n_5543),
.B(n_5446),
.Y(n_6482)
);

AND2x2_ASAP7_75t_L g6483 ( 
.A(n_6019),
.B(n_5128),
.Y(n_6483)
);

NOR2xp33_ASAP7_75t_L g6484 ( 
.A(n_5312),
.B(n_4676),
.Y(n_6484)
);

O2A1O1Ixp33_ASAP7_75t_L g6485 ( 
.A1(n_5231),
.A2(n_5119),
.B(n_4697),
.C(n_4700),
.Y(n_6485)
);

A2O1A1Ixp33_ASAP7_75t_L g6486 ( 
.A1(n_5893),
.A2(n_4886),
.B(n_4738),
.C(n_4570),
.Y(n_6486)
);

BUFx6f_ASAP7_75t_L g6487 ( 
.A(n_6008),
.Y(n_6487)
);

OR2x6_ASAP7_75t_L g6488 ( 
.A(n_5582),
.B(n_4527),
.Y(n_6488)
);

INVx2_ASAP7_75t_L g6489 ( 
.A(n_5985),
.Y(n_6489)
);

INVx2_ASAP7_75t_L g6490 ( 
.A(n_5985),
.Y(n_6490)
);

OAI21xp5_ASAP7_75t_L g6491 ( 
.A1(n_5310),
.A2(n_5119),
.B(n_5115),
.Y(n_6491)
);

NOR2xp33_ASAP7_75t_L g6492 ( 
.A(n_5336),
.B(n_5089),
.Y(n_6492)
);

OAI21x1_ASAP7_75t_L g6493 ( 
.A1(n_5613),
.A2(n_5164),
.B(n_5843),
.Y(n_6493)
);

OAI21x1_ASAP7_75t_SL g6494 ( 
.A1(n_5524),
.A2(n_4998),
.B(n_4994),
.Y(n_6494)
);

OA21x2_ASAP7_75t_L g6495 ( 
.A1(n_5477),
.A2(n_5132),
.B(n_5026),
.Y(n_6495)
);

INVx2_ASAP7_75t_L g6496 ( 
.A(n_6029),
.Y(n_6496)
);

OAI21x1_ASAP7_75t_L g6497 ( 
.A1(n_5843),
.A2(n_5968),
.B(n_5957),
.Y(n_6497)
);

BUFx2_ASAP7_75t_L g6498 ( 
.A(n_6019),
.Y(n_6498)
);

INVx2_ASAP7_75t_L g6499 ( 
.A(n_6029),
.Y(n_6499)
);

INVx1_ASAP7_75t_SL g6500 ( 
.A(n_5378),
.Y(n_6500)
);

INVx1_ASAP7_75t_L g6501 ( 
.A(n_5581),
.Y(n_6501)
);

INVxp67_ASAP7_75t_SL g6502 ( 
.A(n_5736),
.Y(n_6502)
);

OA21x2_ASAP7_75t_L g6503 ( 
.A1(n_5477),
.A2(n_5132),
.B(n_5026),
.Y(n_6503)
);

NAND2x1p5_ASAP7_75t_L g6504 ( 
.A(n_6008),
.B(n_4886),
.Y(n_6504)
);

AOI221xp5_ASAP7_75t_L g6505 ( 
.A1(n_5294),
.A2(n_4640),
.B1(n_4413),
.B2(n_4435),
.C(n_4429),
.Y(n_6505)
);

INVx1_ASAP7_75t_L g6506 ( 
.A(n_5599),
.Y(n_6506)
);

INVx2_ASAP7_75t_L g6507 ( 
.A(n_6029),
.Y(n_6507)
);

OA21x2_ASAP7_75t_L g6508 ( 
.A1(n_5771),
.A2(n_5567),
.B(n_5682),
.Y(n_6508)
);

BUFx4f_ASAP7_75t_L g6509 ( 
.A(n_5171),
.Y(n_6509)
);

AND2x2_ASAP7_75t_L g6510 ( 
.A(n_6019),
.B(n_5128),
.Y(n_6510)
);

INVx1_ASAP7_75t_L g6511 ( 
.A(n_5599),
.Y(n_6511)
);

O2A1O1Ixp33_ASAP7_75t_SL g6512 ( 
.A1(n_5442),
.A2(n_4998),
.B(n_5013),
.C(n_4994),
.Y(n_6512)
);

BUFx8_ASAP7_75t_SL g6513 ( 
.A(n_5286),
.Y(n_6513)
);

AO21x2_ASAP7_75t_L g6514 ( 
.A1(n_5738),
.A2(n_5954),
.B(n_5300),
.Y(n_6514)
);

INVx1_ASAP7_75t_L g6515 ( 
.A(n_5601),
.Y(n_6515)
);

INVx1_ASAP7_75t_L g6516 ( 
.A(n_5601),
.Y(n_6516)
);

INVx1_ASAP7_75t_L g6517 ( 
.A(n_5630),
.Y(n_6517)
);

OA21x2_ASAP7_75t_L g6518 ( 
.A1(n_5771),
.A2(n_5936),
.B(n_5559),
.Y(n_6518)
);

NAND2xp5_ASAP7_75t_SL g6519 ( 
.A(n_5897),
.B(n_4886),
.Y(n_6519)
);

OAI21xp5_ASAP7_75t_L g6520 ( 
.A1(n_5797),
.A2(n_5115),
.B(n_4651),
.Y(n_6520)
);

AOI22xp33_ASAP7_75t_SL g6521 ( 
.A1(n_5950),
.A2(n_4886),
.B1(n_5141),
.B2(n_5136),
.Y(n_6521)
);

INVx1_ASAP7_75t_L g6522 ( 
.A(n_5630),
.Y(n_6522)
);

AND2x2_ASAP7_75t_L g6523 ( 
.A(n_6019),
.B(n_5128),
.Y(n_6523)
);

HB1xp67_ASAP7_75t_L g6524 ( 
.A(n_5149),
.Y(n_6524)
);

OAI22xp5_ASAP7_75t_L g6525 ( 
.A1(n_5897),
.A2(n_4868),
.B1(n_4663),
.B2(n_5013),
.Y(n_6525)
);

AOI21xp5_ASAP7_75t_L g6526 ( 
.A1(n_5740),
.A2(n_5733),
.B(n_5341),
.Y(n_6526)
);

INVx2_ASAP7_75t_L g6527 ( 
.A(n_6029),
.Y(n_6527)
);

AND2x4_ASAP7_75t_L g6528 ( 
.A(n_6008),
.B(n_4886),
.Y(n_6528)
);

INVx2_ASAP7_75t_L g6529 ( 
.A(n_5806),
.Y(n_6529)
);

INVx2_ASAP7_75t_L g6530 ( 
.A(n_5806),
.Y(n_6530)
);

AO31x2_ASAP7_75t_L g6531 ( 
.A1(n_5886),
.A2(n_4888),
.A3(n_4892),
.B(n_4870),
.Y(n_6531)
);

INVx1_ASAP7_75t_L g6532 ( 
.A(n_5653),
.Y(n_6532)
);

CKINVDCx5p33_ASAP7_75t_R g6533 ( 
.A(n_6006),
.Y(n_6533)
);

OR2x6_ASAP7_75t_L g6534 ( 
.A(n_5552),
.B(n_4527),
.Y(n_6534)
);

INVx1_ASAP7_75t_L g6535 ( 
.A(n_5653),
.Y(n_6535)
);

AND2x4_ASAP7_75t_L g6536 ( 
.A(n_5264),
.B(n_4886),
.Y(n_6536)
);

INVx2_ASAP7_75t_L g6537 ( 
.A(n_5806),
.Y(n_6537)
);

OAI21xp5_ASAP7_75t_L g6538 ( 
.A1(n_5456),
.A2(n_4914),
.B(n_4913),
.Y(n_6538)
);

AND2x4_ASAP7_75t_L g6539 ( 
.A(n_5264),
.B(n_5143),
.Y(n_6539)
);

AOI22xp33_ASAP7_75t_L g6540 ( 
.A1(n_5513),
.A2(n_4775),
.B1(n_4741),
.B2(n_5099),
.Y(n_6540)
);

BUFx3_ASAP7_75t_L g6541 ( 
.A(n_5940),
.Y(n_6541)
);

AND2x2_ASAP7_75t_L g6542 ( 
.A(n_6019),
.B(n_5575),
.Y(n_6542)
);

INVx1_ASAP7_75t_L g6543 ( 
.A(n_5657),
.Y(n_6543)
);

BUFx6f_ASAP7_75t_L g6544 ( 
.A(n_5965),
.Y(n_6544)
);

INVx2_ASAP7_75t_L g6545 ( 
.A(n_5806),
.Y(n_6545)
);

OAI22xp33_ASAP7_75t_L g6546 ( 
.A1(n_5489),
.A2(n_4766),
.B1(n_4857),
.B2(n_4769),
.Y(n_6546)
);

INVx1_ASAP7_75t_L g6547 ( 
.A(n_5657),
.Y(n_6547)
);

NAND2xp5_ASAP7_75t_L g6548 ( 
.A(n_5175),
.B(n_4437),
.Y(n_6548)
);

NAND2x1p5_ASAP7_75t_L g6549 ( 
.A(n_5756),
.B(n_5143),
.Y(n_6549)
);

OAI22xp33_ASAP7_75t_L g6550 ( 
.A1(n_5489),
.A2(n_4766),
.B1(n_4857),
.B2(n_4769),
.Y(n_6550)
);

BUFx2_ASAP7_75t_L g6551 ( 
.A(n_5537),
.Y(n_6551)
);

INVx1_ASAP7_75t_L g6552 ( 
.A(n_5667),
.Y(n_6552)
);

INVx4_ASAP7_75t_SL g6553 ( 
.A(n_5228),
.Y(n_6553)
);

BUFx12f_ASAP7_75t_L g6554 ( 
.A(n_5212),
.Y(n_6554)
);

AND2x2_ASAP7_75t_L g6555 ( 
.A(n_5575),
.B(n_5128),
.Y(n_6555)
);

OAI22xp33_ASAP7_75t_L g6556 ( 
.A1(n_5497),
.A2(n_4775),
.B1(n_4741),
.B2(n_5143),
.Y(n_6556)
);

NOR2xp33_ASAP7_75t_SL g6557 ( 
.A(n_5147),
.B(n_5143),
.Y(n_6557)
);

BUFx2_ASAP7_75t_L g6558 ( 
.A(n_5537),
.Y(n_6558)
);

AND2x2_ASAP7_75t_L g6559 ( 
.A(n_5605),
.B(n_4975),
.Y(n_6559)
);

A2O1A1Ixp33_ASAP7_75t_L g6560 ( 
.A1(n_5893),
.A2(n_5143),
.B(n_4880),
.C(n_4775),
.Y(n_6560)
);

AND2x2_ASAP7_75t_L g6561 ( 
.A(n_5605),
.B(n_4975),
.Y(n_6561)
);

INVx1_ASAP7_75t_L g6562 ( 
.A(n_5667),
.Y(n_6562)
);

INVx1_ASAP7_75t_L g6563 ( 
.A(n_5671),
.Y(n_6563)
);

CKINVDCx16_ASAP7_75t_R g6564 ( 
.A(n_5439),
.Y(n_6564)
);

AOI21xp5_ASAP7_75t_L g6565 ( 
.A1(n_5740),
.A2(n_5141),
.B(n_5136),
.Y(n_6565)
);

NAND2xp5_ASAP7_75t_L g6566 ( 
.A(n_5175),
.B(n_4437),
.Y(n_6566)
);

INVx2_ASAP7_75t_L g6567 ( 
.A(n_5806),
.Y(n_6567)
);

INVx2_ASAP7_75t_L g6568 ( 
.A(n_5806),
.Y(n_6568)
);

NOR2xp33_ASAP7_75t_L g6569 ( 
.A(n_5336),
.B(n_5089),
.Y(n_6569)
);

INVx1_ASAP7_75t_L g6570 ( 
.A(n_5671),
.Y(n_6570)
);

AO21x1_ASAP7_75t_L g6571 ( 
.A1(n_5674),
.A2(n_5024),
.B(n_5021),
.Y(n_6571)
);

INVx2_ASAP7_75t_L g6572 ( 
.A(n_5167),
.Y(n_6572)
);

NAND2xp5_ASAP7_75t_SL g6573 ( 
.A(n_5897),
.B(n_5143),
.Y(n_6573)
);

OR2x6_ASAP7_75t_L g6574 ( 
.A(n_5552),
.B(n_4954),
.Y(n_6574)
);

INVx1_ASAP7_75t_L g6575 ( 
.A(n_5672),
.Y(n_6575)
);

OR2x6_ASAP7_75t_L g6576 ( 
.A(n_5552),
.B(n_4954),
.Y(n_6576)
);

NOR2xp33_ASAP7_75t_L g6577 ( 
.A(n_5388),
.B(n_5089),
.Y(n_6577)
);

A2O1A1Ixp33_ASAP7_75t_L g6578 ( 
.A1(n_5513),
.A2(n_4880),
.B(n_4775),
.C(n_4741),
.Y(n_6578)
);

INVx1_ASAP7_75t_L g6579 ( 
.A(n_5672),
.Y(n_6579)
);

INVx1_ASAP7_75t_L g6580 ( 
.A(n_5673),
.Y(n_6580)
);

OAI21x1_ASAP7_75t_L g6581 ( 
.A1(n_5826),
.A2(n_5827),
.B(n_5560),
.Y(n_6581)
);

NAND2xp5_ASAP7_75t_L g6582 ( 
.A(n_5207),
.B(n_4437),
.Y(n_6582)
);

NAND2xp5_ASAP7_75t_L g6583 ( 
.A(n_5253),
.B(n_4437),
.Y(n_6583)
);

CKINVDCx6p67_ASAP7_75t_R g6584 ( 
.A(n_5199),
.Y(n_6584)
);

BUFx2_ASAP7_75t_L g6585 ( 
.A(n_5537),
.Y(n_6585)
);

INVx1_ASAP7_75t_L g6586 ( 
.A(n_5673),
.Y(n_6586)
);

AO21x1_ASAP7_75t_L g6587 ( 
.A1(n_5674),
.A2(n_5024),
.B(n_5021),
.Y(n_6587)
);

AOI22xp33_ASAP7_75t_L g6588 ( 
.A1(n_5395),
.A2(n_5255),
.B1(n_5401),
.B2(n_5683),
.Y(n_6588)
);

INVx4_ASAP7_75t_SL g6589 ( 
.A(n_5228),
.Y(n_6589)
);

OAI221xp5_ASAP7_75t_L g6590 ( 
.A1(n_5407),
.A2(n_4640),
.B1(n_4913),
.B2(n_4928),
.C(n_4914),
.Y(n_6590)
);

AOI21xp33_ASAP7_75t_L g6591 ( 
.A1(n_5640),
.A2(n_5083),
.B(n_5074),
.Y(n_6591)
);

AO32x2_ASAP7_75t_L g6592 ( 
.A1(n_5958),
.A2(n_4636),
.A3(n_4815),
.B1(n_4639),
.B2(n_4631),
.Y(n_6592)
);

OR2x6_ASAP7_75t_L g6593 ( 
.A(n_5552),
.B(n_5004),
.Y(n_6593)
);

AND2x4_ASAP7_75t_L g6594 ( 
.A(n_5264),
.B(n_4496),
.Y(n_6594)
);

AND2x2_ASAP7_75t_L g6595 ( 
.A(n_5932),
.B(n_4975),
.Y(n_6595)
);

INVx2_ASAP7_75t_L g6596 ( 
.A(n_5167),
.Y(n_6596)
);

AND2x2_ASAP7_75t_L g6597 ( 
.A(n_5932),
.B(n_4975),
.Y(n_6597)
);

NOR2xp33_ASAP7_75t_L g6598 ( 
.A(n_5388),
.B(n_5089),
.Y(n_6598)
);

NAND2xp5_ASAP7_75t_L g6599 ( 
.A(n_5490),
.B(n_4437),
.Y(n_6599)
);

BUFx3_ASAP7_75t_L g6600 ( 
.A(n_5940),
.Y(n_6600)
);

OAI21xp5_ASAP7_75t_L g6601 ( 
.A1(n_5456),
.A2(n_4939),
.B(n_4928),
.Y(n_6601)
);

OAI21xp5_ASAP7_75t_L g6602 ( 
.A1(n_5248),
.A2(n_4944),
.B(n_4939),
.Y(n_6602)
);

INVx2_ASAP7_75t_L g6603 ( 
.A(n_5167),
.Y(n_6603)
);

INVx1_ASAP7_75t_SL g6604 ( 
.A(n_5380),
.Y(n_6604)
);

OR2x2_ASAP7_75t_L g6605 ( 
.A(n_6013),
.B(n_4976),
.Y(n_6605)
);

NAND2xp5_ASAP7_75t_L g6606 ( 
.A(n_5490),
.B(n_4437),
.Y(n_6606)
);

OA21x2_ASAP7_75t_L g6607 ( 
.A1(n_5596),
.A2(n_5052),
.B(n_5051),
.Y(n_6607)
);

OR2x6_ASAP7_75t_L g6608 ( 
.A(n_5552),
.B(n_5004),
.Y(n_6608)
);

OA21x2_ASAP7_75t_L g6609 ( 
.A1(n_5772),
.A2(n_5052),
.B(n_5051),
.Y(n_6609)
);

NAND2xp5_ASAP7_75t_L g6610 ( 
.A(n_5577),
.B(n_4437),
.Y(n_6610)
);

AOI22xp5_ASAP7_75t_L g6611 ( 
.A1(n_5497),
.A2(n_3009),
.B1(n_3014),
.B2(n_4880),
.Y(n_6611)
);

INVxp67_ASAP7_75t_SL g6612 ( 
.A(n_5235),
.Y(n_6612)
);

OAI21x1_ASAP7_75t_SL g6613 ( 
.A1(n_5524),
.A2(n_5032),
.B(n_4873),
.Y(n_6613)
);

AOI21x1_ASAP7_75t_L g6614 ( 
.A1(n_5463),
.A2(n_4671),
.B(n_4598),
.Y(n_6614)
);

INVx1_ASAP7_75t_L g6615 ( 
.A(n_5680),
.Y(n_6615)
);

INVx2_ASAP7_75t_SL g6616 ( 
.A(n_5556),
.Y(n_6616)
);

INVx1_ASAP7_75t_L g6617 ( 
.A(n_5680),
.Y(n_6617)
);

AND2x4_ASAP7_75t_L g6618 ( 
.A(n_5264),
.B(n_4619),
.Y(n_6618)
);

AND2x4_ASAP7_75t_L g6619 ( 
.A(n_5264),
.B(n_4619),
.Y(n_6619)
);

NAND2xp33_ASAP7_75t_SL g6620 ( 
.A(n_5199),
.B(n_4619),
.Y(n_6620)
);

AND2x2_ASAP7_75t_L g6621 ( 
.A(n_5493),
.B(n_5539),
.Y(n_6621)
);

INVx2_ASAP7_75t_L g6622 ( 
.A(n_5185),
.Y(n_6622)
);

INVx2_ASAP7_75t_L g6623 ( 
.A(n_5185),
.Y(n_6623)
);

INVx2_ASAP7_75t_L g6624 ( 
.A(n_5185),
.Y(n_6624)
);

AOI21xp5_ASAP7_75t_L g6625 ( 
.A1(n_5341),
.A2(n_5281),
.B(n_5325),
.Y(n_6625)
);

HB1xp67_ASAP7_75t_L g6626 ( 
.A(n_5351),
.Y(n_6626)
);

OA21x2_ASAP7_75t_L g6627 ( 
.A1(n_5772),
.A2(n_5052),
.B(n_5051),
.Y(n_6627)
);

AND2x4_ASAP7_75t_L g6628 ( 
.A(n_5706),
.B(n_4619),
.Y(n_6628)
);

AO21x2_ASAP7_75t_L g6629 ( 
.A1(n_5749),
.A2(n_5018),
.B(n_5008),
.Y(n_6629)
);

AO31x2_ASAP7_75t_L g6630 ( 
.A1(n_5966),
.A2(n_5982),
.A3(n_5931),
.B(n_5531),
.Y(n_6630)
);

HB1xp67_ASAP7_75t_L g6631 ( 
.A(n_5451),
.Y(n_6631)
);

CKINVDCx5p33_ASAP7_75t_R g6632 ( 
.A(n_5375),
.Y(n_6632)
);

OAI21x1_ASAP7_75t_L g6633 ( 
.A1(n_5978),
.A2(n_5463),
.B(n_5382),
.Y(n_6633)
);

AOI22xp33_ASAP7_75t_L g6634 ( 
.A1(n_5401),
.A2(n_4741),
.B1(n_4880),
.B2(n_4410),
.Y(n_6634)
);

INVx1_ASAP7_75t_SL g6635 ( 
.A(n_5380),
.Y(n_6635)
);

INVx1_ASAP7_75t_L g6636 ( 
.A(n_5693),
.Y(n_6636)
);

CKINVDCx11_ASAP7_75t_R g6637 ( 
.A(n_5251),
.Y(n_6637)
);

INVx1_ASAP7_75t_L g6638 ( 
.A(n_5693),
.Y(n_6638)
);

AND2x2_ASAP7_75t_L g6639 ( 
.A(n_5493),
.B(n_4976),
.Y(n_6639)
);

AO21x2_ASAP7_75t_L g6640 ( 
.A1(n_5721),
.A2(n_5018),
.B(n_5008),
.Y(n_6640)
);

HB1xp67_ASAP7_75t_L g6641 ( 
.A(n_5727),
.Y(n_6641)
);

O2A1O1Ixp33_ASAP7_75t_L g6642 ( 
.A1(n_5413),
.A2(n_4663),
.B(n_4946),
.C(n_4944),
.Y(n_6642)
);

O2A1O1Ixp33_ASAP7_75t_SL g6643 ( 
.A1(n_5431),
.A2(n_5032),
.B(n_5083),
.C(n_5074),
.Y(n_6643)
);

OAI21x1_ASAP7_75t_L g6644 ( 
.A1(n_5346),
.A2(n_5621),
.B(n_5616),
.Y(n_6644)
);

OAI21x1_ASAP7_75t_L g6645 ( 
.A1(n_5616),
.A2(n_5621),
.B(n_5397),
.Y(n_6645)
);

INVx1_ASAP7_75t_L g6646 ( 
.A(n_5709),
.Y(n_6646)
);

AND2x4_ASAP7_75t_L g6647 ( 
.A(n_5706),
.B(n_6026),
.Y(n_6647)
);

INVx2_ASAP7_75t_L g6648 ( 
.A(n_5211),
.Y(n_6648)
);

INVx1_ASAP7_75t_L g6649 ( 
.A(n_5709),
.Y(n_6649)
);

OAI21x1_ASAP7_75t_L g6650 ( 
.A1(n_5350),
.A2(n_5397),
.B(n_5518),
.Y(n_6650)
);

AOI21xp5_ASAP7_75t_L g6651 ( 
.A1(n_5651),
.A2(n_5141),
.B(n_5136),
.Y(n_6651)
);

OAI221xp5_ASAP7_75t_L g6652 ( 
.A1(n_5416),
.A2(n_4946),
.B1(n_4919),
.B2(n_4859),
.C(n_4844),
.Y(n_6652)
);

INVx4_ASAP7_75t_L g6653 ( 
.A(n_5834),
.Y(n_6653)
);

INVx1_ASAP7_75t_L g6654 ( 
.A(n_5717),
.Y(n_6654)
);

OR2x2_ASAP7_75t_L g6655 ( 
.A(n_6013),
.B(n_4976),
.Y(n_6655)
);

OR2x2_ASAP7_75t_L g6656 ( 
.A(n_6013),
.B(n_4976),
.Y(n_6656)
);

OAI21xp5_ASAP7_75t_L g6657 ( 
.A1(n_5248),
.A2(n_4415),
.B(n_4410),
.Y(n_6657)
);

CKINVDCx11_ASAP7_75t_R g6658 ( 
.A(n_5251),
.Y(n_6658)
);

INVx3_ASAP7_75t_L g6659 ( 
.A(n_5556),
.Y(n_6659)
);

INVx3_ASAP7_75t_SL g6660 ( 
.A(n_5251),
.Y(n_6660)
);

BUFx6f_ASAP7_75t_L g6661 ( 
.A(n_5965),
.Y(n_6661)
);

AOI21x1_ASAP7_75t_L g6662 ( 
.A1(n_5389),
.A2(n_4671),
.B(n_4598),
.Y(n_6662)
);

INVxp67_ASAP7_75t_L g6663 ( 
.A(n_5526),
.Y(n_6663)
);

NAND3xp33_ASAP7_75t_L g6664 ( 
.A(n_5460),
.B(n_4413),
.C(n_4409),
.Y(n_6664)
);

INVx1_ASAP7_75t_SL g6665 ( 
.A(n_5464),
.Y(n_6665)
);

INVx1_ASAP7_75t_L g6666 ( 
.A(n_5717),
.Y(n_6666)
);

OR2x2_ASAP7_75t_L g6667 ( 
.A(n_6013),
.B(n_4976),
.Y(n_6667)
);

INVx1_ASAP7_75t_L g6668 ( 
.A(n_5730),
.Y(n_6668)
);

OR2x2_ASAP7_75t_L g6669 ( 
.A(n_6013),
.B(n_4976),
.Y(n_6669)
);

NAND2xp5_ASAP7_75t_L g6670 ( 
.A(n_5577),
.B(n_4437),
.Y(n_6670)
);

BUFx3_ASAP7_75t_L g6671 ( 
.A(n_5940),
.Y(n_6671)
);

CKINVDCx5p33_ASAP7_75t_R g6672 ( 
.A(n_5375),
.Y(n_6672)
);

INVx2_ASAP7_75t_L g6673 ( 
.A(n_5211),
.Y(n_6673)
);

AOI221xp5_ASAP7_75t_L g6674 ( 
.A1(n_5636),
.A2(n_4435),
.B1(n_4450),
.B2(n_4429),
.C(n_4409),
.Y(n_6674)
);

NOR2xp33_ASAP7_75t_L g6675 ( 
.A(n_5453),
.B(n_5089),
.Y(n_6675)
);

HB1xp67_ASAP7_75t_L g6676 ( 
.A(n_5727),
.Y(n_6676)
);

NAND2xp5_ASAP7_75t_L g6677 ( 
.A(n_5628),
.B(n_4580),
.Y(n_6677)
);

AOI21x1_ASAP7_75t_L g6678 ( 
.A1(n_5389),
.A2(n_4671),
.B(n_4598),
.Y(n_6678)
);

OA21x2_ASAP7_75t_L g6679 ( 
.A1(n_5917),
.A2(n_5056),
.B(n_5054),
.Y(n_6679)
);

NAND2xp5_ASAP7_75t_L g6680 ( 
.A(n_5628),
.B(n_4580),
.Y(n_6680)
);

INVx1_ASAP7_75t_L g6681 ( 
.A(n_5730),
.Y(n_6681)
);

AOI21xp33_ASAP7_75t_SL g6682 ( 
.A1(n_5319),
.A2(n_5104),
.B(n_5095),
.Y(n_6682)
);

AOI22xp33_ASAP7_75t_L g6683 ( 
.A1(n_5770),
.A2(n_5528),
.B1(n_5992),
.B2(n_5421),
.Y(n_6683)
);

INVx1_ASAP7_75t_L g6684 ( 
.A(n_5739),
.Y(n_6684)
);

AOI21x1_ASAP7_75t_L g6685 ( 
.A1(n_5849),
.A2(n_4671),
.B(n_4598),
.Y(n_6685)
);

OAI22xp5_ASAP7_75t_L g6686 ( 
.A1(n_5992),
.A2(n_4868),
.B1(n_4459),
.B2(n_4461),
.Y(n_6686)
);

OAI21x1_ASAP7_75t_L g6687 ( 
.A1(n_5819),
.A2(n_5067),
.B(n_4908),
.Y(n_6687)
);

INVx1_ASAP7_75t_L g6688 ( 
.A(n_5739),
.Y(n_6688)
);

INVx2_ASAP7_75t_SL g6689 ( 
.A(n_5556),
.Y(n_6689)
);

INVx1_ASAP7_75t_L g6690 ( 
.A(n_5746),
.Y(n_6690)
);

BUFx2_ASAP7_75t_L g6691 ( 
.A(n_5642),
.Y(n_6691)
);

INVx2_ASAP7_75t_L g6692 ( 
.A(n_5211),
.Y(n_6692)
);

OR2x2_ASAP7_75t_L g6693 ( 
.A(n_5333),
.B(n_4976),
.Y(n_6693)
);

OAI21x1_ASAP7_75t_L g6694 ( 
.A1(n_5779),
.A2(n_5815),
.B(n_5417),
.Y(n_6694)
);

OAI221xp5_ASAP7_75t_L g6695 ( 
.A1(n_5647),
.A2(n_4919),
.B1(n_4963),
.B2(n_4859),
.C(n_4844),
.Y(n_6695)
);

OA21x2_ASAP7_75t_L g6696 ( 
.A1(n_5917),
.A2(n_5056),
.B(n_5054),
.Y(n_6696)
);

CKINVDCx5p33_ASAP7_75t_R g6697 ( 
.A(n_5654),
.Y(n_6697)
);

OAI21xp5_ASAP7_75t_L g6698 ( 
.A1(n_5669),
.A2(n_4415),
.B(n_4410),
.Y(n_6698)
);

OAI21xp5_ASAP7_75t_L g6699 ( 
.A1(n_5669),
.A2(n_4456),
.B(n_4415),
.Y(n_6699)
);

CKINVDCx20_ASAP7_75t_R g6700 ( 
.A(n_5629),
.Y(n_6700)
);

BUFx3_ASAP7_75t_L g6701 ( 
.A(n_5811),
.Y(n_6701)
);

NAND2x1_ASAP7_75t_L g6702 ( 
.A(n_5645),
.B(n_4767),
.Y(n_6702)
);

INVx2_ASAP7_75t_L g6703 ( 
.A(n_5226),
.Y(n_6703)
);

AOI22xp33_ASAP7_75t_L g6704 ( 
.A1(n_5528),
.A2(n_4741),
.B1(n_4880),
.B2(n_4456),
.Y(n_6704)
);

OAI21x1_ASAP7_75t_L g6705 ( 
.A1(n_5778),
.A2(n_5067),
.B(n_4908),
.Y(n_6705)
);

INVxp67_ASAP7_75t_L g6706 ( 
.A(n_5555),
.Y(n_6706)
);

NAND2xp5_ASAP7_75t_L g6707 ( 
.A(n_5638),
.B(n_4580),
.Y(n_6707)
);

O2A1O1Ixp5_ASAP7_75t_L g6708 ( 
.A1(n_5203),
.A2(n_5090),
.B(n_4483),
.C(n_4509),
.Y(n_6708)
);

OAI21x1_ASAP7_75t_L g6709 ( 
.A1(n_5533),
.A2(n_5067),
.B(n_4908),
.Y(n_6709)
);

OA21x2_ASAP7_75t_L g6710 ( 
.A1(n_5631),
.A2(n_5056),
.B(n_5054),
.Y(n_6710)
);

OAI21x1_ASAP7_75t_L g6711 ( 
.A1(n_5533),
.A2(n_5067),
.B(n_4912),
.Y(n_6711)
);

NOR2xp33_ASAP7_75t_L g6712 ( 
.A(n_5453),
.B(n_5090),
.Y(n_6712)
);

AOI22xp33_ASAP7_75t_L g6713 ( 
.A1(n_5409),
.A2(n_4456),
.B1(n_4587),
.B2(n_4542),
.Y(n_6713)
);

INVx1_ASAP7_75t_L g6714 ( 
.A(n_5746),
.Y(n_6714)
);

AOI21xp5_ASAP7_75t_L g6715 ( 
.A1(n_5651),
.A2(n_5141),
.B(n_4767),
.Y(n_6715)
);

BUFx2_ASAP7_75t_L g6716 ( 
.A(n_5678),
.Y(n_6716)
);

INVx6_ASAP7_75t_SL g6717 ( 
.A(n_5811),
.Y(n_6717)
);

INVx1_ASAP7_75t_L g6718 ( 
.A(n_5747),
.Y(n_6718)
);

INVx1_ASAP7_75t_L g6719 ( 
.A(n_5747),
.Y(n_6719)
);

OAI21x1_ASAP7_75t_L g6720 ( 
.A1(n_5370),
.A2(n_5381),
.B(n_5376),
.Y(n_6720)
);

OAI22xp5_ASAP7_75t_L g6721 ( 
.A1(n_5785),
.A2(n_4459),
.B1(n_4461),
.B2(n_4450),
.Y(n_6721)
);

INVx1_ASAP7_75t_L g6722 ( 
.A(n_5788),
.Y(n_6722)
);

AND2x4_ASAP7_75t_L g6723 ( 
.A(n_5706),
.B(n_6026),
.Y(n_6723)
);

BUFx3_ASAP7_75t_L g6724 ( 
.A(n_5951),
.Y(n_6724)
);

AND2x2_ASAP7_75t_L g6725 ( 
.A(n_5539),
.B(n_4976),
.Y(n_6725)
);

OAI22xp5_ASAP7_75t_L g6726 ( 
.A1(n_5792),
.A2(n_4467),
.B1(n_4475),
.B2(n_4466),
.Y(n_6726)
);

AOI22xp33_ASAP7_75t_L g6727 ( 
.A1(n_5409),
.A2(n_4542),
.B1(n_4589),
.B2(n_4587),
.Y(n_6727)
);

BUFx6f_ASAP7_75t_L g6728 ( 
.A(n_5965),
.Y(n_6728)
);

INVx2_ASAP7_75t_SL g6729 ( 
.A(n_5556),
.Y(n_6729)
);

OAI21x1_ASAP7_75t_L g6730 ( 
.A1(n_5614),
.A2(n_4912),
.B(n_4896),
.Y(n_6730)
);

OR2x2_ASAP7_75t_L g6731 ( 
.A(n_5333),
.B(n_4894),
.Y(n_6731)
);

NOR2xp67_ASAP7_75t_L g6732 ( 
.A(n_5580),
.B(n_5411),
.Y(n_6732)
);

OAI21x1_ASAP7_75t_L g6733 ( 
.A1(n_5614),
.A2(n_4912),
.B(n_4896),
.Y(n_6733)
);

INVx6_ASAP7_75t_L g6734 ( 
.A(n_5951),
.Y(n_6734)
);

OAI21x1_ASAP7_75t_L g6735 ( 
.A1(n_5614),
.A2(n_4920),
.B(n_4896),
.Y(n_6735)
);

OAI21xp5_ASAP7_75t_L g6736 ( 
.A1(n_5151),
.A2(n_4587),
.B(n_4542),
.Y(n_6736)
);

BUFx2_ASAP7_75t_L g6737 ( 
.A(n_5580),
.Y(n_6737)
);

NAND2xp5_ASAP7_75t_L g6738 ( 
.A(n_5638),
.B(n_4580),
.Y(n_6738)
);

AND2x4_ASAP7_75t_L g6739 ( 
.A(n_5706),
.B(n_4619),
.Y(n_6739)
);

INVx2_ASAP7_75t_L g6740 ( 
.A(n_5226),
.Y(n_6740)
);

INVx2_ASAP7_75t_L g6741 ( 
.A(n_5226),
.Y(n_6741)
);

INVx3_ASAP7_75t_L g6742 ( 
.A(n_5556),
.Y(n_6742)
);

NOR2x1_ASAP7_75t_R g6743 ( 
.A(n_5286),
.B(n_5324),
.Y(n_6743)
);

NAND3xp33_ASAP7_75t_L g6744 ( 
.A(n_5460),
.B(n_4467),
.C(n_4466),
.Y(n_6744)
);

AND2x4_ASAP7_75t_L g6745 ( 
.A(n_5706),
.B(n_4619),
.Y(n_6745)
);

NAND2xp5_ASAP7_75t_L g6746 ( 
.A(n_5832),
.B(n_4580),
.Y(n_6746)
);

OAI21x1_ASAP7_75t_L g6747 ( 
.A1(n_5766),
.A2(n_4923),
.B(n_4920),
.Y(n_6747)
);

INVx1_ASAP7_75t_L g6748 ( 
.A(n_5788),
.Y(n_6748)
);

OAI21x1_ASAP7_75t_L g6749 ( 
.A1(n_5829),
.A2(n_5859),
.B(n_5842),
.Y(n_6749)
);

AOI22xp33_ASAP7_75t_SL g6750 ( 
.A1(n_5636),
.A2(n_5141),
.B1(n_5091),
.B2(n_4698),
.Y(n_6750)
);

CKINVDCx5p33_ASAP7_75t_R g6751 ( 
.A(n_5776),
.Y(n_6751)
);

AND2x4_ASAP7_75t_L g6752 ( 
.A(n_6026),
.B(n_4619),
.Y(n_6752)
);

CKINVDCx5p33_ASAP7_75t_R g6753 ( 
.A(n_5212),
.Y(n_6753)
);

NAND2xp5_ASAP7_75t_L g6754 ( 
.A(n_5677),
.B(n_4580),
.Y(n_6754)
);

O2A1O1Ixp33_ASAP7_75t_SL g6755 ( 
.A1(n_5757),
.A2(n_5085),
.B(n_4859),
.C(n_4919),
.Y(n_6755)
);

OAI22xp33_ASAP7_75t_L g6756 ( 
.A1(n_6017),
.A2(n_4484),
.B1(n_4492),
.B2(n_4475),
.Y(n_6756)
);

OAI22xp5_ASAP7_75t_L g6757 ( 
.A1(n_5326),
.A2(n_4492),
.B1(n_4503),
.B2(n_4484),
.Y(n_6757)
);

AOI22xp33_ASAP7_75t_L g6758 ( 
.A1(n_5421),
.A2(n_4589),
.B1(n_4600),
.B2(n_3598),
.Y(n_6758)
);

NAND2x1p5_ASAP7_75t_L g6759 ( 
.A(n_5411),
.B(n_4767),
.Y(n_6759)
);

AND2x2_ASAP7_75t_L g6760 ( 
.A(n_5564),
.B(n_4894),
.Y(n_6760)
);

HB1xp67_ASAP7_75t_L g6761 ( 
.A(n_5802),
.Y(n_6761)
);

INVx1_ASAP7_75t_L g6762 ( 
.A(n_5793),
.Y(n_6762)
);

INVx2_ASAP7_75t_L g6763 ( 
.A(n_5275),
.Y(n_6763)
);

INVx1_ASAP7_75t_L g6764 ( 
.A(n_5793),
.Y(n_6764)
);

INVx1_ASAP7_75t_L g6765 ( 
.A(n_5814),
.Y(n_6765)
);

INVx1_ASAP7_75t_L g6766 ( 
.A(n_5814),
.Y(n_6766)
);

CKINVDCx20_ASAP7_75t_R g6767 ( 
.A(n_5959),
.Y(n_6767)
);

HB1xp67_ASAP7_75t_L g6768 ( 
.A(n_5802),
.Y(n_6768)
);

BUFx2_ASAP7_75t_L g6769 ( 
.A(n_5612),
.Y(n_6769)
);

INVx2_ASAP7_75t_SL g6770 ( 
.A(n_5556),
.Y(n_6770)
);

NAND2xp5_ASAP7_75t_L g6771 ( 
.A(n_5686),
.B(n_4580),
.Y(n_6771)
);

NAND2x1p5_ASAP7_75t_L g6772 ( 
.A(n_5423),
.B(n_4767),
.Y(n_6772)
);

INVx2_ASAP7_75t_L g6773 ( 
.A(n_5275),
.Y(n_6773)
);

OA21x2_ASAP7_75t_L g6774 ( 
.A1(n_5631),
.A2(n_4931),
.B(n_4926),
.Y(n_6774)
);

OAI21x1_ASAP7_75t_SL g6775 ( 
.A1(n_5586),
.A2(n_4873),
.B(n_4872),
.Y(n_6775)
);

BUFx2_ASAP7_75t_L g6776 ( 
.A(n_5612),
.Y(n_6776)
);

AO21x1_ASAP7_75t_L g6777 ( 
.A1(n_5807),
.A2(n_5085),
.B(n_4872),
.Y(n_6777)
);

NOR2x1_ASAP7_75t_L g6778 ( 
.A(n_5468),
.B(n_5486),
.Y(n_6778)
);

BUFx2_ASAP7_75t_L g6779 ( 
.A(n_5385),
.Y(n_6779)
);

OA21x2_ASAP7_75t_L g6780 ( 
.A1(n_5647),
.A2(n_5100),
.B(n_5093),
.Y(n_6780)
);

AOI22xp5_ASAP7_75t_L g6781 ( 
.A1(n_6017),
.A2(n_3598),
.B1(n_4600),
.B2(n_4589),
.Y(n_6781)
);

AOI21xp5_ASAP7_75t_L g6782 ( 
.A1(n_5877),
.A2(n_5468),
.B(n_5486),
.Y(n_6782)
);

INVx2_ASAP7_75t_L g6783 ( 
.A(n_5275),
.Y(n_6783)
);

INVx2_ASAP7_75t_L g6784 ( 
.A(n_5339),
.Y(n_6784)
);

INVx6_ASAP7_75t_L g6785 ( 
.A(n_5951),
.Y(n_6785)
);

INVx2_ASAP7_75t_L g6786 ( 
.A(n_5339),
.Y(n_6786)
);

NAND2x1p5_ASAP7_75t_L g6787 ( 
.A(n_5423),
.B(n_4767),
.Y(n_6787)
);

AOI21x1_ASAP7_75t_L g6788 ( 
.A1(n_5849),
.A2(n_4671),
.B(n_4598),
.Y(n_6788)
);

INVx2_ASAP7_75t_L g6789 ( 
.A(n_5339),
.Y(n_6789)
);

OR2x6_ASAP7_75t_L g6790 ( 
.A(n_5645),
.B(n_5048),
.Y(n_6790)
);

AND2x2_ASAP7_75t_L g6791 ( 
.A(n_5564),
.B(n_4894),
.Y(n_6791)
);

NAND3xp33_ASAP7_75t_SL g6792 ( 
.A(n_5438),
.B(n_5107),
.C(n_4600),
.Y(n_6792)
);

AOI22xp5_ASAP7_75t_L g6793 ( 
.A1(n_5780),
.A2(n_5090),
.B1(n_4743),
.B2(n_4867),
.Y(n_6793)
);

INVx1_ASAP7_75t_L g6794 ( 
.A(n_5825),
.Y(n_6794)
);

INVx1_ASAP7_75t_L g6795 ( 
.A(n_5825),
.Y(n_6795)
);

BUFx3_ASAP7_75t_L g6796 ( 
.A(n_5951),
.Y(n_6796)
);

INVx2_ASAP7_75t_L g6797 ( 
.A(n_5340),
.Y(n_6797)
);

AO21x2_ASAP7_75t_L g6798 ( 
.A1(n_5721),
.A2(n_5053),
.B(n_5031),
.Y(n_6798)
);

OAI22xp33_ASAP7_75t_L g6799 ( 
.A1(n_5470),
.A2(n_4504),
.B1(n_4529),
.B2(n_4503),
.Y(n_6799)
);

AOI22xp33_ASAP7_75t_L g6800 ( 
.A1(n_5942),
.A2(n_4878),
.B1(n_4855),
.B2(n_4743),
.Y(n_6800)
);

CKINVDCx5p33_ASAP7_75t_R g6801 ( 
.A(n_5212),
.Y(n_6801)
);

AND2x4_ASAP7_75t_SL g6802 ( 
.A(n_5318),
.B(n_3844),
.Y(n_6802)
);

BUFx3_ASAP7_75t_L g6803 ( 
.A(n_5179),
.Y(n_6803)
);

INVx1_ASAP7_75t_L g6804 ( 
.A(n_5833),
.Y(n_6804)
);

AND2x4_ASAP7_75t_L g6805 ( 
.A(n_6026),
.B(n_4619),
.Y(n_6805)
);

AO31x2_ASAP7_75t_L g6806 ( 
.A1(n_6365),
.A2(n_5586),
.A3(n_5369),
.B(n_5437),
.Y(n_6806)
);

AOI21xp5_ASAP7_75t_L g6807 ( 
.A1(n_6625),
.A2(n_5877),
.B(n_5882),
.Y(n_6807)
);

OAI21xp5_ASAP7_75t_L g6808 ( 
.A1(n_6625),
.A2(n_5210),
.B(n_5332),
.Y(n_6808)
);

INVx1_ASAP7_75t_L g6809 ( 
.A(n_6037),
.Y(n_6809)
);

AOI21xp5_ASAP7_75t_L g6810 ( 
.A1(n_6133),
.A2(n_5889),
.B(n_5884),
.Y(n_6810)
);

AO21x2_ASAP7_75t_L g6811 ( 
.A1(n_6196),
.A2(n_5590),
.B(n_5566),
.Y(n_6811)
);

HB1xp67_ASAP7_75t_L g6812 ( 
.A(n_6524),
.Y(n_6812)
);

INVx1_ASAP7_75t_L g6813 ( 
.A(n_6037),
.Y(n_6813)
);

AND2x4_ASAP7_75t_L g6814 ( 
.A(n_6128),
.B(n_6026),
.Y(n_6814)
);

AO31x2_ASAP7_75t_L g6815 ( 
.A1(n_6365),
.A2(n_6292),
.A3(n_6587),
.B(n_6571),
.Y(n_6815)
);

AOI21xp5_ASAP7_75t_L g6816 ( 
.A1(n_6133),
.A2(n_5498),
.B(n_5794),
.Y(n_6816)
);

NOR2xp67_ASAP7_75t_SL g6817 ( 
.A(n_6089),
.B(n_5324),
.Y(n_6817)
);

AND2x4_ASAP7_75t_L g6818 ( 
.A(n_6128),
.B(n_5445),
.Y(n_6818)
);

HB1xp67_ASAP7_75t_L g6819 ( 
.A(n_6524),
.Y(n_6819)
);

OR2x2_ASAP7_75t_L g6820 ( 
.A(n_6070),
.B(n_5333),
.Y(n_6820)
);

INVx3_ASAP7_75t_L g6821 ( 
.A(n_6038),
.Y(n_6821)
);

AO31x2_ASAP7_75t_L g6822 ( 
.A1(n_6365),
.A2(n_5369),
.A3(n_5722),
.B(n_5705),
.Y(n_6822)
);

NAND2x1p5_ASAP7_75t_L g6823 ( 
.A(n_6778),
.B(n_5853),
.Y(n_6823)
);

AND2x4_ASAP7_75t_L g6824 ( 
.A(n_6128),
.B(n_5445),
.Y(n_6824)
);

OAI21x1_ASAP7_75t_L g6825 ( 
.A1(n_6685),
.A2(n_5938),
.B(n_5675),
.Y(n_6825)
);

AO31x2_ASAP7_75t_L g6826 ( 
.A1(n_6292),
.A2(n_5722),
.A3(n_5392),
.B(n_5405),
.Y(n_6826)
);

INVx1_ASAP7_75t_L g6827 ( 
.A(n_6037),
.Y(n_6827)
);

AND2x2_ASAP7_75t_L g6828 ( 
.A(n_6621),
.B(n_6018),
.Y(n_6828)
);

OA21x2_ASAP7_75t_L g6829 ( 
.A1(n_6715),
.A2(n_5590),
.B(n_5566),
.Y(n_6829)
);

OAI21x1_ASAP7_75t_L g6830 ( 
.A1(n_6685),
.A2(n_5938),
.B(n_5675),
.Y(n_6830)
);

INVx1_ASAP7_75t_L g6831 ( 
.A(n_6059),
.Y(n_6831)
);

AOI21xp5_ASAP7_75t_L g6832 ( 
.A1(n_6120),
.A2(n_5652),
.B(n_5737),
.Y(n_6832)
);

INVx1_ASAP7_75t_L g6833 ( 
.A(n_6059),
.Y(n_6833)
);

INVx4_ASAP7_75t_L g6834 ( 
.A(n_6089),
.Y(n_6834)
);

INVx2_ASAP7_75t_L g6835 ( 
.A(n_6284),
.Y(n_6835)
);

INVx2_ASAP7_75t_L g6836 ( 
.A(n_6284),
.Y(n_6836)
);

INVx1_ASAP7_75t_L g6837 ( 
.A(n_6059),
.Y(n_6837)
);

NAND2xp5_ASAP7_75t_L g6838 ( 
.A(n_6215),
.B(n_5844),
.Y(n_6838)
);

INVx1_ASAP7_75t_L g6839 ( 
.A(n_6067),
.Y(n_6839)
);

INVx6_ASAP7_75t_L g6840 ( 
.A(n_6039),
.Y(n_6840)
);

NAND2xp5_ASAP7_75t_L g6841 ( 
.A(n_6215),
.B(n_5847),
.Y(n_6841)
);

AND2x2_ASAP7_75t_L g6842 ( 
.A(n_6621),
.B(n_6018),
.Y(n_6842)
);

INVx3_ASAP7_75t_L g6843 ( 
.A(n_6038),
.Y(n_6843)
);

AOI21xp5_ASAP7_75t_L g6844 ( 
.A1(n_6120),
.A2(n_5690),
.B(n_5926),
.Y(n_6844)
);

AND2x2_ASAP7_75t_L g6845 ( 
.A(n_6621),
.B(n_6014),
.Y(n_6845)
);

INVx2_ASAP7_75t_L g6846 ( 
.A(n_6284),
.Y(n_6846)
);

NOR2xp33_ASAP7_75t_L g6847 ( 
.A(n_6189),
.B(n_5324),
.Y(n_6847)
);

INVx2_ASAP7_75t_SL g6848 ( 
.A(n_6452),
.Y(n_6848)
);

OAI21x1_ASAP7_75t_L g6849 ( 
.A1(n_6685),
.A2(n_6788),
.B(n_6702),
.Y(n_6849)
);

NAND2xp5_ASAP7_75t_L g6850 ( 
.A(n_6160),
.B(n_5465),
.Y(n_6850)
);

AOI21xp5_ASAP7_75t_L g6851 ( 
.A1(n_6238),
.A2(n_5960),
.B(n_5315),
.Y(n_6851)
);

NAND2xp5_ASAP7_75t_L g6852 ( 
.A(n_6160),
.B(n_5465),
.Y(n_6852)
);

AND2x2_ASAP7_75t_L g6853 ( 
.A(n_6355),
.B(n_6014),
.Y(n_6853)
);

INVx1_ASAP7_75t_L g6854 ( 
.A(n_6067),
.Y(n_6854)
);

AOI21xp5_ASAP7_75t_L g6855 ( 
.A1(n_6238),
.A2(n_5989),
.B(n_5731),
.Y(n_6855)
);

INVx1_ASAP7_75t_L g6856 ( 
.A(n_6067),
.Y(n_6856)
);

OAI21x1_ASAP7_75t_L g6857 ( 
.A1(n_6788),
.A2(n_5688),
.B(n_5676),
.Y(n_6857)
);

BUFx2_ASAP7_75t_L g6858 ( 
.A(n_6743),
.Y(n_6858)
);

OR2x2_ASAP7_75t_L g6859 ( 
.A(n_6070),
.B(n_5333),
.Y(n_6859)
);

AOI21xp33_ASAP7_75t_L g6860 ( 
.A1(n_6123),
.A2(n_5708),
.B(n_5665),
.Y(n_6860)
);

OAI21x1_ASAP7_75t_L g6861 ( 
.A1(n_6788),
.A2(n_5688),
.B(n_5676),
.Y(n_6861)
);

AOI21xp33_ASAP7_75t_SL g6862 ( 
.A1(n_6533),
.A2(n_5412),
.B(n_5239),
.Y(n_6862)
);

INVx1_ASAP7_75t_L g6863 ( 
.A(n_6075),
.Y(n_6863)
);

OA21x2_ASAP7_75t_L g6864 ( 
.A1(n_6715),
.A2(n_5361),
.B(n_5506),
.Y(n_6864)
);

AOI21xp33_ASAP7_75t_SL g6865 ( 
.A1(n_6533),
.A2(n_5454),
.B(n_5261),
.Y(n_6865)
);

AO21x2_ASAP7_75t_L g6866 ( 
.A1(n_6196),
.A2(n_6502),
.B(n_6074),
.Y(n_6866)
);

INVx1_ASAP7_75t_L g6867 ( 
.A(n_6075),
.Y(n_6867)
);

INVx2_ASAP7_75t_L g6868 ( 
.A(n_6284),
.Y(n_6868)
);

CKINVDCx11_ASAP7_75t_R g6869 ( 
.A(n_6131),
.Y(n_6869)
);

OA21x2_ASAP7_75t_L g6870 ( 
.A1(n_6066),
.A2(n_5506),
.B(n_5554),
.Y(n_6870)
);

OR2x2_ASAP7_75t_L g6871 ( 
.A(n_6246),
.B(n_5333),
.Y(n_6871)
);

NAND2xp5_ASAP7_75t_L g6872 ( 
.A(n_6213),
.B(n_5433),
.Y(n_6872)
);

BUFx2_ASAP7_75t_L g6873 ( 
.A(n_6743),
.Y(n_6873)
);

AO31x2_ASAP7_75t_L g6874 ( 
.A1(n_6292),
.A2(n_5725),
.A3(n_5696),
.B(n_5525),
.Y(n_6874)
);

OAI21x1_ASAP7_75t_L g6875 ( 
.A1(n_6702),
.A2(n_5659),
.B(n_5929),
.Y(n_6875)
);

INVx2_ASAP7_75t_L g6876 ( 
.A(n_6294),
.Y(n_6876)
);

AO22x2_ASAP7_75t_L g6877 ( 
.A1(n_6066),
.A2(n_5997),
.B1(n_5610),
.B2(n_5544),
.Y(n_6877)
);

OAI21x1_ASAP7_75t_SL g6878 ( 
.A1(n_6782),
.A2(n_5222),
.B(n_5209),
.Y(n_6878)
);

OAI21x1_ASAP7_75t_L g6879 ( 
.A1(n_6702),
.A2(n_5659),
.B(n_5929),
.Y(n_6879)
);

INVx1_ASAP7_75t_L g6880 ( 
.A(n_6075),
.Y(n_6880)
);

AND2x4_ASAP7_75t_L g6881 ( 
.A(n_6128),
.B(n_6198),
.Y(n_6881)
);

INVx2_ASAP7_75t_SL g6882 ( 
.A(n_6452),
.Y(n_6882)
);

HB1xp67_ASAP7_75t_L g6883 ( 
.A(n_6626),
.Y(n_6883)
);

OAI21x1_ASAP7_75t_L g6884 ( 
.A1(n_6782),
.A2(n_5930),
.B(n_5933),
.Y(n_6884)
);

OAI21xp5_ASAP7_75t_L g6885 ( 
.A1(n_6123),
.A2(n_6371),
.B(n_6436),
.Y(n_6885)
);

BUFx12f_ASAP7_75t_L g6886 ( 
.A(n_6126),
.Y(n_6886)
);

INVx2_ASAP7_75t_L g6887 ( 
.A(n_6294),
.Y(n_6887)
);

NOR2xp33_ASAP7_75t_L g6888 ( 
.A(n_6189),
.B(n_5335),
.Y(n_6888)
);

INVx2_ASAP7_75t_L g6889 ( 
.A(n_6294),
.Y(n_6889)
);

BUFx6f_ASAP7_75t_L g6890 ( 
.A(n_6126),
.Y(n_6890)
);

AND2x4_ASAP7_75t_SL g6891 ( 
.A(n_6189),
.B(n_5209),
.Y(n_6891)
);

NAND2xp5_ASAP7_75t_L g6892 ( 
.A(n_6213),
.B(n_5433),
.Y(n_6892)
);

INVx1_ASAP7_75t_L g6893 ( 
.A(n_6099),
.Y(n_6893)
);

NOR2xp33_ASAP7_75t_L g6894 ( 
.A(n_6062),
.B(n_5335),
.Y(n_6894)
);

NAND2xp5_ASAP7_75t_L g6895 ( 
.A(n_6082),
.B(n_5406),
.Y(n_6895)
);

AOI21xp5_ASAP7_75t_L g6896 ( 
.A1(n_6055),
.A2(n_5751),
.B(n_5816),
.Y(n_6896)
);

INVx1_ASAP7_75t_L g6897 ( 
.A(n_6099),
.Y(n_6897)
);

NAND2xp5_ASAP7_75t_L g6898 ( 
.A(n_6082),
.B(n_5406),
.Y(n_6898)
);

INVx2_ASAP7_75t_SL g6899 ( 
.A(n_6647),
.Y(n_6899)
);

AO31x2_ASAP7_75t_L g6900 ( 
.A1(n_6571),
.A2(n_5514),
.A3(n_5444),
.B(n_5997),
.Y(n_6900)
);

NAND2x1p5_ASAP7_75t_L g6901 ( 
.A(n_6778),
.B(n_5853),
.Y(n_6901)
);

OAI21x1_ASAP7_75t_L g6902 ( 
.A1(n_6057),
.A2(n_5930),
.B(n_5933),
.Y(n_6902)
);

NAND2xp5_ASAP7_75t_L g6903 ( 
.A(n_6088),
.B(n_5918),
.Y(n_6903)
);

AOI21xp5_ASAP7_75t_L g6904 ( 
.A1(n_6055),
.A2(n_5270),
.B(n_5331),
.Y(n_6904)
);

INVx1_ASAP7_75t_L g6905 ( 
.A(n_6099),
.Y(n_6905)
);

AO21x2_ASAP7_75t_L g6906 ( 
.A1(n_6074),
.A2(n_5721),
.B(n_5874),
.Y(n_6906)
);

AOI21xp5_ASAP7_75t_L g6907 ( 
.A1(n_6085),
.A2(n_5328),
.B(n_5609),
.Y(n_6907)
);

AND2x2_ASAP7_75t_L g6908 ( 
.A(n_6355),
.B(n_5445),
.Y(n_6908)
);

OAI21x1_ASAP7_75t_L g6909 ( 
.A1(n_6057),
.A2(n_5933),
.B(n_5860),
.Y(n_6909)
);

OAI21x1_ASAP7_75t_L g6910 ( 
.A1(n_6057),
.A2(n_5933),
.B(n_5870),
.Y(n_6910)
);

AOI21xp5_ASAP7_75t_L g6911 ( 
.A1(n_6085),
.A2(n_5820),
.B(n_5858),
.Y(n_6911)
);

NAND2xp5_ASAP7_75t_L g6912 ( 
.A(n_6088),
.B(n_5918),
.Y(n_6912)
);

INVx2_ASAP7_75t_L g6913 ( 
.A(n_6294),
.Y(n_6913)
);

INVx1_ASAP7_75t_L g6914 ( 
.A(n_6102),
.Y(n_6914)
);

OAI21x1_ASAP7_75t_L g6915 ( 
.A1(n_6662),
.A2(n_5848),
.B(n_5549),
.Y(n_6915)
);

INVx3_ASAP7_75t_L g6916 ( 
.A(n_6038),
.Y(n_6916)
);

NAND2x1p5_ASAP7_75t_L g6917 ( 
.A(n_6509),
.B(n_5503),
.Y(n_6917)
);

HB1xp67_ASAP7_75t_L g6918 ( 
.A(n_6626),
.Y(n_6918)
);

AND2x2_ASAP7_75t_L g6919 ( 
.A(n_6355),
.B(n_5445),
.Y(n_6919)
);

HB1xp67_ASAP7_75t_L g6920 ( 
.A(n_6631),
.Y(n_6920)
);

INVx2_ASAP7_75t_L g6921 ( 
.A(n_6386),
.Y(n_6921)
);

OAI21xp5_ASAP7_75t_L g6922 ( 
.A1(n_6371),
.A2(n_5195),
.B(n_5729),
.Y(n_6922)
);

OAI21xp5_ASAP7_75t_L g6923 ( 
.A1(n_6436),
.A2(n_5774),
.B(n_5670),
.Y(n_6923)
);

BUFx2_ASAP7_75t_L g6924 ( 
.A(n_6647),
.Y(n_6924)
);

HB1xp67_ASAP7_75t_L g6925 ( 
.A(n_6631),
.Y(n_6925)
);

AND2x4_ASAP7_75t_L g6926 ( 
.A(n_6128),
.B(n_5426),
.Y(n_6926)
);

OAI21x1_ASAP7_75t_L g6927 ( 
.A1(n_6662),
.A2(n_5549),
.B(n_5658),
.Y(n_6927)
);

INVx1_ASAP7_75t_L g6928 ( 
.A(n_6102),
.Y(n_6928)
);

AOI21xp5_ASAP7_75t_L g6929 ( 
.A1(n_6035),
.A2(n_5171),
.B(n_5972),
.Y(n_6929)
);

AOI21xp5_ASAP7_75t_L g6930 ( 
.A1(n_6035),
.A2(n_5171),
.B(n_6011),
.Y(n_6930)
);

NAND2x1p5_ASAP7_75t_L g6931 ( 
.A(n_6509),
.B(n_5503),
.Y(n_6931)
);

INVx2_ASAP7_75t_SL g6932 ( 
.A(n_6647),
.Y(n_6932)
);

AOI21x1_ASAP7_75t_L g6933 ( 
.A1(n_6260),
.A2(n_5896),
.B(n_5874),
.Y(n_6933)
);

BUFx2_ASAP7_75t_L g6934 ( 
.A(n_6647),
.Y(n_6934)
);

OA21x2_ASAP7_75t_L g6935 ( 
.A1(n_6502),
.A2(n_5561),
.B(n_5554),
.Y(n_6935)
);

OA21x2_ASAP7_75t_L g6936 ( 
.A1(n_6651),
.A2(n_5563),
.B(n_5561),
.Y(n_6936)
);

AOI22xp33_ASAP7_75t_L g6937 ( 
.A1(n_6683),
.A2(n_5443),
.B1(n_5666),
.B2(n_5569),
.Y(n_6937)
);

INVx1_ASAP7_75t_L g6938 ( 
.A(n_6102),
.Y(n_6938)
);

INVxp33_ASAP7_75t_L g6939 ( 
.A(n_6109),
.Y(n_6939)
);

OAI21xp5_ASAP7_75t_L g6940 ( 
.A1(n_6343),
.A2(n_5670),
.B(n_5434),
.Y(n_6940)
);

INVx1_ASAP7_75t_L g6941 ( 
.A(n_6116),
.Y(n_6941)
);

NAND2xp5_ASAP7_75t_L g6942 ( 
.A(n_6195),
.B(n_5866),
.Y(n_6942)
);

AOI22xp5_ASAP7_75t_L g6943 ( 
.A1(n_6683),
.A2(n_5780),
.B1(n_5470),
.B2(n_5754),
.Y(n_6943)
);

AOI21xp5_ASAP7_75t_L g6944 ( 
.A1(n_6526),
.A2(n_5910),
.B(n_5572),
.Y(n_6944)
);

INVx6_ASAP7_75t_L g6945 ( 
.A(n_6039),
.Y(n_6945)
);

AOI21x1_ASAP7_75t_L g6946 ( 
.A1(n_6260),
.A2(n_5896),
.B(n_5386),
.Y(n_6946)
);

OA21x2_ASAP7_75t_L g6947 ( 
.A1(n_6651),
.A2(n_5563),
.B(n_5426),
.Y(n_6947)
);

AND2x4_ASAP7_75t_L g6948 ( 
.A(n_6128),
.B(n_5684),
.Y(n_6948)
);

BUFx6f_ASAP7_75t_SL g6949 ( 
.A(n_6269),
.Y(n_6949)
);

OAI21x1_ASAP7_75t_L g6950 ( 
.A1(n_6662),
.A2(n_5549),
.B(n_5658),
.Y(n_6950)
);

NAND2xp5_ASAP7_75t_L g6951 ( 
.A(n_6195),
.B(n_5866),
.Y(n_6951)
);

HB1xp67_ASAP7_75t_L g6952 ( 
.A(n_6641),
.Y(n_6952)
);

A2O1A1Ixp33_ASAP7_75t_L g6953 ( 
.A1(n_6642),
.A2(n_5830),
.B(n_5438),
.C(n_5482),
.Y(n_6953)
);

BUFx12f_ASAP7_75t_L g6954 ( 
.A(n_6457),
.Y(n_6954)
);

OAI21x1_ASAP7_75t_L g6955 ( 
.A1(n_6678),
.A2(n_5549),
.B(n_5943),
.Y(n_6955)
);

CKINVDCx11_ASAP7_75t_R g6956 ( 
.A(n_6131),
.Y(n_6956)
);

OAI21x1_ASAP7_75t_L g6957 ( 
.A1(n_6678),
.A2(n_5943),
.B(n_5952),
.Y(n_6957)
);

NAND2x1p5_ASAP7_75t_L g6958 ( 
.A(n_6509),
.B(n_5400),
.Y(n_6958)
);

AO21x2_ASAP7_75t_L g6959 ( 
.A1(n_6526),
.A2(n_5721),
.B(n_5544),
.Y(n_6959)
);

BUFx3_ASAP7_75t_L g6960 ( 
.A(n_6089),
.Y(n_6960)
);

OR2x2_ASAP7_75t_L g6961 ( 
.A(n_6246),
.B(n_5333),
.Y(n_6961)
);

OAI21x1_ASAP7_75t_L g6962 ( 
.A1(n_6678),
.A2(n_5943),
.B(n_5952),
.Y(n_6962)
);

INVx1_ASAP7_75t_L g6963 ( 
.A(n_6116),
.Y(n_6963)
);

INVx2_ASAP7_75t_L g6964 ( 
.A(n_6305),
.Y(n_6964)
);

AOI21xp5_ASAP7_75t_L g6965 ( 
.A1(n_6200),
.A2(n_5574),
.B(n_5557),
.Y(n_6965)
);

NAND2xp5_ASAP7_75t_L g6966 ( 
.A(n_6470),
.B(n_5474),
.Y(n_6966)
);

INVx2_ASAP7_75t_SL g6967 ( 
.A(n_6647),
.Y(n_6967)
);

AOI21xp33_ASAP7_75t_L g6968 ( 
.A1(n_6200),
.A2(n_5274),
.B(n_5273),
.Y(n_6968)
);

OA21x2_ASAP7_75t_L g6969 ( 
.A1(n_6565),
.A2(n_5632),
.B(n_5644),
.Y(n_6969)
);

INVx2_ASAP7_75t_L g6970 ( 
.A(n_6305),
.Y(n_6970)
);

INVx2_ASAP7_75t_L g6971 ( 
.A(n_6305),
.Y(n_6971)
);

AOI21xp5_ASAP7_75t_L g6972 ( 
.A1(n_6150),
.A2(n_5622),
.B(n_5762),
.Y(n_6972)
);

OR2x6_ASAP7_75t_L g6973 ( 
.A(n_6150),
.B(n_5179),
.Y(n_6973)
);

AND2x4_ASAP7_75t_L g6974 ( 
.A(n_6128),
.B(n_5684),
.Y(n_6974)
);

NOR2xp33_ASAP7_75t_L g6975 ( 
.A(n_6062),
.B(n_5335),
.Y(n_6975)
);

AND2x4_ASAP7_75t_L g6976 ( 
.A(n_6198),
.B(n_5684),
.Y(n_6976)
);

BUFx12f_ASAP7_75t_L g6977 ( 
.A(n_6457),
.Y(n_6977)
);

HB1xp67_ASAP7_75t_L g6978 ( 
.A(n_6641),
.Y(n_6978)
);

INVx3_ASAP7_75t_L g6979 ( 
.A(n_6038),
.Y(n_6979)
);

HB1xp67_ASAP7_75t_L g6980 ( 
.A(n_6676),
.Y(n_6980)
);

OR2x2_ASAP7_75t_L g6981 ( 
.A(n_6246),
.B(n_5343),
.Y(n_6981)
);

INVx1_ASAP7_75t_L g6982 ( 
.A(n_6116),
.Y(n_6982)
);

AOI21xp5_ASAP7_75t_L g6983 ( 
.A1(n_6158),
.A2(n_5800),
.B(n_5147),
.Y(n_6983)
);

CKINVDCx16_ASAP7_75t_R g6984 ( 
.A(n_6109),
.Y(n_6984)
);

BUFx3_ASAP7_75t_L g6985 ( 
.A(n_6089),
.Y(n_6985)
);

INVx1_ASAP7_75t_L g6986 ( 
.A(n_6125),
.Y(n_6986)
);

INVx2_ASAP7_75t_L g6987 ( 
.A(n_6305),
.Y(n_6987)
);

INVx1_ASAP7_75t_L g6988 ( 
.A(n_6125),
.Y(n_6988)
);

OAI21x1_ASAP7_75t_L g6989 ( 
.A1(n_6418),
.A2(n_5943),
.B(n_5952),
.Y(n_6989)
);

INVx2_ASAP7_75t_L g6990 ( 
.A(n_6310),
.Y(n_6990)
);

AOI21xp5_ASAP7_75t_L g6991 ( 
.A1(n_6158),
.A2(n_5813),
.B(n_5434),
.Y(n_6991)
);

INVx2_ASAP7_75t_L g6992 ( 
.A(n_6310),
.Y(n_6992)
);

INVx1_ASAP7_75t_L g6993 ( 
.A(n_6125),
.Y(n_6993)
);

INVx1_ASAP7_75t_L g6994 ( 
.A(n_6127),
.Y(n_6994)
);

OA21x2_ASAP7_75t_L g6995 ( 
.A1(n_6565),
.A2(n_5632),
.B(n_5644),
.Y(n_6995)
);

A2O1A1Ixp33_ASAP7_75t_L g6996 ( 
.A1(n_6642),
.A2(n_5578),
.B(n_5562),
.C(n_5480),
.Y(n_6996)
);

INVx2_ASAP7_75t_L g6997 ( 
.A(n_6310),
.Y(n_6997)
);

OR2x2_ASAP7_75t_L g6998 ( 
.A(n_6299),
.B(n_5343),
.Y(n_6998)
);

CKINVDCx16_ASAP7_75t_R g6999 ( 
.A(n_6469),
.Y(n_6999)
);

OA21x2_ASAP7_75t_L g7000 ( 
.A1(n_6056),
.A2(n_5487),
.B(n_5713),
.Y(n_7000)
);

AOI21x1_ASAP7_75t_L g7001 ( 
.A1(n_6260),
.A2(n_5386),
.B(n_5464),
.Y(n_7001)
);

INVxp67_ASAP7_75t_SL g7002 ( 
.A(n_6777),
.Y(n_7002)
);

A2O1A1Ixp33_ASAP7_75t_L g7003 ( 
.A1(n_6485),
.A2(n_5419),
.B(n_5450),
.C(n_5942),
.Y(n_7003)
);

AO31x2_ASAP7_75t_L g7004 ( 
.A1(n_6571),
.A2(n_5863),
.A3(n_5865),
.B(n_5655),
.Y(n_7004)
);

INVx1_ASAP7_75t_L g7005 ( 
.A(n_6127),
.Y(n_7005)
);

AND2x2_ASAP7_75t_L g7006 ( 
.A(n_6410),
.B(n_6769),
.Y(n_7006)
);

NOR2x1_ASAP7_75t_SL g7007 ( 
.A(n_6792),
.B(n_5385),
.Y(n_7007)
);

A2O1A1Ixp33_ASAP7_75t_L g7008 ( 
.A1(n_6485),
.A2(n_6374),
.B(n_6505),
.C(n_6343),
.Y(n_7008)
);

NOR2xp33_ASAP7_75t_L g7009 ( 
.A(n_6062),
.B(n_5427),
.Y(n_7009)
);

OAI21x1_ASAP7_75t_L g7010 ( 
.A1(n_6418),
.A2(n_5980),
.B(n_5719),
.Y(n_7010)
);

BUFx12f_ASAP7_75t_L g7011 ( 
.A(n_6637),
.Y(n_7011)
);

NAND2xp5_ASAP7_75t_L g7012 ( 
.A(n_6470),
.B(n_5474),
.Y(n_7012)
);

BUFx2_ASAP7_75t_L g7013 ( 
.A(n_6647),
.Y(n_7013)
);

AOI21x1_ASAP7_75t_L g7014 ( 
.A1(n_6444),
.A2(n_5583),
.B(n_5475),
.Y(n_7014)
);

INVx2_ASAP7_75t_SL g7015 ( 
.A(n_6723),
.Y(n_7015)
);

NAND2xp5_ASAP7_75t_L g7016 ( 
.A(n_6484),
.B(n_5894),
.Y(n_7016)
);

AND2x2_ASAP7_75t_L g7017 ( 
.A(n_6410),
.B(n_6769),
.Y(n_7017)
);

OAI21x1_ASAP7_75t_L g7018 ( 
.A1(n_6418),
.A2(n_5980),
.B(n_5719),
.Y(n_7018)
);

OAI21x1_ASAP7_75t_L g7019 ( 
.A1(n_6459),
.A2(n_5980),
.B(n_5969),
.Y(n_7019)
);

OAI21x1_ASAP7_75t_L g7020 ( 
.A1(n_6459),
.A2(n_5969),
.B(n_5964),
.Y(n_7020)
);

AOI21xp5_ASAP7_75t_L g7021 ( 
.A1(n_6509),
.A2(n_5419),
.B(n_5999),
.Y(n_7021)
);

OR2x2_ASAP7_75t_L g7022 ( 
.A(n_6299),
.B(n_6369),
.Y(n_7022)
);

INVx2_ASAP7_75t_L g7023 ( 
.A(n_6310),
.Y(n_7023)
);

OAI21xp5_ASAP7_75t_SL g7024 ( 
.A1(n_6588),
.A2(n_5329),
.B(n_5750),
.Y(n_7024)
);

AND2x2_ASAP7_75t_L g7025 ( 
.A(n_6410),
.B(n_5892),
.Y(n_7025)
);

OAI21x1_ASAP7_75t_L g7026 ( 
.A1(n_6459),
.A2(n_5973),
.B(n_5964),
.Y(n_7026)
);

NAND2xp5_ASAP7_75t_L g7027 ( 
.A(n_6484),
.B(n_5894),
.Y(n_7027)
);

NAND2xp5_ASAP7_75t_L g7028 ( 
.A(n_6492),
.B(n_5529),
.Y(n_7028)
);

AND2x2_ASAP7_75t_L g7029 ( 
.A(n_6769),
.B(n_5901),
.Y(n_7029)
);

AOI21x1_ASAP7_75t_L g7030 ( 
.A1(n_6444),
.A2(n_5583),
.B(n_5475),
.Y(n_7030)
);

OAI21x1_ASAP7_75t_L g7031 ( 
.A1(n_6056),
.A2(n_5973),
.B(n_5298),
.Y(n_7031)
);

AOI22xp33_ASAP7_75t_L g7032 ( 
.A1(n_6588),
.A2(n_6428),
.B1(n_6151),
.B2(n_6300),
.Y(n_7032)
);

AOI22xp5_ASAP7_75t_L g7033 ( 
.A1(n_6428),
.A2(n_5750),
.B1(n_5754),
.B2(n_6024),
.Y(n_7033)
);

AO31x2_ASAP7_75t_L g7034 ( 
.A1(n_6587),
.A2(n_6303),
.A3(n_6777),
.B(n_6434),
.Y(n_7034)
);

AND2x2_ASAP7_75t_L g7035 ( 
.A(n_6776),
.B(n_5913),
.Y(n_7035)
);

AO31x2_ASAP7_75t_L g7036 ( 
.A1(n_6587),
.A2(n_5863),
.A3(n_5865),
.B(n_5655),
.Y(n_7036)
);

BUFx6f_ASAP7_75t_L g7037 ( 
.A(n_6554),
.Y(n_7037)
);

NAND2xp5_ASAP7_75t_L g7038 ( 
.A(n_6492),
.B(n_5529),
.Y(n_7038)
);

AOI21x1_ASAP7_75t_L g7039 ( 
.A1(n_6052),
.A2(n_5649),
.B(n_5608),
.Y(n_7039)
);

AOI21xp5_ASAP7_75t_L g7040 ( 
.A1(n_6509),
.A2(n_6094),
.B(n_6374),
.Y(n_7040)
);

INVx1_ASAP7_75t_L g7041 ( 
.A(n_6127),
.Y(n_7041)
);

OAI21x1_ASAP7_75t_L g7042 ( 
.A1(n_6056),
.A2(n_5298),
.B(n_5663),
.Y(n_7042)
);

OA21x2_ASAP7_75t_L g7043 ( 
.A1(n_6063),
.A2(n_5714),
.B(n_5713),
.Y(n_7043)
);

OAI21x1_ASAP7_75t_L g7044 ( 
.A1(n_6068),
.A2(n_5298),
.B(n_5663),
.Y(n_7044)
);

AOI21xp5_ASAP7_75t_L g7045 ( 
.A1(n_6094),
.A2(n_6000),
.B(n_5999),
.Y(n_7045)
);

INVx4_ASAP7_75t_SL g7046 ( 
.A(n_6660),
.Y(n_7046)
);

NAND2x1p5_ASAP7_75t_L g7047 ( 
.A(n_6573),
.B(n_5400),
.Y(n_7047)
);

AOI21xp5_ASAP7_75t_L g7048 ( 
.A1(n_6218),
.A2(n_6000),
.B(n_5591),
.Y(n_7048)
);

OAI21xp5_ASAP7_75t_L g7049 ( 
.A1(n_6095),
.A2(n_5641),
.B(n_5510),
.Y(n_7049)
);

OR2x6_ASAP7_75t_L g7050 ( 
.A(n_6239),
.B(n_5179),
.Y(n_7050)
);

OAI221xp5_ASAP7_75t_L g7051 ( 
.A1(n_6095),
.A2(n_6117),
.B1(n_6146),
.B2(n_6249),
.C(n_6239),
.Y(n_7051)
);

OAI21xp5_ASAP7_75t_L g7052 ( 
.A1(n_6117),
.A2(n_5510),
.B(n_5495),
.Y(n_7052)
);

AOI21x1_ASAP7_75t_L g7053 ( 
.A1(n_6052),
.A2(n_5649),
.B(n_5608),
.Y(n_7053)
);

BUFx12f_ASAP7_75t_L g7054 ( 
.A(n_6637),
.Y(n_7054)
);

AND2x4_ASAP7_75t_L g7055 ( 
.A(n_6198),
.B(n_5684),
.Y(n_7055)
);

OAI21x1_ASAP7_75t_L g7056 ( 
.A1(n_6068),
.A2(n_5298),
.B(n_5242),
.Y(n_7056)
);

INVx2_ASAP7_75t_L g7057 ( 
.A(n_6640),
.Y(n_7057)
);

AOI21x1_ASAP7_75t_L g7058 ( 
.A1(n_6115),
.A2(n_6301),
.B(n_6270),
.Y(n_7058)
);

HB1xp67_ASAP7_75t_L g7059 ( 
.A(n_6676),
.Y(n_7059)
);

NAND2xp5_ASAP7_75t_L g7060 ( 
.A(n_6569),
.B(n_5546),
.Y(n_7060)
);

AO21x1_ASAP7_75t_L g7061 ( 
.A1(n_6114),
.A2(n_5522),
.B(n_5507),
.Y(n_7061)
);

AO21x2_ASAP7_75t_L g7062 ( 
.A1(n_6212),
.A2(n_5496),
.B(n_5637),
.Y(n_7062)
);

OA21x2_ASAP7_75t_L g7063 ( 
.A1(n_6063),
.A2(n_5714),
.B(n_5716),
.Y(n_7063)
);

OA21x2_ASAP7_75t_L g7064 ( 
.A1(n_6063),
.A2(n_5716),
.B(n_5661),
.Y(n_7064)
);

INVx1_ASAP7_75t_L g7065 ( 
.A(n_6132),
.Y(n_7065)
);

INVx4_ASAP7_75t_SL g7066 ( 
.A(n_6660),
.Y(n_7066)
);

OA21x2_ASAP7_75t_L g7067 ( 
.A1(n_6064),
.A2(n_6060),
.B(n_6493),
.Y(n_7067)
);

AOI21xp5_ASAP7_75t_L g7068 ( 
.A1(n_6218),
.A2(n_5591),
.B(n_5624),
.Y(n_7068)
);

INVx1_ASAP7_75t_L g7069 ( 
.A(n_6132),
.Y(n_7069)
);

BUFx2_ASAP7_75t_L g7070 ( 
.A(n_6723),
.Y(n_7070)
);

AND2x4_ASAP7_75t_L g7071 ( 
.A(n_6198),
.B(n_5684),
.Y(n_7071)
);

NOR2x1_ASAP7_75t_SL g7072 ( 
.A(n_6792),
.B(n_6333),
.Y(n_7072)
);

BUFx6f_ASAP7_75t_L g7073 ( 
.A(n_6554),
.Y(n_7073)
);

NAND2xp5_ASAP7_75t_L g7074 ( 
.A(n_6569),
.B(n_6674),
.Y(n_7074)
);

INVx1_ASAP7_75t_L g7075 ( 
.A(n_6132),
.Y(n_7075)
);

INVx1_ASAP7_75t_L g7076 ( 
.A(n_6143),
.Y(n_7076)
);

OAI21x1_ASAP7_75t_L g7077 ( 
.A1(n_6068),
.A2(n_5242),
.B(n_5189),
.Y(n_7077)
);

A2O1A1Ixp33_ASAP7_75t_L g7078 ( 
.A1(n_6505),
.A2(n_5427),
.B(n_6020),
.C(n_5293),
.Y(n_7078)
);

AND2x2_ASAP7_75t_L g7079 ( 
.A(n_6776),
.B(n_6737),
.Y(n_7079)
);

INVx2_ASAP7_75t_L g7080 ( 
.A(n_6640),
.Y(n_7080)
);

INVx1_ASAP7_75t_L g7081 ( 
.A(n_6143),
.Y(n_7081)
);

OAI21x1_ASAP7_75t_L g7082 ( 
.A1(n_6068),
.A2(n_5242),
.B(n_5189),
.Y(n_7082)
);

INVx2_ASAP7_75t_L g7083 ( 
.A(n_6640),
.Y(n_7083)
);

INVx1_ASAP7_75t_L g7084 ( 
.A(n_6143),
.Y(n_7084)
);

NAND2xp5_ASAP7_75t_L g7085 ( 
.A(n_6674),
.B(n_5546),
.Y(n_7085)
);

NAND2xp5_ASAP7_75t_L g7086 ( 
.A(n_6477),
.B(n_5548),
.Y(n_7086)
);

INVx1_ASAP7_75t_L g7087 ( 
.A(n_6153),
.Y(n_7087)
);

NOR2x1_ASAP7_75t_SL g7088 ( 
.A(n_6333),
.B(n_5385),
.Y(n_7088)
);

INVx2_ASAP7_75t_L g7089 ( 
.A(n_6386),
.Y(n_7089)
);

OAI21x1_ASAP7_75t_L g7090 ( 
.A1(n_6068),
.A2(n_5242),
.B(n_5189),
.Y(n_7090)
);

OR2x2_ASAP7_75t_L g7091 ( 
.A(n_6299),
.B(n_5343),
.Y(n_7091)
);

AND2x4_ASAP7_75t_L g7092 ( 
.A(n_6198),
.B(n_5761),
.Y(n_7092)
);

AOI21xp5_ASAP7_75t_L g7093 ( 
.A1(n_6046),
.A2(n_5635),
.B(n_5627),
.Y(n_7093)
);

NAND2xp5_ASAP7_75t_L g7094 ( 
.A(n_6477),
.B(n_5548),
.Y(n_7094)
);

NAND2xp5_ASAP7_75t_L g7095 ( 
.A(n_6092),
.B(n_6105),
.Y(n_7095)
);

OAI21x1_ASAP7_75t_L g7096 ( 
.A1(n_6073),
.A2(n_6183),
.B(n_6134),
.Y(n_7096)
);

INVx1_ASAP7_75t_L g7097 ( 
.A(n_6153),
.Y(n_7097)
);

OAI21x1_ASAP7_75t_L g7098 ( 
.A1(n_6073),
.A2(n_5304),
.B(n_5189),
.Y(n_7098)
);

INVx1_ASAP7_75t_L g7099 ( 
.A(n_6153),
.Y(n_7099)
);

OAI21x1_ASAP7_75t_L g7100 ( 
.A1(n_6073),
.A2(n_5357),
.B(n_5304),
.Y(n_7100)
);

NAND2xp5_ASAP7_75t_L g7101 ( 
.A(n_6092),
.B(n_5570),
.Y(n_7101)
);

INVx2_ASAP7_75t_L g7102 ( 
.A(n_6640),
.Y(n_7102)
);

NAND2xp5_ASAP7_75t_L g7103 ( 
.A(n_6105),
.B(n_5570),
.Y(n_7103)
);

NAND2xp5_ASAP7_75t_L g7104 ( 
.A(n_6149),
.B(n_5478),
.Y(n_7104)
);

OAI21x1_ASAP7_75t_L g7105 ( 
.A1(n_6073),
.A2(n_5357),
.B(n_5304),
.Y(n_7105)
);

INVx1_ASAP7_75t_L g7106 ( 
.A(n_6157),
.Y(n_7106)
);

OAI21x1_ASAP7_75t_L g7107 ( 
.A1(n_6073),
.A2(n_5357),
.B(n_5304),
.Y(n_7107)
);

BUFx3_ASAP7_75t_L g7108 ( 
.A(n_6554),
.Y(n_7108)
);

INVx2_ASAP7_75t_L g7109 ( 
.A(n_6386),
.Y(n_7109)
);

AO21x2_ASAP7_75t_L g7110 ( 
.A1(n_6212),
.A2(n_5496),
.B(n_5637),
.Y(n_7110)
);

AOI21xp5_ASAP7_75t_L g7111 ( 
.A1(n_6046),
.A2(n_6156),
.B(n_6249),
.Y(n_7111)
);

HB1xp67_ASAP7_75t_L g7112 ( 
.A(n_6761),
.Y(n_7112)
);

OAI21xp5_ASAP7_75t_L g7113 ( 
.A1(n_6402),
.A2(n_5495),
.B(n_5241),
.Y(n_7113)
);

AOI21xp5_ASAP7_75t_L g7114 ( 
.A1(n_6156),
.A2(n_6300),
.B(n_6230),
.Y(n_7114)
);

OAI21x1_ASAP7_75t_SL g7115 ( 
.A1(n_6777),
.A2(n_6447),
.B(n_6396),
.Y(n_7115)
);

AO31x2_ASAP7_75t_L g7116 ( 
.A1(n_6303),
.A2(n_5661),
.A3(n_5707),
.B(n_5697),
.Y(n_7116)
);

OAI21x1_ASAP7_75t_L g7117 ( 
.A1(n_6134),
.A2(n_5359),
.B(n_5357),
.Y(n_7117)
);

NAND2xp5_ASAP7_75t_L g7118 ( 
.A(n_6149),
.B(n_5478),
.Y(n_7118)
);

BUFx2_ASAP7_75t_R g7119 ( 
.A(n_6513),
.Y(n_7119)
);

A2O1A1Ixp33_ASAP7_75t_L g7120 ( 
.A1(n_6425),
.A2(n_5427),
.B(n_6020),
.C(n_5720),
.Y(n_7120)
);

AO21x2_ASAP7_75t_L g7121 ( 
.A1(n_6096),
.A2(n_5637),
.B(n_5911),
.Y(n_7121)
);

AO21x2_ASAP7_75t_L g7122 ( 
.A1(n_6096),
.A2(n_5637),
.B(n_5963),
.Y(n_7122)
);

AND2x2_ASAP7_75t_L g7123 ( 
.A(n_6776),
.B(n_5305),
.Y(n_7123)
);

BUFx3_ASAP7_75t_L g7124 ( 
.A(n_6554),
.Y(n_7124)
);

CKINVDCx11_ASAP7_75t_R g7125 ( 
.A(n_6242),
.Y(n_7125)
);

BUFx8_ASAP7_75t_L g7126 ( 
.A(n_6062),
.Y(n_7126)
);

AND2x2_ASAP7_75t_L g7127 ( 
.A(n_6737),
.B(n_5305),
.Y(n_7127)
);

INVx2_ASAP7_75t_L g7128 ( 
.A(n_6640),
.Y(n_7128)
);

INVx1_ASAP7_75t_L g7129 ( 
.A(n_6157),
.Y(n_7129)
);

OAI21xp5_ASAP7_75t_L g7130 ( 
.A1(n_6402),
.A2(n_5681),
.B(n_5297),
.Y(n_7130)
);

NAND2xp5_ASAP7_75t_L g7131 ( 
.A(n_6161),
.B(n_5485),
.Y(n_7131)
);

OAI21x1_ASAP7_75t_L g7132 ( 
.A1(n_6134),
.A2(n_5516),
.B(n_5359),
.Y(n_7132)
);

OAI21x1_ASAP7_75t_L g7133 ( 
.A1(n_6134),
.A2(n_5516),
.B(n_5359),
.Y(n_7133)
);

AO31x2_ASAP7_75t_L g7134 ( 
.A1(n_6434),
.A2(n_5707),
.A3(n_5734),
.B(n_5697),
.Y(n_7134)
);

OAI21x1_ASAP7_75t_L g7135 ( 
.A1(n_6134),
.A2(n_5516),
.B(n_5359),
.Y(n_7135)
);

NAND2xp5_ASAP7_75t_L g7136 ( 
.A(n_6161),
.B(n_5485),
.Y(n_7136)
);

OAI21x1_ASAP7_75t_L g7137 ( 
.A1(n_6183),
.A2(n_5604),
.B(n_5516),
.Y(n_7137)
);

AOI21x1_ASAP7_75t_L g7138 ( 
.A1(n_6115),
.A2(n_5753),
.B(n_5734),
.Y(n_7138)
);

NAND2xp5_ASAP7_75t_L g7139 ( 
.A(n_6180),
.B(n_5854),
.Y(n_7139)
);

INVx2_ASAP7_75t_L g7140 ( 
.A(n_6798),
.Y(n_7140)
);

AOI21xp33_ASAP7_75t_L g7141 ( 
.A1(n_6054),
.A2(n_5274),
.B(n_5273),
.Y(n_7141)
);

INVx3_ASAP7_75t_L g7142 ( 
.A(n_6038),
.Y(n_7142)
);

OA21x2_ASAP7_75t_L g7143 ( 
.A1(n_6064),
.A2(n_6005),
.B(n_5946),
.Y(n_7143)
);

AOI21x1_ASAP7_75t_L g7144 ( 
.A1(n_6270),
.A2(n_5789),
.B(n_5753),
.Y(n_7144)
);

AO21x2_ASAP7_75t_L g7145 ( 
.A1(n_6096),
.A2(n_5715),
.B(n_5752),
.Y(n_7145)
);

INVx1_ASAP7_75t_L g7146 ( 
.A(n_6157),
.Y(n_7146)
);

INVx1_ASAP7_75t_L g7147 ( 
.A(n_6163),
.Y(n_7147)
);

BUFx4f_ASAP7_75t_SL g7148 ( 
.A(n_6242),
.Y(n_7148)
);

NAND2xp5_ASAP7_75t_L g7149 ( 
.A(n_6180),
.B(n_5854),
.Y(n_7149)
);

AOI21xp5_ASAP7_75t_L g7150 ( 
.A1(n_6230),
.A2(n_6130),
.B(n_6757),
.Y(n_7150)
);

AND2x2_ASAP7_75t_L g7151 ( 
.A(n_6737),
.B(n_5391),
.Y(n_7151)
);

AOI22xp33_ASAP7_75t_L g7152 ( 
.A1(n_6151),
.A2(n_6054),
.B1(n_6269),
.B2(n_6032),
.Y(n_7152)
);

OA21x2_ASAP7_75t_L g7153 ( 
.A1(n_6064),
.A2(n_6060),
.B(n_6493),
.Y(n_7153)
);

BUFx8_ASAP7_75t_L g7154 ( 
.A(n_6204),
.Y(n_7154)
);

NAND2xp5_ASAP7_75t_L g7155 ( 
.A(n_6211),
.B(n_5511),
.Y(n_7155)
);

INVx1_ASAP7_75t_L g7156 ( 
.A(n_6163),
.Y(n_7156)
);

BUFx3_ASAP7_75t_L g7157 ( 
.A(n_6469),
.Y(n_7157)
);

INVx1_ASAP7_75t_L g7158 ( 
.A(n_6163),
.Y(n_7158)
);

AND2x2_ASAP7_75t_L g7159 ( 
.A(n_6334),
.B(n_5391),
.Y(n_7159)
);

INVx2_ASAP7_75t_L g7160 ( 
.A(n_6798),
.Y(n_7160)
);

INVx1_ASAP7_75t_L g7161 ( 
.A(n_6171),
.Y(n_7161)
);

BUFx2_ASAP7_75t_L g7162 ( 
.A(n_6723),
.Y(n_7162)
);

OAI22xp5_ASAP7_75t_L g7163 ( 
.A1(n_6032),
.A2(n_5681),
.B1(n_5967),
.B2(n_5536),
.Y(n_7163)
);

NAND2xp5_ASAP7_75t_L g7164 ( 
.A(n_6211),
.B(n_5511),
.Y(n_7164)
);

AO21x2_ASAP7_75t_L g7165 ( 
.A1(n_6754),
.A2(n_5752),
.B(n_5921),
.Y(n_7165)
);

INVx1_ASAP7_75t_L g7166 ( 
.A(n_6171),
.Y(n_7166)
);

NAND2xp5_ASAP7_75t_L g7167 ( 
.A(n_6425),
.B(n_5527),
.Y(n_7167)
);

OA21x2_ASAP7_75t_L g7168 ( 
.A1(n_6060),
.A2(n_6005),
.B(n_5946),
.Y(n_7168)
);

AOI211xp5_ASAP7_75t_SL g7169 ( 
.A1(n_6370),
.A2(n_6023),
.B(n_5790),
.C(n_5791),
.Y(n_7169)
);

INVx2_ASAP7_75t_L g7170 ( 
.A(n_6798),
.Y(n_7170)
);

OAI22xp33_ASAP7_75t_L g7171 ( 
.A1(n_6334),
.A2(n_6010),
.B1(n_5953),
.B2(n_5783),
.Y(n_7171)
);

INVx2_ASAP7_75t_L g7172 ( 
.A(n_6798),
.Y(n_7172)
);

AND2x2_ASAP7_75t_L g7173 ( 
.A(n_6377),
.B(n_5418),
.Y(n_7173)
);

AND2x4_ASAP7_75t_L g7174 ( 
.A(n_6198),
.B(n_5761),
.Y(n_7174)
);

AO21x2_ASAP7_75t_L g7175 ( 
.A1(n_6754),
.A2(n_5921),
.B(n_5307),
.Y(n_7175)
);

AO31x2_ASAP7_75t_L g7176 ( 
.A1(n_6318),
.A2(n_5803),
.A3(n_5924),
.B(n_5789),
.Y(n_7176)
);

INVx2_ASAP7_75t_L g7177 ( 
.A(n_6798),
.Y(n_7177)
);

INVx3_ASAP7_75t_L g7178 ( 
.A(n_6038),
.Y(n_7178)
);

OAI21x1_ASAP7_75t_L g7179 ( 
.A1(n_6183),
.A2(n_5643),
.B(n_5604),
.Y(n_7179)
);

AOI21x1_ASAP7_75t_L g7180 ( 
.A1(n_6301),
.A2(n_6391),
.B(n_6389),
.Y(n_7180)
);

INVx3_ASAP7_75t_L g7181 ( 
.A(n_6038),
.Y(n_7181)
);

INVx1_ASAP7_75t_L g7182 ( 
.A(n_6171),
.Y(n_7182)
);

OAI21x1_ASAP7_75t_L g7183 ( 
.A1(n_6183),
.A2(n_5643),
.B(n_5604),
.Y(n_7183)
);

INVx1_ASAP7_75t_L g7184 ( 
.A(n_6177),
.Y(n_7184)
);

OAI21x1_ASAP7_75t_L g7185 ( 
.A1(n_6183),
.A2(n_5643),
.B(n_5604),
.Y(n_7185)
);

INVx1_ASAP7_75t_L g7186 ( 
.A(n_6177),
.Y(n_7186)
);

INVx2_ASAP7_75t_L g7187 ( 
.A(n_6386),
.Y(n_7187)
);

OAI21x1_ASAP7_75t_L g7188 ( 
.A1(n_6233),
.A2(n_5735),
.B(n_5643),
.Y(n_7188)
);

INVx1_ASAP7_75t_L g7189 ( 
.A(n_6177),
.Y(n_7189)
);

AOI21xp5_ASAP7_75t_L g7190 ( 
.A1(n_6130),
.A2(n_6022),
.B(n_5767),
.Y(n_7190)
);

INVx2_ASAP7_75t_L g7191 ( 
.A(n_6406),
.Y(n_7191)
);

OAI21xp5_ASAP7_75t_L g7192 ( 
.A1(n_6146),
.A2(n_5573),
.B(n_5712),
.Y(n_7192)
);

NOR2xp33_ASAP7_75t_L g7193 ( 
.A(n_6168),
.B(n_5256),
.Y(n_7193)
);

INVx1_ASAP7_75t_L g7194 ( 
.A(n_6179),
.Y(n_7194)
);

INVx1_ASAP7_75t_L g7195 ( 
.A(n_6179),
.Y(n_7195)
);

INVx2_ASAP7_75t_L g7196 ( 
.A(n_6406),
.Y(n_7196)
);

AOI21xp5_ASAP7_75t_L g7197 ( 
.A1(n_6757),
.A2(n_6022),
.B(n_5200),
.Y(n_7197)
);

AO31x2_ASAP7_75t_L g7198 ( 
.A1(n_6318),
.A2(n_5924),
.A3(n_5803),
.B(n_5836),
.Y(n_7198)
);

INVx1_ASAP7_75t_L g7199 ( 
.A(n_6179),
.Y(n_7199)
);

NOR2x1_ASAP7_75t_SL g7200 ( 
.A(n_6333),
.B(n_5385),
.Y(n_7200)
);

BUFx2_ASAP7_75t_L g7201 ( 
.A(n_6723),
.Y(n_7201)
);

OAI21x1_ASAP7_75t_L g7202 ( 
.A1(n_6233),
.A2(n_5768),
.B(n_5735),
.Y(n_7202)
);

AO21x2_ASAP7_75t_L g7203 ( 
.A1(n_6771),
.A2(n_5921),
.B(n_5307),
.Y(n_7203)
);

BUFx8_ASAP7_75t_L g7204 ( 
.A(n_6204),
.Y(n_7204)
);

HB1xp67_ASAP7_75t_L g7205 ( 
.A(n_6761),
.Y(n_7205)
);

AO21x2_ASAP7_75t_L g7206 ( 
.A1(n_6771),
.A2(n_5921),
.B(n_5307),
.Y(n_7206)
);

AND2x2_ASAP7_75t_L g7207 ( 
.A(n_6377),
.B(n_5418),
.Y(n_7207)
);

INVx1_ASAP7_75t_L g7208 ( 
.A(n_6186),
.Y(n_7208)
);

NAND2xp5_ASAP7_75t_L g7209 ( 
.A(n_6030),
.B(n_5527),
.Y(n_7209)
);

AO31x2_ASAP7_75t_L g7210 ( 
.A1(n_6451),
.A2(n_5836),
.A3(n_5861),
.B(n_5833),
.Y(n_7210)
);

INVx4_ASAP7_75t_L g7211 ( 
.A(n_6168),
.Y(n_7211)
);

OAI21x1_ASAP7_75t_L g7212 ( 
.A1(n_6233),
.A2(n_5768),
.B(n_5735),
.Y(n_7212)
);

INVx1_ASAP7_75t_L g7213 ( 
.A(n_6186),
.Y(n_7213)
);

BUFx8_ASAP7_75t_L g7214 ( 
.A(n_6427),
.Y(n_7214)
);

AOI21xp5_ASAP7_75t_L g7215 ( 
.A1(n_6137),
.A2(n_6022),
.B(n_5200),
.Y(n_7215)
);

INVx2_ASAP7_75t_L g7216 ( 
.A(n_6314),
.Y(n_7216)
);

OAI21x1_ASAP7_75t_L g7217 ( 
.A1(n_6233),
.A2(n_5768),
.B(n_5735),
.Y(n_7217)
);

OAI21x1_ASAP7_75t_L g7218 ( 
.A1(n_6233),
.A2(n_5846),
.B(n_5768),
.Y(n_7218)
);

OAI21x1_ASAP7_75t_L g7219 ( 
.A1(n_6397),
.A2(n_5850),
.B(n_5846),
.Y(n_7219)
);

OAI21x1_ASAP7_75t_L g7220 ( 
.A1(n_6397),
.A2(n_5850),
.B(n_5846),
.Y(n_7220)
);

NAND2xp5_ASAP7_75t_L g7221 ( 
.A(n_6030),
.B(n_6021),
.Y(n_7221)
);

OAI21x1_ASAP7_75t_L g7222 ( 
.A1(n_6397),
.A2(n_5850),
.B(n_5846),
.Y(n_7222)
);

NAND2xp5_ASAP7_75t_L g7223 ( 
.A(n_6221),
.B(n_6021),
.Y(n_7223)
);

INVx2_ASAP7_75t_L g7224 ( 
.A(n_6406),
.Y(n_7224)
);

INVx1_ASAP7_75t_L g7225 ( 
.A(n_6186),
.Y(n_7225)
);

INVx3_ASAP7_75t_L g7226 ( 
.A(n_6038),
.Y(n_7226)
);

OA21x2_ASAP7_75t_L g7227 ( 
.A1(n_6493),
.A2(n_5949),
.B(n_5945),
.Y(n_7227)
);

INVx3_ASAP7_75t_L g7228 ( 
.A(n_6040),
.Y(n_7228)
);

OAI21x1_ASAP7_75t_L g7229 ( 
.A1(n_6397),
.A2(n_6474),
.B(n_6458),
.Y(n_7229)
);

CKINVDCx5p33_ASAP7_75t_R g7230 ( 
.A(n_6368),
.Y(n_7230)
);

AO31x2_ASAP7_75t_L g7231 ( 
.A1(n_6451),
.A2(n_5867),
.A3(n_5868),
.B(n_5861),
.Y(n_7231)
);

INVx1_ASAP7_75t_L g7232 ( 
.A(n_6192),
.Y(n_7232)
);

INVx2_ASAP7_75t_L g7233 ( 
.A(n_6314),
.Y(n_7233)
);

INVx2_ASAP7_75t_L g7234 ( 
.A(n_6314),
.Y(n_7234)
);

INVx2_ASAP7_75t_L g7235 ( 
.A(n_6314),
.Y(n_7235)
);

INVx1_ASAP7_75t_L g7236 ( 
.A(n_6192),
.Y(n_7236)
);

OAI21x1_ASAP7_75t_L g7237 ( 
.A1(n_6397),
.A2(n_5879),
.B(n_5850),
.Y(n_7237)
);

INVx5_ASAP7_75t_L g7238 ( 
.A(n_6040),
.Y(n_7238)
);

NAND2xp5_ASAP7_75t_L g7239 ( 
.A(n_6221),
.B(n_5758),
.Y(n_7239)
);

INVx1_ASAP7_75t_L g7240 ( 
.A(n_6192),
.Y(n_7240)
);

NOR2xp33_ASAP7_75t_L g7241 ( 
.A(n_6427),
.B(n_6584),
.Y(n_7241)
);

AND2x4_ASAP7_75t_L g7242 ( 
.A(n_6198),
.B(n_5761),
.Y(n_7242)
);

INVx2_ASAP7_75t_L g7243 ( 
.A(n_6315),
.Y(n_7243)
);

NAND2xp5_ASAP7_75t_L g7244 ( 
.A(n_6675),
.B(n_5758),
.Y(n_7244)
);

INVx1_ASAP7_75t_L g7245 ( 
.A(n_6199),
.Y(n_7245)
);

INVx1_ASAP7_75t_L g7246 ( 
.A(n_6199),
.Y(n_7246)
);

OAI21x1_ASAP7_75t_L g7247 ( 
.A1(n_6458),
.A2(n_5891),
.B(n_5879),
.Y(n_7247)
);

INVx1_ASAP7_75t_L g7248 ( 
.A(n_6199),
.Y(n_7248)
);

OAI21xp5_ASAP7_75t_L g7249 ( 
.A1(n_6295),
.A2(n_5492),
.B(n_5698),
.Y(n_7249)
);

CKINVDCx5p33_ASAP7_75t_R g7250 ( 
.A(n_6368),
.Y(n_7250)
);

NAND2xp5_ASAP7_75t_L g7251 ( 
.A(n_6675),
.B(n_5483),
.Y(n_7251)
);

NOR2xp33_ASAP7_75t_L g7252 ( 
.A(n_6584),
.B(n_5256),
.Y(n_7252)
);

OAI21x1_ASAP7_75t_L g7253 ( 
.A1(n_6458),
.A2(n_5891),
.B(n_5879),
.Y(n_7253)
);

INVx2_ASAP7_75t_L g7254 ( 
.A(n_6315),
.Y(n_7254)
);

NAND2x1p5_ASAP7_75t_L g7255 ( 
.A(n_6573),
.B(n_5400),
.Y(n_7255)
);

OA21x2_ASAP7_75t_L g7256 ( 
.A1(n_6086),
.A2(n_5949),
.B(n_5945),
.Y(n_7256)
);

NAND2xp5_ASAP7_75t_L g7257 ( 
.A(n_6712),
.B(n_5483),
.Y(n_7257)
);

OA21x2_ASAP7_75t_L g7258 ( 
.A1(n_6086),
.A2(n_5974),
.B(n_5955),
.Y(n_7258)
);

OAI21x1_ASAP7_75t_L g7259 ( 
.A1(n_6458),
.A2(n_5891),
.B(n_5879),
.Y(n_7259)
);

INVx1_ASAP7_75t_L g7260 ( 
.A(n_6223),
.Y(n_7260)
);

A2O1A1Ixp33_ASAP7_75t_L g7261 ( 
.A1(n_6453),
.A2(n_5720),
.B(n_5279),
.C(n_6015),
.Y(n_7261)
);

INVx2_ASAP7_75t_L g7262 ( 
.A(n_6315),
.Y(n_7262)
);

INVx1_ASAP7_75t_L g7263 ( 
.A(n_6223),
.Y(n_7263)
);

INVx1_ASAP7_75t_L g7264 ( 
.A(n_6223),
.Y(n_7264)
);

INVx1_ASAP7_75t_L g7265 ( 
.A(n_6226),
.Y(n_7265)
);

INVx2_ASAP7_75t_L g7266 ( 
.A(n_6315),
.Y(n_7266)
);

INVx1_ASAP7_75t_L g7267 ( 
.A(n_6226),
.Y(n_7267)
);

AOI21xp5_ASAP7_75t_L g7268 ( 
.A1(n_6137),
.A2(n_6022),
.B(n_5200),
.Y(n_7268)
);

HB1xp67_ASAP7_75t_L g7269 ( 
.A(n_6768),
.Y(n_7269)
);

INVx1_ASAP7_75t_L g7270 ( 
.A(n_6226),
.Y(n_7270)
);

AO31x2_ASAP7_75t_L g7271 ( 
.A1(n_6122),
.A2(n_6148),
.A3(n_6107),
.B(n_6295),
.Y(n_7271)
);

INVx1_ASAP7_75t_L g7272 ( 
.A(n_6229),
.Y(n_7272)
);

NOR2x1_ASAP7_75t_SL g7273 ( 
.A(n_6228),
.B(n_5385),
.Y(n_7273)
);

INVx1_ASAP7_75t_L g7274 ( 
.A(n_6229),
.Y(n_7274)
);

AOI21x1_ASAP7_75t_L g7275 ( 
.A1(n_6389),
.A2(n_5352),
.B(n_5340),
.Y(n_7275)
);

OA21x2_ASAP7_75t_L g7276 ( 
.A1(n_6086),
.A2(n_6248),
.B(n_6247),
.Y(n_7276)
);

INVx1_ASAP7_75t_L g7277 ( 
.A(n_6229),
.Y(n_7277)
);

INVx2_ASAP7_75t_L g7278 ( 
.A(n_6316),
.Y(n_7278)
);

NAND2x1p5_ASAP7_75t_L g7279 ( 
.A(n_6508),
.B(n_5400),
.Y(n_7279)
);

AND2x2_ASAP7_75t_L g7280 ( 
.A(n_6377),
.B(n_6378),
.Y(n_7280)
);

BUFx2_ASAP7_75t_L g7281 ( 
.A(n_6723),
.Y(n_7281)
);

HB1xp67_ASAP7_75t_L g7282 ( 
.A(n_6768),
.Y(n_7282)
);

OAI21x1_ASAP7_75t_L g7283 ( 
.A1(n_6458),
.A2(n_6016),
.B(n_5891),
.Y(n_7283)
);

AO21x2_ASAP7_75t_L g7284 ( 
.A1(n_6347),
.A2(n_5307),
.B(n_5955),
.Y(n_7284)
);

INVx1_ASAP7_75t_L g7285 ( 
.A(n_6252),
.Y(n_7285)
);

INVx1_ASAP7_75t_L g7286 ( 
.A(n_6252),
.Y(n_7286)
);

OAI22xp5_ASAP7_75t_L g7287 ( 
.A1(n_6564),
.A2(n_5975),
.B1(n_6010),
.B2(n_5953),
.Y(n_7287)
);

HB1xp67_ASAP7_75t_L g7288 ( 
.A(n_6663),
.Y(n_7288)
);

OA21x2_ASAP7_75t_L g7289 ( 
.A1(n_6247),
.A2(n_5981),
.B(n_5974),
.Y(n_7289)
);

NAND2xp5_ASAP7_75t_L g7290 ( 
.A(n_6712),
.B(n_5796),
.Y(n_7290)
);

OAI21x1_ASAP7_75t_L g7291 ( 
.A1(n_6474),
.A2(n_6016),
.B(n_5984),
.Y(n_7291)
);

INVx2_ASAP7_75t_L g7292 ( 
.A(n_6406),
.Y(n_7292)
);

AOI21xp5_ASAP7_75t_L g7293 ( 
.A1(n_6137),
.A2(n_5200),
.B(n_5809),
.Y(n_7293)
);

OAI21x1_ASAP7_75t_L g7294 ( 
.A1(n_6474),
.A2(n_6016),
.B(n_5984),
.Y(n_7294)
);

OAI21x1_ASAP7_75t_SL g7295 ( 
.A1(n_6396),
.A2(n_5222),
.B(n_5209),
.Y(n_7295)
);

NOR2xp33_ASAP7_75t_L g7296 ( 
.A(n_6584),
.B(n_5256),
.Y(n_7296)
);

AOI21xp5_ASAP7_75t_L g7297 ( 
.A1(n_6137),
.A2(n_5200),
.B(n_5818),
.Y(n_7297)
);

INVx1_ASAP7_75t_L g7298 ( 
.A(n_6252),
.Y(n_7298)
);

CKINVDCx5p33_ASAP7_75t_R g7299 ( 
.A(n_6335),
.Y(n_7299)
);

NAND2xp5_ASAP7_75t_L g7300 ( 
.A(n_6577),
.B(n_5862),
.Y(n_7300)
);

INVx1_ASAP7_75t_L g7301 ( 
.A(n_6267),
.Y(n_7301)
);

CKINVDCx20_ASAP7_75t_R g7302 ( 
.A(n_6700),
.Y(n_7302)
);

OAI21x1_ASAP7_75t_L g7303 ( 
.A1(n_6474),
.A2(n_6016),
.B(n_5993),
.Y(n_7303)
);

INVx6_ASAP7_75t_L g7304 ( 
.A(n_6039),
.Y(n_7304)
);

OAI21xp5_ASAP7_75t_L g7305 ( 
.A1(n_6478),
.A2(n_6256),
.B(n_6538),
.Y(n_7305)
);

INVx1_ASAP7_75t_L g7306 ( 
.A(n_6267),
.Y(n_7306)
);

INVx3_ASAP7_75t_L g7307 ( 
.A(n_6040),
.Y(n_7307)
);

AO31x2_ASAP7_75t_L g7308 ( 
.A1(n_6122),
.A2(n_5868),
.A3(n_5872),
.B(n_5867),
.Y(n_7308)
);

OAI21x1_ASAP7_75t_L g7309 ( 
.A1(n_6474),
.A2(n_5993),
.B(n_5976),
.Y(n_7309)
);

AOI21xp5_ASAP7_75t_L g7310 ( 
.A1(n_6137),
.A2(n_5194),
.B(n_6004),
.Y(n_7310)
);

AO21x1_ASAP7_75t_L g7311 ( 
.A1(n_6114),
.A2(n_5222),
.B(n_5209),
.Y(n_7311)
);

INVx3_ASAP7_75t_L g7312 ( 
.A(n_6040),
.Y(n_7312)
);

INVx2_ASAP7_75t_L g7313 ( 
.A(n_6316),
.Y(n_7313)
);

NAND2xp5_ASAP7_75t_L g7314 ( 
.A(n_6577),
.B(n_5538),
.Y(n_7314)
);

INVx2_ASAP7_75t_L g7315 ( 
.A(n_6316),
.Y(n_7315)
);

INVx2_ASAP7_75t_L g7316 ( 
.A(n_6316),
.Y(n_7316)
);

AO21x2_ASAP7_75t_L g7317 ( 
.A1(n_6347),
.A2(n_5981),
.B(n_5250),
.Y(n_7317)
);

AND2x2_ASAP7_75t_L g7318 ( 
.A(n_6377),
.B(n_5625),
.Y(n_7318)
);

AOI22xp33_ASAP7_75t_L g7319 ( 
.A1(n_6269),
.A2(n_5876),
.B1(n_5915),
.B2(n_5856),
.Y(n_7319)
);

OAI21x1_ASAP7_75t_SL g7320 ( 
.A1(n_6396),
.A2(n_5222),
.B(n_5193),
.Y(n_7320)
);

AO21x2_ASAP7_75t_L g7321 ( 
.A1(n_6313),
.A2(n_5250),
.B(n_5225),
.Y(n_7321)
);

BUFx2_ASAP7_75t_L g7322 ( 
.A(n_6723),
.Y(n_7322)
);

BUFx8_ASAP7_75t_L g7323 ( 
.A(n_6051),
.Y(n_7323)
);

INVx4_ASAP7_75t_L g7324 ( 
.A(n_6182),
.Y(n_7324)
);

NAND2xp5_ASAP7_75t_L g7325 ( 
.A(n_6598),
.B(n_5538),
.Y(n_7325)
);

AND2x4_ASAP7_75t_L g7326 ( 
.A(n_6272),
.B(n_5761),
.Y(n_7326)
);

AOI21xp5_ASAP7_75t_L g7327 ( 
.A1(n_6182),
.A2(n_5194),
.B(n_5821),
.Y(n_7327)
);

OA21x2_ASAP7_75t_L g7328 ( 
.A1(n_6247),
.A2(n_5702),
.B(n_5700),
.Y(n_7328)
);

BUFx2_ASAP7_75t_L g7329 ( 
.A(n_6717),
.Y(n_7329)
);

AO31x2_ASAP7_75t_L g7330 ( 
.A1(n_6148),
.A2(n_5934),
.A3(n_5941),
.B(n_5872),
.Y(n_7330)
);

AND2x4_ASAP7_75t_L g7331 ( 
.A(n_6272),
.B(n_5851),
.Y(n_7331)
);

OAI21xp5_ASAP7_75t_L g7332 ( 
.A1(n_6478),
.A2(n_5194),
.B(n_5695),
.Y(n_7332)
);

NAND2xp5_ASAP7_75t_L g7333 ( 
.A(n_6598),
.B(n_5619),
.Y(n_7333)
);

AO31x2_ASAP7_75t_L g7334 ( 
.A1(n_6107),
.A2(n_5941),
.A3(n_5947),
.B(n_5934),
.Y(n_7334)
);

AO21x2_ASAP7_75t_L g7335 ( 
.A1(n_6313),
.A2(n_5265),
.B(n_5225),
.Y(n_7335)
);

BUFx10_ASAP7_75t_L g7336 ( 
.A(n_6753),
.Y(n_7336)
);

OR2x6_ASAP7_75t_SL g7337 ( 
.A(n_6632),
.B(n_5588),
.Y(n_7337)
);

AOI21x1_ASAP7_75t_L g7338 ( 
.A1(n_6391),
.A2(n_5352),
.B(n_5340),
.Y(n_7338)
);

BUFx2_ASAP7_75t_L g7339 ( 
.A(n_6717),
.Y(n_7339)
);

AND2x4_ASAP7_75t_L g7340 ( 
.A(n_6272),
.B(n_5851),
.Y(n_7340)
);

AO21x2_ASAP7_75t_L g7341 ( 
.A1(n_6520),
.A2(n_5266),
.B(n_5265),
.Y(n_7341)
);

OAI21x1_ASAP7_75t_L g7342 ( 
.A1(n_6504),
.A2(n_5976),
.B(n_5995),
.Y(n_7342)
);

AO21x2_ASAP7_75t_L g7343 ( 
.A1(n_6520),
.A2(n_6202),
.B(n_6331),
.Y(n_7343)
);

OAI22xp5_ASAP7_75t_L g7344 ( 
.A1(n_6564),
.A2(n_5711),
.B1(n_5998),
.B2(n_5986),
.Y(n_7344)
);

INVx3_ASAP7_75t_L g7345 ( 
.A(n_6040),
.Y(n_7345)
);

AOI21xp5_ASAP7_75t_L g7346 ( 
.A1(n_6182),
.A2(n_5821),
.B(n_5808),
.Y(n_7346)
);

AOI22xp33_ASAP7_75t_L g7347 ( 
.A1(n_6269),
.A2(n_5915),
.B1(n_5876),
.B2(n_5291),
.Y(n_7347)
);

NAND2xp5_ASAP7_75t_L g7348 ( 
.A(n_6538),
.B(n_5619),
.Y(n_7348)
);

NAND2xp5_ASAP7_75t_L g7349 ( 
.A(n_6601),
.B(n_5571),
.Y(n_7349)
);

AO21x2_ASAP7_75t_L g7350 ( 
.A1(n_6202),
.A2(n_5266),
.B(n_5900),
.Y(n_7350)
);

INVx1_ASAP7_75t_L g7351 ( 
.A(n_6267),
.Y(n_7351)
);

AND2x4_ASAP7_75t_L g7352 ( 
.A(n_6272),
.B(n_5851),
.Y(n_7352)
);

AOI22xp5_ASAP7_75t_L g7353 ( 
.A1(n_6342),
.A2(n_5781),
.B1(n_5828),
.B2(n_5783),
.Y(n_7353)
);

AO21x2_ASAP7_75t_L g7354 ( 
.A1(n_6331),
.A2(n_5905),
.B(n_5900),
.Y(n_7354)
);

NAND2xp5_ASAP7_75t_L g7355 ( 
.A(n_6601),
.B(n_5571),
.Y(n_7355)
);

OAI21x1_ASAP7_75t_L g7356 ( 
.A1(n_6504),
.A2(n_5995),
.B(n_5148),
.Y(n_7356)
);

INVx2_ASAP7_75t_L g7357 ( 
.A(n_6352),
.Y(n_7357)
);

OA21x2_ASAP7_75t_L g7358 ( 
.A1(n_6248),
.A2(n_5403),
.B(n_5905),
.Y(n_7358)
);

OR2x2_ASAP7_75t_L g7359 ( 
.A(n_6369),
.B(n_6330),
.Y(n_7359)
);

NOR2x1_ASAP7_75t_SL g7360 ( 
.A(n_6228),
.B(n_6340),
.Y(n_7360)
);

INVx1_ASAP7_75t_L g7361 ( 
.A(n_6275),
.Y(n_7361)
);

INVx1_ASAP7_75t_L g7362 ( 
.A(n_6275),
.Y(n_7362)
);

XOR2xp5_ASAP7_75t_L g7363 ( 
.A(n_6700),
.B(n_5512),
.Y(n_7363)
);

INVx1_ASAP7_75t_L g7364 ( 
.A(n_6275),
.Y(n_7364)
);

INVx1_ASAP7_75t_L g7365 ( 
.A(n_6279),
.Y(n_7365)
);

AO31x2_ASAP7_75t_L g7366 ( 
.A1(n_6185),
.A2(n_5971),
.A3(n_5979),
.B(n_5947),
.Y(n_7366)
);

INVx1_ASAP7_75t_L g7367 ( 
.A(n_6279),
.Y(n_7367)
);

NAND2xp5_ASAP7_75t_L g7368 ( 
.A(n_6256),
.B(n_5576),
.Y(n_7368)
);

OR2x2_ASAP7_75t_L g7369 ( 
.A(n_6369),
.B(n_5343),
.Y(n_7369)
);

AND2x2_ASAP7_75t_L g7370 ( 
.A(n_6377),
.B(n_5625),
.Y(n_7370)
);

AOI21x1_ASAP7_75t_L g7371 ( 
.A1(n_6392),
.A2(n_5377),
.B(n_5352),
.Y(n_7371)
);

AO21x2_ASAP7_75t_L g7372 ( 
.A1(n_6331),
.A2(n_5979),
.B(n_5971),
.Y(n_7372)
);

NAND2xp5_ASAP7_75t_L g7373 ( 
.A(n_6413),
.B(n_5576),
.Y(n_7373)
);

NAND2xp5_ASAP7_75t_L g7374 ( 
.A(n_6413),
.B(n_5181),
.Y(n_7374)
);

INVx1_ASAP7_75t_L g7375 ( 
.A(n_6279),
.Y(n_7375)
);

NOR2xp33_ASAP7_75t_L g7376 ( 
.A(n_6658),
.B(n_5256),
.Y(n_7376)
);

INVx1_ASAP7_75t_L g7377 ( 
.A(n_6282),
.Y(n_7377)
);

OAI22xp5_ASAP7_75t_L g7378 ( 
.A1(n_6138),
.A2(n_5711),
.B1(n_5279),
.B2(n_5835),
.Y(n_7378)
);

OAI21x1_ASAP7_75t_L g7379 ( 
.A1(n_6504),
.A2(n_5148),
.B(n_5467),
.Y(n_7379)
);

HB1xp67_ASAP7_75t_L g7380 ( 
.A(n_6663),
.Y(n_7380)
);

HB1xp67_ASAP7_75t_L g7381 ( 
.A(n_6706),
.Y(n_7381)
);

AOI21xp5_ASAP7_75t_L g7382 ( 
.A1(n_6182),
.A2(n_5804),
.B(n_5845),
.Y(n_7382)
);

A2O1A1Ixp33_ASAP7_75t_L g7383 ( 
.A1(n_6453),
.A2(n_5279),
.B(n_5881),
.C(n_5880),
.Y(n_7383)
);

AOI21xp5_ASAP7_75t_L g7384 ( 
.A1(n_6182),
.A2(n_5895),
.B(n_5864),
.Y(n_7384)
);

NAND2x1p5_ASAP7_75t_L g7385 ( 
.A(n_6508),
.B(n_5148),
.Y(n_7385)
);

NOR2xp33_ASAP7_75t_L g7386 ( 
.A(n_6658),
.B(n_5668),
.Y(n_7386)
);

INVx1_ASAP7_75t_L g7387 ( 
.A(n_6282),
.Y(n_7387)
);

OAI21xp5_ASAP7_75t_L g7388 ( 
.A1(n_6460),
.A2(n_5466),
.B(n_5484),
.Y(n_7388)
);

OAI21x1_ASAP7_75t_L g7389 ( 
.A1(n_6504),
.A2(n_5148),
.B(n_5467),
.Y(n_7389)
);

INVx1_ASAP7_75t_SL g7390 ( 
.A(n_6660),
.Y(n_7390)
);

INVx1_ASAP7_75t_L g7391 ( 
.A(n_6282),
.Y(n_7391)
);

AOI21xp5_ASAP7_75t_L g7392 ( 
.A1(n_6442),
.A2(n_5899),
.B(n_5983),
.Y(n_7392)
);

INVx3_ASAP7_75t_L g7393 ( 
.A(n_6040),
.Y(n_7393)
);

NAND2xp5_ASAP7_75t_L g7394 ( 
.A(n_6439),
.B(n_5181),
.Y(n_7394)
);

AO31x2_ASAP7_75t_L g7395 ( 
.A1(n_6185),
.A2(n_6025),
.A3(n_6027),
.B(n_5996),
.Y(n_7395)
);

INVx3_ASAP7_75t_L g7396 ( 
.A(n_6040),
.Y(n_7396)
);

AO21x2_ASAP7_75t_L g7397 ( 
.A1(n_6166),
.A2(n_6025),
.B(n_5996),
.Y(n_7397)
);

INVx1_ASAP7_75t_L g7398 ( 
.A(n_6291),
.Y(n_7398)
);

AND2x4_ASAP7_75t_L g7399 ( 
.A(n_6272),
.B(n_5851),
.Y(n_7399)
);

NAND2xp5_ASAP7_75t_L g7400 ( 
.A(n_6439),
.B(n_5246),
.Y(n_7400)
);

NOR2xp33_ASAP7_75t_R g7401 ( 
.A(n_6697),
.B(n_5512),
.Y(n_7401)
);

NAND2xp5_ASAP7_75t_L g7402 ( 
.A(n_6466),
.B(n_5246),
.Y(n_7402)
);

AOI21xp5_ASAP7_75t_L g7403 ( 
.A1(n_6442),
.A2(n_5987),
.B(n_5907),
.Y(n_7403)
);

AO21x2_ASAP7_75t_L g7404 ( 
.A1(n_6166),
.A2(n_6408),
.B(n_6353),
.Y(n_7404)
);

INVx1_ASAP7_75t_L g7405 ( 
.A(n_6291),
.Y(n_7405)
);

NOR2xp33_ASAP7_75t_L g7406 ( 
.A(n_6753),
.B(n_5668),
.Y(n_7406)
);

OAI21x1_ASAP7_75t_L g7407 ( 
.A1(n_6504),
.A2(n_5467),
.B(n_5799),
.Y(n_7407)
);

INVx1_ASAP7_75t_L g7408 ( 
.A(n_6291),
.Y(n_7408)
);

BUFx3_ASAP7_75t_L g7409 ( 
.A(n_6513),
.Y(n_7409)
);

A2O1A1Ixp33_ASAP7_75t_L g7410 ( 
.A1(n_6736),
.A2(n_5881),
.B(n_5937),
.C(n_5880),
.Y(n_7410)
);

OAI21xp5_ASAP7_75t_L g7411 ( 
.A1(n_6460),
.A2(n_6342),
.B(n_6356),
.Y(n_7411)
);

INVx1_ASAP7_75t_L g7412 ( 
.A(n_6302),
.Y(n_7412)
);

OAI21x1_ASAP7_75t_SL g7413 ( 
.A1(n_6447),
.A2(n_5223),
.B(n_5193),
.Y(n_7413)
);

OAI21xp5_ASAP7_75t_L g7414 ( 
.A1(n_6356),
.A2(n_5466),
.B(n_5589),
.Y(n_7414)
);

AOI21xp5_ASAP7_75t_L g7415 ( 
.A1(n_6643),
.A2(n_5594),
.B(n_5592),
.Y(n_7415)
);

OR2x2_ASAP7_75t_L g7416 ( 
.A(n_6330),
.B(n_5343),
.Y(n_7416)
);

AOI21xp5_ASAP7_75t_L g7417 ( 
.A1(n_6643),
.A2(n_5623),
.B(n_5600),
.Y(n_7417)
);

INVx1_ASAP7_75t_L g7418 ( 
.A(n_6302),
.Y(n_7418)
);

INVx1_ASAP7_75t_L g7419 ( 
.A(n_6302),
.Y(n_7419)
);

INVx1_ASAP7_75t_SL g7420 ( 
.A(n_6660),
.Y(n_7420)
);

AOI21xp5_ASAP7_75t_L g7421 ( 
.A1(n_6370),
.A2(n_6009),
.B(n_6007),
.Y(n_7421)
);

NAND2xp5_ASAP7_75t_L g7422 ( 
.A(n_6466),
.B(n_5633),
.Y(n_7422)
);

AND2x2_ASAP7_75t_L g7423 ( 
.A(n_6378),
.B(n_5728),
.Y(n_7423)
);

NAND2xp33_ASAP7_75t_L g7424 ( 
.A(n_6801),
.B(n_5228),
.Y(n_7424)
);

A2O1A1Ixp33_ASAP7_75t_L g7425 ( 
.A1(n_6736),
.A2(n_5937),
.B(n_5773),
.C(n_5823),
.Y(n_7425)
);

NAND2xp5_ASAP7_75t_L g7426 ( 
.A(n_6448),
.B(n_5699),
.Y(n_7426)
);

AOI21xp33_ASAP7_75t_SL g7427 ( 
.A1(n_6632),
.A2(n_5617),
.B(n_5606),
.Y(n_7427)
);

AOI21xp5_ASAP7_75t_L g7428 ( 
.A1(n_6290),
.A2(n_5823),
.B(n_5773),
.Y(n_7428)
);

OAI22xp5_ASAP7_75t_L g7429 ( 
.A1(n_6138),
.A2(n_5835),
.B1(n_5781),
.B2(n_5741),
.Y(n_7429)
);

AND2x4_ASAP7_75t_L g7430 ( 
.A(n_6272),
.B(n_5928),
.Y(n_7430)
);

INVx2_ASAP7_75t_L g7431 ( 
.A(n_6352),
.Y(n_7431)
);

AND2x4_ASAP7_75t_L g7432 ( 
.A(n_6272),
.B(n_5928),
.Y(n_7432)
);

BUFx6f_ASAP7_75t_L g7433 ( 
.A(n_6040),
.Y(n_7433)
);

BUFx6f_ASAP7_75t_L g7434 ( 
.A(n_6042),
.Y(n_7434)
);

INVx1_ASAP7_75t_L g7435 ( 
.A(n_6304),
.Y(n_7435)
);

OA21x2_ASAP7_75t_L g7436 ( 
.A1(n_6248),
.A2(n_6273),
.B(n_6147),
.Y(n_7436)
);

AOI22xp5_ASAP7_75t_L g7437 ( 
.A1(n_6043),
.A2(n_6219),
.B1(n_6053),
.B2(n_6398),
.Y(n_7437)
);

AOI22xp5_ASAP7_75t_L g7438 ( 
.A1(n_6043),
.A2(n_5828),
.B1(n_5915),
.B2(n_5876),
.Y(n_7438)
);

OAI21x1_ASAP7_75t_L g7439 ( 
.A1(n_6549),
.A2(n_5799),
.B(n_5394),
.Y(n_7439)
);

INVx1_ASAP7_75t_L g7440 ( 
.A(n_6304),
.Y(n_7440)
);

NAND2xp5_ASAP7_75t_L g7441 ( 
.A(n_6448),
.B(n_5906),
.Y(n_7441)
);

AOI21xp5_ASAP7_75t_L g7442 ( 
.A1(n_6290),
.A2(n_6519),
.B(n_6578),
.Y(n_7442)
);

BUFx6f_ASAP7_75t_L g7443 ( 
.A(n_6042),
.Y(n_7443)
);

AO31x2_ASAP7_75t_L g7444 ( 
.A1(n_6083),
.A2(n_6560),
.A3(n_6449),
.B(n_6691),
.Y(n_7444)
);

A2O1A1Ixp33_ASAP7_75t_L g7445 ( 
.A1(n_6280),
.A2(n_5904),
.B(n_5935),
.C(n_5403),
.Y(n_7445)
);

AOI21xp5_ASAP7_75t_L g7446 ( 
.A1(n_6519),
.A2(n_6578),
.B(n_6508),
.Y(n_7446)
);

AOI21xp5_ASAP7_75t_L g7447 ( 
.A1(n_6508),
.A2(n_5798),
.B(n_5795),
.Y(n_7447)
);

INVx1_ASAP7_75t_L g7448 ( 
.A(n_6304),
.Y(n_7448)
);

INVx2_ASAP7_75t_L g7449 ( 
.A(n_6352),
.Y(n_7449)
);

INVx1_ASAP7_75t_L g7450 ( 
.A(n_6309),
.Y(n_7450)
);

NAND2xp5_ASAP7_75t_L g7451 ( 
.A(n_6081),
.B(n_5906),
.Y(n_7451)
);

HB1xp67_ASAP7_75t_L g7452 ( 
.A(n_6706),
.Y(n_7452)
);

AOI21xp5_ASAP7_75t_L g7453 ( 
.A1(n_6508),
.A2(n_5530),
.B(n_5603),
.Y(n_7453)
);

OAI21x1_ASAP7_75t_L g7454 ( 
.A1(n_6549),
.A2(n_5799),
.B(n_5394),
.Y(n_7454)
);

AND2x4_ASAP7_75t_L g7455 ( 
.A(n_6446),
.B(n_5928),
.Y(n_7455)
);

AOI22xp5_ASAP7_75t_L g7456 ( 
.A1(n_6219),
.A2(n_5530),
.B1(n_5228),
.B2(n_5323),
.Y(n_7456)
);

CKINVDCx6p67_ASAP7_75t_R g7457 ( 
.A(n_6269),
.Y(n_7457)
);

AOI22xp33_ASAP7_75t_L g7458 ( 
.A1(n_6112),
.A2(n_5291),
.B1(n_5545),
.B2(n_5323),
.Y(n_7458)
);

AND2x2_ASAP7_75t_L g7459 ( 
.A(n_6378),
.B(n_5728),
.Y(n_7459)
);

INVx1_ASAP7_75t_L g7460 ( 
.A(n_6309),
.Y(n_7460)
);

AOI21xp5_ASAP7_75t_L g7461 ( 
.A1(n_6508),
.A2(n_6280),
.B(n_6590),
.Y(n_7461)
);

OAI21x1_ASAP7_75t_L g7462 ( 
.A1(n_6549),
.A2(n_5799),
.B(n_5394),
.Y(n_7462)
);

INVx3_ASAP7_75t_L g7463 ( 
.A(n_6042),
.Y(n_7463)
);

BUFx6f_ASAP7_75t_L g7464 ( 
.A(n_6042),
.Y(n_7464)
);

AOI21xp5_ASAP7_75t_L g7465 ( 
.A1(n_6590),
.A2(n_5603),
.B(n_5650),
.Y(n_7465)
);

NAND2x1p5_ASAP7_75t_L g7466 ( 
.A(n_6042),
.B(n_5215),
.Y(n_7466)
);

BUFx8_ASAP7_75t_L g7467 ( 
.A(n_6051),
.Y(n_7467)
);

INVx1_ASAP7_75t_L g7468 ( 
.A(n_6309),
.Y(n_7468)
);

OA21x2_ASAP7_75t_L g7469 ( 
.A1(n_6273),
.A2(n_5197),
.B(n_5176),
.Y(n_7469)
);

BUFx6f_ASAP7_75t_L g7470 ( 
.A(n_6042),
.Y(n_7470)
);

OA21x2_ASAP7_75t_L g7471 ( 
.A1(n_6273),
.A2(n_5197),
.B(n_5176),
.Y(n_7471)
);

INVx1_ASAP7_75t_L g7472 ( 
.A(n_6321),
.Y(n_7472)
);

AOI21xp5_ASAP7_75t_L g7473 ( 
.A1(n_6686),
.A2(n_5650),
.B(n_5215),
.Y(n_7473)
);

OAI21xp5_ASAP7_75t_L g7474 ( 
.A1(n_6356),
.A2(n_5660),
.B(n_5648),
.Y(n_7474)
);

BUFx3_ASAP7_75t_L g7475 ( 
.A(n_6801),
.Y(n_7475)
);

AO21x1_ASAP7_75t_SL g7476 ( 
.A1(n_6288),
.A2(n_5857),
.B(n_5871),
.Y(n_7476)
);

OAI21xp5_ASAP7_75t_L g7477 ( 
.A1(n_6286),
.A2(n_6463),
.B(n_6521),
.Y(n_7477)
);

OA21x2_ASAP7_75t_L g7478 ( 
.A1(n_6147),
.A2(n_5229),
.B(n_5206),
.Y(n_7478)
);

OA21x2_ASAP7_75t_L g7479 ( 
.A1(n_6147),
.A2(n_5229),
.B(n_5206),
.Y(n_7479)
);

OAI21x1_ASAP7_75t_L g7480 ( 
.A1(n_6549),
.A2(n_5414),
.B(n_5377),
.Y(n_7480)
);

AO31x2_ASAP7_75t_L g7481 ( 
.A1(n_6083),
.A2(n_6027),
.A3(n_5244),
.B(n_5268),
.Y(n_7481)
);

OAI21x1_ASAP7_75t_L g7482 ( 
.A1(n_6549),
.A2(n_5414),
.B(n_5377),
.Y(n_7482)
);

INVx1_ASAP7_75t_L g7483 ( 
.A(n_6321),
.Y(n_7483)
);

INVx1_ASAP7_75t_L g7484 ( 
.A(n_6321),
.Y(n_7484)
);

AOI21xp5_ASAP7_75t_L g7485 ( 
.A1(n_6686),
.A2(n_5215),
.B(n_5763),
.Y(n_7485)
);

OR2x2_ASAP7_75t_L g7486 ( 
.A(n_6332),
.B(n_6336),
.Y(n_7486)
);

INVx2_ASAP7_75t_L g7487 ( 
.A(n_6352),
.Y(n_7487)
);

INVx1_ASAP7_75t_L g7488 ( 
.A(n_6323),
.Y(n_7488)
);

NAND2xp5_ASAP7_75t_L g7489 ( 
.A(n_6081),
.B(n_5840),
.Y(n_7489)
);

NOR2xp33_ASAP7_75t_L g7490 ( 
.A(n_6672),
.B(n_6140),
.Y(n_7490)
);

AO21x2_ASAP7_75t_L g7491 ( 
.A1(n_6408),
.A2(n_6353),
.B(n_6514),
.Y(n_7491)
);

NAND2xp5_ASAP7_75t_L g7492 ( 
.A(n_6205),
.B(n_5840),
.Y(n_7492)
);

NAND2xp5_ASAP7_75t_SL g7493 ( 
.A(n_6672),
.B(n_5223),
.Y(n_7493)
);

NAND2xp5_ASAP7_75t_L g7494 ( 
.A(n_6205),
.B(n_5810),
.Y(n_7494)
);

OAI21x1_ASAP7_75t_L g7495 ( 
.A1(n_6464),
.A2(n_5420),
.B(n_5414),
.Y(n_7495)
);

AO21x2_ASAP7_75t_L g7496 ( 
.A1(n_6353),
.A2(n_5244),
.B(n_5230),
.Y(n_7496)
);

NOR2x1_ASAP7_75t_R g7497 ( 
.A(n_6033),
.B(n_5512),
.Y(n_7497)
);

INVx1_ASAP7_75t_L g7498 ( 
.A(n_6323),
.Y(n_7498)
);

NAND2xp5_ASAP7_75t_L g7499 ( 
.A(n_6417),
.B(n_5810),
.Y(n_7499)
);

INVx1_ASAP7_75t_L g7500 ( 
.A(n_6323),
.Y(n_7500)
);

AOI21xp5_ASAP7_75t_L g7501 ( 
.A1(n_6486),
.A2(n_5215),
.B(n_5763),
.Y(n_7501)
);

OAI21xp5_ASAP7_75t_L g7502 ( 
.A1(n_6286),
.A2(n_5660),
.B(n_5648),
.Y(n_7502)
);

INVx1_ASAP7_75t_L g7503 ( 
.A(n_6337),
.Y(n_7503)
);

OAI22xp5_ASAP7_75t_L g7504 ( 
.A1(n_6540),
.A2(n_5741),
.B1(n_6003),
.B2(n_5323),
.Y(n_7504)
);

BUFx3_ASAP7_75t_L g7505 ( 
.A(n_6051),
.Y(n_7505)
);

OAI21x1_ASAP7_75t_L g7506 ( 
.A1(n_6464),
.A2(n_5430),
.B(n_5420),
.Y(n_7506)
);

OR2x2_ASAP7_75t_L g7507 ( 
.A(n_6332),
.B(n_5343),
.Y(n_7507)
);

BUFx6f_ASAP7_75t_L g7508 ( 
.A(n_6042),
.Y(n_7508)
);

OAI21x1_ASAP7_75t_L g7509 ( 
.A1(n_6464),
.A2(n_5430),
.B(n_5420),
.Y(n_7509)
);

A2O1A1Ixp33_ASAP7_75t_L g7510 ( 
.A1(n_6732),
.A2(n_5994),
.B(n_6012),
.C(n_5857),
.Y(n_7510)
);

BUFx8_ASAP7_75t_L g7511 ( 
.A(n_6051),
.Y(n_7511)
);

INVx2_ASAP7_75t_L g7512 ( 
.A(n_6462),
.Y(n_7512)
);

HB1xp67_ASAP7_75t_L g7513 ( 
.A(n_6612),
.Y(n_7513)
);

OA21x2_ASAP7_75t_L g7514 ( 
.A1(n_6274),
.A2(n_5268),
.B(n_5230),
.Y(n_7514)
);

INVx1_ASAP7_75t_L g7515 ( 
.A(n_6337),
.Y(n_7515)
);

NAND2xp5_ASAP7_75t_L g7516 ( 
.A(n_6417),
.B(n_5838),
.Y(n_7516)
);

OA21x2_ASAP7_75t_L g7517 ( 
.A1(n_6274),
.A2(n_5269),
.B(n_5430),
.Y(n_7517)
);

AO31x2_ASAP7_75t_L g7518 ( 
.A1(n_6560),
.A2(n_5269),
.A3(n_5501),
.B(n_5471),
.Y(n_7518)
);

AOI21xp5_ASAP7_75t_L g7519 ( 
.A1(n_6486),
.A2(n_5763),
.B(n_5540),
.Y(n_7519)
);

OAI21x1_ASAP7_75t_L g7520 ( 
.A1(n_6614),
.A2(n_5501),
.B(n_5471),
.Y(n_7520)
);

AND2x4_ASAP7_75t_L g7521 ( 
.A(n_6446),
.B(n_6553),
.Y(n_7521)
);

INVx1_ASAP7_75t_L g7522 ( 
.A(n_6337),
.Y(n_7522)
);

CKINVDCx20_ASAP7_75t_R g7523 ( 
.A(n_6767),
.Y(n_7523)
);

INVx1_ASAP7_75t_L g7524 ( 
.A(n_6350),
.Y(n_7524)
);

INVx2_ASAP7_75t_L g7525 ( 
.A(n_6462),
.Y(n_7525)
);

OAI21x1_ASAP7_75t_L g7526 ( 
.A1(n_6614),
.A2(n_5501),
.B(n_5471),
.Y(n_7526)
);

INVx1_ASAP7_75t_L g7527 ( 
.A(n_6350),
.Y(n_7527)
);

BUFx2_ASAP7_75t_L g7528 ( 
.A(n_6717),
.Y(n_7528)
);

OR2x2_ASAP7_75t_L g7529 ( 
.A(n_6336),
.B(n_5368),
.Y(n_7529)
);

A2O1A1Ixp33_ASAP7_75t_L g7530 ( 
.A1(n_6732),
.A2(n_5878),
.B(n_5875),
.C(n_5602),
.Y(n_7530)
);

NAND2xp5_ASAP7_75t_L g7531 ( 
.A(n_6591),
.B(n_5838),
.Y(n_7531)
);

OR2x2_ASAP7_75t_L g7532 ( 
.A(n_6357),
.B(n_5368),
.Y(n_7532)
);

OAI21x1_ASAP7_75t_L g7533 ( 
.A1(n_6614),
.A2(n_5585),
.B(n_5547),
.Y(n_7533)
);

AOI21x1_ASAP7_75t_L g7534 ( 
.A1(n_6392),
.A2(n_5585),
.B(n_5547),
.Y(n_7534)
);

OAI21x1_ASAP7_75t_L g7535 ( 
.A1(n_6408),
.A2(n_5585),
.B(n_5547),
.Y(n_7535)
);

OAI21x1_ASAP7_75t_L g7536 ( 
.A1(n_6581),
.A2(n_6283),
.B(n_6287),
.Y(n_7536)
);

BUFx6f_ASAP7_75t_L g7537 ( 
.A(n_6042),
.Y(n_7537)
);

INVx2_ASAP7_75t_L g7538 ( 
.A(n_6462),
.Y(n_7538)
);

CKINVDCx20_ASAP7_75t_R g7539 ( 
.A(n_6767),
.Y(n_7539)
);

INVx2_ASAP7_75t_SL g7540 ( 
.A(n_6803),
.Y(n_7540)
);

AOI21xp5_ASAP7_75t_L g7541 ( 
.A1(n_6755),
.A2(n_5763),
.B(n_5540),
.Y(n_7541)
);

INVx2_ASAP7_75t_SL g7542 ( 
.A(n_6803),
.Y(n_7542)
);

OR2x6_ASAP7_75t_L g7543 ( 
.A(n_6790),
.B(n_5291),
.Y(n_7543)
);

AOI21xp5_ASAP7_75t_L g7544 ( 
.A1(n_6755),
.A2(n_5763),
.B(n_5540),
.Y(n_7544)
);

BUFx2_ASAP7_75t_L g7545 ( 
.A(n_6717),
.Y(n_7545)
);

INVx6_ASAP7_75t_L g7546 ( 
.A(n_6039),
.Y(n_7546)
);

INVx1_ASAP7_75t_L g7547 ( 
.A(n_6350),
.Y(n_7547)
);

INVx2_ASAP7_75t_L g7548 ( 
.A(n_6462),
.Y(n_7548)
);

OR2x2_ASAP7_75t_L g7549 ( 
.A(n_6357),
.B(n_5368),
.Y(n_7549)
);

NAND2xp5_ASAP7_75t_L g7550 ( 
.A(n_6591),
.B(n_5368),
.Y(n_7550)
);

NAND2xp5_ASAP7_75t_L g7551 ( 
.A(n_6351),
.B(n_5368),
.Y(n_7551)
);

AOI21xp5_ASAP7_75t_L g7552 ( 
.A1(n_6721),
.A2(n_5323),
.B(n_5291),
.Y(n_7552)
);

NAND3xp33_ASAP7_75t_L g7553 ( 
.A(n_6521),
.B(n_5502),
.C(n_5744),
.Y(n_7553)
);

NAND2xp5_ASAP7_75t_L g7554 ( 
.A(n_6351),
.B(n_5368),
.Y(n_7554)
);

INVx1_ASAP7_75t_L g7555 ( 
.A(n_6362),
.Y(n_7555)
);

BUFx3_ASAP7_75t_L g7556 ( 
.A(n_6071),
.Y(n_7556)
);

NAND2xp5_ASAP7_75t_L g7557 ( 
.A(n_6358),
.B(n_5396),
.Y(n_7557)
);

AOI22xp33_ASAP7_75t_SL g7558 ( 
.A1(n_6112),
.A2(n_5741),
.B1(n_5923),
.B2(n_5545),
.Y(n_7558)
);

OAI21x1_ASAP7_75t_L g7559 ( 
.A1(n_6581),
.A2(n_5634),
.B(n_5615),
.Y(n_7559)
);

NAND2xp5_ASAP7_75t_L g7560 ( 
.A(n_6358),
.B(n_5396),
.Y(n_7560)
);

OAI21x1_ASAP7_75t_L g7561 ( 
.A1(n_6581),
.A2(n_5634),
.B(n_5615),
.Y(n_7561)
);

OA21x2_ASAP7_75t_L g7562 ( 
.A1(n_6274),
.A2(n_5634),
.B(n_5615),
.Y(n_7562)
);

AND2x4_ASAP7_75t_L g7563 ( 
.A(n_6446),
.B(n_5928),
.Y(n_7563)
);

AOI21x1_ASAP7_75t_L g7564 ( 
.A1(n_6416),
.A2(n_5703),
.B(n_5679),
.Y(n_7564)
);

AND2x2_ASAP7_75t_L g7565 ( 
.A(n_6378),
.B(n_5191),
.Y(n_7565)
);

AOI21x1_ASAP7_75t_L g7566 ( 
.A1(n_6416),
.A2(n_5703),
.B(n_5679),
.Y(n_7566)
);

AO31x2_ASAP7_75t_L g7567 ( 
.A1(n_6449),
.A2(n_5679),
.A3(n_5748),
.B(n_5703),
.Y(n_7567)
);

OR2x2_ASAP7_75t_L g7568 ( 
.A(n_6243),
.B(n_5396),
.Y(n_7568)
);

NAND2x1p5_ASAP7_75t_L g7569 ( 
.A(n_6076),
.B(n_5545),
.Y(n_7569)
);

NAND3xp33_ASAP7_75t_L g7570 ( 
.A(n_6231),
.B(n_5502),
.C(n_5744),
.Y(n_7570)
);

AO31x2_ASAP7_75t_L g7571 ( 
.A1(n_6691),
.A2(n_5748),
.A3(n_5831),
.B(n_5786),
.Y(n_7571)
);

AND2x4_ASAP7_75t_L g7572 ( 
.A(n_6446),
.B(n_5191),
.Y(n_7572)
);

A2O1A1Ixp33_ASAP7_75t_L g7573 ( 
.A1(n_6463),
.A2(n_5602),
.B(n_5499),
.C(n_6003),
.Y(n_7573)
);

AOI21xp5_ASAP7_75t_L g7574 ( 
.A1(n_6721),
.A2(n_5923),
.B(n_5545),
.Y(n_7574)
);

CKINVDCx5p33_ASAP7_75t_R g7575 ( 
.A(n_6335),
.Y(n_7575)
);

NAND2x1p5_ASAP7_75t_L g7576 ( 
.A(n_6076),
.B(n_5923),
.Y(n_7576)
);

AOI21x1_ASAP7_75t_L g7577 ( 
.A1(n_6691),
.A2(n_5786),
.B(n_5748),
.Y(n_7577)
);

INVx1_ASAP7_75t_L g7578 ( 
.A(n_6362),
.Y(n_7578)
);

OR2x2_ASAP7_75t_L g7579 ( 
.A(n_6243),
.B(n_5396),
.Y(n_7579)
);

INVx1_ASAP7_75t_L g7580 ( 
.A(n_6362),
.Y(n_7580)
);

NOR2x1_ASAP7_75t_SL g7581 ( 
.A(n_6340),
.B(n_5579),
.Y(n_7581)
);

OA21x2_ASAP7_75t_L g7582 ( 
.A1(n_6283),
.A2(n_5831),
.B(n_5786),
.Y(n_7582)
);

AND2x2_ASAP7_75t_L g7583 ( 
.A(n_6378),
.B(n_5191),
.Y(n_7583)
);

NAND2x1p5_ASAP7_75t_L g7584 ( 
.A(n_6076),
.B(n_5923),
.Y(n_7584)
);

NAND2xp5_ASAP7_75t_L g7585 ( 
.A(n_6799),
.B(n_5396),
.Y(n_7585)
);

INVx2_ASAP7_75t_L g7586 ( 
.A(n_6479),
.Y(n_7586)
);

OAI21x1_ASAP7_75t_L g7587 ( 
.A1(n_6283),
.A2(n_5852),
.B(n_5831),
.Y(n_7587)
);

INVx2_ASAP7_75t_L g7588 ( 
.A(n_6479),
.Y(n_7588)
);

INVx1_ASAP7_75t_L g7589 ( 
.A(n_6364),
.Y(n_7589)
);

INVx2_ASAP7_75t_L g7590 ( 
.A(n_6479),
.Y(n_7590)
);

NAND2x1p5_ASAP7_75t_L g7591 ( 
.A(n_6076),
.B(n_4675),
.Y(n_7591)
);

INVx2_ASAP7_75t_L g7592 ( 
.A(n_6415),
.Y(n_7592)
);

AOI21x1_ASAP7_75t_L g7593 ( 
.A1(n_6716),
.A2(n_5898),
.B(n_5852),
.Y(n_7593)
);

AND2x4_ASAP7_75t_L g7594 ( 
.A(n_6446),
.B(n_5191),
.Y(n_7594)
);

INVx1_ASAP7_75t_L g7595 ( 
.A(n_6364),
.Y(n_7595)
);

INVx2_ASAP7_75t_L g7596 ( 
.A(n_6415),
.Y(n_7596)
);

AOI22x1_ASAP7_75t_L g7597 ( 
.A1(n_6112),
.A2(n_5606),
.B1(n_5617),
.B2(n_5499),
.Y(n_7597)
);

INVx1_ASAP7_75t_L g7598 ( 
.A(n_6364),
.Y(n_7598)
);

HB1xp67_ASAP7_75t_L g7599 ( 
.A(n_6612),
.Y(n_7599)
);

INVx1_ASAP7_75t_L g7600 ( 
.A(n_6366),
.Y(n_7600)
);

OR2x2_ASAP7_75t_L g7601 ( 
.A(n_6395),
.B(n_6254),
.Y(n_7601)
);

INVx2_ASAP7_75t_L g7602 ( 
.A(n_6415),
.Y(n_7602)
);

AOI21xp5_ASAP7_75t_L g7603 ( 
.A1(n_6726),
.A2(n_5873),
.B(n_5871),
.Y(n_7603)
);

AOI22xp33_ASAP7_75t_SL g7604 ( 
.A1(n_6112),
.A2(n_5741),
.B1(n_5308),
.B2(n_5366),
.Y(n_7604)
);

NAND2xp5_ASAP7_75t_L g7605 ( 
.A(n_6799),
.B(n_6756),
.Y(n_7605)
);

OA21x2_ASAP7_75t_L g7606 ( 
.A1(n_6287),
.A2(n_5898),
.B(n_5852),
.Y(n_7606)
);

BUFx6f_ASAP7_75t_L g7607 ( 
.A(n_6076),
.Y(n_7607)
);

INVx4_ASAP7_75t_L g7608 ( 
.A(n_6079),
.Y(n_7608)
);

OAI21x1_ASAP7_75t_L g7609 ( 
.A1(n_6287),
.A2(n_5920),
.B(n_5898),
.Y(n_7609)
);

NAND2xp5_ASAP7_75t_L g7610 ( 
.A(n_6756),
.B(n_5396),
.Y(n_7610)
);

AND2x4_ASAP7_75t_L g7611 ( 
.A(n_6446),
.B(n_5308),
.Y(n_7611)
);

AOI21xp5_ASAP7_75t_L g7612 ( 
.A1(n_6726),
.A2(n_5888),
.B(n_5873),
.Y(n_7612)
);

AOI21x1_ASAP7_75t_L g7613 ( 
.A1(n_6716),
.A2(n_5925),
.B(n_5920),
.Y(n_7613)
);

AND2x4_ASAP7_75t_L g7614 ( 
.A(n_6446),
.B(n_5308),
.Y(n_7614)
);

OAI21xp33_ASAP7_75t_SL g7615 ( 
.A1(n_6345),
.A2(n_5452),
.B(n_5691),
.Y(n_7615)
);

OAI21x1_ASAP7_75t_L g7616 ( 
.A1(n_6124),
.A2(n_5925),
.B(n_5920),
.Y(n_7616)
);

AND2x2_ASAP7_75t_L g7617 ( 
.A(n_6407),
.B(n_5308),
.Y(n_7617)
);

AO31x2_ASAP7_75t_L g7618 ( 
.A1(n_6716),
.A2(n_5948),
.A3(n_6001),
.B(n_5925),
.Y(n_7618)
);

AO21x2_ASAP7_75t_L g7619 ( 
.A1(n_6514),
.A2(n_5888),
.B(n_5948),
.Y(n_7619)
);

NAND2xp5_ASAP7_75t_L g7620 ( 
.A(n_6254),
.B(n_5182),
.Y(n_7620)
);

INVx2_ASAP7_75t_L g7621 ( 
.A(n_6479),
.Y(n_7621)
);

AND2x4_ASAP7_75t_L g7622 ( 
.A(n_6553),
.B(n_5313),
.Y(n_7622)
);

INVx2_ASAP7_75t_L g7623 ( 
.A(n_6489),
.Y(n_7623)
);

AOI22xp33_ASAP7_75t_L g7624 ( 
.A1(n_6112),
.A2(n_5090),
.B1(n_5366),
.B2(n_5313),
.Y(n_7624)
);

OAI22xp5_ASAP7_75t_L g7625 ( 
.A1(n_6540),
.A2(n_5741),
.B1(n_6003),
.B2(n_5617),
.Y(n_7625)
);

OAI21xp5_ASAP7_75t_L g7626 ( 
.A1(n_6694),
.A2(n_5692),
.B(n_5687),
.Y(n_7626)
);

AND2x4_ASAP7_75t_L g7627 ( 
.A(n_6553),
.B(n_5313),
.Y(n_7627)
);

AOI21x1_ASAP7_75t_L g7628 ( 
.A1(n_6498),
.A2(n_6001),
.B(n_5948),
.Y(n_7628)
);

INVx1_ASAP7_75t_L g7629 ( 
.A(n_6366),
.Y(n_7629)
);

AOI22xp33_ASAP7_75t_L g7630 ( 
.A1(n_7032),
.A2(n_6432),
.B1(n_6142),
.B2(n_6403),
.Y(n_7630)
);

OAI22xp5_ASAP7_75t_L g7631 ( 
.A1(n_7008),
.A2(n_6053),
.B1(n_6288),
.B2(n_6398),
.Y(n_7631)
);

NAND2xp5_ASAP7_75t_L g7632 ( 
.A(n_7113),
.B(n_6306),
.Y(n_7632)
);

OAI22x1_ASAP7_75t_SL g7633 ( 
.A1(n_6848),
.A2(n_6140),
.B1(n_6359),
.B2(n_6697),
.Y(n_7633)
);

AOI22xp5_ASAP7_75t_L g7634 ( 
.A1(n_6885),
.A2(n_6255),
.B1(n_6481),
.B2(n_6306),
.Y(n_7634)
);

OAI22xp33_ASAP7_75t_L g7635 ( 
.A1(n_7437),
.A2(n_6285),
.B1(n_6176),
.B2(n_6049),
.Y(n_7635)
);

AND2x2_ASAP7_75t_L g7636 ( 
.A(n_6924),
.B(n_6555),
.Y(n_7636)
);

BUFx2_ASAP7_75t_L g7637 ( 
.A(n_7497),
.Y(n_7637)
);

OAI22xp5_ASAP7_75t_L g7638 ( 
.A1(n_7152),
.A2(n_6403),
.B1(n_6424),
.B2(n_6190),
.Y(n_7638)
);

AOI22xp33_ASAP7_75t_SL g7639 ( 
.A1(n_7051),
.A2(n_7093),
.B1(n_7049),
.B2(n_6851),
.Y(n_7639)
);

BUFx8_ASAP7_75t_L g7640 ( 
.A(n_6890),
.Y(n_7640)
);

AND2x2_ASAP7_75t_L g7641 ( 
.A(n_6924),
.B(n_6555),
.Y(n_7641)
);

AOI22xp33_ASAP7_75t_L g7642 ( 
.A1(n_7068),
.A2(n_6432),
.B1(n_6142),
.B2(n_6167),
.Y(n_7642)
);

CKINVDCx20_ASAP7_75t_R g7643 ( 
.A(n_7125),
.Y(n_7643)
);

HB1xp67_ASAP7_75t_L g7644 ( 
.A(n_6812),
.Y(n_7644)
);

AOI22xp33_ASAP7_75t_SL g7645 ( 
.A1(n_7305),
.A2(n_6167),
.B1(n_6432),
.B2(n_6467),
.Y(n_7645)
);

AOI22xp33_ASAP7_75t_L g7646 ( 
.A1(n_7045),
.A2(n_6167),
.B1(n_6255),
.B2(n_6704),
.Y(n_7646)
);

INVx3_ASAP7_75t_L g7647 ( 
.A(n_6881),
.Y(n_7647)
);

AOI22xp33_ASAP7_75t_L g7648 ( 
.A1(n_7048),
.A2(n_6704),
.B1(n_6348),
.B2(n_6481),
.Y(n_7648)
);

INVx4_ASAP7_75t_L g7649 ( 
.A(n_6890),
.Y(n_7649)
);

AOI222xp33_ASAP7_75t_L g7650 ( 
.A1(n_7052),
.A2(n_6090),
.B1(n_6084),
.B2(n_6525),
.C1(n_6231),
.C2(n_6491),
.Y(n_7650)
);

OAI222xp33_ASAP7_75t_L g7651 ( 
.A1(n_7437),
.A2(n_6727),
.B1(n_6713),
.B2(n_6348),
.C1(n_6781),
.C2(n_6695),
.Y(n_7651)
);

OAI22xp5_ASAP7_75t_L g7652 ( 
.A1(n_6984),
.A2(n_6424),
.B1(n_6190),
.B2(n_6206),
.Y(n_7652)
);

NOR2xp33_ASAP7_75t_L g7653 ( 
.A(n_6984),
.B(n_6359),
.Y(n_7653)
);

OAI22xp5_ASAP7_75t_L g7654 ( 
.A1(n_7078),
.A2(n_6206),
.B1(n_6078),
.B2(n_6758),
.Y(n_7654)
);

AOI22xp33_ASAP7_75t_L g7655 ( 
.A1(n_7040),
.A2(n_6514),
.B1(n_6634),
.B2(n_6467),
.Y(n_7655)
);

OAI21xp5_ASAP7_75t_SL g7656 ( 
.A1(n_6810),
.A2(n_6750),
.B(n_6078),
.Y(n_7656)
);

OR2x6_ASAP7_75t_L g7657 ( 
.A(n_7415),
.B(n_6079),
.Y(n_7657)
);

AOI22xp33_ASAP7_75t_L g7658 ( 
.A1(n_7114),
.A2(n_7150),
.B1(n_7249),
.B2(n_7192),
.Y(n_7658)
);

INVx1_ASAP7_75t_L g7659 ( 
.A(n_6809),
.Y(n_7659)
);

AOI22xp33_ASAP7_75t_L g7660 ( 
.A1(n_6808),
.A2(n_6514),
.B1(n_6634),
.B2(n_6467),
.Y(n_7660)
);

INVxp67_ASAP7_75t_L g7661 ( 
.A(n_7154),
.Y(n_7661)
);

INVx2_ASAP7_75t_L g7662 ( 
.A(n_7372),
.Y(n_7662)
);

OAI22xp5_ASAP7_75t_L g7663 ( 
.A1(n_6896),
.A2(n_6758),
.B1(n_6781),
.B2(n_6159),
.Y(n_7663)
);

INVx2_ASAP7_75t_L g7664 ( 
.A(n_7372),
.Y(n_7664)
);

AOI22xp33_ASAP7_75t_L g7665 ( 
.A1(n_7465),
.A2(n_6940),
.B1(n_7477),
.B2(n_7388),
.Y(n_7665)
);

AOI22xp33_ASAP7_75t_L g7666 ( 
.A1(n_6907),
.A2(n_6514),
.B1(n_6296),
.B2(n_6090),
.Y(n_7666)
);

AOI22xp33_ASAP7_75t_SL g7667 ( 
.A1(n_6807),
.A2(n_6387),
.B1(n_6399),
.B2(n_6380),
.Y(n_7667)
);

AOI22xp33_ASAP7_75t_SL g7668 ( 
.A1(n_7072),
.A2(n_6387),
.B1(n_6399),
.B2(n_6380),
.Y(n_7668)
);

AOI22xp33_ASAP7_75t_L g7669 ( 
.A1(n_6904),
.A2(n_6296),
.B1(n_6084),
.B2(n_6159),
.Y(n_7669)
);

BUFx12f_ASAP7_75t_L g7670 ( 
.A(n_7154),
.Y(n_7670)
);

CKINVDCx5p33_ASAP7_75t_R g7671 ( 
.A(n_6869),
.Y(n_7671)
);

OAI22xp5_ASAP7_75t_L g7672 ( 
.A1(n_6844),
.A2(n_6375),
.B1(n_6454),
.B2(n_6404),
.Y(n_7672)
);

INVx2_ASAP7_75t_SL g7673 ( 
.A(n_7238),
.Y(n_7673)
);

CKINVDCx5p33_ASAP7_75t_R g7674 ( 
.A(n_6956),
.Y(n_7674)
);

BUFx12f_ASAP7_75t_L g7675 ( 
.A(n_7154),
.Y(n_7675)
);

AOI22xp33_ASAP7_75t_L g7676 ( 
.A1(n_7348),
.A2(n_6296),
.B1(n_6803),
.B2(n_6699),
.Y(n_7676)
);

INVx1_ASAP7_75t_SL g7677 ( 
.A(n_7119),
.Y(n_7677)
);

INVx4_ASAP7_75t_L g7678 ( 
.A(n_6890),
.Y(n_7678)
);

NOR2xp33_ASAP7_75t_L g7679 ( 
.A(n_6939),
.B(n_6751),
.Y(n_7679)
);

INVx1_ASAP7_75t_L g7680 ( 
.A(n_6809),
.Y(n_7680)
);

AND2x2_ASAP7_75t_L g7681 ( 
.A(n_6934),
.B(n_6555),
.Y(n_7681)
);

NOR2x1_ASAP7_75t_R g7682 ( 
.A(n_6886),
.B(n_6033),
.Y(n_7682)
);

AND2x2_ASAP7_75t_L g7683 ( 
.A(n_6934),
.B(n_6542),
.Y(n_7683)
);

OAI21xp5_ASAP7_75t_SL g7684 ( 
.A1(n_6929),
.A2(n_6750),
.B(n_6727),
.Y(n_7684)
);

OAI22xp5_ASAP7_75t_L g7685 ( 
.A1(n_7456),
.A2(n_6375),
.B1(n_6454),
.B2(n_6404),
.Y(n_7685)
);

AOI22xp33_ASAP7_75t_SL g7686 ( 
.A1(n_7072),
.A2(n_6387),
.B1(n_6399),
.B2(n_6380),
.Y(n_7686)
);

AOI22xp33_ASAP7_75t_L g7687 ( 
.A1(n_7141),
.A2(n_6296),
.B1(n_6803),
.B2(n_6699),
.Y(n_7687)
);

OAI22xp5_ASAP7_75t_L g7688 ( 
.A1(n_7456),
.A2(n_6420),
.B1(n_6713),
.B2(n_6611),
.Y(n_7688)
);

AOI22xp33_ASAP7_75t_L g7689 ( 
.A1(n_7605),
.A2(n_6296),
.B1(n_6698),
.B2(n_6488),
.Y(n_7689)
);

INVx6_ASAP7_75t_L g7690 ( 
.A(n_7126),
.Y(n_7690)
);

AOI22xp33_ASAP7_75t_L g7691 ( 
.A1(n_7111),
.A2(n_6698),
.B1(n_6488),
.B2(n_6340),
.Y(n_7691)
);

INVx1_ASAP7_75t_L g7692 ( 
.A(n_6813),
.Y(n_7692)
);

OAI22xp5_ASAP7_75t_L g7693 ( 
.A1(n_6937),
.A2(n_6420),
.B1(n_6611),
.B2(n_6793),
.Y(n_7693)
);

OAI21xp5_ASAP7_75t_SL g7694 ( 
.A1(n_6930),
.A2(n_6456),
.B(n_6483),
.Y(n_7694)
);

AOI21xp5_ASAP7_75t_L g7695 ( 
.A1(n_7417),
.A2(n_6620),
.B(n_6491),
.Y(n_7695)
);

AOI22xp33_ASAP7_75t_L g7696 ( 
.A1(n_6911),
.A2(n_6488),
.B1(n_6340),
.B2(n_6551),
.Y(n_7696)
);

OAI22xp5_ASAP7_75t_L g7697 ( 
.A1(n_7353),
.A2(n_6793),
.B1(n_6800),
.B2(n_6695),
.Y(n_7697)
);

INVx1_ASAP7_75t_L g7698 ( 
.A(n_6813),
.Y(n_7698)
);

OAI22xp5_ASAP7_75t_L g7699 ( 
.A1(n_7353),
.A2(n_6800),
.B1(n_6071),
.B2(n_6136),
.Y(n_7699)
);

AOI22xp33_ASAP7_75t_SL g7700 ( 
.A1(n_7002),
.A2(n_6354),
.B1(n_6345),
.B2(n_6518),
.Y(n_7700)
);

AND2x2_ASAP7_75t_L g7701 ( 
.A(n_7013),
.B(n_6542),
.Y(n_7701)
);

OAI22xp33_ASAP7_75t_L g7702 ( 
.A1(n_6943),
.A2(n_6285),
.B1(n_6049),
.B2(n_6176),
.Y(n_7702)
);

BUFx4f_ASAP7_75t_SL g7703 ( 
.A(n_6886),
.Y(n_7703)
);

OAI22xp33_ASAP7_75t_L g7704 ( 
.A1(n_6943),
.A2(n_7074),
.B1(n_7024),
.B2(n_7033),
.Y(n_7704)
);

AOI22xp33_ASAP7_75t_SL g7705 ( 
.A1(n_7411),
.A2(n_6354),
.B1(n_6345),
.B2(n_6518),
.Y(n_7705)
);

OAI21xp5_ASAP7_75t_SL g7706 ( 
.A1(n_7024),
.A2(n_6456),
.B(n_6483),
.Y(n_7706)
);

INVx1_ASAP7_75t_L g7707 ( 
.A(n_6827),
.Y(n_7707)
);

CKINVDCx5p33_ASAP7_75t_R g7708 ( 
.A(n_7154),
.Y(n_7708)
);

HB1xp67_ASAP7_75t_L g7709 ( 
.A(n_6819),
.Y(n_7709)
);

AOI22xp33_ASAP7_75t_L g7710 ( 
.A1(n_7061),
.A2(n_6488),
.B1(n_6340),
.B2(n_6551),
.Y(n_7710)
);

CKINVDCx5p33_ASAP7_75t_R g7711 ( 
.A(n_7204),
.Y(n_7711)
);

INVx1_ASAP7_75t_L g7712 ( 
.A(n_6827),
.Y(n_7712)
);

AND2x2_ASAP7_75t_L g7713 ( 
.A(n_7013),
.B(n_6542),
.Y(n_7713)
);

AOI22xp5_ASAP7_75t_L g7714 ( 
.A1(n_7061),
.A2(n_6556),
.B1(n_6620),
.B2(n_6550),
.Y(n_7714)
);

AOI22xp33_ASAP7_75t_L g7715 ( 
.A1(n_6855),
.A2(n_6488),
.B1(n_6340),
.B2(n_6551),
.Y(n_7715)
);

AOI22xp33_ASAP7_75t_L g7716 ( 
.A1(n_7453),
.A2(n_6488),
.B1(n_6340),
.B2(n_6558),
.Y(n_7716)
);

INVx2_ASAP7_75t_L g7717 ( 
.A(n_7372),
.Y(n_7717)
);

AOI22xp33_ASAP7_75t_L g7718 ( 
.A1(n_6991),
.A2(n_6488),
.B1(n_6585),
.B2(n_6558),
.Y(n_7718)
);

INVx1_ASAP7_75t_L g7719 ( 
.A(n_6831),
.Y(n_7719)
);

BUFx12f_ASAP7_75t_L g7720 ( 
.A(n_7204),
.Y(n_7720)
);

AOI22xp33_ASAP7_75t_L g7721 ( 
.A1(n_7429),
.A2(n_7461),
.B1(n_6972),
.B2(n_7332),
.Y(n_7721)
);

NOR2xp33_ASAP7_75t_L g7722 ( 
.A(n_6890),
.B(n_6751),
.Y(n_7722)
);

BUFx6f_ASAP7_75t_L g7723 ( 
.A(n_6890),
.Y(n_7723)
);

AOI22xp33_ASAP7_75t_L g7724 ( 
.A1(n_6944),
.A2(n_6585),
.B1(n_6558),
.B2(n_6103),
.Y(n_7724)
);

NAND3xp33_ASAP7_75t_L g7725 ( 
.A(n_7003),
.B(n_6518),
.C(n_6297),
.Y(n_7725)
);

OAI22xp5_ASAP7_75t_L g7726 ( 
.A1(n_6996),
.A2(n_6071),
.B1(n_6136),
.B2(n_6091),
.Y(n_7726)
);

CKINVDCx5p33_ASAP7_75t_R g7727 ( 
.A(n_7204),
.Y(n_7727)
);

AOI22xp33_ASAP7_75t_L g7728 ( 
.A1(n_6923),
.A2(n_6585),
.B1(n_6103),
.B2(n_6033),
.Y(n_7728)
);

NOR2xp67_ASAP7_75t_L g7729 ( 
.A(n_7238),
.B(n_6407),
.Y(n_7729)
);

AOI22xp5_ASAP7_75t_L g7730 ( 
.A1(n_6858),
.A2(n_6556),
.B1(n_6550),
.B2(n_6546),
.Y(n_7730)
);

OAI22xp33_ASAP7_75t_L g7731 ( 
.A1(n_7033),
.A2(n_6308),
.B1(n_6557),
.B2(n_6546),
.Y(n_7731)
);

OAI22xp33_ASAP7_75t_L g7732 ( 
.A1(n_7438),
.A2(n_6308),
.B1(n_6557),
.B2(n_6790),
.Y(n_7732)
);

OAI222xp33_ASAP7_75t_L g7733 ( 
.A1(n_7344),
.A2(n_6652),
.B1(n_6354),
.B2(n_6731),
.C1(n_6525),
.C2(n_6693),
.Y(n_7733)
);

BUFx12f_ASAP7_75t_L g7734 ( 
.A(n_7204),
.Y(n_7734)
);

CKINVDCx11_ASAP7_75t_R g7735 ( 
.A(n_6954),
.Y(n_7735)
);

OAI22xp5_ASAP7_75t_L g7736 ( 
.A1(n_6953),
.A2(n_6071),
.B1(n_6136),
.B2(n_6091),
.Y(n_7736)
);

OAI22xp5_ASAP7_75t_L g7737 ( 
.A1(n_7120),
.A2(n_6091),
.B1(n_6141),
.B2(n_6136),
.Y(n_7737)
);

INVx1_ASAP7_75t_L g7738 ( 
.A(n_6831),
.Y(n_7738)
);

INVx1_ASAP7_75t_L g7739 ( 
.A(n_6833),
.Y(n_7739)
);

INVx2_ASAP7_75t_L g7740 ( 
.A(n_7618),
.Y(n_7740)
);

INVx2_ASAP7_75t_L g7741 ( 
.A(n_7618),
.Y(n_7741)
);

INVx2_ASAP7_75t_SL g7742 ( 
.A(n_7238),
.Y(n_7742)
);

OAI22xp5_ASAP7_75t_L g7743 ( 
.A1(n_7445),
.A2(n_6091),
.B1(n_6227),
.B2(n_6141),
.Y(n_7743)
);

NAND2xp5_ASAP7_75t_L g7744 ( 
.A(n_6895),
.B(n_6898),
.Y(n_7744)
);

OAI22xp33_ASAP7_75t_L g7745 ( 
.A1(n_7438),
.A2(n_7516),
.B1(n_7499),
.B2(n_7085),
.Y(n_7745)
);

OAI21xp33_ASAP7_75t_L g7746 ( 
.A1(n_7414),
.A2(n_6510),
.B(n_6483),
.Y(n_7746)
);

INVx1_ASAP7_75t_L g7747 ( 
.A(n_6833),
.Y(n_7747)
);

NAND3xp33_ASAP7_75t_L g7748 ( 
.A(n_7473),
.B(n_6518),
.C(n_6297),
.Y(n_7748)
);

AOI22xp5_ASAP7_75t_L g7749 ( 
.A1(n_6858),
.A2(n_6790),
.B1(n_6523),
.B2(n_6510),
.Y(n_7749)
);

AOI222xp33_ASAP7_75t_L g7750 ( 
.A1(n_7502),
.A2(n_6523),
.B1(n_6510),
.B2(n_6744),
.C1(n_6664),
.C2(n_6253),
.Y(n_7750)
);

OAI222xp33_ASAP7_75t_L g7751 ( 
.A1(n_7378),
.A2(n_6652),
.B1(n_6731),
.B2(n_6693),
.C1(n_6293),
.C2(n_6087),
.Y(n_7751)
);

INVxp67_ASAP7_75t_L g7752 ( 
.A(n_7214),
.Y(n_7752)
);

AOI22xp33_ASAP7_75t_L g7753 ( 
.A1(n_6922),
.A2(n_6983),
.B1(n_6973),
.B2(n_7171),
.Y(n_7753)
);

INVx1_ASAP7_75t_L g7754 ( 
.A(n_6837),
.Y(n_7754)
);

BUFx3_ASAP7_75t_L g7755 ( 
.A(n_6954),
.Y(n_7755)
);

AOI22xp5_ASAP7_75t_L g7756 ( 
.A1(n_6873),
.A2(n_6790),
.B1(n_6523),
.B2(n_6253),
.Y(n_7756)
);

AOI222xp33_ASAP7_75t_L g7757 ( 
.A1(n_7610),
.A2(n_6664),
.B1(n_6744),
.B2(n_6325),
.C1(n_6395),
.C2(n_6657),
.Y(n_7757)
);

INVx3_ASAP7_75t_L g7758 ( 
.A(n_6881),
.Y(n_7758)
);

CKINVDCx6p67_ASAP7_75t_R g7759 ( 
.A(n_6977),
.Y(n_7759)
);

OAI22xp5_ASAP7_75t_L g7760 ( 
.A1(n_7410),
.A2(n_6227),
.B1(n_6232),
.B2(n_6141),
.Y(n_7760)
);

BUFx6f_ASAP7_75t_L g7761 ( 
.A(n_7409),
.Y(n_7761)
);

OAI22xp5_ASAP7_75t_L g7762 ( 
.A1(n_7383),
.A2(n_6227),
.B1(n_6232),
.B2(n_6141),
.Y(n_7762)
);

AOI22xp33_ASAP7_75t_L g7763 ( 
.A1(n_6973),
.A2(n_6103),
.B1(n_6033),
.B2(n_6058),
.Y(n_7763)
);

INVx2_ASAP7_75t_L g7764 ( 
.A(n_7571),
.Y(n_7764)
);

OAI21xp5_ASAP7_75t_L g7765 ( 
.A1(n_6816),
.A2(n_6694),
.B(n_6650),
.Y(n_7765)
);

INVxp67_ASAP7_75t_L g7766 ( 
.A(n_7214),
.Y(n_7766)
);

AOI222xp33_ASAP7_75t_L g7767 ( 
.A1(n_7585),
.A2(n_6325),
.B1(n_6657),
.B2(n_6602),
.C1(n_6498),
.C2(n_6566),
.Y(n_7767)
);

OAI22xp5_ASAP7_75t_SL g7768 ( 
.A1(n_6977),
.A2(n_7011),
.B1(n_7054),
.B2(n_6999),
.Y(n_7768)
);

INVx1_ASAP7_75t_L g7769 ( 
.A(n_6837),
.Y(n_7769)
);

INVx1_ASAP7_75t_L g7770 ( 
.A(n_6839),
.Y(n_7770)
);

AOI22xp5_ASAP7_75t_L g7771 ( 
.A1(n_6873),
.A2(n_6790),
.B1(n_6411),
.B2(n_6734),
.Y(n_7771)
);

INVx1_ASAP7_75t_SL g7772 ( 
.A(n_7157),
.Y(n_7772)
);

NOR2xp33_ASAP7_75t_L g7773 ( 
.A(n_7211),
.B(n_6033),
.Y(n_7773)
);

AOI22xp33_ASAP7_75t_L g7774 ( 
.A1(n_6973),
.A2(n_6103),
.B1(n_6058),
.B2(n_6437),
.Y(n_7774)
);

OAI21xp33_ASAP7_75t_L g7775 ( 
.A1(n_7425),
.A2(n_6731),
.B(n_6693),
.Y(n_7775)
);

INVx1_ASAP7_75t_SL g7776 ( 
.A(n_7157),
.Y(n_7776)
);

OAI22xp5_ASAP7_75t_L g7777 ( 
.A1(n_7261),
.A2(n_6227),
.B1(n_6240),
.B2(n_6232),
.Y(n_7777)
);

OAI22xp5_ASAP7_75t_L g7778 ( 
.A1(n_6832),
.A2(n_7510),
.B1(n_7337),
.B2(n_7530),
.Y(n_7778)
);

OR2x2_ASAP7_75t_L g7779 ( 
.A(n_7317),
.B(n_6582),
.Y(n_7779)
);

BUFx4f_ASAP7_75t_SL g7780 ( 
.A(n_7011),
.Y(n_7780)
);

AOI22xp33_ASAP7_75t_L g7781 ( 
.A1(n_6973),
.A2(n_6103),
.B1(n_6058),
.B2(n_6437),
.Y(n_7781)
);

BUFx3_ASAP7_75t_L g7782 ( 
.A(n_7054),
.Y(n_7782)
);

AOI22xp33_ASAP7_75t_L g7783 ( 
.A1(n_6973),
.A2(n_6653),
.B1(n_6437),
.B2(n_6518),
.Y(n_7783)
);

AOI22xp33_ASAP7_75t_SL g7784 ( 
.A1(n_7214),
.A2(n_7007),
.B1(n_7273),
.B2(n_6870),
.Y(n_7784)
);

CKINVDCx20_ASAP7_75t_R g7785 ( 
.A(n_7148),
.Y(n_7785)
);

INVx1_ASAP7_75t_L g7786 ( 
.A(n_6839),
.Y(n_7786)
);

INVx1_ASAP7_75t_L g7787 ( 
.A(n_6854),
.Y(n_7787)
);

OAI22xp5_ASAP7_75t_L g7788 ( 
.A1(n_7337),
.A2(n_6240),
.B1(n_6268),
.B2(n_6232),
.Y(n_7788)
);

INVx5_ASAP7_75t_L g7789 ( 
.A(n_7433),
.Y(n_7789)
);

AND2x2_ASAP7_75t_L g7790 ( 
.A(n_7070),
.B(n_6407),
.Y(n_7790)
);

INVx1_ASAP7_75t_L g7791 ( 
.A(n_6854),
.Y(n_7791)
);

AOI22xp33_ASAP7_75t_L g7792 ( 
.A1(n_7163),
.A2(n_6653),
.B1(n_6437),
.B2(n_6518),
.Y(n_7792)
);

AOI22xp33_ASAP7_75t_L g7793 ( 
.A1(n_7476),
.A2(n_6653),
.B1(n_6437),
.B2(n_6339),
.Y(n_7793)
);

BUFx6f_ASAP7_75t_L g7794 ( 
.A(n_7409),
.Y(n_7794)
);

INVx1_ASAP7_75t_L g7795 ( 
.A(n_6856),
.Y(n_7795)
);

AOI22xp33_ASAP7_75t_L g7796 ( 
.A1(n_7476),
.A2(n_6653),
.B1(n_6339),
.B2(n_6319),
.Y(n_7796)
);

OAI21xp33_ASAP7_75t_L g7797 ( 
.A1(n_6877),
.A2(n_6473),
.B(n_6393),
.Y(n_7797)
);

OAI21xp33_ASAP7_75t_L g7798 ( 
.A1(n_6877),
.A2(n_6473),
.B(n_6393),
.Y(n_7798)
);

INVx2_ASAP7_75t_L g7799 ( 
.A(n_7571),
.Y(n_7799)
);

AOI22xp33_ASAP7_75t_L g7800 ( 
.A1(n_7050),
.A2(n_6653),
.B1(n_6339),
.B2(n_6319),
.Y(n_7800)
);

AOI222xp33_ASAP7_75t_L g7801 ( 
.A1(n_7349),
.A2(n_6602),
.B1(n_6498),
.B2(n_6548),
.C1(n_6566),
.C2(n_6597),
.Y(n_7801)
);

AOI22xp33_ASAP7_75t_L g7802 ( 
.A1(n_7050),
.A2(n_6319),
.B1(n_6431),
.B2(n_6790),
.Y(n_7802)
);

INVx2_ASAP7_75t_L g7803 ( 
.A(n_7571),
.Y(n_7803)
);

INVx1_ASAP7_75t_L g7804 ( 
.A(n_6856),
.Y(n_7804)
);

OAI22xp5_ASAP7_75t_L g7805 ( 
.A1(n_7553),
.A2(n_6268),
.B1(n_6341),
.B2(n_6240),
.Y(n_7805)
);

AOI222xp33_ASAP7_75t_L g7806 ( 
.A1(n_7355),
.A2(n_6548),
.B1(n_6595),
.B2(n_6597),
.C1(n_6445),
.C2(n_6760),
.Y(n_7806)
);

AOI22xp33_ASAP7_75t_L g7807 ( 
.A1(n_7050),
.A2(n_6319),
.B1(n_6431),
.B2(n_6790),
.Y(n_7807)
);

INVx1_ASAP7_75t_SL g7808 ( 
.A(n_7157),
.Y(n_7808)
);

INVx2_ASAP7_75t_L g7809 ( 
.A(n_7571),
.Y(n_7809)
);

OAI22xp33_ASAP7_75t_L g7810 ( 
.A1(n_6965),
.A2(n_7167),
.B1(n_7325),
.B2(n_7314),
.Y(n_7810)
);

OAI22xp33_ASAP7_75t_SL g7811 ( 
.A1(n_6823),
.A2(n_6087),
.B1(n_6250),
.B2(n_6178),
.Y(n_7811)
);

AOI22xp33_ASAP7_75t_L g7812 ( 
.A1(n_7050),
.A2(n_6319),
.B1(n_6431),
.B2(n_6494),
.Y(n_7812)
);

OR2x2_ASAP7_75t_L g7813 ( 
.A(n_7317),
.B(n_6582),
.Y(n_7813)
);

INVx1_ASAP7_75t_L g7814 ( 
.A(n_6863),
.Y(n_7814)
);

BUFx6f_ASAP7_75t_SL g7815 ( 
.A(n_7409),
.Y(n_7815)
);

INVx4_ASAP7_75t_SL g7816 ( 
.A(n_6949),
.Y(n_7816)
);

AOI22xp33_ASAP7_75t_L g7817 ( 
.A1(n_7050),
.A2(n_6319),
.B1(n_6494),
.B2(n_6613),
.Y(n_7817)
);

HB1xp67_ASAP7_75t_L g7818 ( 
.A(n_6883),
.Y(n_7818)
);

AOI222xp33_ASAP7_75t_L g7819 ( 
.A1(n_7086),
.A2(n_6597),
.B1(n_6595),
.B2(n_6445),
.C1(n_6791),
.C2(n_6760),
.Y(n_7819)
);

NOR2xp67_ASAP7_75t_SL g7820 ( 
.A(n_7037),
.B(n_6240),
.Y(n_7820)
);

BUFx12f_ASAP7_75t_L g7821 ( 
.A(n_7214),
.Y(n_7821)
);

AOI22xp33_ASAP7_75t_L g7822 ( 
.A1(n_6840),
.A2(n_6319),
.B1(n_6494),
.B2(n_6613),
.Y(n_7822)
);

BUFx3_ASAP7_75t_L g7823 ( 
.A(n_7126),
.Y(n_7823)
);

AOI22xp33_ASAP7_75t_L g7824 ( 
.A1(n_6840),
.A2(n_6613),
.B1(n_6775),
.B2(n_6268),
.Y(n_7824)
);

BUFx4f_ASAP7_75t_SL g7825 ( 
.A(n_7302),
.Y(n_7825)
);

CKINVDCx5p33_ASAP7_75t_R g7826 ( 
.A(n_6999),
.Y(n_7826)
);

OAI22xp5_ASAP7_75t_SL g7827 ( 
.A1(n_6848),
.A2(n_6268),
.B1(n_6394),
.B2(n_6341),
.Y(n_7827)
);

INVx1_ASAP7_75t_L g7828 ( 
.A(n_6863),
.Y(n_7828)
);

HB1xp67_ASAP7_75t_L g7829 ( 
.A(n_6918),
.Y(n_7829)
);

AOI22xp33_ASAP7_75t_L g7830 ( 
.A1(n_6840),
.A2(n_6775),
.B1(n_6341),
.B2(n_6422),
.Y(n_7830)
);

AOI22xp33_ASAP7_75t_L g7831 ( 
.A1(n_6840),
.A2(n_6775),
.B1(n_6341),
.B2(n_6422),
.Y(n_7831)
);

BUFx12f_ASAP7_75t_L g7832 ( 
.A(n_7126),
.Y(n_7832)
);

OAI22xp33_ASAP7_75t_L g7833 ( 
.A1(n_7333),
.A2(n_6422),
.B1(n_6472),
.B2(n_6394),
.Y(n_7833)
);

NAND3xp33_ASAP7_75t_L g7834 ( 
.A(n_6870),
.B(n_6289),
.C(n_6110),
.Y(n_7834)
);

OAI22xp5_ASAP7_75t_SL g7835 ( 
.A1(n_6882),
.A2(n_6394),
.B1(n_6472),
.B2(n_6422),
.Y(n_7835)
);

BUFx3_ASAP7_75t_L g7836 ( 
.A(n_7126),
.Y(n_7836)
);

AOI22xp33_ASAP7_75t_L g7837 ( 
.A1(n_6945),
.A2(n_6394),
.B1(n_6541),
.B2(n_6472),
.Y(n_7837)
);

OAI22xp5_ASAP7_75t_L g7838 ( 
.A1(n_7553),
.A2(n_6541),
.B1(n_6600),
.B2(n_6472),
.Y(n_7838)
);

AOI22xp33_ASAP7_75t_L g7839 ( 
.A1(n_6945),
.A2(n_6541),
.B1(n_6671),
.B2(n_6600),
.Y(n_7839)
);

OAI22xp33_ASAP7_75t_L g7840 ( 
.A1(n_7094),
.A2(n_6600),
.B1(n_6671),
.B2(n_6541),
.Y(n_7840)
);

INVx1_ASAP7_75t_L g7841 ( 
.A(n_6867),
.Y(n_7841)
);

AOI22xp33_ASAP7_75t_SL g7842 ( 
.A1(n_7007),
.A2(n_6661),
.B1(n_6728),
.B2(n_6544),
.Y(n_7842)
);

AOI22xp33_ASAP7_75t_SL g7843 ( 
.A1(n_7273),
.A2(n_6661),
.B1(n_6728),
.B2(n_6544),
.Y(n_7843)
);

AOI22xp33_ASAP7_75t_L g7844 ( 
.A1(n_6945),
.A2(n_6600),
.B1(n_6671),
.B2(n_6079),
.Y(n_7844)
);

OAI21xp5_ASAP7_75t_SL g7845 ( 
.A1(n_6862),
.A2(n_6682),
.B(n_6536),
.Y(n_7845)
);

OAI21xp5_ASAP7_75t_SL g7846 ( 
.A1(n_6862),
.A2(n_6682),
.B(n_6536),
.Y(n_7846)
);

NOR2xp33_ASAP7_75t_SL g7847 ( 
.A(n_7497),
.B(n_7241),
.Y(n_7847)
);

AOI22xp33_ASAP7_75t_L g7848 ( 
.A1(n_6945),
.A2(n_6671),
.B1(n_6079),
.B2(n_6534),
.Y(n_7848)
);

AOI22xp33_ASAP7_75t_L g7849 ( 
.A1(n_7304),
.A2(n_6079),
.B1(n_6534),
.B2(n_6281),
.Y(n_7849)
);

OAI22xp5_ASAP7_75t_L g7850 ( 
.A1(n_6882),
.A2(n_6087),
.B1(n_6250),
.B2(n_6178),
.Y(n_7850)
);

AOI22xp33_ASAP7_75t_L g7851 ( 
.A1(n_7304),
.A2(n_6079),
.B1(n_6534),
.B2(n_6281),
.Y(n_7851)
);

AOI22xp33_ASAP7_75t_L g7852 ( 
.A1(n_7304),
.A2(n_6079),
.B1(n_6534),
.B2(n_6281),
.Y(n_7852)
);

OAI21xp5_ASAP7_75t_SL g7853 ( 
.A1(n_7446),
.A2(n_6536),
.B(n_6779),
.Y(n_7853)
);

NAND2xp5_ASAP7_75t_L g7854 ( 
.A(n_6850),
.B(n_6595),
.Y(n_7854)
);

AOI22xp33_ASAP7_75t_SL g7855 ( 
.A1(n_6870),
.A2(n_6661),
.B1(n_6728),
.B2(n_6544),
.Y(n_7855)
);

INVx1_ASAP7_75t_L g7856 ( 
.A(n_6867),
.Y(n_7856)
);

BUFx6f_ASAP7_75t_L g7857 ( 
.A(n_7037),
.Y(n_7857)
);

NAND2xp5_ASAP7_75t_L g7858 ( 
.A(n_6852),
.B(n_6599),
.Y(n_7858)
);

OAI21xp5_ASAP7_75t_SL g7859 ( 
.A1(n_7428),
.A2(n_6536),
.B(n_6779),
.Y(n_7859)
);

AOI22xp33_ASAP7_75t_L g7860 ( 
.A1(n_7304),
.A2(n_6534),
.B1(n_6281),
.B2(n_6039),
.Y(n_7860)
);

AOI22xp33_ASAP7_75t_L g7861 ( 
.A1(n_7546),
.A2(n_6534),
.B1(n_6281),
.B2(n_6039),
.Y(n_7861)
);

OAI21xp5_ASAP7_75t_SL g7862 ( 
.A1(n_7021),
.A2(n_7442),
.B(n_7319),
.Y(n_7862)
);

INVx2_ASAP7_75t_L g7863 ( 
.A(n_7571),
.Y(n_7863)
);

CKINVDCx11_ASAP7_75t_R g7864 ( 
.A(n_7336),
.Y(n_7864)
);

INVx2_ASAP7_75t_L g7865 ( 
.A(n_7571),
.Y(n_7865)
);

AOI222xp33_ASAP7_75t_L g7866 ( 
.A1(n_7570),
.A2(n_6445),
.B1(n_6791),
.B2(n_6760),
.C1(n_6725),
.C2(n_6639),
.Y(n_7866)
);

BUFx2_ASAP7_75t_L g7867 ( 
.A(n_6881),
.Y(n_7867)
);

INVx2_ASAP7_75t_L g7868 ( 
.A(n_7618),
.Y(n_7868)
);

INVx1_ASAP7_75t_L g7869 ( 
.A(n_6880),
.Y(n_7869)
);

AOI22xp33_ASAP7_75t_L g7870 ( 
.A1(n_7546),
.A2(n_6534),
.B1(n_6104),
.B2(n_6388),
.Y(n_7870)
);

NAND2xp5_ASAP7_75t_L g7871 ( 
.A(n_6942),
.B(n_6599),
.Y(n_7871)
);

NAND2xp5_ASAP7_75t_L g7872 ( 
.A(n_6951),
.B(n_6606),
.Y(n_7872)
);

AOI22xp33_ASAP7_75t_L g7873 ( 
.A1(n_7546),
.A2(n_6104),
.B1(n_6388),
.B2(n_6574),
.Y(n_7873)
);

BUFx4f_ASAP7_75t_SL g7874 ( 
.A(n_7523),
.Y(n_7874)
);

AOI22xp33_ASAP7_75t_L g7875 ( 
.A1(n_7546),
.A2(n_6104),
.B1(n_6388),
.B2(n_6574),
.Y(n_7875)
);

INVx1_ASAP7_75t_L g7876 ( 
.A(n_6880),
.Y(n_7876)
);

INVx2_ASAP7_75t_L g7877 ( 
.A(n_7618),
.Y(n_7877)
);

NOR2xp33_ASAP7_75t_L g7878 ( 
.A(n_7211),
.B(n_6407),
.Y(n_7878)
);

AOI22xp33_ASAP7_75t_L g7879 ( 
.A1(n_7324),
.A2(n_6949),
.B1(n_6968),
.B2(n_6870),
.Y(n_7879)
);

NAND2xp5_ASAP7_75t_L g7880 ( 
.A(n_6903),
.B(n_6606),
.Y(n_7880)
);

AOI22xp33_ASAP7_75t_SL g7881 ( 
.A1(n_7360),
.A2(n_6661),
.B1(n_6728),
.B2(n_6544),
.Y(n_7881)
);

OAI22xp5_ASAP7_75t_L g7882 ( 
.A1(n_7573),
.A2(n_6178),
.B1(n_6293),
.B2(n_6250),
.Y(n_7882)
);

AOI22xp33_ASAP7_75t_SL g7883 ( 
.A1(n_7360),
.A2(n_6935),
.B1(n_6949),
.B2(n_6877),
.Y(n_7883)
);

AOI22xp33_ASAP7_75t_L g7884 ( 
.A1(n_7324),
.A2(n_6104),
.B1(n_6388),
.B2(n_6574),
.Y(n_7884)
);

AOI22xp33_ASAP7_75t_L g7885 ( 
.A1(n_7324),
.A2(n_6104),
.B1(n_6388),
.B2(n_6574),
.Y(n_7885)
);

OAI22xp5_ASAP7_75t_L g7886 ( 
.A1(n_7604),
.A2(n_6293),
.B1(n_6411),
.B2(n_6145),
.Y(n_7886)
);

INVx1_ASAP7_75t_L g7887 ( 
.A(n_6893),
.Y(n_7887)
);

INVx1_ASAP7_75t_L g7888 ( 
.A(n_6893),
.Y(n_7888)
);

BUFx6f_ASAP7_75t_L g7889 ( 
.A(n_7037),
.Y(n_7889)
);

BUFx3_ASAP7_75t_L g7890 ( 
.A(n_7475),
.Y(n_7890)
);

OAI22xp5_ASAP7_75t_L g7891 ( 
.A1(n_6823),
.A2(n_6901),
.B1(n_7570),
.B2(n_7624),
.Y(n_7891)
);

INVx1_ASAP7_75t_L g7892 ( 
.A(n_6897),
.Y(n_7892)
);

AOI22xp33_ASAP7_75t_L g7893 ( 
.A1(n_7324),
.A2(n_6104),
.B1(n_6388),
.B2(n_6574),
.Y(n_7893)
);

OAI21xp33_ASAP7_75t_L g7894 ( 
.A1(n_6877),
.A2(n_6605),
.B(n_6405),
.Y(n_7894)
);

AND2x2_ASAP7_75t_L g7895 ( 
.A(n_7070),
.B(n_6407),
.Y(n_7895)
);

INVx2_ASAP7_75t_L g7896 ( 
.A(n_7618),
.Y(n_7896)
);

INVx2_ASAP7_75t_L g7897 ( 
.A(n_7618),
.Y(n_7897)
);

HB1xp67_ASAP7_75t_L g7898 ( 
.A(n_6920),
.Y(n_7898)
);

OAI22xp5_ASAP7_75t_L g7899 ( 
.A1(n_6823),
.A2(n_6411),
.B1(n_6734),
.B2(n_6145),
.Y(n_7899)
);

OR2x2_ASAP7_75t_L g7900 ( 
.A(n_7317),
.B(n_7330),
.Y(n_7900)
);

NOR2xp33_ASAP7_75t_L g7901 ( 
.A(n_7211),
.B(n_6435),
.Y(n_7901)
);

INVx2_ASAP7_75t_SL g7902 ( 
.A(n_7238),
.Y(n_7902)
);

AOI22xp33_ASAP7_75t_SL g7903 ( 
.A1(n_6935),
.A2(n_6661),
.B1(n_6728),
.B2(n_6544),
.Y(n_7903)
);

AOI22xp33_ASAP7_75t_L g7904 ( 
.A1(n_7287),
.A2(n_6576),
.B1(n_6593),
.B2(n_6574),
.Y(n_7904)
);

AOI22xp33_ASAP7_75t_L g7905 ( 
.A1(n_6834),
.A2(n_6576),
.B1(n_6593),
.B2(n_6574),
.Y(n_7905)
);

AND2x2_ASAP7_75t_L g7906 ( 
.A(n_7162),
.B(n_6435),
.Y(n_7906)
);

AOI22xp33_ASAP7_75t_L g7907 ( 
.A1(n_6834),
.A2(n_6593),
.B1(n_6608),
.B2(n_6576),
.Y(n_7907)
);

INVx2_ASAP7_75t_SL g7908 ( 
.A(n_7238),
.Y(n_7908)
);

INVx1_ASAP7_75t_L g7909 ( 
.A(n_6897),
.Y(n_7909)
);

BUFx6f_ASAP7_75t_L g7910 ( 
.A(n_7037),
.Y(n_7910)
);

INVx1_ASAP7_75t_L g7911 ( 
.A(n_6905),
.Y(n_7911)
);

BUFx6f_ASAP7_75t_L g7912 ( 
.A(n_7037),
.Y(n_7912)
);

BUFx5_ASAP7_75t_L g7913 ( 
.A(n_7505),
.Y(n_7913)
);

AOI22xp33_ASAP7_75t_L g7914 ( 
.A1(n_6834),
.A2(n_6593),
.B1(n_6608),
.B2(n_6576),
.Y(n_7914)
);

AND2x2_ASAP7_75t_L g7915 ( 
.A(n_7162),
.B(n_6435),
.Y(n_7915)
);

AOI22xp33_ASAP7_75t_L g7916 ( 
.A1(n_6834),
.A2(n_6593),
.B1(n_6608),
.B2(n_6576),
.Y(n_7916)
);

AOI222xp33_ASAP7_75t_L g7917 ( 
.A1(n_7368),
.A2(n_6445),
.B1(n_6791),
.B2(n_6639),
.C1(n_6725),
.C2(n_6583),
.Y(n_7917)
);

INVx2_ASAP7_75t_L g7918 ( 
.A(n_7577),
.Y(n_7918)
);

OAI21xp5_ASAP7_75t_SL g7919 ( 
.A1(n_7382),
.A2(n_7403),
.B(n_7297),
.Y(n_7919)
);

INVx2_ASAP7_75t_L g7920 ( 
.A(n_7577),
.Y(n_7920)
);

AOI22xp33_ASAP7_75t_L g7921 ( 
.A1(n_6960),
.A2(n_6593),
.B1(n_6608),
.B2(n_6576),
.Y(n_7921)
);

NAND2xp5_ASAP7_75t_L g7922 ( 
.A(n_6912),
.B(n_6610),
.Y(n_7922)
);

INVx1_ASAP7_75t_L g7923 ( 
.A(n_6905),
.Y(n_7923)
);

NAND2xp5_ASAP7_75t_L g7924 ( 
.A(n_6872),
.B(n_6610),
.Y(n_7924)
);

AOI22xp33_ASAP7_75t_L g7925 ( 
.A1(n_6960),
.A2(n_6593),
.B1(n_6608),
.B2(n_6576),
.Y(n_7925)
);

INVx1_ASAP7_75t_L g7926 ( 
.A(n_6914),
.Y(n_7926)
);

OAI22xp5_ASAP7_75t_L g7927 ( 
.A1(n_6901),
.A2(n_7551),
.B1(n_7557),
.B2(n_7554),
.Y(n_7927)
);

OAI22xp5_ASAP7_75t_L g7928 ( 
.A1(n_6901),
.A2(n_6411),
.B1(n_6734),
.B2(n_6145),
.Y(n_7928)
);

OAI21xp5_ASAP7_75t_SL g7929 ( 
.A1(n_7293),
.A2(n_6536),
.B(n_6779),
.Y(n_7929)
);

INVx1_ASAP7_75t_L g7930 ( 
.A(n_6914),
.Y(n_7930)
);

INVx2_ASAP7_75t_L g7931 ( 
.A(n_7593),
.Y(n_7931)
);

INVxp67_ASAP7_75t_SL g7932 ( 
.A(n_7311),
.Y(n_7932)
);

AOI22xp5_ASAP7_75t_L g7933 ( 
.A1(n_7390),
.A2(n_6411),
.B1(n_6734),
.B2(n_6145),
.Y(n_7933)
);

INVx1_ASAP7_75t_L g7934 ( 
.A(n_6928),
.Y(n_7934)
);

AOI22xp33_ASAP7_75t_SL g7935 ( 
.A1(n_6935),
.A2(n_6661),
.B1(n_6728),
.B2(n_6544),
.Y(n_7935)
);

INVx1_ASAP7_75t_L g7936 ( 
.A(n_6928),
.Y(n_7936)
);

INVx2_ASAP7_75t_L g7937 ( 
.A(n_7593),
.Y(n_7937)
);

BUFx6f_ASAP7_75t_L g7938 ( 
.A(n_7073),
.Y(n_7938)
);

AOI22xp33_ASAP7_75t_SL g7939 ( 
.A1(n_6935),
.A2(n_6661),
.B1(n_6728),
.B2(n_6544),
.Y(n_7939)
);

OAI22xp5_ASAP7_75t_L g7940 ( 
.A1(n_7560),
.A2(n_6411),
.B1(n_6734),
.B2(n_6145),
.Y(n_7940)
);

OAI22xp5_ASAP7_75t_L g7941 ( 
.A1(n_6892),
.A2(n_6411),
.B1(n_6734),
.B2(n_6145),
.Y(n_7941)
);

INVx2_ASAP7_75t_L g7942 ( 
.A(n_7613),
.Y(n_7942)
);

OR2x2_ASAP7_75t_L g7943 ( 
.A(n_7330),
.B(n_6583),
.Y(n_7943)
);

AOI22xp33_ASAP7_75t_L g7944 ( 
.A1(n_6960),
.A2(n_6608),
.B1(n_6108),
.B2(n_6145),
.Y(n_7944)
);

AOI22xp33_ASAP7_75t_L g7945 ( 
.A1(n_6985),
.A2(n_6608),
.B1(n_6108),
.B2(n_6734),
.Y(n_7945)
);

NAND2xp5_ASAP7_75t_L g7946 ( 
.A(n_7426),
.B(n_6670),
.Y(n_7946)
);

HB1xp67_ASAP7_75t_L g7947 ( 
.A(n_6925),
.Y(n_7947)
);

OAI21xp5_ASAP7_75t_SL g7948 ( 
.A1(n_7197),
.A2(n_7190),
.B(n_7558),
.Y(n_7948)
);

AOI22xp33_ASAP7_75t_SL g7949 ( 
.A1(n_6866),
.A2(n_6661),
.B1(n_6728),
.B2(n_6544),
.Y(n_7949)
);

AOI22xp5_ASAP7_75t_L g7950 ( 
.A1(n_7420),
.A2(n_7424),
.B1(n_7504),
.B2(n_7505),
.Y(n_7950)
);

INVx3_ASAP7_75t_L g7951 ( 
.A(n_6881),
.Y(n_7951)
);

INVx1_ASAP7_75t_L g7952 ( 
.A(n_6938),
.Y(n_7952)
);

OAI22xp5_ASAP7_75t_L g7953 ( 
.A1(n_7505),
.A2(n_7556),
.B1(n_6888),
.B2(n_6847),
.Y(n_7953)
);

AOI22xp5_ASAP7_75t_L g7954 ( 
.A1(n_7556),
.A2(n_6785),
.B1(n_6536),
.B2(n_6111),
.Y(n_7954)
);

INVx1_ASAP7_75t_L g7955 ( 
.A(n_6938),
.Y(n_7955)
);

AOI22xp33_ASAP7_75t_SL g7956 ( 
.A1(n_6866),
.A2(n_7130),
.B1(n_6936),
.B2(n_7088),
.Y(n_7956)
);

AND2x2_ASAP7_75t_L g7957 ( 
.A(n_7201),
.B(n_6435),
.Y(n_7957)
);

BUFx12f_ASAP7_75t_L g7958 ( 
.A(n_7211),
.Y(n_7958)
);

AOI22xp33_ASAP7_75t_SL g7959 ( 
.A1(n_6866),
.A2(n_6144),
.B1(n_6187),
.B2(n_6165),
.Y(n_7959)
);

CKINVDCx5p33_ASAP7_75t_R g7960 ( 
.A(n_7230),
.Y(n_7960)
);

AOI22xp33_ASAP7_75t_SL g7961 ( 
.A1(n_6936),
.A2(n_6144),
.B1(n_6187),
.B2(n_6165),
.Y(n_7961)
);

AOI22xp5_ASAP7_75t_L g7962 ( 
.A1(n_7556),
.A2(n_6785),
.B1(n_6111),
.B2(n_6245),
.Y(n_7962)
);

INVx1_ASAP7_75t_L g7963 ( 
.A(n_6941),
.Y(n_7963)
);

AOI22xp33_ASAP7_75t_L g7964 ( 
.A1(n_6985),
.A2(n_7108),
.B1(n_7124),
.B2(n_6860),
.Y(n_7964)
);

AOI22xp33_ASAP7_75t_L g7965 ( 
.A1(n_6985),
.A2(n_6108),
.B1(n_6785),
.B2(n_6289),
.Y(n_7965)
);

AOI22xp33_ASAP7_75t_SL g7966 ( 
.A1(n_6936),
.A2(n_6144),
.B1(n_6187),
.B2(n_6165),
.Y(n_7966)
);

OAI22xp5_ASAP7_75t_L g7967 ( 
.A1(n_7347),
.A2(n_6785),
.B1(n_6111),
.B2(n_6245),
.Y(n_7967)
);

OAI22xp5_ASAP7_75t_L g7968 ( 
.A1(n_7458),
.A2(n_6785),
.B1(n_6111),
.B2(n_6245),
.Y(n_7968)
);

OAI222xp33_ASAP7_75t_L g7969 ( 
.A1(n_7014),
.A2(n_6656),
.B1(n_6605),
.B2(n_6667),
.C1(n_6655),
.C2(n_6405),
.Y(n_7969)
);

AOI22xp33_ASAP7_75t_L g7970 ( 
.A1(n_7108),
.A2(n_6108),
.B1(n_6785),
.B2(n_6289),
.Y(n_7970)
);

OAI22xp33_ASAP7_75t_L g7971 ( 
.A1(n_7169),
.A2(n_7550),
.B1(n_7441),
.B2(n_7457),
.Y(n_7971)
);

AOI22xp33_ASAP7_75t_L g7972 ( 
.A1(n_7108),
.A2(n_6108),
.B1(n_6785),
.B2(n_6289),
.Y(n_7972)
);

BUFx4f_ASAP7_75t_SL g7973 ( 
.A(n_7539),
.Y(n_7973)
);

AND2x2_ASAP7_75t_L g7974 ( 
.A(n_7201),
.B(n_6435),
.Y(n_7974)
);

INVx1_ASAP7_75t_L g7975 ( 
.A(n_6941),
.Y(n_7975)
);

HB1xp67_ASAP7_75t_L g7976 ( 
.A(n_7288),
.Y(n_7976)
);

INVx1_ASAP7_75t_L g7977 ( 
.A(n_6963),
.Y(n_7977)
);

OAI21xp5_ASAP7_75t_SL g7978 ( 
.A1(n_7485),
.A2(n_6655),
.B(n_6405),
.Y(n_7978)
);

AOI22xp33_ASAP7_75t_L g7979 ( 
.A1(n_7124),
.A2(n_6289),
.B1(n_6111),
.B2(n_6245),
.Y(n_7979)
);

AOI22xp33_ASAP7_75t_L g7980 ( 
.A1(n_7124),
.A2(n_6289),
.B1(n_6245),
.B2(n_6036),
.Y(n_7980)
);

NAND2xp5_ASAP7_75t_L g7981 ( 
.A(n_7603),
.B(n_6670),
.Y(n_7981)
);

AOI22xp33_ASAP7_75t_L g7982 ( 
.A1(n_7625),
.A2(n_6320),
.B1(n_6036),
.B2(n_5313),
.Y(n_7982)
);

AOI22xp33_ASAP7_75t_L g7983 ( 
.A1(n_7457),
.A2(n_6320),
.B1(n_6036),
.B2(n_5366),
.Y(n_7983)
);

AOI22xp33_ASAP7_75t_L g7984 ( 
.A1(n_7073),
.A2(n_6320),
.B1(n_6036),
.B2(n_5366),
.Y(n_7984)
);

AOI22xp33_ASAP7_75t_SL g7985 ( 
.A1(n_6936),
.A2(n_6220),
.B1(n_6298),
.B2(n_6278),
.Y(n_7985)
);

AOI22xp33_ASAP7_75t_SL g7986 ( 
.A1(n_7088),
.A2(n_6220),
.B1(n_6298),
.B2(n_6278),
.Y(n_7986)
);

BUFx2_ASAP7_75t_L g7987 ( 
.A(n_7521),
.Y(n_7987)
);

AOI22xp33_ASAP7_75t_L g7988 ( 
.A1(n_7073),
.A2(n_6320),
.B1(n_6036),
.B2(n_5371),
.Y(n_7988)
);

OR2x2_ASAP7_75t_L g7989 ( 
.A(n_7330),
.B(n_6746),
.Y(n_7989)
);

AOI22xp33_ASAP7_75t_L g7990 ( 
.A1(n_7073),
.A2(n_6320),
.B1(n_5371),
.B2(n_6276),
.Y(n_7990)
);

AND2x4_ASAP7_75t_L g7991 ( 
.A(n_7046),
.B(n_6553),
.Y(n_7991)
);

OAI21xp33_ASAP7_75t_L g7992 ( 
.A1(n_7447),
.A2(n_6655),
.B(n_6605),
.Y(n_7992)
);

AOI22xp33_ASAP7_75t_L g7993 ( 
.A1(n_7073),
.A2(n_5371),
.B1(n_6276),
.B2(n_6257),
.Y(n_7993)
);

AND2x2_ASAP7_75t_L g7994 ( 
.A(n_7281),
.B(n_6220),
.Y(n_7994)
);

AOI22xp33_ASAP7_75t_L g7995 ( 
.A1(n_7608),
.A2(n_5371),
.B1(n_6276),
.B2(n_6257),
.Y(n_7995)
);

OAI22xp5_ASAP7_75t_L g7996 ( 
.A1(n_6838),
.A2(n_6667),
.B1(n_6669),
.B2(n_6656),
.Y(n_7996)
);

HB1xp67_ASAP7_75t_L g7997 ( 
.A(n_7380),
.Y(n_7997)
);

CKINVDCx5p33_ASAP7_75t_R g7998 ( 
.A(n_7250),
.Y(n_7998)
);

AOI22xp33_ASAP7_75t_L g7999 ( 
.A1(n_7608),
.A2(n_6257),
.B1(n_6276),
.B2(n_6701),
.Y(n_7999)
);

INVx1_ASAP7_75t_L g8000 ( 
.A(n_6963),
.Y(n_8000)
);

AOI22xp33_ASAP7_75t_SL g8001 ( 
.A1(n_7200),
.A2(n_6298),
.B1(n_6278),
.B2(n_6447),
.Y(n_8001)
);

AOI21xp5_ASAP7_75t_L g8002 ( 
.A1(n_7346),
.A2(n_6512),
.B(n_6694),
.Y(n_8002)
);

OAI21xp5_ASAP7_75t_SL g8003 ( 
.A1(n_7310),
.A2(n_6667),
.B(n_6656),
.Y(n_8003)
);

OAI22xp33_ASAP7_75t_L g8004 ( 
.A1(n_7014),
.A2(n_6669),
.B1(n_5606),
.B2(n_6382),
.Y(n_8004)
);

AOI22xp33_ASAP7_75t_L g8005 ( 
.A1(n_7608),
.A2(n_6257),
.B1(n_6276),
.B2(n_6701),
.Y(n_8005)
);

OAI21xp5_ASAP7_75t_SL g8006 ( 
.A1(n_7392),
.A2(n_6669),
.B(n_6173),
.Y(n_8006)
);

AOI22xp33_ASAP7_75t_L g8007 ( 
.A1(n_7608),
.A2(n_6257),
.B1(n_6724),
.B2(n_6701),
.Y(n_8007)
);

CKINVDCx5p33_ASAP7_75t_R g8008 ( 
.A(n_7299),
.Y(n_8008)
);

OAI21xp5_ASAP7_75t_L g8009 ( 
.A1(n_7541),
.A2(n_6650),
.B(n_6708),
.Y(n_8009)
);

AOI22xp33_ASAP7_75t_L g8010 ( 
.A1(n_7311),
.A2(n_6701),
.B1(n_6796),
.B2(n_6724),
.Y(n_8010)
);

OAI21xp5_ASAP7_75t_SL g8011 ( 
.A1(n_6865),
.A2(n_6173),
.B(n_6164),
.Y(n_8011)
);

AOI22xp33_ASAP7_75t_SL g8012 ( 
.A1(n_7200),
.A2(n_6725),
.B1(n_6639),
.B2(n_6650),
.Y(n_8012)
);

AND2x2_ASAP7_75t_L g8013 ( 
.A(n_7281),
.B(n_6559),
.Y(n_8013)
);

INVx5_ASAP7_75t_L g8014 ( 
.A(n_7433),
.Y(n_8014)
);

NAND2xp5_ASAP7_75t_L g8015 ( 
.A(n_7612),
.B(n_6072),
.Y(n_8015)
);

AND2x2_ASAP7_75t_L g8016 ( 
.A(n_7322),
.B(n_6559),
.Y(n_8016)
);

CKINVDCx5p33_ASAP7_75t_R g8017 ( 
.A(n_7575),
.Y(n_8017)
);

AOI22xp33_ASAP7_75t_SL g8018 ( 
.A1(n_7159),
.A2(n_6774),
.B1(n_6710),
.B2(n_6780),
.Y(n_8018)
);

NOR2xp33_ASAP7_75t_L g8019 ( 
.A(n_7475),
.B(n_6512),
.Y(n_8019)
);

NAND2xp5_ASAP7_75t_L g8020 ( 
.A(n_6966),
.B(n_6072),
.Y(n_8020)
);

AOI22xp33_ASAP7_75t_L g8021 ( 
.A1(n_7159),
.A2(n_6724),
.B1(n_6796),
.B2(n_5090),
.Y(n_8021)
);

INVx1_ASAP7_75t_L g8022 ( 
.A(n_6982),
.Y(n_8022)
);

OAI22xp5_ASAP7_75t_L g8023 ( 
.A1(n_6841),
.A2(n_6796),
.B1(n_6724),
.B2(n_6618),
.Y(n_8023)
);

AOI22xp5_ASAP7_75t_L g8024 ( 
.A1(n_6817),
.A2(n_6539),
.B1(n_6618),
.B2(n_6594),
.Y(n_8024)
);

HB1xp67_ASAP7_75t_L g8025 ( 
.A(n_7381),
.Y(n_8025)
);

BUFx2_ASAP7_75t_L g8026 ( 
.A(n_7521),
.Y(n_8026)
);

INVx1_ASAP7_75t_L g8027 ( 
.A(n_6982),
.Y(n_8027)
);

INVx2_ASAP7_75t_L g8028 ( 
.A(n_7613),
.Y(n_8028)
);

INVx1_ASAP7_75t_L g8029 ( 
.A(n_6986),
.Y(n_8029)
);

INVxp67_ASAP7_75t_L g8030 ( 
.A(n_7452),
.Y(n_8030)
);

CKINVDCx11_ASAP7_75t_R g8031 ( 
.A(n_7336),
.Y(n_8031)
);

INVx1_ASAP7_75t_SL g8032 ( 
.A(n_7401),
.Y(n_8032)
);

AOI22xp33_ASAP7_75t_SL g8033 ( 
.A1(n_6947),
.A2(n_6774),
.B1(n_6710),
.B2(n_6780),
.Y(n_8033)
);

INVx2_ASAP7_75t_L g8034 ( 
.A(n_7496),
.Y(n_8034)
);

AOI22xp33_ASAP7_75t_SL g8035 ( 
.A1(n_6947),
.A2(n_6774),
.B1(n_6710),
.B2(n_6780),
.Y(n_8035)
);

OAI222xp33_ASAP7_75t_L g8036 ( 
.A1(n_7030),
.A2(n_6561),
.B1(n_6559),
.B2(n_6772),
.C1(n_6787),
.C2(n_6759),
.Y(n_8036)
);

INVx1_ASAP7_75t_L g8037 ( 
.A(n_6986),
.Y(n_8037)
);

INVx5_ASAP7_75t_SL g8038 ( 
.A(n_7433),
.Y(n_8038)
);

OAI22xp5_ASAP7_75t_L g8039 ( 
.A1(n_7252),
.A2(n_6796),
.B1(n_6618),
.B2(n_6619),
.Y(n_8039)
);

INVx2_ASAP7_75t_L g8040 ( 
.A(n_7496),
.Y(n_8040)
);

INVx5_ASAP7_75t_L g8041 ( 
.A(n_7433),
.Y(n_8041)
);

HB1xp67_ASAP7_75t_SL g8042 ( 
.A(n_7323),
.Y(n_8042)
);

AOI222xp33_ASAP7_75t_L g8043 ( 
.A1(n_7531),
.A2(n_6746),
.B1(n_6738),
.B2(n_6680),
.C1(n_6707),
.C2(n_6677),
.Y(n_8043)
);

BUFx12f_ASAP7_75t_L g8044 ( 
.A(n_7336),
.Y(n_8044)
);

OAI222xp33_ASAP7_75t_L g8045 ( 
.A1(n_7030),
.A2(n_6561),
.B1(n_6787),
.B2(n_6772),
.C1(n_6759),
.C2(n_6400),
.Y(n_8045)
);

AOI222xp33_ASAP7_75t_L g8046 ( 
.A1(n_7626),
.A2(n_6738),
.B1(n_6680),
.B2(n_6707),
.C1(n_6677),
.C2(n_6031),
.Y(n_8046)
);

AOI22xp33_ASAP7_75t_L g8047 ( 
.A1(n_7323),
.A2(n_4743),
.B1(n_4867),
.B2(n_4777),
.Y(n_8047)
);

AOI22xp33_ASAP7_75t_L g8048 ( 
.A1(n_7323),
.A2(n_4743),
.B1(n_4867),
.B2(n_4777),
.Y(n_8048)
);

AOI22xp33_ASAP7_75t_L g8049 ( 
.A1(n_7323),
.A2(n_4743),
.B1(n_4867),
.B2(n_4777),
.Y(n_8049)
);

OAI22xp5_ASAP7_75t_L g8050 ( 
.A1(n_7296),
.A2(n_6618),
.B1(n_6619),
.B2(n_6594),
.Y(n_8050)
);

OAI22xp5_ASAP7_75t_L g8051 ( 
.A1(n_7363),
.A2(n_6618),
.B1(n_6619),
.B2(n_6594),
.Y(n_8051)
);

OAI22xp5_ASAP7_75t_L g8052 ( 
.A1(n_7363),
.A2(n_6618),
.B1(n_6619),
.B2(n_6594),
.Y(n_8052)
);

INVx3_ASAP7_75t_L g8053 ( 
.A(n_7521),
.Y(n_8053)
);

OAI22xp5_ASAP7_75t_L g8054 ( 
.A1(n_7012),
.A2(n_6619),
.B1(n_6628),
.B2(n_6594),
.Y(n_8054)
);

AOI22xp33_ASAP7_75t_L g8055 ( 
.A1(n_7467),
.A2(n_4777),
.B1(n_4867),
.B2(n_6720),
.Y(n_8055)
);

INVx1_ASAP7_75t_L g8056 ( 
.A(n_6988),
.Y(n_8056)
);

OAI22xp5_ASAP7_75t_L g8057 ( 
.A1(n_7493),
.A2(n_6619),
.B1(n_6628),
.B2(n_6594),
.Y(n_8057)
);

INVx2_ASAP7_75t_L g8058 ( 
.A(n_7496),
.Y(n_8058)
);

INVx2_ASAP7_75t_SL g8059 ( 
.A(n_7238),
.Y(n_8059)
);

AOI22xp33_ASAP7_75t_L g8060 ( 
.A1(n_7467),
.A2(n_4777),
.B1(n_6720),
.B2(n_6110),
.Y(n_8060)
);

AOI22xp33_ASAP7_75t_L g8061 ( 
.A1(n_7467),
.A2(n_6720),
.B1(n_6110),
.B2(n_5091),
.Y(n_8061)
);

OAI21xp33_ASAP7_75t_L g8062 ( 
.A1(n_7501),
.A2(n_6561),
.B(n_6121),
.Y(n_8062)
);

OAI222xp33_ASAP7_75t_L g8063 ( 
.A1(n_6817),
.A2(n_6772),
.B1(n_6787),
.B2(n_6759),
.C1(n_6400),
.C2(n_6234),
.Y(n_8063)
);

INVx3_ASAP7_75t_L g8064 ( 
.A(n_7521),
.Y(n_8064)
);

AOI22xp33_ASAP7_75t_L g8065 ( 
.A1(n_7467),
.A2(n_6110),
.B1(n_5091),
.B2(n_4698),
.Y(n_8065)
);

AOI22xp33_ASAP7_75t_L g8066 ( 
.A1(n_7511),
.A2(n_6110),
.B1(n_5091),
.B2(n_4698),
.Y(n_8066)
);

NAND2xp5_ASAP7_75t_L g8067 ( 
.A(n_7060),
.B(n_6121),
.Y(n_8067)
);

INVx1_ASAP7_75t_SL g8068 ( 
.A(n_7475),
.Y(n_8068)
);

BUFx2_ASAP7_75t_L g8069 ( 
.A(n_7046),
.Y(n_8069)
);

NAND2xp5_ASAP7_75t_L g8070 ( 
.A(n_7028),
.B(n_6214),
.Y(n_8070)
);

AOI22xp33_ASAP7_75t_SL g8071 ( 
.A1(n_6947),
.A2(n_6774),
.B1(n_6710),
.B2(n_6780),
.Y(n_8071)
);

OAI21xp33_ASAP7_75t_L g8072 ( 
.A1(n_7385),
.A2(n_6173),
.B(n_6497),
.Y(n_8072)
);

AOI22xp33_ASAP7_75t_L g8073 ( 
.A1(n_7511),
.A2(n_7597),
.B1(n_6894),
.B2(n_7009),
.Y(n_8073)
);

INVx2_ASAP7_75t_L g8074 ( 
.A(n_7628),
.Y(n_8074)
);

AOI22xp33_ASAP7_75t_L g8075 ( 
.A1(n_7511),
.A2(n_7597),
.B1(n_6975),
.B2(n_6948),
.Y(n_8075)
);

NAND2xp5_ASAP7_75t_L g8076 ( 
.A(n_7038),
.B(n_6214),
.Y(n_8076)
);

INVx3_ASAP7_75t_L g8077 ( 
.A(n_7397),
.Y(n_8077)
);

INVx2_ASAP7_75t_L g8078 ( 
.A(n_7628),
.Y(n_8078)
);

OAI21xp5_ASAP7_75t_SL g8079 ( 
.A1(n_6865),
.A2(n_6164),
.B(n_6152),
.Y(n_8079)
);

OAI22xp5_ASAP7_75t_L g8080 ( 
.A1(n_7385),
.A2(n_6739),
.B1(n_6745),
.B2(n_6628),
.Y(n_8080)
);

INVx1_ASAP7_75t_L g8081 ( 
.A(n_6988),
.Y(n_8081)
);

HB1xp67_ASAP7_75t_L g8082 ( 
.A(n_7513),
.Y(n_8082)
);

AND2x2_ASAP7_75t_L g8083 ( 
.A(n_7322),
.B(n_6818),
.Y(n_8083)
);

INVx2_ASAP7_75t_L g8084 ( 
.A(n_6906),
.Y(n_8084)
);

AOI22xp33_ASAP7_75t_L g8085 ( 
.A1(n_7511),
.A2(n_6110),
.B1(n_5091),
.B2(n_4698),
.Y(n_8085)
);

BUFx2_ASAP7_75t_L g8086 ( 
.A(n_7046),
.Y(n_8086)
);

BUFx12f_ASAP7_75t_L g8087 ( 
.A(n_7336),
.Y(n_8087)
);

CKINVDCx5p33_ASAP7_75t_R g8088 ( 
.A(n_7490),
.Y(n_8088)
);

BUFx3_ASAP7_75t_L g8089 ( 
.A(n_7376),
.Y(n_8089)
);

AOI222xp33_ASAP7_75t_L g8090 ( 
.A1(n_7474),
.A2(n_6031),
.B1(n_6041),
.B2(n_6113),
.C1(n_6100),
.C2(n_6050),
.Y(n_8090)
);

HB1xp67_ASAP7_75t_SL g8091 ( 
.A(n_7193),
.Y(n_8091)
);

AOI22xp33_ASAP7_75t_L g8092 ( 
.A1(n_6948),
.A2(n_5091),
.B1(n_4698),
.B2(n_6717),
.Y(n_8092)
);

INVx4_ASAP7_75t_SL g8093 ( 
.A(n_6815),
.Y(n_8093)
);

AOI22xp33_ASAP7_75t_L g8094 ( 
.A1(n_6948),
.A2(n_6976),
.B1(n_7055),
.B2(n_6974),
.Y(n_8094)
);

AOI22xp33_ASAP7_75t_L g8095 ( 
.A1(n_6948),
.A2(n_5091),
.B1(n_4698),
.B2(n_6717),
.Y(n_8095)
);

AOI22xp33_ASAP7_75t_L g8096 ( 
.A1(n_6974),
.A2(n_5091),
.B1(n_4698),
.B2(n_6780),
.Y(n_8096)
);

NAND2xp5_ASAP7_75t_L g8097 ( 
.A(n_7290),
.B(n_6214),
.Y(n_8097)
);

INVx1_ASAP7_75t_L g8098 ( 
.A(n_6993),
.Y(n_8098)
);

INVxp67_ASAP7_75t_SL g8099 ( 
.A(n_7599),
.Y(n_8099)
);

INVx1_ASAP7_75t_L g8100 ( 
.A(n_6993),
.Y(n_8100)
);

BUFx6f_ASAP7_75t_L g8101 ( 
.A(n_7433),
.Y(n_8101)
);

AOI22xp33_ASAP7_75t_SL g8102 ( 
.A1(n_6947),
.A2(n_6710),
.B1(n_6774),
.B2(n_6780),
.Y(n_8102)
);

OAI21xp33_ASAP7_75t_L g8103 ( 
.A1(n_7385),
.A2(n_7421),
.B(n_7223),
.Y(n_8103)
);

AOI22xp33_ASAP7_75t_L g8104 ( 
.A1(n_6974),
.A2(n_5091),
.B1(n_4698),
.B2(n_6539),
.Y(n_8104)
);

OAI22xp5_ASAP7_75t_L g8105 ( 
.A1(n_6891),
.A2(n_6739),
.B1(n_6745),
.B2(n_6628),
.Y(n_8105)
);

INVx5_ASAP7_75t_SL g8106 ( 
.A(n_7434),
.Y(n_8106)
);

AND2x2_ASAP7_75t_L g8107 ( 
.A(n_6818),
.B(n_6553),
.Y(n_8107)
);

AOI22xp33_ASAP7_75t_L g8108 ( 
.A1(n_6974),
.A2(n_7055),
.B1(n_7071),
.B2(n_6976),
.Y(n_8108)
);

AOI22xp33_ASAP7_75t_L g8109 ( 
.A1(n_6976),
.A2(n_5091),
.B1(n_4698),
.B2(n_6539),
.Y(n_8109)
);

AOI22xp33_ASAP7_75t_SL g8110 ( 
.A1(n_6864),
.A2(n_6710),
.B1(n_6774),
.B2(n_6208),
.Y(n_8110)
);

BUFx4f_ASAP7_75t_SL g8111 ( 
.A(n_7434),
.Y(n_8111)
);

AOI22xp33_ASAP7_75t_L g8112 ( 
.A1(n_6976),
.A2(n_5091),
.B1(n_4698),
.B2(n_6539),
.Y(n_8112)
);

BUFx2_ASAP7_75t_L g8113 ( 
.A(n_7046),
.Y(n_8113)
);

NAND2xp5_ASAP7_75t_L g8114 ( 
.A(n_7300),
.B(n_7373),
.Y(n_8114)
);

CKINVDCx20_ASAP7_75t_R g8115 ( 
.A(n_7386),
.Y(n_8115)
);

INVx2_ASAP7_75t_L g8116 ( 
.A(n_6906),
.Y(n_8116)
);

BUFx2_ASAP7_75t_L g8117 ( 
.A(n_7046),
.Y(n_8117)
);

INVx2_ASAP7_75t_L g8118 ( 
.A(n_6906),
.Y(n_8118)
);

INVx1_ASAP7_75t_L g8119 ( 
.A(n_6994),
.Y(n_8119)
);

AOI22xp33_ASAP7_75t_L g8120 ( 
.A1(n_7055),
.A2(n_5091),
.B1(n_4698),
.B2(n_6539),
.Y(n_8120)
);

AOI22xp33_ASAP7_75t_SL g8121 ( 
.A1(n_6864),
.A2(n_6208),
.B1(n_6101),
.B2(n_6076),
.Y(n_8121)
);

OAI22xp5_ASAP7_75t_L g8122 ( 
.A1(n_6891),
.A2(n_6739),
.B1(n_6745),
.B2(n_6628),
.Y(n_8122)
);

OAI21xp5_ASAP7_75t_SL g8123 ( 
.A1(n_7384),
.A2(n_6164),
.B(n_6152),
.Y(n_8123)
);

INVx2_ASAP7_75t_SL g8124 ( 
.A(n_6891),
.Y(n_8124)
);

AND2x4_ASAP7_75t_L g8125 ( 
.A(n_7066),
.B(n_6553),
.Y(n_8125)
);

AND2x2_ASAP7_75t_L g8126 ( 
.A(n_6818),
.B(n_6553),
.Y(n_8126)
);

OAI21xp5_ASAP7_75t_SL g8127 ( 
.A1(n_7327),
.A2(n_6164),
.B(n_6152),
.Y(n_8127)
);

AOI22xp33_ASAP7_75t_L g8128 ( 
.A1(n_7055),
.A2(n_4698),
.B1(n_6539),
.B2(n_6164),
.Y(n_8128)
);

INVx2_ASAP7_75t_L g8129 ( 
.A(n_7478),
.Y(n_8129)
);

NAND2xp5_ASAP7_75t_L g8130 ( 
.A(n_7489),
.B(n_6214),
.Y(n_8130)
);

HB1xp67_ASAP7_75t_L g8131 ( 
.A(n_6853),
.Y(n_8131)
);

AOI22xp33_ASAP7_75t_L g8132 ( 
.A1(n_7071),
.A2(n_6164),
.B1(n_6193),
.B2(n_6152),
.Y(n_8132)
);

NAND3xp33_ASAP7_75t_L g8133 ( 
.A(n_6864),
.B(n_6708),
.C(n_6265),
.Y(n_8133)
);

INVx2_ASAP7_75t_L g8134 ( 
.A(n_7478),
.Y(n_8134)
);

AOI22xp33_ASAP7_75t_L g8135 ( 
.A1(n_7071),
.A2(n_6193),
.B1(n_6376),
.B2(n_6152),
.Y(n_8135)
);

AND2x2_ASAP7_75t_SL g8136 ( 
.A(n_6864),
.B(n_6926),
.Y(n_8136)
);

HB1xp67_ASAP7_75t_L g8137 ( 
.A(n_6853),
.Y(n_8137)
);

INVx2_ASAP7_75t_L g8138 ( 
.A(n_7478),
.Y(n_8138)
);

INVx1_ASAP7_75t_L g8139 ( 
.A(n_6994),
.Y(n_8139)
);

AOI22xp33_ASAP7_75t_SL g8140 ( 
.A1(n_6811),
.A2(n_6208),
.B1(n_6101),
.B2(n_6076),
.Y(n_8140)
);

OAI22xp5_ASAP7_75t_L g8141 ( 
.A1(n_7016),
.A2(n_6739),
.B1(n_6745),
.B2(n_6628),
.Y(n_8141)
);

AND2x2_ASAP7_75t_L g8142 ( 
.A(n_6818),
.B(n_6589),
.Y(n_8142)
);

INVx1_ASAP7_75t_L g8143 ( 
.A(n_7005),
.Y(n_8143)
);

INVx1_ASAP7_75t_L g8144 ( 
.A(n_7005),
.Y(n_8144)
);

AOI22xp33_ASAP7_75t_L g8145 ( 
.A1(n_7071),
.A2(n_6193),
.B1(n_6376),
.B2(n_6152),
.Y(n_8145)
);

INVx1_ASAP7_75t_L g8146 ( 
.A(n_7041),
.Y(n_8146)
);

AND2x2_ASAP7_75t_L g8147 ( 
.A(n_6824),
.B(n_6589),
.Y(n_8147)
);

BUFx6f_ASAP7_75t_L g8148 ( 
.A(n_7434),
.Y(n_8148)
);

INVx1_ASAP7_75t_L g8149 ( 
.A(n_7041),
.Y(n_8149)
);

AOI22xp33_ASAP7_75t_L g8150 ( 
.A1(n_7127),
.A2(n_6376),
.B1(n_6423),
.B2(n_6193),
.Y(n_8150)
);

AOI22xp33_ASAP7_75t_SL g8151 ( 
.A1(n_6811),
.A2(n_6101),
.B1(n_6266),
.B2(n_6076),
.Y(n_8151)
);

OAI22xp5_ASAP7_75t_L g8152 ( 
.A1(n_7027),
.A2(n_6745),
.B1(n_6752),
.B2(n_6739),
.Y(n_8152)
);

AOI22xp33_ASAP7_75t_L g8153 ( 
.A1(n_7127),
.A2(n_6193),
.B1(n_6423),
.B2(n_6376),
.Y(n_8153)
);

AOI22xp33_ASAP7_75t_L g8154 ( 
.A1(n_7151),
.A2(n_6193),
.B1(n_6423),
.B2(n_6376),
.Y(n_8154)
);

INVx2_ASAP7_75t_L g8155 ( 
.A(n_7478),
.Y(n_8155)
);

INVx2_ASAP7_75t_SL g8156 ( 
.A(n_7434),
.Y(n_8156)
);

AOI22xp5_ASAP7_75t_SL g8157 ( 
.A1(n_7329),
.A2(n_6266),
.B1(n_6277),
.B2(n_6101),
.Y(n_8157)
);

INVx2_ASAP7_75t_L g8158 ( 
.A(n_7479),
.Y(n_8158)
);

INVx1_ASAP7_75t_L g8159 ( 
.A(n_7065),
.Y(n_8159)
);

OAI21xp5_ASAP7_75t_L g8160 ( 
.A1(n_7544),
.A2(n_6497),
.B(n_6482),
.Y(n_8160)
);

INVx1_ASAP7_75t_L g8161 ( 
.A(n_7065),
.Y(n_8161)
);

AOI22xp33_ASAP7_75t_L g8162 ( 
.A1(n_7151),
.A2(n_6423),
.B1(n_6426),
.B2(n_6376),
.Y(n_8162)
);

INVx1_ASAP7_75t_L g8163 ( 
.A(n_7069),
.Y(n_8163)
);

HB1xp67_ASAP7_75t_L g8164 ( 
.A(n_7006),
.Y(n_8164)
);

AOI22xp33_ASAP7_75t_SL g8165 ( 
.A1(n_6811),
.A2(n_6266),
.B1(n_6277),
.B2(n_6101),
.Y(n_8165)
);

NAND2xp5_ASAP7_75t_L g8166 ( 
.A(n_7494),
.B(n_6214),
.Y(n_8166)
);

NOR2xp33_ASAP7_75t_L g8167 ( 
.A(n_7406),
.B(n_6234),
.Y(n_8167)
);

AOI22xp33_ASAP7_75t_L g8168 ( 
.A1(n_6814),
.A2(n_6426),
.B1(n_6528),
.B2(n_6423),
.Y(n_8168)
);

AOI22xp33_ASAP7_75t_L g8169 ( 
.A1(n_6814),
.A2(n_7350),
.B1(n_6926),
.B2(n_7145),
.Y(n_8169)
);

NOR2xp33_ASAP7_75t_L g8170 ( 
.A(n_7492),
.B(n_6338),
.Y(n_8170)
);

BUFx3_ASAP7_75t_L g8171 ( 
.A(n_7434),
.Y(n_8171)
);

NAND2xp5_ASAP7_75t_L g8172 ( 
.A(n_7209),
.B(n_6214),
.Y(n_8172)
);

INVx4_ASAP7_75t_L g8173 ( 
.A(n_7066),
.Y(n_8173)
);

AOI22xp33_ASAP7_75t_L g8174 ( 
.A1(n_6814),
.A2(n_6426),
.B1(n_6528),
.B2(n_6423),
.Y(n_8174)
);

AOI22xp33_ASAP7_75t_L g8175 ( 
.A1(n_6814),
.A2(n_6528),
.B1(n_6426),
.B2(n_6266),
.Y(n_8175)
);

INVx2_ASAP7_75t_L g8176 ( 
.A(n_7479),
.Y(n_8176)
);

INVx2_ASAP7_75t_L g8177 ( 
.A(n_7479),
.Y(n_8177)
);

AOI22xp33_ASAP7_75t_SL g8178 ( 
.A1(n_7350),
.A2(n_6266),
.B1(n_6277),
.B2(n_6101),
.Y(n_8178)
);

BUFx6f_ASAP7_75t_L g8179 ( 
.A(n_7443),
.Y(n_8179)
);

OAI22xp5_ASAP7_75t_L g8180 ( 
.A1(n_7519),
.A2(n_6745),
.B1(n_6752),
.B2(n_6739),
.Y(n_8180)
);

AND2x2_ASAP7_75t_L g8181 ( 
.A(n_6824),
.B(n_6589),
.Y(n_8181)
);

INVx4_ASAP7_75t_L g8182 ( 
.A(n_7066),
.Y(n_8182)
);

AND2x2_ASAP7_75t_L g8183 ( 
.A(n_6824),
.B(n_7092),
.Y(n_8183)
);

OAI22xp33_ASAP7_75t_L g8184 ( 
.A1(n_6871),
.A2(n_6101),
.B1(n_6277),
.B2(n_6266),
.Y(n_8184)
);

BUFx4f_ASAP7_75t_SL g8185 ( 
.A(n_7443),
.Y(n_8185)
);

AOI22xp33_ASAP7_75t_L g8186 ( 
.A1(n_7350),
.A2(n_6528),
.B1(n_6426),
.B2(n_6266),
.Y(n_8186)
);

AOI22xp5_ASAP7_75t_L g8187 ( 
.A1(n_6926),
.A2(n_6805),
.B1(n_6752),
.B2(n_6528),
.Y(n_8187)
);

BUFx4f_ASAP7_75t_SL g8188 ( 
.A(n_7443),
.Y(n_8188)
);

INVx1_ASAP7_75t_L g8189 ( 
.A(n_7069),
.Y(n_8189)
);

OAI21xp5_ASAP7_75t_SL g8190 ( 
.A1(n_7215),
.A2(n_6528),
.B(n_6426),
.Y(n_8190)
);

AOI22xp33_ASAP7_75t_L g8191 ( 
.A1(n_6926),
.A2(n_6266),
.B1(n_6277),
.B2(n_6101),
.Y(n_8191)
);

AOI22xp33_ASAP7_75t_L g8192 ( 
.A1(n_7145),
.A2(n_6824),
.B1(n_6959),
.B2(n_7268),
.Y(n_8192)
);

INVx1_ASAP7_75t_L g8193 ( 
.A(n_7075),
.Y(n_8193)
);

INVx5_ASAP7_75t_L g8194 ( 
.A(n_7443),
.Y(n_8194)
);

AOI22xp33_ASAP7_75t_SL g8195 ( 
.A1(n_7581),
.A2(n_6277),
.B1(n_6344),
.B2(n_6328),
.Y(n_8195)
);

AOI22xp33_ASAP7_75t_L g8196 ( 
.A1(n_7145),
.A2(n_6277),
.B1(n_6344),
.B2(n_6328),
.Y(n_8196)
);

AOI22xp33_ASAP7_75t_L g8197 ( 
.A1(n_6959),
.A2(n_7343),
.B1(n_7594),
.B2(n_7572),
.Y(n_8197)
);

AOI22xp33_ASAP7_75t_L g8198 ( 
.A1(n_6959),
.A2(n_6277),
.B1(n_6344),
.B2(n_6328),
.Y(n_8198)
);

INVx1_ASAP7_75t_L g8199 ( 
.A(n_7075),
.Y(n_8199)
);

OAI22xp5_ASAP7_75t_L g8200 ( 
.A1(n_6871),
.A2(n_6752),
.B1(n_6805),
.B2(n_5691),
.Y(n_8200)
);

OAI22xp5_ASAP7_75t_L g8201 ( 
.A1(n_6961),
.A2(n_6752),
.B1(n_6805),
.B2(n_5724),
.Y(n_8201)
);

AND2x2_ASAP7_75t_L g8202 ( 
.A(n_7092),
.B(n_6589),
.Y(n_8202)
);

OAI21xp5_ASAP7_75t_SL g8203 ( 
.A1(n_7427),
.A2(n_6065),
.B(n_6061),
.Y(n_8203)
);

INVx1_ASAP7_75t_L g8204 ( 
.A(n_7076),
.Y(n_8204)
);

AOI22xp33_ASAP7_75t_L g8205 ( 
.A1(n_7343),
.A2(n_6328),
.B1(n_6382),
.B2(n_6344),
.Y(n_8205)
);

AOI21xp33_ASAP7_75t_L g8206 ( 
.A1(n_6878),
.A2(n_6237),
.B(n_6224),
.Y(n_8206)
);

INVx2_ASAP7_75t_L g8207 ( 
.A(n_7479),
.Y(n_8207)
);

BUFx3_ASAP7_75t_L g8208 ( 
.A(n_7443),
.Y(n_8208)
);

CKINVDCx5p33_ASAP7_75t_R g8209 ( 
.A(n_7066),
.Y(n_8209)
);

INVx1_ASAP7_75t_L g8210 ( 
.A(n_7076),
.Y(n_8210)
);

INVx1_ASAP7_75t_L g8211 ( 
.A(n_7081),
.Y(n_8211)
);

OAI22xp33_ASAP7_75t_L g8212 ( 
.A1(n_6961),
.A2(n_6382),
.B1(n_6344),
.B2(n_6328),
.Y(n_8212)
);

INVx1_ASAP7_75t_L g8213 ( 
.A(n_7081),
.Y(n_8213)
);

INVx3_ASAP7_75t_L g8214 ( 
.A(n_7397),
.Y(n_8214)
);

INVx1_ASAP7_75t_L g8215 ( 
.A(n_7084),
.Y(n_8215)
);

AOI22xp33_ASAP7_75t_L g8216 ( 
.A1(n_7343),
.A2(n_6328),
.B1(n_6382),
.B2(n_6344),
.Y(n_8216)
);

OAI21xp33_ASAP7_75t_L g8217 ( 
.A1(n_7221),
.A2(n_6497),
.B(n_6041),
.Y(n_8217)
);

OAI21xp5_ASAP7_75t_SL g8218 ( 
.A1(n_7427),
.A2(n_6065),
.B(n_6061),
.Y(n_8218)
);

OAI21xp33_ASAP7_75t_L g8219 ( 
.A1(n_7079),
.A2(n_6041),
.B(n_6031),
.Y(n_8219)
);

AOI22xp33_ASAP7_75t_SL g8220 ( 
.A1(n_7581),
.A2(n_6328),
.B1(n_6382),
.B2(n_6344),
.Y(n_8220)
);

AND2x4_ASAP7_75t_L g8221 ( 
.A(n_7066),
.B(n_6589),
.Y(n_8221)
);

AOI22xp33_ASAP7_75t_SL g8222 ( 
.A1(n_7006),
.A2(n_6328),
.B1(n_6382),
.B2(n_6344),
.Y(n_8222)
);

AO22x1_ASAP7_75t_L g8223 ( 
.A1(n_7464),
.A2(n_6419),
.B1(n_6487),
.B2(n_6382),
.Y(n_8223)
);

INVx2_ASAP7_75t_L g8224 ( 
.A(n_7469),
.Y(n_8224)
);

INVx3_ASAP7_75t_SL g8225 ( 
.A(n_7464),
.Y(n_8225)
);

AOI22xp33_ASAP7_75t_L g8226 ( 
.A1(n_7572),
.A2(n_6382),
.B1(n_6487),
.B2(n_6419),
.Y(n_8226)
);

AND2x2_ASAP7_75t_L g8227 ( 
.A(n_7092),
.B(n_6589),
.Y(n_8227)
);

OAI22xp5_ASAP7_75t_L g8228 ( 
.A1(n_6981),
.A2(n_7091),
.B1(n_7369),
.B2(n_6998),
.Y(n_8228)
);

INVx1_ASAP7_75t_L g8229 ( 
.A(n_7084),
.Y(n_8229)
);

AOI22xp33_ASAP7_75t_L g8230 ( 
.A1(n_7572),
.A2(n_6419),
.B1(n_6487),
.B2(n_6589),
.Y(n_8230)
);

AOI22xp33_ASAP7_75t_SL g8231 ( 
.A1(n_7017),
.A2(n_6419),
.B1(n_6487),
.B2(n_6174),
.Y(n_8231)
);

OAI22xp33_ASAP7_75t_L g8232 ( 
.A1(n_6981),
.A2(n_6487),
.B1(n_6419),
.B2(n_6235),
.Y(n_8232)
);

INVx1_ASAP7_75t_L g8233 ( 
.A(n_7087),
.Y(n_8233)
);

AOI22xp33_ASAP7_75t_SL g8234 ( 
.A1(n_7017),
.A2(n_6419),
.B1(n_6487),
.B2(n_6174),
.Y(n_8234)
);

INVx1_ASAP7_75t_L g8235 ( 
.A(n_7087),
.Y(n_8235)
);

NOR2xp33_ASAP7_75t_L g8236 ( 
.A(n_7251),
.B(n_6338),
.Y(n_8236)
);

INVx1_ASAP7_75t_L g8237 ( 
.A(n_7097),
.Y(n_8237)
);

BUFx3_ASAP7_75t_L g8238 ( 
.A(n_7464),
.Y(n_8238)
);

OAI21xp5_ASAP7_75t_SL g8239 ( 
.A1(n_7552),
.A2(n_6065),
.B(n_6061),
.Y(n_8239)
);

HB1xp67_ASAP7_75t_L g8240 ( 
.A(n_6952),
.Y(n_8240)
);

OAI21xp33_ASAP7_75t_L g8241 ( 
.A1(n_7079),
.A2(n_6041),
.B(n_6031),
.Y(n_8241)
);

AOI22xp33_ASAP7_75t_L g8242 ( 
.A1(n_7572),
.A2(n_6419),
.B1(n_6487),
.B2(n_6752),
.Y(n_8242)
);

AND2x2_ASAP7_75t_L g8243 ( 
.A(n_7092),
.B(n_6805),
.Y(n_8243)
);

BUFx4f_ASAP7_75t_SL g8244 ( 
.A(n_7464),
.Y(n_8244)
);

AOI22xp5_ASAP7_75t_L g8245 ( 
.A1(n_7174),
.A2(n_6805),
.B1(n_6802),
.B2(n_6061),
.Y(n_8245)
);

AO22x1_ASAP7_75t_L g8246 ( 
.A1(n_7464),
.A2(n_6487),
.B1(n_6419),
.B2(n_6235),
.Y(n_8246)
);

BUFx12f_ASAP7_75t_L g8247 ( 
.A(n_7470),
.Y(n_8247)
);

NAND2xp5_ASAP7_75t_L g8248 ( 
.A(n_7244),
.B(n_6214),
.Y(n_8248)
);

HB1xp67_ASAP7_75t_L g8249 ( 
.A(n_6978),
.Y(n_8249)
);

NAND2xp5_ASAP7_75t_L g8250 ( 
.A(n_7374),
.B(n_6214),
.Y(n_8250)
);

INVx1_ASAP7_75t_L g8251 ( 
.A(n_7097),
.Y(n_8251)
);

OAI222xp33_ASAP7_75t_L g8252 ( 
.A1(n_6998),
.A2(n_6772),
.B1(n_6759),
.B2(n_6787),
.C1(n_6665),
.C2(n_6604),
.Y(n_8252)
);

INVx1_ASAP7_75t_L g8253 ( 
.A(n_7099),
.Y(n_8253)
);

OAI222xp33_ASAP7_75t_L g8254 ( 
.A1(n_7091),
.A2(n_6772),
.B1(n_6759),
.B2(n_6787),
.C1(n_6665),
.C2(n_6604),
.Y(n_8254)
);

AND2x2_ASAP7_75t_L g8255 ( 
.A(n_7174),
.B(n_6805),
.Y(n_8255)
);

AOI22xp33_ASAP7_75t_L g8256 ( 
.A1(n_7594),
.A2(n_6174),
.B1(n_6237),
.B2(n_6224),
.Y(n_8256)
);

AOI22xp33_ASAP7_75t_SL g8257 ( 
.A1(n_7321),
.A2(n_6174),
.B1(n_6203),
.B2(n_6679),
.Y(n_8257)
);

NAND2xp5_ASAP7_75t_L g8258 ( 
.A(n_7394),
.B(n_6263),
.Y(n_8258)
);

OAI21xp5_ASAP7_75t_SL g8259 ( 
.A1(n_7574),
.A2(n_6065),
.B(n_6061),
.Y(n_8259)
);

NAND2xp5_ASAP7_75t_SL g8260 ( 
.A(n_7470),
.B(n_6061),
.Y(n_8260)
);

INVx4_ASAP7_75t_L g8261 ( 
.A(n_7470),
.Y(n_8261)
);

OAI21xp5_ASAP7_75t_SL g8262 ( 
.A1(n_6917),
.A2(n_6065),
.B(n_6802),
.Y(n_8262)
);

AOI22xp33_ASAP7_75t_SL g8263 ( 
.A1(n_7321),
.A2(n_6174),
.B1(n_6203),
.B2(n_6679),
.Y(n_8263)
);

AOI22xp33_ASAP7_75t_L g8264 ( 
.A1(n_7594),
.A2(n_7614),
.B1(n_7622),
.B2(n_7611),
.Y(n_8264)
);

AOI22xp33_ASAP7_75t_SL g8265 ( 
.A1(n_7321),
.A2(n_6203),
.B1(n_6696),
.B2(n_6679),
.Y(n_8265)
);

AND2x2_ASAP7_75t_L g8266 ( 
.A(n_7174),
.B(n_6630),
.Y(n_8266)
);

AOI22xp33_ASAP7_75t_L g8267 ( 
.A1(n_7594),
.A2(n_6237),
.B1(n_6224),
.B2(n_6065),
.Y(n_8267)
);

INVx2_ASAP7_75t_L g8268 ( 
.A(n_7469),
.Y(n_8268)
);

INVx2_ASAP7_75t_L g8269 ( 
.A(n_7469),
.Y(n_8269)
);

OAI22xp5_ASAP7_75t_L g8270 ( 
.A1(n_7369),
.A2(n_5724),
.B1(n_5452),
.B2(n_5970),
.Y(n_8270)
);

NAND2xp5_ASAP7_75t_L g8271 ( 
.A(n_7400),
.B(n_6263),
.Y(n_8271)
);

OAI22xp5_ASAP7_75t_SL g8272 ( 
.A1(n_7569),
.A2(n_6235),
.B1(n_6236),
.B2(n_6181),
.Y(n_8272)
);

AOI22xp33_ASAP7_75t_L g8273 ( 
.A1(n_7611),
.A2(n_7614),
.B1(n_7627),
.B2(n_7622),
.Y(n_8273)
);

OAI22xp5_ASAP7_75t_L g8274 ( 
.A1(n_7257),
.A2(n_5970),
.B1(n_5373),
.B2(n_5387),
.Y(n_8274)
);

AOI22xp33_ASAP7_75t_L g8275 ( 
.A1(n_7611),
.A2(n_6224),
.B1(n_6237),
.B2(n_5970),
.Y(n_8275)
);

CKINVDCx14_ASAP7_75t_R g8276 ( 
.A(n_7329),
.Y(n_8276)
);

NAND2xp5_ASAP7_75t_L g8277 ( 
.A(n_7402),
.B(n_6263),
.Y(n_8277)
);

AOI22xp5_ASAP7_75t_L g8278 ( 
.A1(n_7174),
.A2(n_6802),
.B1(n_5970),
.B2(n_6237),
.Y(n_8278)
);

NAND2xp5_ASAP7_75t_L g8279 ( 
.A(n_7239),
.B(n_6263),
.Y(n_8279)
);

AOI22xp5_ASAP7_75t_L g8280 ( 
.A1(n_7242),
.A2(n_6802),
.B1(n_6224),
.B2(n_6236),
.Y(n_8280)
);

NOR2xp33_ASAP7_75t_L g8281 ( 
.A(n_7451),
.B(n_6500),
.Y(n_8281)
);

OAI21xp5_ASAP7_75t_SL g8282 ( 
.A1(n_6917),
.A2(n_6100),
.B(n_6050),
.Y(n_8282)
);

AOI22xp33_ASAP7_75t_L g8283 ( 
.A1(n_7611),
.A2(n_4679),
.B1(n_6503),
.B2(n_6495),
.Y(n_8283)
);

AOI22xp33_ASAP7_75t_SL g8284 ( 
.A1(n_7335),
.A2(n_6696),
.B1(n_6679),
.B2(n_6495),
.Y(n_8284)
);

HB1xp67_ASAP7_75t_L g8285 ( 
.A(n_6980),
.Y(n_8285)
);

OAI22xp5_ASAP7_75t_L g8286 ( 
.A1(n_6899),
.A2(n_5373),
.B1(n_5387),
.B2(n_5182),
.Y(n_8286)
);

OAI222xp33_ASAP7_75t_L g8287 ( 
.A1(n_6908),
.A2(n_6635),
.B1(n_6500),
.B2(n_6139),
.C1(n_6100),
.C2(n_6113),
.Y(n_8287)
);

AOI22xp33_ASAP7_75t_L g8288 ( 
.A1(n_7614),
.A2(n_4679),
.B1(n_6503),
.B2(n_6495),
.Y(n_8288)
);

OAI21xp5_ASAP7_75t_L g8289 ( 
.A1(n_7279),
.A2(n_6482),
.B(n_6644),
.Y(n_8289)
);

AOI22xp5_ASAP7_75t_L g8290 ( 
.A1(n_7242),
.A2(n_6236),
.B1(n_6317),
.B2(n_6181),
.Y(n_8290)
);

AOI22xp33_ASAP7_75t_L g8291 ( 
.A1(n_7614),
.A2(n_4679),
.B1(n_6503),
.B2(n_6495),
.Y(n_8291)
);

INVx2_ASAP7_75t_L g8292 ( 
.A(n_7469),
.Y(n_8292)
);

AND2x2_ASAP7_75t_L g8293 ( 
.A(n_7242),
.B(n_6630),
.Y(n_8293)
);

OAI21xp5_ASAP7_75t_L g8294 ( 
.A1(n_7279),
.A2(n_6482),
.B(n_6644),
.Y(n_8294)
);

AND2x2_ASAP7_75t_L g8295 ( 
.A(n_7242),
.B(n_6630),
.Y(n_8295)
);

OAI22xp5_ASAP7_75t_L g8296 ( 
.A1(n_6899),
.A2(n_6317),
.B1(n_6346),
.B2(n_6181),
.Y(n_8296)
);

INVx1_ASAP7_75t_L g8297 ( 
.A(n_7099),
.Y(n_8297)
);

AOI22xp33_ASAP7_75t_L g8298 ( 
.A1(n_7622),
.A2(n_6475),
.B1(n_6503),
.B2(n_6495),
.Y(n_8298)
);

BUFx8_ASAP7_75t_L g8299 ( 
.A(n_7339),
.Y(n_8299)
);

AOI21xp5_ASAP7_75t_L g8300 ( 
.A1(n_6878),
.A2(n_6346),
.B(n_6317),
.Y(n_8300)
);

AOI22xp33_ASAP7_75t_L g8301 ( 
.A1(n_7622),
.A2(n_6503),
.B1(n_6495),
.B2(n_6475),
.Y(n_8301)
);

INVx3_ASAP7_75t_L g8302 ( 
.A(n_7397),
.Y(n_8302)
);

AOI22xp33_ASAP7_75t_L g8303 ( 
.A1(n_7627),
.A2(n_6503),
.B1(n_6475),
.B2(n_6191),
.Y(n_8303)
);

AO22x1_ASAP7_75t_L g8304 ( 
.A1(n_7470),
.A2(n_6409),
.B1(n_6461),
.B2(n_6346),
.Y(n_8304)
);

BUFx5_ASAP7_75t_L g8305 ( 
.A(n_7627),
.Y(n_8305)
);

INVx3_ASAP7_75t_L g8306 ( 
.A(n_6933),
.Y(n_8306)
);

AOI22xp33_ASAP7_75t_L g8307 ( 
.A1(n_7627),
.A2(n_6475),
.B1(n_6191),
.B2(n_6461),
.Y(n_8307)
);

INVx1_ASAP7_75t_L g8308 ( 
.A(n_7106),
.Y(n_8308)
);

AND2x2_ASAP7_75t_L g8309 ( 
.A(n_7326),
.B(n_6630),
.Y(n_8309)
);

INVx1_ASAP7_75t_L g8310 ( 
.A(n_7106),
.Y(n_8310)
);

AOI22xp33_ASAP7_75t_SL g8311 ( 
.A1(n_7335),
.A2(n_6679),
.B1(n_6696),
.B2(n_6475),
.Y(n_8311)
);

AOI22xp33_ASAP7_75t_L g8312 ( 
.A1(n_7326),
.A2(n_6475),
.B1(n_6191),
.B2(n_6461),
.Y(n_8312)
);

INVx2_ASAP7_75t_L g8313 ( 
.A(n_7471),
.Y(n_8313)
);

BUFx4f_ASAP7_75t_SL g8314 ( 
.A(n_7470),
.Y(n_8314)
);

AOI221xp5_ASAP7_75t_L g8315 ( 
.A1(n_7335),
.A2(n_6100),
.B1(n_6139),
.B2(n_6113),
.C(n_6050),
.Y(n_8315)
);

INVx2_ASAP7_75t_L g8316 ( 
.A(n_7471),
.Y(n_8316)
);

NAND2xp5_ASAP7_75t_L g8317 ( 
.A(n_7422),
.B(n_6263),
.Y(n_8317)
);

AOI22xp33_ASAP7_75t_L g8318 ( 
.A1(n_7326),
.A2(n_6476),
.B1(n_6409),
.B2(n_5424),
.Y(n_8318)
);

OAI222xp33_ASAP7_75t_L g8319 ( 
.A1(n_6908),
.A2(n_6635),
.B1(n_6050),
.B2(n_6139),
.C1(n_6113),
.C2(n_6476),
.Y(n_8319)
);

HB1xp67_ASAP7_75t_L g8320 ( 
.A(n_7059),
.Y(n_8320)
);

OAI22xp5_ASAP7_75t_L g8321 ( 
.A1(n_6932),
.A2(n_6409),
.B1(n_6476),
.B2(n_6139),
.Y(n_8321)
);

INVx1_ASAP7_75t_L g8322 ( 
.A(n_7129),
.Y(n_8322)
);

AOI22xp33_ASAP7_75t_L g8323 ( 
.A1(n_7326),
.A2(n_5424),
.B1(n_5565),
.B2(n_5318),
.Y(n_8323)
);

CKINVDCx5p33_ASAP7_75t_R g8324 ( 
.A(n_7508),
.Y(n_8324)
);

NOR2xp33_ASAP7_75t_L g8325 ( 
.A(n_7104),
.B(n_6044),
.Y(n_8325)
);

INVx1_ASAP7_75t_L g8326 ( 
.A(n_7129),
.Y(n_8326)
);

HB1xp67_ASAP7_75t_L g8327 ( 
.A(n_7112),
.Y(n_8327)
);

CKINVDCx6p67_ASAP7_75t_R g8328 ( 
.A(n_7508),
.Y(n_8328)
);

AOI22xp33_ASAP7_75t_L g8329 ( 
.A1(n_7331),
.A2(n_5424),
.B1(n_5565),
.B2(n_5318),
.Y(n_8329)
);

BUFx4f_ASAP7_75t_SL g8330 ( 
.A(n_7508),
.Y(n_8330)
);

NOR2xp33_ASAP7_75t_R g8331 ( 
.A(n_7001),
.B(n_6197),
.Y(n_8331)
);

NAND3xp33_ASAP7_75t_L g8332 ( 
.A(n_7328),
.B(n_6265),
.C(n_6225),
.Y(n_8332)
);

INVx1_ASAP7_75t_L g8333 ( 
.A(n_7146),
.Y(n_8333)
);

INVx2_ASAP7_75t_L g8334 ( 
.A(n_8077),
.Y(n_8334)
);

AND2x2_ASAP7_75t_L g8335 ( 
.A(n_7784),
.B(n_6932),
.Y(n_8335)
);

NOR2xp33_ASAP7_75t_L g8336 ( 
.A(n_7661),
.B(n_7339),
.Y(n_8336)
);

BUFx6f_ASAP7_75t_L g8337 ( 
.A(n_7735),
.Y(n_8337)
);

INVx2_ASAP7_75t_L g8338 ( 
.A(n_8077),
.Y(n_8338)
);

HB1xp67_ASAP7_75t_L g8339 ( 
.A(n_8164),
.Y(n_8339)
);

INVx2_ASAP7_75t_L g8340 ( 
.A(n_8077),
.Y(n_8340)
);

BUFx10_ASAP7_75t_L g8341 ( 
.A(n_7815),
.Y(n_8341)
);

AND2x2_ASAP7_75t_L g8342 ( 
.A(n_8136),
.B(n_6967),
.Y(n_8342)
);

INVx2_ASAP7_75t_L g8343 ( 
.A(n_8214),
.Y(n_8343)
);

INVx1_ASAP7_75t_L g8344 ( 
.A(n_7976),
.Y(n_8344)
);

AO21x2_ASAP7_75t_L g8345 ( 
.A1(n_7932),
.A2(n_7765),
.B(n_7725),
.Y(n_8345)
);

INVx2_ASAP7_75t_L g8346 ( 
.A(n_8214),
.Y(n_8346)
);

INVx4_ASAP7_75t_SL g8347 ( 
.A(n_7815),
.Y(n_8347)
);

INVx1_ASAP7_75t_L g8348 ( 
.A(n_7997),
.Y(n_8348)
);

AO21x2_ASAP7_75t_L g8349 ( 
.A1(n_8331),
.A2(n_7115),
.B(n_7413),
.Y(n_8349)
);

INVx1_ASAP7_75t_L g8350 ( 
.A(n_8025),
.Y(n_8350)
);

INVx2_ASAP7_75t_L g8351 ( 
.A(n_8214),
.Y(n_8351)
);

INVx2_ASAP7_75t_L g8352 ( 
.A(n_8302),
.Y(n_8352)
);

INVx2_ASAP7_75t_L g8353 ( 
.A(n_8302),
.Y(n_8353)
);

OA21x2_ASAP7_75t_L g8354 ( 
.A1(n_7665),
.A2(n_7080),
.B(n_7057),
.Y(n_8354)
);

OR2x2_ASAP7_75t_L g8355 ( 
.A(n_8020),
.B(n_8030),
.Y(n_8355)
);

AND2x4_ASAP7_75t_L g8356 ( 
.A(n_8173),
.B(n_6967),
.Y(n_8356)
);

INVx1_ASAP7_75t_SL g8357 ( 
.A(n_7735),
.Y(n_8357)
);

INVx2_ASAP7_75t_L g8358 ( 
.A(n_8302),
.Y(n_8358)
);

OA21x2_ASAP7_75t_L g8359 ( 
.A1(n_7632),
.A2(n_7080),
.B(n_7057),
.Y(n_8359)
);

AND2x2_ASAP7_75t_L g8360 ( 
.A(n_8136),
.B(n_7015),
.Y(n_8360)
);

INVx1_ASAP7_75t_L g8361 ( 
.A(n_7754),
.Y(n_8361)
);

INVx2_ASAP7_75t_L g8362 ( 
.A(n_8093),
.Y(n_8362)
);

OR2x2_ASAP7_75t_L g8363 ( 
.A(n_8067),
.B(n_8015),
.Y(n_8363)
);

INVx2_ASAP7_75t_L g8364 ( 
.A(n_8093),
.Y(n_8364)
);

HB1xp67_ASAP7_75t_L g8365 ( 
.A(n_8131),
.Y(n_8365)
);

INVx2_ASAP7_75t_L g8366 ( 
.A(n_8093),
.Y(n_8366)
);

INVx2_ASAP7_75t_L g8367 ( 
.A(n_8093),
.Y(n_8367)
);

OR2x2_ASAP7_75t_L g8368 ( 
.A(n_8137),
.B(n_7271),
.Y(n_8368)
);

INVx2_ASAP7_75t_L g8369 ( 
.A(n_8101),
.Y(n_8369)
);

INVx3_ASAP7_75t_L g8370 ( 
.A(n_8173),
.Y(n_8370)
);

HB1xp67_ASAP7_75t_L g8371 ( 
.A(n_8082),
.Y(n_8371)
);

OAI21x1_ASAP7_75t_L g8372 ( 
.A1(n_7900),
.A2(n_7115),
.B(n_7053),
.Y(n_8372)
);

NAND2xp5_ASAP7_75t_L g8373 ( 
.A(n_7704),
.B(n_7271),
.Y(n_8373)
);

INVx1_ASAP7_75t_SL g8374 ( 
.A(n_7643),
.Y(n_8374)
);

INVx2_ASAP7_75t_L g8375 ( 
.A(n_8101),
.Y(n_8375)
);

INVx1_ASAP7_75t_L g8376 ( 
.A(n_7754),
.Y(n_8376)
);

AO21x2_ASAP7_75t_L g8377 ( 
.A1(n_8331),
.A2(n_7413),
.B(n_7320),
.Y(n_8377)
);

INVx1_ASAP7_75t_L g8378 ( 
.A(n_7769),
.Y(n_8378)
);

AND2x2_ASAP7_75t_L g8379 ( 
.A(n_8183),
.B(n_7991),
.Y(n_8379)
);

INVx2_ASAP7_75t_L g8380 ( 
.A(n_8101),
.Y(n_8380)
);

INVx3_ASAP7_75t_L g8381 ( 
.A(n_8173),
.Y(n_8381)
);

NOR2xp33_ASAP7_75t_L g8382 ( 
.A(n_7752),
.B(n_7528),
.Y(n_8382)
);

AO21x2_ASAP7_75t_L g8383 ( 
.A1(n_7748),
.A2(n_7320),
.B(n_7295),
.Y(n_8383)
);

INVx2_ASAP7_75t_L g8384 ( 
.A(n_8101),
.Y(n_8384)
);

INVx1_ASAP7_75t_L g8385 ( 
.A(n_7769),
.Y(n_8385)
);

INVx1_ASAP7_75t_L g8386 ( 
.A(n_7770),
.Y(n_8386)
);

AND2x2_ASAP7_75t_L g8387 ( 
.A(n_8183),
.B(n_7015),
.Y(n_8387)
);

AO21x2_ASAP7_75t_L g8388 ( 
.A1(n_8004),
.A2(n_7295),
.B(n_7491),
.Y(n_8388)
);

AND2x2_ASAP7_75t_L g8389 ( 
.A(n_7991),
.B(n_7331),
.Y(n_8389)
);

INVxp67_ASAP7_75t_L g8390 ( 
.A(n_7772),
.Y(n_8390)
);

NAND2xp5_ASAP7_75t_L g8391 ( 
.A(n_7810),
.B(n_7639),
.Y(n_8391)
);

AND2x2_ASAP7_75t_L g8392 ( 
.A(n_7991),
.B(n_7331),
.Y(n_8392)
);

AND2x4_ASAP7_75t_L g8393 ( 
.A(n_8182),
.B(n_7331),
.Y(n_8393)
);

OR2x2_ASAP7_75t_L g8394 ( 
.A(n_7744),
.B(n_7271),
.Y(n_8394)
);

INVx2_ASAP7_75t_L g8395 ( 
.A(n_8101),
.Y(n_8395)
);

NOR2xp33_ASAP7_75t_L g8396 ( 
.A(n_7766),
.B(n_7528),
.Y(n_8396)
);

OR2x2_ASAP7_75t_L g8397 ( 
.A(n_8099),
.B(n_7271),
.Y(n_8397)
);

NAND2xp5_ASAP7_75t_L g8398 ( 
.A(n_7745),
.B(n_7271),
.Y(n_8398)
);

INVx1_ASAP7_75t_L g8399 ( 
.A(n_7770),
.Y(n_8399)
);

INVx2_ASAP7_75t_L g8400 ( 
.A(n_8148),
.Y(n_8400)
);

BUFx2_ASAP7_75t_SL g8401 ( 
.A(n_7643),
.Y(n_8401)
);

INVx2_ASAP7_75t_L g8402 ( 
.A(n_8148),
.Y(n_8402)
);

AND2x4_ASAP7_75t_L g8403 ( 
.A(n_8182),
.B(n_7340),
.Y(n_8403)
);

INVx2_ASAP7_75t_L g8404 ( 
.A(n_8148),
.Y(n_8404)
);

INVx1_ASAP7_75t_L g8405 ( 
.A(n_7909),
.Y(n_8405)
);

AO21x2_ASAP7_75t_L g8406 ( 
.A1(n_7971),
.A2(n_7491),
.B(n_7341),
.Y(n_8406)
);

INVx1_ASAP7_75t_L g8407 ( 
.A(n_7909),
.Y(n_8407)
);

AND2x2_ASAP7_75t_L g8408 ( 
.A(n_8125),
.B(n_7340),
.Y(n_8408)
);

AO21x2_ASAP7_75t_L g8409 ( 
.A1(n_7706),
.A2(n_7491),
.B(n_7341),
.Y(n_8409)
);

INVx1_ASAP7_75t_L g8410 ( 
.A(n_7911),
.Y(n_8410)
);

AND2x2_ASAP7_75t_L g8411 ( 
.A(n_8125),
.B(n_7340),
.Y(n_8411)
);

INVx1_ASAP7_75t_L g8412 ( 
.A(n_7911),
.Y(n_8412)
);

BUFx3_ASAP7_75t_L g8413 ( 
.A(n_7640),
.Y(n_8413)
);

INVx3_ASAP7_75t_L g8414 ( 
.A(n_8182),
.Y(n_8414)
);

HB1xp67_ASAP7_75t_L g8415 ( 
.A(n_7644),
.Y(n_8415)
);

AND2x2_ASAP7_75t_L g8416 ( 
.A(n_8125),
.B(n_7340),
.Y(n_8416)
);

OAI21xp5_ASAP7_75t_L g8417 ( 
.A1(n_7658),
.A2(n_7576),
.B(n_7569),
.Y(n_8417)
);

INVx2_ASAP7_75t_L g8418 ( 
.A(n_8148),
.Y(n_8418)
);

INVx1_ASAP7_75t_L g8419 ( 
.A(n_8022),
.Y(n_8419)
);

INVx1_ASAP7_75t_L g8420 ( 
.A(n_8022),
.Y(n_8420)
);

INVx1_ASAP7_75t_L g8421 ( 
.A(n_8027),
.Y(n_8421)
);

INVx2_ASAP7_75t_L g8422 ( 
.A(n_8148),
.Y(n_8422)
);

NAND2xp5_ASAP7_75t_L g8423 ( 
.A(n_7776),
.B(n_7271),
.Y(n_8423)
);

OA21x2_ASAP7_75t_L g8424 ( 
.A1(n_7694),
.A2(n_7080),
.B(n_7057),
.Y(n_8424)
);

INVx2_ASAP7_75t_L g8425 ( 
.A(n_8179),
.Y(n_8425)
);

BUFx2_ASAP7_75t_L g8426 ( 
.A(n_8044),
.Y(n_8426)
);

NOR2xp33_ASAP7_75t_L g8427 ( 
.A(n_7755),
.B(n_7545),
.Y(n_8427)
);

AO21x1_ASAP7_75t_SL g8428 ( 
.A1(n_7714),
.A2(n_7269),
.B(n_7205),
.Y(n_8428)
);

INVx2_ASAP7_75t_L g8429 ( 
.A(n_8179),
.Y(n_8429)
);

AND2x2_ASAP7_75t_L g8430 ( 
.A(n_8221),
.B(n_7352),
.Y(n_8430)
);

INVx1_ASAP7_75t_L g8431 ( 
.A(n_8027),
.Y(n_8431)
);

AND2x2_ASAP7_75t_L g8432 ( 
.A(n_8221),
.B(n_7352),
.Y(n_8432)
);

INVx1_ASAP7_75t_L g8433 ( 
.A(n_8029),
.Y(n_8433)
);

AND2x2_ASAP7_75t_L g8434 ( 
.A(n_8221),
.B(n_7352),
.Y(n_8434)
);

INVx1_ASAP7_75t_L g8435 ( 
.A(n_8029),
.Y(n_8435)
);

INVx1_ASAP7_75t_SL g8436 ( 
.A(n_7826),
.Y(n_8436)
);

OA21x2_ASAP7_75t_L g8437 ( 
.A1(n_8045),
.A2(n_7102),
.B(n_7083),
.Y(n_8437)
);

INVx2_ASAP7_75t_L g8438 ( 
.A(n_8179),
.Y(n_8438)
);

AO21x2_ASAP7_75t_L g8439 ( 
.A1(n_7729),
.A2(n_7341),
.B(n_7619),
.Y(n_8439)
);

BUFx2_ASAP7_75t_L g8440 ( 
.A(n_8044),
.Y(n_8440)
);

AND2x2_ASAP7_75t_L g8441 ( 
.A(n_8107),
.B(n_7352),
.Y(n_8441)
);

INVx2_ASAP7_75t_SL g8442 ( 
.A(n_7723),
.Y(n_8442)
);

INVx1_ASAP7_75t_L g8443 ( 
.A(n_8037),
.Y(n_8443)
);

INVx1_ASAP7_75t_SL g8444 ( 
.A(n_7826),
.Y(n_8444)
);

INVx2_ASAP7_75t_L g8445 ( 
.A(n_8179),
.Y(n_8445)
);

INVx1_ASAP7_75t_L g8446 ( 
.A(n_8037),
.Y(n_8446)
);

HB1xp67_ASAP7_75t_L g8447 ( 
.A(n_7709),
.Y(n_8447)
);

AO21x2_ASAP7_75t_L g8448 ( 
.A1(n_7751),
.A2(n_7619),
.B(n_7180),
.Y(n_8448)
);

INVx1_ASAP7_75t_L g8449 ( 
.A(n_8139),
.Y(n_8449)
);

INVx2_ASAP7_75t_L g8450 ( 
.A(n_8179),
.Y(n_8450)
);

AND2x2_ASAP7_75t_L g8451 ( 
.A(n_8107),
.B(n_7399),
.Y(n_8451)
);

INVx1_ASAP7_75t_L g8452 ( 
.A(n_8139),
.Y(n_8452)
);

INVx1_ASAP7_75t_L g8453 ( 
.A(n_8159),
.Y(n_8453)
);

INVx1_ASAP7_75t_L g8454 ( 
.A(n_8159),
.Y(n_8454)
);

INVx1_ASAP7_75t_L g8455 ( 
.A(n_8233),
.Y(n_8455)
);

AND2x2_ASAP7_75t_L g8456 ( 
.A(n_8126),
.B(n_7399),
.Y(n_8456)
);

OR2x6_ASAP7_75t_L g8457 ( 
.A(n_7637),
.B(n_7508),
.Y(n_8457)
);

AND2x2_ASAP7_75t_L g8458 ( 
.A(n_8126),
.B(n_7399),
.Y(n_8458)
);

BUFx3_ASAP7_75t_L g8459 ( 
.A(n_7640),
.Y(n_8459)
);

INVx2_ASAP7_75t_L g8460 ( 
.A(n_7683),
.Y(n_8460)
);

INVx1_ASAP7_75t_L g8461 ( 
.A(n_8233),
.Y(n_8461)
);

OR2x2_ASAP7_75t_L g8462 ( 
.A(n_8114),
.B(n_7330),
.Y(n_8462)
);

INVx4_ASAP7_75t_L g8463 ( 
.A(n_7759),
.Y(n_8463)
);

INVx1_ASAP7_75t_L g8464 ( 
.A(n_8235),
.Y(n_8464)
);

INVx2_ASAP7_75t_L g8465 ( 
.A(n_7683),
.Y(n_8465)
);

INVx1_ASAP7_75t_L g8466 ( 
.A(n_8235),
.Y(n_8466)
);

AND2x2_ASAP7_75t_L g8467 ( 
.A(n_8142),
.B(n_7399),
.Y(n_8467)
);

INVx2_ASAP7_75t_L g8468 ( 
.A(n_7701),
.Y(n_8468)
);

BUFx4f_ASAP7_75t_SL g8469 ( 
.A(n_7832),
.Y(n_8469)
);

AOI21xp5_ASAP7_75t_L g8470 ( 
.A1(n_7656),
.A2(n_7284),
.B(n_7619),
.Y(n_8470)
);

AND2x2_ASAP7_75t_L g8471 ( 
.A(n_8142),
.B(n_7430),
.Y(n_8471)
);

OR2x2_ASAP7_75t_L g8472 ( 
.A(n_7818),
.B(n_7330),
.Y(n_8472)
);

INVx1_ASAP7_75t_L g8473 ( 
.A(n_8333),
.Y(n_8473)
);

AND2x2_ASAP7_75t_L g8474 ( 
.A(n_8147),
.B(n_7430),
.Y(n_8474)
);

INVx2_ASAP7_75t_L g8475 ( 
.A(n_7701),
.Y(n_8475)
);

BUFx3_ASAP7_75t_L g8476 ( 
.A(n_7640),
.Y(n_8476)
);

AND2x2_ASAP7_75t_L g8477 ( 
.A(n_8147),
.B(n_7430),
.Y(n_8477)
);

AO21x2_ASAP7_75t_L g8478 ( 
.A1(n_8009),
.A2(n_7180),
.B(n_7058),
.Y(n_8478)
);

BUFx6f_ASAP7_75t_L g8479 ( 
.A(n_7755),
.Y(n_8479)
);

OR2x6_ASAP7_75t_L g8480 ( 
.A(n_7637),
.B(n_7508),
.Y(n_8480)
);

INVx1_ASAP7_75t_L g8481 ( 
.A(n_8333),
.Y(n_8481)
);

AOI22xp33_ASAP7_75t_L g8482 ( 
.A1(n_7721),
.A2(n_7284),
.B1(n_7062),
.B2(n_7110),
.Y(n_8482)
);

INVx2_ASAP7_75t_L g8483 ( 
.A(n_7713),
.Y(n_8483)
);

AND2x2_ASAP7_75t_L g8484 ( 
.A(n_8181),
.B(n_7430),
.Y(n_8484)
);

BUFx3_ASAP7_75t_L g8485 ( 
.A(n_7670),
.Y(n_8485)
);

INVx1_ASAP7_75t_L g8486 ( 
.A(n_7659),
.Y(n_8486)
);

BUFx2_ASAP7_75t_L g8487 ( 
.A(n_8087),
.Y(n_8487)
);

AND2x2_ASAP7_75t_L g8488 ( 
.A(n_8181),
.B(n_7432),
.Y(n_8488)
);

BUFx6f_ASAP7_75t_L g8489 ( 
.A(n_7782),
.Y(n_8489)
);

AND2x2_ASAP7_75t_L g8490 ( 
.A(n_8202),
.B(n_7432),
.Y(n_8490)
);

INVx2_ASAP7_75t_SL g8491 ( 
.A(n_7723),
.Y(n_8491)
);

INVx1_ASAP7_75t_L g8492 ( 
.A(n_7680),
.Y(n_8492)
);

INVx1_ASAP7_75t_L g8493 ( 
.A(n_7692),
.Y(n_8493)
);

BUFx6f_ASAP7_75t_L g8494 ( 
.A(n_7782),
.Y(n_8494)
);

AO21x2_ASAP7_75t_L g8495 ( 
.A1(n_8184),
.A2(n_7058),
.B(n_7083),
.Y(n_8495)
);

INVx1_ASAP7_75t_L g8496 ( 
.A(n_7698),
.Y(n_8496)
);

INVx3_ASAP7_75t_L g8497 ( 
.A(n_7649),
.Y(n_8497)
);

INVx3_ASAP7_75t_L g8498 ( 
.A(n_7649),
.Y(n_8498)
);

AO21x2_ASAP7_75t_L g8499 ( 
.A1(n_8212),
.A2(n_7102),
.B(n_7083),
.Y(n_8499)
);

INVx2_ASAP7_75t_L g8500 ( 
.A(n_7713),
.Y(n_8500)
);

INVx1_ASAP7_75t_L g8501 ( 
.A(n_7707),
.Y(n_8501)
);

HB1xp67_ASAP7_75t_L g8502 ( 
.A(n_7829),
.Y(n_8502)
);

OR2x2_ASAP7_75t_L g8503 ( 
.A(n_7898),
.B(n_7330),
.Y(n_8503)
);

BUFx2_ASAP7_75t_L g8504 ( 
.A(n_8087),
.Y(n_8504)
);

INVx4_ASAP7_75t_L g8505 ( 
.A(n_7759),
.Y(n_8505)
);

INVx2_ASAP7_75t_L g8506 ( 
.A(n_7900),
.Y(n_8506)
);

INVx1_ASAP7_75t_L g8507 ( 
.A(n_7712),
.Y(n_8507)
);

INVx1_ASAP7_75t_L g8508 ( 
.A(n_7719),
.Y(n_8508)
);

OR2x2_ASAP7_75t_L g8509 ( 
.A(n_7947),
.B(n_6822),
.Y(n_8509)
);

HB1xp67_ASAP7_75t_L g8510 ( 
.A(n_8240),
.Y(n_8510)
);

BUFx3_ASAP7_75t_L g8511 ( 
.A(n_7670),
.Y(n_8511)
);

INVxp67_ASAP7_75t_SL g8512 ( 
.A(n_8019),
.Y(n_8512)
);

INVx1_ASAP7_75t_L g8513 ( 
.A(n_7738),
.Y(n_8513)
);

NOR2xp33_ASAP7_75t_SL g8514 ( 
.A(n_7675),
.B(n_7545),
.Y(n_8514)
);

HB1xp67_ASAP7_75t_L g8515 ( 
.A(n_8249),
.Y(n_8515)
);

OR2x2_ASAP7_75t_L g8516 ( 
.A(n_8285),
.B(n_6822),
.Y(n_8516)
);

INVx3_ASAP7_75t_L g8517 ( 
.A(n_7649),
.Y(n_8517)
);

OA21x2_ASAP7_75t_L g8518 ( 
.A1(n_8196),
.A2(n_7128),
.B(n_7102),
.Y(n_8518)
);

INVx1_ASAP7_75t_L g8519 ( 
.A(n_7739),
.Y(n_8519)
);

NOR2xp33_ASAP7_75t_L g8520 ( 
.A(n_7678),
.B(n_7537),
.Y(n_8520)
);

INVx2_ASAP7_75t_SL g8521 ( 
.A(n_7723),
.Y(n_8521)
);

BUFx2_ASAP7_75t_L g8522 ( 
.A(n_7832),
.Y(n_8522)
);

INVx1_ASAP7_75t_L g8523 ( 
.A(n_7747),
.Y(n_8523)
);

INVx1_ASAP7_75t_L g8524 ( 
.A(n_7786),
.Y(n_8524)
);

INVx1_ASAP7_75t_L g8525 ( 
.A(n_7787),
.Y(n_8525)
);

INVx2_ASAP7_75t_L g8526 ( 
.A(n_8171),
.Y(n_8526)
);

OR2x2_ASAP7_75t_L g8527 ( 
.A(n_8320),
.B(n_6822),
.Y(n_8527)
);

INVx1_ASAP7_75t_L g8528 ( 
.A(n_7791),
.Y(n_8528)
);

INVx1_ASAP7_75t_L g8529 ( 
.A(n_7795),
.Y(n_8529)
);

INVx1_ASAP7_75t_L g8530 ( 
.A(n_7804),
.Y(n_8530)
);

INVx1_ASAP7_75t_L g8531 ( 
.A(n_7814),
.Y(n_8531)
);

INVx2_ASAP7_75t_L g8532 ( 
.A(n_8171),
.Y(n_8532)
);

INVx1_ASAP7_75t_L g8533 ( 
.A(n_7828),
.Y(n_8533)
);

INVx2_ASAP7_75t_L g8534 ( 
.A(n_8208),
.Y(n_8534)
);

AO21x2_ASAP7_75t_L g8535 ( 
.A1(n_8036),
.A2(n_7140),
.B(n_7128),
.Y(n_8535)
);

OAI21x1_ASAP7_75t_L g8536 ( 
.A1(n_8306),
.A2(n_7053),
.B(n_7039),
.Y(n_8536)
);

HB1xp67_ASAP7_75t_L g8537 ( 
.A(n_8327),
.Y(n_8537)
);

OAI33xp33_ASAP7_75t_L g8538 ( 
.A1(n_7778),
.A2(n_7529),
.A3(n_7549),
.B1(n_7532),
.B2(n_7507),
.B3(n_7416),
.Y(n_8538)
);

AND2x2_ASAP7_75t_L g8539 ( 
.A(n_8202),
.B(n_7432),
.Y(n_8539)
);

AND2x2_ASAP7_75t_L g8540 ( 
.A(n_8227),
.B(n_7647),
.Y(n_8540)
);

AND2x4_ASAP7_75t_L g8541 ( 
.A(n_7867),
.B(n_7432),
.Y(n_8541)
);

INVx1_ASAP7_75t_L g8542 ( 
.A(n_7841),
.Y(n_8542)
);

AOI22xp33_ASAP7_75t_L g8543 ( 
.A1(n_7654),
.A2(n_7284),
.B1(n_7062),
.B2(n_7110),
.Y(n_8543)
);

INVx1_ASAP7_75t_L g8544 ( 
.A(n_7856),
.Y(n_8544)
);

OR2x6_ASAP7_75t_L g8545 ( 
.A(n_8069),
.B(n_8086),
.Y(n_8545)
);

OR2x6_ASAP7_75t_L g8546 ( 
.A(n_8069),
.B(n_7537),
.Y(n_8546)
);

INVx1_ASAP7_75t_L g8547 ( 
.A(n_7869),
.Y(n_8547)
);

AND2x2_ASAP7_75t_L g8548 ( 
.A(n_8227),
.B(n_7455),
.Y(n_8548)
);

INVx1_ASAP7_75t_L g8549 ( 
.A(n_7876),
.Y(n_8549)
);

BUFx2_ASAP7_75t_L g8550 ( 
.A(n_7675),
.Y(n_8550)
);

INVx2_ASAP7_75t_L g8551 ( 
.A(n_8208),
.Y(n_8551)
);

BUFx3_ASAP7_75t_L g8552 ( 
.A(n_7720),
.Y(n_8552)
);

BUFx2_ASAP7_75t_L g8553 ( 
.A(n_7720),
.Y(n_8553)
);

INVx1_ASAP7_75t_L g8554 ( 
.A(n_7887),
.Y(n_8554)
);

OR2x2_ASAP7_75t_L g8555 ( 
.A(n_7981),
.B(n_6815),
.Y(n_8555)
);

HB1xp67_ASAP7_75t_L g8556 ( 
.A(n_7808),
.Y(n_8556)
);

INVx1_ASAP7_75t_L g8557 ( 
.A(n_7888),
.Y(n_8557)
);

BUFx3_ASAP7_75t_L g8558 ( 
.A(n_7734),
.Y(n_8558)
);

INVx3_ASAP7_75t_L g8559 ( 
.A(n_7678),
.Y(n_8559)
);

INVx2_ASAP7_75t_L g8560 ( 
.A(n_8238),
.Y(n_8560)
);

OAI21xp5_ASAP7_75t_L g8561 ( 
.A1(n_7753),
.A2(n_7576),
.B(n_7569),
.Y(n_8561)
);

AO21x2_ASAP7_75t_L g8562 ( 
.A1(n_7797),
.A2(n_7140),
.B(n_7128),
.Y(n_8562)
);

INVx2_ASAP7_75t_L g8563 ( 
.A(n_8238),
.Y(n_8563)
);

AND2x2_ASAP7_75t_L g8564 ( 
.A(n_7647),
.B(n_7758),
.Y(n_8564)
);

NAND2xp5_ASAP7_75t_L g8565 ( 
.A(n_8068),
.B(n_7123),
.Y(n_8565)
);

INVx2_ASAP7_75t_L g8566 ( 
.A(n_7994),
.Y(n_8566)
);

INVx1_ASAP7_75t_L g8567 ( 
.A(n_7892),
.Y(n_8567)
);

INVx2_ASAP7_75t_L g8568 ( 
.A(n_7994),
.Y(n_8568)
);

INVx1_ASAP7_75t_L g8569 ( 
.A(n_7923),
.Y(n_8569)
);

AO21x2_ASAP7_75t_L g8570 ( 
.A1(n_7798),
.A2(n_7160),
.B(n_7140),
.Y(n_8570)
);

AO21x2_ASAP7_75t_L g8571 ( 
.A1(n_8011),
.A2(n_7170),
.B(n_7160),
.Y(n_8571)
);

INVx2_ASAP7_75t_L g8572 ( 
.A(n_7790),
.Y(n_8572)
);

AND2x2_ASAP7_75t_L g8573 ( 
.A(n_7647),
.B(n_7455),
.Y(n_8573)
);

AND2x2_ASAP7_75t_L g8574 ( 
.A(n_7758),
.B(n_7455),
.Y(n_8574)
);

INVx2_ASAP7_75t_L g8575 ( 
.A(n_7790),
.Y(n_8575)
);

NAND2xp5_ASAP7_75t_L g8576 ( 
.A(n_7634),
.B(n_7123),
.Y(n_8576)
);

INVx2_ASAP7_75t_SL g8577 ( 
.A(n_7723),
.Y(n_8577)
);

BUFx2_ASAP7_75t_L g8578 ( 
.A(n_7734),
.Y(n_8578)
);

INVx2_ASAP7_75t_L g8579 ( 
.A(n_7895),
.Y(n_8579)
);

INVx2_ASAP7_75t_L g8580 ( 
.A(n_7895),
.Y(n_8580)
);

INVx1_ASAP7_75t_L g8581 ( 
.A(n_7926),
.Y(n_8581)
);

OR2x2_ASAP7_75t_L g8582 ( 
.A(n_7854),
.B(n_6822),
.Y(n_8582)
);

INVx2_ASAP7_75t_L g8583 ( 
.A(n_7906),
.Y(n_8583)
);

INVx1_ASAP7_75t_L g8584 ( 
.A(n_7930),
.Y(n_8584)
);

INVx2_ASAP7_75t_L g8585 ( 
.A(n_7906),
.Y(n_8585)
);

INVx2_ASAP7_75t_L g8586 ( 
.A(n_7915),
.Y(n_8586)
);

INVx1_ASAP7_75t_L g8587 ( 
.A(n_7934),
.Y(n_8587)
);

INVx2_ASAP7_75t_L g8588 ( 
.A(n_7915),
.Y(n_8588)
);

INVx2_ASAP7_75t_L g8589 ( 
.A(n_7957),
.Y(n_8589)
);

AO21x2_ASAP7_75t_L g8590 ( 
.A1(n_7894),
.A2(n_8002),
.B(n_7664),
.Y(n_8590)
);

OA21x2_ASAP7_75t_L g8591 ( 
.A1(n_8332),
.A2(n_7170),
.B(n_7160),
.Y(n_8591)
);

BUFx3_ASAP7_75t_L g8592 ( 
.A(n_7821),
.Y(n_8592)
);

INVx1_ASAP7_75t_L g8593 ( 
.A(n_7936),
.Y(n_8593)
);

AND2x2_ASAP7_75t_L g8594 ( 
.A(n_7758),
.B(n_7951),
.Y(n_8594)
);

INVx5_ASAP7_75t_L g8595 ( 
.A(n_7723),
.Y(n_8595)
);

HB1xp67_ASAP7_75t_L g8596 ( 
.A(n_7867),
.Y(n_8596)
);

INVx2_ASAP7_75t_L g8597 ( 
.A(n_7957),
.Y(n_8597)
);

INVx1_ASAP7_75t_L g8598 ( 
.A(n_7952),
.Y(n_8598)
);

INVx1_ASAP7_75t_L g8599 ( 
.A(n_7955),
.Y(n_8599)
);

INVx2_ASAP7_75t_L g8600 ( 
.A(n_7974),
.Y(n_8600)
);

BUFx2_ASAP7_75t_L g8601 ( 
.A(n_7821),
.Y(n_8601)
);

INVx2_ASAP7_75t_L g8602 ( 
.A(n_7974),
.Y(n_8602)
);

AO21x2_ASAP7_75t_L g8603 ( 
.A1(n_7662),
.A2(n_7172),
.B(n_7170),
.Y(n_8603)
);

INVx1_ASAP7_75t_L g8604 ( 
.A(n_7963),
.Y(n_8604)
);

INVx2_ASAP7_75t_L g8605 ( 
.A(n_8261),
.Y(n_8605)
);

INVxp67_ASAP7_75t_SL g8606 ( 
.A(n_7761),
.Y(n_8606)
);

INVx2_ASAP7_75t_L g8607 ( 
.A(n_8261),
.Y(n_8607)
);

INVx1_ASAP7_75t_L g8608 ( 
.A(n_7975),
.Y(n_8608)
);

NOR3xp33_ASAP7_75t_L g8609 ( 
.A(n_7736),
.B(n_6843),
.C(n_6821),
.Y(n_8609)
);

INVx1_ASAP7_75t_L g8610 ( 
.A(n_7977),
.Y(n_8610)
);

OR2x2_ASAP7_75t_L g8611 ( 
.A(n_8097),
.B(n_6822),
.Y(n_8611)
);

BUFx3_ASAP7_75t_L g8612 ( 
.A(n_7703),
.Y(n_8612)
);

INVx3_ASAP7_75t_L g8613 ( 
.A(n_7678),
.Y(n_8613)
);

INVx2_ASAP7_75t_L g8614 ( 
.A(n_8261),
.Y(n_8614)
);

INVx2_ASAP7_75t_L g8615 ( 
.A(n_7913),
.Y(n_8615)
);

AND2x2_ASAP7_75t_L g8616 ( 
.A(n_7951),
.B(n_7455),
.Y(n_8616)
);

INVx1_ASAP7_75t_L g8617 ( 
.A(n_8000),
.Y(n_8617)
);

NAND2xp5_ASAP7_75t_L g8618 ( 
.A(n_7964),
.B(n_7366),
.Y(n_8618)
);

INVx1_ASAP7_75t_L g8619 ( 
.A(n_8056),
.Y(n_8619)
);

INVxp67_ASAP7_75t_SL g8620 ( 
.A(n_7761),
.Y(n_8620)
);

INVx1_ASAP7_75t_L g8621 ( 
.A(n_8081),
.Y(n_8621)
);

INVx1_ASAP7_75t_L g8622 ( 
.A(n_8098),
.Y(n_8622)
);

INVx2_ASAP7_75t_L g8623 ( 
.A(n_7913),
.Y(n_8623)
);

BUFx3_ASAP7_75t_L g8624 ( 
.A(n_7780),
.Y(n_8624)
);

INVx1_ASAP7_75t_SL g8625 ( 
.A(n_7708),
.Y(n_8625)
);

INVx2_ASAP7_75t_L g8626 ( 
.A(n_7913),
.Y(n_8626)
);

INVx1_ASAP7_75t_L g8627 ( 
.A(n_8100),
.Y(n_8627)
);

BUFx6f_ASAP7_75t_L g8628 ( 
.A(n_7761),
.Y(n_8628)
);

AND2x2_ASAP7_75t_L g8629 ( 
.A(n_7951),
.B(n_7563),
.Y(n_8629)
);

INVx1_ASAP7_75t_L g8630 ( 
.A(n_8119),
.Y(n_8630)
);

OR2x2_ASAP7_75t_L g8631 ( 
.A(n_7858),
.B(n_6815),
.Y(n_8631)
);

AO21x2_ASAP7_75t_L g8632 ( 
.A1(n_7662),
.A2(n_7177),
.B(n_7172),
.Y(n_8632)
);

AND2x2_ASAP7_75t_L g8633 ( 
.A(n_8053),
.B(n_7563),
.Y(n_8633)
);

INVx1_ASAP7_75t_L g8634 ( 
.A(n_8143),
.Y(n_8634)
);

AND2x4_ASAP7_75t_L g8635 ( 
.A(n_7987),
.B(n_7563),
.Y(n_8635)
);

BUFx6f_ASAP7_75t_L g8636 ( 
.A(n_7761),
.Y(n_8636)
);

AND2x2_ASAP7_75t_L g8637 ( 
.A(n_8053),
.B(n_7563),
.Y(n_8637)
);

OR2x2_ASAP7_75t_L g8638 ( 
.A(n_7871),
.B(n_6822),
.Y(n_8638)
);

AND2x4_ASAP7_75t_L g8639 ( 
.A(n_7987),
.B(n_6815),
.Y(n_8639)
);

INVx2_ASAP7_75t_L g8640 ( 
.A(n_7913),
.Y(n_8640)
);

HB1xp67_ASAP7_75t_L g8641 ( 
.A(n_8026),
.Y(n_8641)
);

INVx1_ASAP7_75t_L g8642 ( 
.A(n_8144),
.Y(n_8642)
);

INVx1_ASAP7_75t_L g8643 ( 
.A(n_8146),
.Y(n_8643)
);

OR2x6_ASAP7_75t_L g8644 ( 
.A(n_8086),
.B(n_7537),
.Y(n_8644)
);

INVx2_ASAP7_75t_L g8645 ( 
.A(n_7913),
.Y(n_8645)
);

INVx2_ASAP7_75t_L g8646 ( 
.A(n_7913),
.Y(n_8646)
);

INVx2_ASAP7_75t_SL g8647 ( 
.A(n_7789),
.Y(n_8647)
);

INVx4_ASAP7_75t_L g8648 ( 
.A(n_7958),
.Y(n_8648)
);

NAND2xp5_ASAP7_75t_L g8649 ( 
.A(n_7631),
.B(n_7366),
.Y(n_8649)
);

INVx3_ASAP7_75t_L g8650 ( 
.A(n_7761),
.Y(n_8650)
);

NAND2xp5_ASAP7_75t_L g8651 ( 
.A(n_7757),
.B(n_7366),
.Y(n_8651)
);

BUFx3_ASAP7_75t_L g8652 ( 
.A(n_7794),
.Y(n_8652)
);

HB1xp67_ASAP7_75t_L g8653 ( 
.A(n_8026),
.Y(n_8653)
);

HB1xp67_ASAP7_75t_L g8654 ( 
.A(n_7890),
.Y(n_8654)
);

INVx2_ASAP7_75t_L g8655 ( 
.A(n_7913),
.Y(n_8655)
);

AND2x2_ASAP7_75t_L g8656 ( 
.A(n_8053),
.B(n_6919),
.Y(n_8656)
);

BUFx6f_ASAP7_75t_L g8657 ( 
.A(n_7794),
.Y(n_8657)
);

INVx1_ASAP7_75t_L g8658 ( 
.A(n_8149),
.Y(n_8658)
);

INVx2_ASAP7_75t_L g8659 ( 
.A(n_7789),
.Y(n_8659)
);

INVx3_ASAP7_75t_L g8660 ( 
.A(n_7794),
.Y(n_8660)
);

INVx2_ASAP7_75t_L g8661 ( 
.A(n_7789),
.Y(n_8661)
);

AND2x2_ASAP7_75t_L g8662 ( 
.A(n_8064),
.B(n_6919),
.Y(n_8662)
);

INVx4_ASAP7_75t_L g8663 ( 
.A(n_7958),
.Y(n_8663)
);

INVx1_ASAP7_75t_L g8664 ( 
.A(n_8161),
.Y(n_8664)
);

INVx1_ASAP7_75t_L g8665 ( 
.A(n_8163),
.Y(n_8665)
);

INVx2_ASAP7_75t_L g8666 ( 
.A(n_7789),
.Y(n_8666)
);

INVx1_ASAP7_75t_L g8667 ( 
.A(n_8189),
.Y(n_8667)
);

AND2x2_ASAP7_75t_L g8668 ( 
.A(n_8064),
.B(n_7444),
.Y(n_8668)
);

AND2x4_ASAP7_75t_L g8669 ( 
.A(n_8113),
.B(n_6815),
.Y(n_8669)
);

AND2x2_ASAP7_75t_L g8670 ( 
.A(n_8064),
.B(n_8243),
.Y(n_8670)
);

INVx1_ASAP7_75t_L g8671 ( 
.A(n_8193),
.Y(n_8671)
);

AO21x2_ASAP7_75t_L g8672 ( 
.A1(n_7664),
.A2(n_7177),
.B(n_7172),
.Y(n_8672)
);

INVx1_ASAP7_75t_L g8673 ( 
.A(n_8199),
.Y(n_8673)
);

CKINVDCx20_ASAP7_75t_R g8674 ( 
.A(n_7785),
.Y(n_8674)
);

INVx3_ASAP7_75t_L g8675 ( 
.A(n_7794),
.Y(n_8675)
);

OR2x2_ASAP7_75t_L g8676 ( 
.A(n_7872),
.B(n_7366),
.Y(n_8676)
);

INVx1_ASAP7_75t_L g8677 ( 
.A(n_8204),
.Y(n_8677)
);

INVx2_ASAP7_75t_L g8678 ( 
.A(n_7789),
.Y(n_8678)
);

AND2x2_ASAP7_75t_L g8679 ( 
.A(n_8243),
.B(n_7444),
.Y(n_8679)
);

INVx2_ASAP7_75t_L g8680 ( 
.A(n_8014),
.Y(n_8680)
);

INVx1_ASAP7_75t_L g8681 ( 
.A(n_8210),
.Y(n_8681)
);

BUFx2_ASAP7_75t_L g8682 ( 
.A(n_8299),
.Y(n_8682)
);

INVx2_ASAP7_75t_L g8683 ( 
.A(n_8014),
.Y(n_8683)
);

INVx2_ASAP7_75t_L g8684 ( 
.A(n_8014),
.Y(n_8684)
);

AND2x2_ASAP7_75t_L g8685 ( 
.A(n_8255),
.B(n_7444),
.Y(n_8685)
);

BUFx2_ASAP7_75t_L g8686 ( 
.A(n_8299),
.Y(n_8686)
);

INVx2_ASAP7_75t_L g8687 ( 
.A(n_8014),
.Y(n_8687)
);

AND2x2_ASAP7_75t_L g8688 ( 
.A(n_8255),
.B(n_7444),
.Y(n_8688)
);

OR2x2_ASAP7_75t_L g8689 ( 
.A(n_7880),
.B(n_7366),
.Y(n_8689)
);

INVx1_ASAP7_75t_L g8690 ( 
.A(n_8211),
.Y(n_8690)
);

AND2x2_ASAP7_75t_L g8691 ( 
.A(n_8083),
.B(n_7444),
.Y(n_8691)
);

INVx2_ASAP7_75t_L g8692 ( 
.A(n_8014),
.Y(n_8692)
);

AOI21xp5_ASAP7_75t_SL g8693 ( 
.A1(n_7682),
.A2(n_6815),
.B(n_7576),
.Y(n_8693)
);

AOI22xp5_ASAP7_75t_L g8694 ( 
.A1(n_7762),
.A2(n_7543),
.B1(n_7000),
.B2(n_7110),
.Y(n_8694)
);

NAND2xp5_ASAP7_75t_SL g8695 ( 
.A(n_7635),
.B(n_7537),
.Y(n_8695)
);

BUFx2_ASAP7_75t_L g8696 ( 
.A(n_8299),
.Y(n_8696)
);

AND2x2_ASAP7_75t_L g8697 ( 
.A(n_8083),
.B(n_7444),
.Y(n_8697)
);

INVx1_ASAP7_75t_L g8698 ( 
.A(n_8213),
.Y(n_8698)
);

HB1xp67_ASAP7_75t_L g8699 ( 
.A(n_7890),
.Y(n_8699)
);

INVx1_ASAP7_75t_L g8700 ( 
.A(n_8215),
.Y(n_8700)
);

OAI21x1_ASAP7_75t_L g8701 ( 
.A1(n_8306),
.A2(n_7138),
.B(n_7039),
.Y(n_8701)
);

INVx3_ASAP7_75t_L g8702 ( 
.A(n_7794),
.Y(n_8702)
);

OR2x2_ASAP7_75t_L g8703 ( 
.A(n_7922),
.B(n_7366),
.Y(n_8703)
);

INVx1_ASAP7_75t_L g8704 ( 
.A(n_8229),
.Y(n_8704)
);

OA21x2_ASAP7_75t_L g8705 ( 
.A1(n_7834),
.A2(n_7177),
.B(n_6849),
.Y(n_8705)
);

INVxp33_ASAP7_75t_L g8706 ( 
.A(n_7768),
.Y(n_8706)
);

BUFx2_ASAP7_75t_L g8707 ( 
.A(n_8209),
.Y(n_8707)
);

INVx1_ASAP7_75t_L g8708 ( 
.A(n_8237),
.Y(n_8708)
);

AOI22xp33_ASAP7_75t_L g8709 ( 
.A1(n_7638),
.A2(n_7062),
.B1(n_7328),
.B2(n_7121),
.Y(n_8709)
);

INVx1_ASAP7_75t_L g8710 ( 
.A(n_8251),
.Y(n_8710)
);

INVx1_ASAP7_75t_L g8711 ( 
.A(n_8253),
.Y(n_8711)
);

INVx1_ASAP7_75t_L g8712 ( 
.A(n_8297),
.Y(n_8712)
);

BUFx6f_ASAP7_75t_L g8713 ( 
.A(n_7857),
.Y(n_8713)
);

INVx1_ASAP7_75t_SL g8714 ( 
.A(n_7708),
.Y(n_8714)
);

INVx1_ASAP7_75t_L g8715 ( 
.A(n_8308),
.Y(n_8715)
);

BUFx3_ASAP7_75t_L g8716 ( 
.A(n_7671),
.Y(n_8716)
);

AND2x2_ASAP7_75t_L g8717 ( 
.A(n_8222),
.B(n_7540),
.Y(n_8717)
);

INVx2_ASAP7_75t_L g8718 ( 
.A(n_8041),
.Y(n_8718)
);

INVx2_ASAP7_75t_L g8719 ( 
.A(n_8041),
.Y(n_8719)
);

BUFx2_ASAP7_75t_L g8720 ( 
.A(n_8209),
.Y(n_8720)
);

AO21x2_ASAP7_75t_L g8721 ( 
.A1(n_7717),
.A2(n_6849),
.B(n_7138),
.Y(n_8721)
);

AO21x2_ASAP7_75t_L g8722 ( 
.A1(n_7717),
.A2(n_7144),
.B(n_7536),
.Y(n_8722)
);

NAND2xp5_ASAP7_75t_L g8723 ( 
.A(n_7792),
.B(n_7395),
.Y(n_8723)
);

BUFx2_ASAP7_75t_L g8724 ( 
.A(n_8113),
.Y(n_8724)
);

AOI33xp33_ASAP7_75t_L g8725 ( 
.A1(n_7666),
.A2(n_7705),
.A3(n_7700),
.B1(n_7879),
.B2(n_7687),
.B3(n_7645),
.Y(n_8725)
);

NAND2xp5_ASAP7_75t_L g8726 ( 
.A(n_7750),
.B(n_7395),
.Y(n_8726)
);

AND2x2_ASAP7_75t_L g8727 ( 
.A(n_8276),
.B(n_7540),
.Y(n_8727)
);

INVx1_ASAP7_75t_L g8728 ( 
.A(n_8310),
.Y(n_8728)
);

NAND2xp5_ASAP7_75t_L g8729 ( 
.A(n_7767),
.B(n_7395),
.Y(n_8729)
);

INVx2_ASAP7_75t_L g8730 ( 
.A(n_8041),
.Y(n_8730)
);

OA21x2_ASAP7_75t_L g8731 ( 
.A1(n_8289),
.A2(n_7536),
.B(n_6955),
.Y(n_8731)
);

INVx1_ASAP7_75t_L g8732 ( 
.A(n_8322),
.Y(n_8732)
);

OR2x6_ASAP7_75t_L g8733 ( 
.A(n_8117),
.B(n_7690),
.Y(n_8733)
);

INVx2_ASAP7_75t_L g8734 ( 
.A(n_8041),
.Y(n_8734)
);

BUFx2_ASAP7_75t_L g8735 ( 
.A(n_8117),
.Y(n_8735)
);

INVx1_ASAP7_75t_L g8736 ( 
.A(n_8326),
.Y(n_8736)
);

OR2x2_ASAP7_75t_L g8737 ( 
.A(n_7924),
.B(n_7395),
.Y(n_8737)
);

AND2x2_ASAP7_75t_L g8738 ( 
.A(n_8276),
.B(n_7542),
.Y(n_8738)
);

AND2x2_ASAP7_75t_L g8739 ( 
.A(n_7883),
.B(n_7542),
.Y(n_8739)
);

INVx2_ASAP7_75t_L g8740 ( 
.A(n_8041),
.Y(n_8740)
);

INVx2_ASAP7_75t_L g8741 ( 
.A(n_8194),
.Y(n_8741)
);

AND2x2_ASAP7_75t_L g8742 ( 
.A(n_8157),
.B(n_7537),
.Y(n_8742)
);

AND2x4_ASAP7_75t_L g8743 ( 
.A(n_7816),
.B(n_6821),
.Y(n_8743)
);

HB1xp67_ASAP7_75t_L g8744 ( 
.A(n_8156),
.Y(n_8744)
);

NAND2xp5_ASAP7_75t_L g8745 ( 
.A(n_7630),
.B(n_7395),
.Y(n_8745)
);

INVxp67_ASAP7_75t_L g8746 ( 
.A(n_7815),
.Y(n_8746)
);

AND2x2_ASAP7_75t_L g8747 ( 
.A(n_8124),
.B(n_7607),
.Y(n_8747)
);

AND2x2_ASAP7_75t_L g8748 ( 
.A(n_8124),
.B(n_7607),
.Y(n_8748)
);

INVx1_ASAP7_75t_L g8749 ( 
.A(n_8156),
.Y(n_8749)
);

OAI21x1_ASAP7_75t_L g8750 ( 
.A1(n_8306),
.A2(n_7144),
.B(n_6933),
.Y(n_8750)
);

INVx1_ASAP7_75t_L g8751 ( 
.A(n_8325),
.Y(n_8751)
);

INVx11_ASAP7_75t_L g8752 ( 
.A(n_8247),
.Y(n_8752)
);

AOI21x1_ASAP7_75t_L g8753 ( 
.A1(n_8223),
.A2(n_7282),
.B(n_7001),
.Y(n_8753)
);

HB1xp67_ASAP7_75t_L g8754 ( 
.A(n_7636),
.Y(n_8754)
);

AND2x4_ASAP7_75t_L g8755 ( 
.A(n_7816),
.B(n_8194),
.Y(n_8755)
);

OR2x2_ASAP7_75t_L g8756 ( 
.A(n_7805),
.B(n_7395),
.Y(n_8756)
);

AND2x2_ASAP7_75t_L g8757 ( 
.A(n_7636),
.B(n_7607),
.Y(n_8757)
);

OR2x2_ASAP7_75t_L g8758 ( 
.A(n_7838),
.B(n_7095),
.Y(n_8758)
);

AO21x2_ASAP7_75t_L g8759 ( 
.A1(n_8034),
.A2(n_7354),
.B(n_7122),
.Y(n_8759)
);

AND2x4_ASAP7_75t_L g8760 ( 
.A(n_7816),
.B(n_6821),
.Y(n_8760)
);

AO21x2_ASAP7_75t_L g8761 ( 
.A1(n_8034),
.A2(n_7354),
.B(n_7122),
.Y(n_8761)
);

BUFx6f_ASAP7_75t_L g8762 ( 
.A(n_7857),
.Y(n_8762)
);

HB1xp67_ASAP7_75t_L g8763 ( 
.A(n_7641),
.Y(n_8763)
);

NAND2xp5_ASAP7_75t_SL g8764 ( 
.A(n_7702),
.B(n_7650),
.Y(n_8764)
);

INVx1_ASAP7_75t_L g8765 ( 
.A(n_8040),
.Y(n_8765)
);

AO21x2_ASAP7_75t_L g8766 ( 
.A1(n_8040),
.A2(n_7354),
.B(n_7122),
.Y(n_8766)
);

INVx1_ASAP7_75t_L g8767 ( 
.A(n_8058),
.Y(n_8767)
);

INVx2_ASAP7_75t_L g8768 ( 
.A(n_8194),
.Y(n_8768)
);

INVx1_ASAP7_75t_L g8769 ( 
.A(n_8058),
.Y(n_8769)
);

NAND2xp5_ASAP7_75t_L g8770 ( 
.A(n_8170),
.B(n_6845),
.Y(n_8770)
);

AO21x2_ASAP7_75t_L g8771 ( 
.A1(n_8287),
.A2(n_7121),
.B(n_7404),
.Y(n_8771)
);

BUFx2_ASAP7_75t_L g8772 ( 
.A(n_7711),
.Y(n_8772)
);

AOI31xp33_ASAP7_75t_L g8773 ( 
.A1(n_7726),
.A2(n_7584),
.A3(n_6931),
.B(n_6917),
.Y(n_8773)
);

INVx2_ASAP7_75t_SL g8774 ( 
.A(n_8194),
.Y(n_8774)
);

AND2x2_ASAP7_75t_L g8775 ( 
.A(n_7641),
.B(n_7607),
.Y(n_8775)
);

OA21x2_ASAP7_75t_L g8776 ( 
.A1(n_8294),
.A2(n_6955),
.B(n_7216),
.Y(n_8776)
);

OAI21x1_ASAP7_75t_L g8777 ( 
.A1(n_8010),
.A2(n_7229),
.B(n_7096),
.Y(n_8777)
);

AND2x4_ASAP7_75t_L g8778 ( 
.A(n_7816),
.B(n_6821),
.Y(n_8778)
);

INVxp67_ASAP7_75t_SL g8779 ( 
.A(n_7633),
.Y(n_8779)
);

OR2x2_ASAP7_75t_L g8780 ( 
.A(n_7946),
.B(n_7620),
.Y(n_8780)
);

HB1xp67_ASAP7_75t_L g8781 ( 
.A(n_7681),
.Y(n_8781)
);

INVx2_ASAP7_75t_L g8782 ( 
.A(n_8194),
.Y(n_8782)
);

OAI21x1_ASAP7_75t_L g8783 ( 
.A1(n_8300),
.A2(n_7229),
.B(n_7096),
.Y(n_8783)
);

AND2x2_ASAP7_75t_L g8784 ( 
.A(n_7681),
.B(n_7607),
.Y(n_8784)
);

HB1xp67_ASAP7_75t_L g8785 ( 
.A(n_7673),
.Y(n_8785)
);

INVx2_ASAP7_75t_L g8786 ( 
.A(n_7673),
.Y(n_8786)
);

INVx2_ASAP7_75t_L g8787 ( 
.A(n_7742),
.Y(n_8787)
);

INVx2_ASAP7_75t_L g8788 ( 
.A(n_7742),
.Y(n_8788)
);

HB1xp67_ASAP7_75t_L g8789 ( 
.A(n_7902),
.Y(n_8789)
);

OR2x6_ASAP7_75t_L g8790 ( 
.A(n_7690),
.B(n_7584),
.Y(n_8790)
);

INVx1_ASAP7_75t_L g8791 ( 
.A(n_8328),
.Y(n_8791)
);

INVx2_ASAP7_75t_SL g8792 ( 
.A(n_7690),
.Y(n_8792)
);

INVx1_ASAP7_75t_L g8793 ( 
.A(n_8328),
.Y(n_8793)
);

INVx2_ASAP7_75t_L g8794 ( 
.A(n_7902),
.Y(n_8794)
);

AND2x2_ASAP7_75t_L g8795 ( 
.A(n_8264),
.B(n_6828),
.Y(n_8795)
);

INVx1_ASAP7_75t_L g8796 ( 
.A(n_7908),
.Y(n_8796)
);

INVx1_ASAP7_75t_L g8797 ( 
.A(n_7908),
.Y(n_8797)
);

BUFx6f_ASAP7_75t_L g8798 ( 
.A(n_7857),
.Y(n_8798)
);

INVx1_ASAP7_75t_L g8799 ( 
.A(n_8059),
.Y(n_8799)
);

INVx1_ASAP7_75t_L g8800 ( 
.A(n_8059),
.Y(n_8800)
);

AO21x2_ASAP7_75t_L g8801 ( 
.A1(n_8160),
.A2(n_7121),
.B(n_7404),
.Y(n_8801)
);

INVx1_ASAP7_75t_L g8802 ( 
.A(n_8129),
.Y(n_8802)
);

AND2x2_ASAP7_75t_L g8803 ( 
.A(n_8273),
.B(n_6828),
.Y(n_8803)
);

INVx1_ASAP7_75t_L g8804 ( 
.A(n_8129),
.Y(n_8804)
);

INVx2_ASAP7_75t_L g8805 ( 
.A(n_7918),
.Y(n_8805)
);

NAND2xp5_ASAP7_75t_SL g8806 ( 
.A(n_7956),
.B(n_7584),
.Y(n_8806)
);

INVx2_ASAP7_75t_SL g8807 ( 
.A(n_7690),
.Y(n_8807)
);

INVx1_ASAP7_75t_L g8808 ( 
.A(n_8134),
.Y(n_8808)
);

OAI22xp5_ASAP7_75t_L g8809 ( 
.A1(n_7669),
.A2(n_6931),
.B1(n_7507),
.B2(n_7416),
.Y(n_8809)
);

INVx3_ASAP7_75t_SL g8810 ( 
.A(n_7711),
.Y(n_8810)
);

AO21x2_ASAP7_75t_L g8811 ( 
.A1(n_7891),
.A2(n_7404),
.B(n_6836),
.Y(n_8811)
);

HB1xp67_ASAP7_75t_L g8812 ( 
.A(n_8013),
.Y(n_8812)
);

OA21x2_ASAP7_75t_L g8813 ( 
.A1(n_7733),
.A2(n_7233),
.B(n_7216),
.Y(n_8813)
);

AND2x4_ASAP7_75t_L g8814 ( 
.A(n_8089),
.B(n_6843),
.Y(n_8814)
);

INVx2_ASAP7_75t_L g8815 ( 
.A(n_7918),
.Y(n_8815)
);

OAI21xp5_ASAP7_75t_L g8816 ( 
.A1(n_7862),
.A2(n_7279),
.B(n_7466),
.Y(n_8816)
);

INVx2_ASAP7_75t_SL g8817 ( 
.A(n_8305),
.Y(n_8817)
);

HB1xp67_ASAP7_75t_L g8818 ( 
.A(n_8013),
.Y(n_8818)
);

AND2x4_ASAP7_75t_L g8819 ( 
.A(n_8089),
.B(n_6843),
.Y(n_8819)
);

OA21x2_ASAP7_75t_L g8820 ( 
.A1(n_8205),
.A2(n_7233),
.B(n_7216),
.Y(n_8820)
);

NAND2xp5_ASAP7_75t_L g8821 ( 
.A(n_8236),
.B(n_6845),
.Y(n_8821)
);

INVx2_ASAP7_75t_L g8822 ( 
.A(n_7920),
.Y(n_8822)
);

OR2x6_ASAP7_75t_L g8823 ( 
.A(n_8223),
.B(n_6843),
.Y(n_8823)
);

NAND2xp5_ASAP7_75t_L g8824 ( 
.A(n_7660),
.B(n_7308),
.Y(n_8824)
);

INVxp67_ASAP7_75t_L g8825 ( 
.A(n_8042),
.Y(n_8825)
);

AOI21xp5_ASAP7_75t_SL g8826 ( 
.A1(n_7777),
.A2(n_7063),
.B(n_7043),
.Y(n_8826)
);

OA21x2_ASAP7_75t_L g8827 ( 
.A1(n_8216),
.A2(n_7234),
.B(n_7233),
.Y(n_8827)
);

HB1xp67_ASAP7_75t_L g8828 ( 
.A(n_8016),
.Y(n_8828)
);

BUFx2_ASAP7_75t_L g8829 ( 
.A(n_7727),
.Y(n_8829)
);

BUFx6f_ASAP7_75t_L g8830 ( 
.A(n_7857),
.Y(n_8830)
);

INVx2_ASAP7_75t_SL g8831 ( 
.A(n_8305),
.Y(n_8831)
);

HB1xp67_ASAP7_75t_L g8832 ( 
.A(n_8016),
.Y(n_8832)
);

INVx1_ASAP7_75t_L g8833 ( 
.A(n_8134),
.Y(n_8833)
);

AND2x4_ASAP7_75t_L g8834 ( 
.A(n_8024),
.B(n_6916),
.Y(n_8834)
);

BUFx2_ASAP7_75t_L g8835 ( 
.A(n_7727),
.Y(n_8835)
);

HB1xp67_ASAP7_75t_L g8836 ( 
.A(n_8324),
.Y(n_8836)
);

NAND2xp5_ASAP7_75t_L g8837 ( 
.A(n_7801),
.B(n_8103),
.Y(n_8837)
);

INVx1_ASAP7_75t_L g8838 ( 
.A(n_8138),
.Y(n_8838)
);

INVx1_ASAP7_75t_L g8839 ( 
.A(n_8138),
.Y(n_8839)
);

BUFx2_ASAP7_75t_L g8840 ( 
.A(n_7823),
.Y(n_8840)
);

OA21x2_ASAP7_75t_L g8841 ( 
.A1(n_8198),
.A2(n_7235),
.B(n_7234),
.Y(n_8841)
);

AO21x2_ASAP7_75t_L g8842 ( 
.A1(n_8232),
.A2(n_6836),
.B(n_6835),
.Y(n_8842)
);

NAND2xp5_ASAP7_75t_L g8843 ( 
.A(n_8043),
.B(n_7308),
.Y(n_8843)
);

OAI21xp5_ASAP7_75t_SL g8844 ( 
.A1(n_7919),
.A2(n_6931),
.B(n_7466),
.Y(n_8844)
);

INVx1_ASAP7_75t_L g8845 ( 
.A(n_8155),
.Y(n_8845)
);

OR2x2_ASAP7_75t_L g8846 ( 
.A(n_8070),
.B(n_7481),
.Y(n_8846)
);

NAND2xp5_ASAP7_75t_L g8847 ( 
.A(n_8032),
.B(n_7308),
.Y(n_8847)
);

INVx1_ASAP7_75t_L g8848 ( 
.A(n_8155),
.Y(n_8848)
);

INVx2_ASAP7_75t_L g8849 ( 
.A(n_7920),
.Y(n_8849)
);

AO21x2_ASAP7_75t_L g8850 ( 
.A1(n_8063),
.A2(n_6836),
.B(n_6835),
.Y(n_8850)
);

INVx2_ASAP7_75t_L g8851 ( 
.A(n_7931),
.Y(n_8851)
);

OR2x2_ASAP7_75t_L g8852 ( 
.A(n_7699),
.B(n_7693),
.Y(n_8852)
);

AO21x2_ASAP7_75t_L g8853 ( 
.A1(n_7695),
.A2(n_6846),
.B(n_6835),
.Y(n_8853)
);

INVx1_ASAP7_75t_L g8854 ( 
.A(n_8158),
.Y(n_8854)
);

AND2x4_ASAP7_75t_L g8855 ( 
.A(n_8187),
.B(n_8094),
.Y(n_8855)
);

AO21x2_ASAP7_75t_L g8856 ( 
.A1(n_8319),
.A2(n_6868),
.B(n_6846),
.Y(n_8856)
);

OA21x2_ASAP7_75t_L g8857 ( 
.A1(n_8158),
.A2(n_7235),
.B(n_7234),
.Y(n_8857)
);

INVx2_ASAP7_75t_L g8858 ( 
.A(n_7931),
.Y(n_8858)
);

INVx1_ASAP7_75t_L g8859 ( 
.A(n_8176),
.Y(n_8859)
);

INVx2_ASAP7_75t_L g8860 ( 
.A(n_7937),
.Y(n_8860)
);

AOI21x1_ASAP7_75t_L g8861 ( 
.A1(n_8246),
.A2(n_6946),
.B(n_7025),
.Y(n_8861)
);

INVx1_ASAP7_75t_L g8862 ( 
.A(n_8176),
.Y(n_8862)
);

AND2x2_ASAP7_75t_L g8863 ( 
.A(n_8305),
.B(n_6842),
.Y(n_8863)
);

INVx1_ASAP7_75t_L g8864 ( 
.A(n_8177),
.Y(n_8864)
);

AND2x2_ASAP7_75t_L g8865 ( 
.A(n_8305),
.B(n_7881),
.Y(n_8865)
);

INVx3_ASAP7_75t_L g8866 ( 
.A(n_8247),
.Y(n_8866)
);

NAND2xp5_ASAP7_75t_L g8867 ( 
.A(n_7652),
.B(n_7308),
.Y(n_8867)
);

AO21x2_ASAP7_75t_L g8868 ( 
.A1(n_8252),
.A2(n_6868),
.B(n_6846),
.Y(n_8868)
);

INVx2_ASAP7_75t_L g8869 ( 
.A(n_7937),
.Y(n_8869)
);

INVx2_ASAP7_75t_L g8870 ( 
.A(n_7942),
.Y(n_8870)
);

INVx4_ASAP7_75t_L g8871 ( 
.A(n_7857),
.Y(n_8871)
);

INVx2_ASAP7_75t_L g8872 ( 
.A(n_7942),
.Y(n_8872)
);

INVx1_ASAP7_75t_L g8873 ( 
.A(n_8177),
.Y(n_8873)
);

AO21x2_ASAP7_75t_L g8874 ( 
.A1(n_8254),
.A2(n_6876),
.B(n_6868),
.Y(n_8874)
);

INVx2_ASAP7_75t_L g8875 ( 
.A(n_8028),
.Y(n_8875)
);

NAND2xp5_ASAP7_75t_L g8876 ( 
.A(n_7724),
.B(n_7308),
.Y(n_8876)
);

AND2x2_ASAP7_75t_L g8877 ( 
.A(n_8305),
.B(n_6842),
.Y(n_8877)
);

INVx2_ASAP7_75t_L g8878 ( 
.A(n_8028),
.Y(n_8878)
);

NOR2xp33_ASAP7_75t_L g8879 ( 
.A(n_7677),
.B(n_6916),
.Y(n_8879)
);

HB1xp67_ASAP7_75t_L g8880 ( 
.A(n_8324),
.Y(n_8880)
);

AND2x4_ASAP7_75t_L g8881 ( 
.A(n_8108),
.B(n_6916),
.Y(n_8881)
);

AND2x2_ASAP7_75t_L g8882 ( 
.A(n_8305),
.B(n_6806),
.Y(n_8882)
);

NAND2xp5_ASAP7_75t_L g8883 ( 
.A(n_7672),
.B(n_7308),
.Y(n_8883)
);

INVx1_ASAP7_75t_L g8884 ( 
.A(n_8207),
.Y(n_8884)
);

AND2x2_ASAP7_75t_L g8885 ( 
.A(n_8305),
.B(n_6806),
.Y(n_8885)
);

HB1xp67_ASAP7_75t_L g8886 ( 
.A(n_7889),
.Y(n_8886)
);

INVx1_ASAP7_75t_L g8887 ( 
.A(n_8207),
.Y(n_8887)
);

INVx2_ASAP7_75t_SL g8888 ( 
.A(n_7889),
.Y(n_8888)
);

INVx2_ASAP7_75t_L g8889 ( 
.A(n_8084),
.Y(n_8889)
);

BUFx2_ASAP7_75t_L g8890 ( 
.A(n_7823),
.Y(n_8890)
);

INVx2_ASAP7_75t_L g8891 ( 
.A(n_8084),
.Y(n_8891)
);

INVx1_ASAP7_75t_L g8892 ( 
.A(n_8224),
.Y(n_8892)
);

INVx2_ASAP7_75t_L g8893 ( 
.A(n_8116),
.Y(n_8893)
);

AND2x2_ASAP7_75t_L g8894 ( 
.A(n_8230),
.B(n_6806),
.Y(n_8894)
);

AO22x1_ASAP7_75t_L g8895 ( 
.A1(n_7737),
.A2(n_6979),
.B1(n_7142),
.B2(n_6916),
.Y(n_8895)
);

AND2x2_ASAP7_75t_L g8896 ( 
.A(n_8038),
.B(n_6806),
.Y(n_8896)
);

AO21x2_ASAP7_75t_L g8897 ( 
.A1(n_8116),
.A2(n_6887),
.B(n_6876),
.Y(n_8897)
);

NAND2xp5_ASAP7_75t_L g8898 ( 
.A(n_7676),
.B(n_7029),
.Y(n_8898)
);

INVx2_ASAP7_75t_L g8899 ( 
.A(n_8118),
.Y(n_8899)
);

BUFx2_ASAP7_75t_L g8900 ( 
.A(n_7836),
.Y(n_8900)
);

AND2x4_ASAP7_75t_L g8901 ( 
.A(n_8245),
.B(n_6979),
.Y(n_8901)
);

AO21x2_ASAP7_75t_L g8902 ( 
.A1(n_8118),
.A2(n_6887),
.B(n_6876),
.Y(n_8902)
);

AND2x2_ASAP7_75t_L g8903 ( 
.A(n_8038),
.B(n_6806),
.Y(n_8903)
);

INVx1_ASAP7_75t_L g8904 ( 
.A(n_8224),
.Y(n_8904)
);

INVx1_ASAP7_75t_L g8905 ( 
.A(n_8268),
.Y(n_8905)
);

OR2x2_ASAP7_75t_L g8906 ( 
.A(n_7850),
.B(n_6826),
.Y(n_8906)
);

AO21x2_ASAP7_75t_L g8907 ( 
.A1(n_8006),
.A2(n_6889),
.B(n_6887),
.Y(n_8907)
);

INVx1_ASAP7_75t_L g8908 ( 
.A(n_8268),
.Y(n_8908)
);

INVx1_ASAP7_75t_L g8909 ( 
.A(n_8269),
.Y(n_8909)
);

INVx2_ASAP7_75t_L g8910 ( 
.A(n_8074),
.Y(n_8910)
);

OA21x2_ASAP7_75t_L g8911 ( 
.A1(n_8269),
.A2(n_7243),
.B(n_7235),
.Y(n_8911)
);

INVx2_ASAP7_75t_L g8912 ( 
.A(n_8074),
.Y(n_8912)
);

OR2x2_ASAP7_75t_L g8913 ( 
.A(n_7953),
.B(n_6826),
.Y(n_8913)
);

OAI21xp5_ASAP7_75t_L g8914 ( 
.A1(n_7760),
.A2(n_7466),
.B(n_7042),
.Y(n_8914)
);

OR2x6_ASAP7_75t_L g8915 ( 
.A(n_7889),
.B(n_7307),
.Y(n_8915)
);

AND2x2_ASAP7_75t_L g8916 ( 
.A(n_8038),
.B(n_6806),
.Y(n_8916)
);

INVx3_ASAP7_75t_L g8917 ( 
.A(n_8038),
.Y(n_8917)
);

INVx1_ASAP7_75t_L g8918 ( 
.A(n_8292),
.Y(n_8918)
);

INVx1_ASAP7_75t_L g8919 ( 
.A(n_8292),
.Y(n_8919)
);

INVx1_ASAP7_75t_L g8920 ( 
.A(n_8313),
.Y(n_8920)
);

AO21x2_ASAP7_75t_L g8921 ( 
.A1(n_7853),
.A2(n_6964),
.B(n_6889),
.Y(n_8921)
);

NOR2xp67_ASAP7_75t_R g8922 ( 
.A(n_8682),
.B(n_7836),
.Y(n_8922)
);

INVx1_ASAP7_75t_L g8923 ( 
.A(n_8596),
.Y(n_8923)
);

HB1xp67_ASAP7_75t_L g8924 ( 
.A(n_8641),
.Y(n_8924)
);

AND2x2_ASAP7_75t_L g8925 ( 
.A(n_8379),
.B(n_7847),
.Y(n_8925)
);

INVx2_ASAP7_75t_L g8926 ( 
.A(n_8545),
.Y(n_8926)
);

AND2x2_ASAP7_75t_L g8927 ( 
.A(n_8379),
.B(n_7653),
.Y(n_8927)
);

AND2x2_ASAP7_75t_L g8928 ( 
.A(n_8436),
.B(n_8075),
.Y(n_8928)
);

BUFx6f_ASAP7_75t_L g8929 ( 
.A(n_8337),
.Y(n_8929)
);

INVx1_ASAP7_75t_L g8930 ( 
.A(n_8653),
.Y(n_8930)
);

AND2x2_ASAP7_75t_L g8931 ( 
.A(n_8444),
.B(n_7773),
.Y(n_8931)
);

AND2x2_ASAP7_75t_L g8932 ( 
.A(n_8686),
.B(n_8073),
.Y(n_8932)
);

OAI22xp33_ASAP7_75t_L g8933 ( 
.A1(n_8373),
.A2(n_7730),
.B1(n_7684),
.B2(n_7743),
.Y(n_8933)
);

AND2x2_ASAP7_75t_L g8934 ( 
.A(n_8696),
.B(n_7864),
.Y(n_8934)
);

NAND2xp5_ASAP7_75t_L g8935 ( 
.A(n_8556),
.B(n_7889),
.Y(n_8935)
);

INVx1_ASAP7_75t_L g8936 ( 
.A(n_8339),
.Y(n_8936)
);

INVx1_ASAP7_75t_L g8937 ( 
.A(n_8365),
.Y(n_8937)
);

INVx2_ASAP7_75t_L g8938 ( 
.A(n_8545),
.Y(n_8938)
);

INVx1_ASAP7_75t_L g8939 ( 
.A(n_8361),
.Y(n_8939)
);

NAND2xp5_ASAP7_75t_L g8940 ( 
.A(n_8390),
.B(n_8606),
.Y(n_8940)
);

AOI211xp5_ASAP7_75t_L g8941 ( 
.A1(n_8764),
.A2(n_7948),
.B(n_7840),
.C(n_7833),
.Y(n_8941)
);

INVx1_ASAP7_75t_L g8942 ( 
.A(n_8376),
.Y(n_8942)
);

INVx2_ASAP7_75t_L g8943 ( 
.A(n_8545),
.Y(n_8943)
);

INVx2_ASAP7_75t_L g8944 ( 
.A(n_8545),
.Y(n_8944)
);

INVx2_ASAP7_75t_L g8945 ( 
.A(n_8628),
.Y(n_8945)
);

INVx1_ASAP7_75t_L g8946 ( 
.A(n_8378),
.Y(n_8946)
);

OR2x2_ASAP7_75t_L g8947 ( 
.A(n_8565),
.B(n_7728),
.Y(n_8947)
);

AND2x2_ASAP7_75t_L g8948 ( 
.A(n_8441),
.B(n_7864),
.Y(n_8948)
);

NOR2xp33_ASAP7_75t_R g8949 ( 
.A(n_8337),
.B(n_8031),
.Y(n_8949)
);

INVx2_ASAP7_75t_L g8950 ( 
.A(n_8628),
.Y(n_8950)
);

AND2x2_ASAP7_75t_L g8951 ( 
.A(n_8441),
.B(n_8031),
.Y(n_8951)
);

INVx1_ASAP7_75t_L g8952 ( 
.A(n_8385),
.Y(n_8952)
);

AND2x2_ASAP7_75t_L g8953 ( 
.A(n_8451),
.B(n_7820),
.Y(n_8953)
);

AND2x2_ASAP7_75t_L g8954 ( 
.A(n_8451),
.B(n_8456),
.Y(n_8954)
);

INVx1_ASAP7_75t_L g8955 ( 
.A(n_8386),
.Y(n_8955)
);

AND2x2_ASAP7_75t_L g8956 ( 
.A(n_8456),
.B(n_7820),
.Y(n_8956)
);

OR2x2_ASAP7_75t_L g8957 ( 
.A(n_8344),
.B(n_7788),
.Y(n_8957)
);

OR2x2_ASAP7_75t_L g8958 ( 
.A(n_8348),
.B(n_8051),
.Y(n_8958)
);

INVx1_ASAP7_75t_L g8959 ( 
.A(n_8399),
.Y(n_8959)
);

INVx2_ASAP7_75t_L g8960 ( 
.A(n_8628),
.Y(n_8960)
);

AND2x2_ASAP7_75t_L g8961 ( 
.A(n_8458),
.B(n_7878),
.Y(n_8961)
);

HB1xp67_ASAP7_75t_L g8962 ( 
.A(n_8415),
.Y(n_8962)
);

INVx1_ASAP7_75t_L g8963 ( 
.A(n_8405),
.Y(n_8963)
);

INVx2_ASAP7_75t_L g8964 ( 
.A(n_8628),
.Y(n_8964)
);

INVx1_ASAP7_75t_L g8965 ( 
.A(n_8407),
.Y(n_8965)
);

INVx3_ASAP7_75t_L g8966 ( 
.A(n_8716),
.Y(n_8966)
);

INVx1_ASAP7_75t_L g8967 ( 
.A(n_8410),
.Y(n_8967)
);

HB1xp67_ASAP7_75t_L g8968 ( 
.A(n_8447),
.Y(n_8968)
);

INVx2_ASAP7_75t_L g8969 ( 
.A(n_8636),
.Y(n_8969)
);

INVx2_ASAP7_75t_L g8970 ( 
.A(n_8636),
.Y(n_8970)
);

AND2x2_ASAP7_75t_L g8971 ( 
.A(n_8458),
.B(n_7901),
.Y(n_8971)
);

INVx1_ASAP7_75t_L g8972 ( 
.A(n_8412),
.Y(n_8972)
);

HB1xp67_ASAP7_75t_L g8973 ( 
.A(n_8502),
.Y(n_8973)
);

INVx1_ASAP7_75t_L g8974 ( 
.A(n_8419),
.Y(n_8974)
);

INVx2_ASAP7_75t_SL g8975 ( 
.A(n_8595),
.Y(n_8975)
);

INVx3_ASAP7_75t_L g8976 ( 
.A(n_8716),
.Y(n_8976)
);

INVx1_ASAP7_75t_L g8977 ( 
.A(n_8420),
.Y(n_8977)
);

INVx1_ASAP7_75t_L g8978 ( 
.A(n_8421),
.Y(n_8978)
);

INVx1_ASAP7_75t_L g8979 ( 
.A(n_8431),
.Y(n_8979)
);

AND2x2_ASAP7_75t_L g8980 ( 
.A(n_8467),
.B(n_7889),
.Y(n_8980)
);

AOI22xp33_ASAP7_75t_L g8981 ( 
.A1(n_8764),
.A2(n_8391),
.B1(n_8837),
.B2(n_8852),
.Y(n_8981)
);

INVx2_ASAP7_75t_L g8982 ( 
.A(n_8636),
.Y(n_8982)
);

NOR2xp33_ASAP7_75t_R g8983 ( 
.A(n_8337),
.B(n_7671),
.Y(n_8983)
);

INVx1_ASAP7_75t_L g8984 ( 
.A(n_8433),
.Y(n_8984)
);

INVx1_ASAP7_75t_L g8985 ( 
.A(n_8435),
.Y(n_8985)
);

AND2x2_ASAP7_75t_L g8986 ( 
.A(n_8467),
.B(n_7910),
.Y(n_8986)
);

AND2x2_ASAP7_75t_L g8987 ( 
.A(n_8471),
.B(n_7910),
.Y(n_8987)
);

INVx2_ASAP7_75t_L g8988 ( 
.A(n_8636),
.Y(n_8988)
);

AND2x2_ASAP7_75t_L g8989 ( 
.A(n_8471),
.B(n_7910),
.Y(n_8989)
);

AND2x2_ASAP7_75t_L g8990 ( 
.A(n_8474),
.B(n_7910),
.Y(n_8990)
);

OAI22xp5_ASAP7_75t_L g8991 ( 
.A1(n_8398),
.A2(n_7646),
.B1(n_7655),
.B2(n_7668),
.Y(n_8991)
);

NAND2xp5_ASAP7_75t_L g8992 ( 
.A(n_8620),
.B(n_7910),
.Y(n_8992)
);

HB1xp67_ASAP7_75t_L g8993 ( 
.A(n_8510),
.Y(n_8993)
);

INVx1_ASAP7_75t_L g8994 ( 
.A(n_8443),
.Y(n_8994)
);

INVx1_ASAP7_75t_L g8995 ( 
.A(n_8446),
.Y(n_8995)
);

INVx3_ASAP7_75t_L g8996 ( 
.A(n_8541),
.Y(n_8996)
);

AOI222xp33_ASAP7_75t_L g8997 ( 
.A1(n_8651),
.A2(n_7775),
.B1(n_8062),
.B2(n_7651),
.C1(n_7746),
.C2(n_7697),
.Y(n_8997)
);

AND2x2_ASAP7_75t_L g8998 ( 
.A(n_8474),
.B(n_7912),
.Y(n_8998)
);

OR2x2_ASAP7_75t_L g8999 ( 
.A(n_8350),
.B(n_8052),
.Y(n_8999)
);

AND2x2_ASAP7_75t_L g9000 ( 
.A(n_8477),
.B(n_8484),
.Y(n_9000)
);

INVx1_ASAP7_75t_L g9001 ( 
.A(n_8449),
.Y(n_9001)
);

HB1xp67_ASAP7_75t_L g9002 ( 
.A(n_8515),
.Y(n_9002)
);

OR2x2_ASAP7_75t_L g9003 ( 
.A(n_8355),
.B(n_7642),
.Y(n_9003)
);

INVx1_ASAP7_75t_L g9004 ( 
.A(n_8452),
.Y(n_9004)
);

INVx1_ASAP7_75t_L g9005 ( 
.A(n_8453),
.Y(n_9005)
);

INVx1_ASAP7_75t_L g9006 ( 
.A(n_8454),
.Y(n_9006)
);

INVxp67_ASAP7_75t_SL g9007 ( 
.A(n_8813),
.Y(n_9007)
);

INVx3_ASAP7_75t_L g9008 ( 
.A(n_8541),
.Y(n_9008)
);

AND2x2_ASAP7_75t_L g9009 ( 
.A(n_8477),
.B(n_8484),
.Y(n_9009)
);

INVx1_ASAP7_75t_L g9010 ( 
.A(n_8455),
.Y(n_9010)
);

OAI21x1_ASAP7_75t_L g9011 ( 
.A1(n_8861),
.A2(n_8169),
.B(n_8197),
.Y(n_9011)
);

INVx2_ASAP7_75t_L g9012 ( 
.A(n_8657),
.Y(n_9012)
);

INVx2_ASAP7_75t_L g9013 ( 
.A(n_8657),
.Y(n_9013)
);

INVx1_ASAP7_75t_L g9014 ( 
.A(n_8461),
.Y(n_9014)
);

INVx1_ASAP7_75t_L g9015 ( 
.A(n_8464),
.Y(n_9015)
);

AND2x2_ASAP7_75t_L g9016 ( 
.A(n_8488),
.B(n_7912),
.Y(n_9016)
);

INVx1_ASAP7_75t_L g9017 ( 
.A(n_8466),
.Y(n_9017)
);

INVx2_ASAP7_75t_L g9018 ( 
.A(n_8657),
.Y(n_9018)
);

OA21x2_ASAP7_75t_L g9019 ( 
.A1(n_8536),
.A2(n_8315),
.B(n_8313),
.Y(n_9019)
);

INVx1_ASAP7_75t_L g9020 ( 
.A(n_8473),
.Y(n_9020)
);

INVx2_ASAP7_75t_SL g9021 ( 
.A(n_8341),
.Y(n_9021)
);

INVx3_ASAP7_75t_L g9022 ( 
.A(n_8541),
.Y(n_9022)
);

BUFx2_ASAP7_75t_L g9023 ( 
.A(n_8772),
.Y(n_9023)
);

INVx2_ASAP7_75t_L g9024 ( 
.A(n_8657),
.Y(n_9024)
);

INVx1_ASAP7_75t_L g9025 ( 
.A(n_8481),
.Y(n_9025)
);

NOR4xp25_ASAP7_75t_SL g9026 ( 
.A(n_8806),
.B(n_7846),
.C(n_7845),
.D(n_8079),
.Y(n_9026)
);

NAND2xp5_ASAP7_75t_L g9027 ( 
.A(n_8654),
.B(n_7912),
.Y(n_9027)
);

INVx1_ASAP7_75t_L g9028 ( 
.A(n_8371),
.Y(n_9028)
);

INVx2_ASAP7_75t_SL g9029 ( 
.A(n_8595),
.Y(n_9029)
);

INVx1_ASAP7_75t_L g9030 ( 
.A(n_8537),
.Y(n_9030)
);

BUFx2_ASAP7_75t_L g9031 ( 
.A(n_8829),
.Y(n_9031)
);

INVx1_ASAP7_75t_SL g9032 ( 
.A(n_8401),
.Y(n_9032)
);

INVxp67_ASAP7_75t_SL g9033 ( 
.A(n_8813),
.Y(n_9033)
);

AND2x2_ASAP7_75t_L g9034 ( 
.A(n_8488),
.B(n_7912),
.Y(n_9034)
);

HB1xp67_ASAP7_75t_L g9035 ( 
.A(n_8724),
.Y(n_9035)
);

INVx2_ASAP7_75t_L g9036 ( 
.A(n_8564),
.Y(n_9036)
);

INVx5_ASAP7_75t_L g9037 ( 
.A(n_8337),
.Y(n_9037)
);

INVx2_ASAP7_75t_L g9038 ( 
.A(n_8564),
.Y(n_9038)
);

NAND2xp5_ASAP7_75t_L g9039 ( 
.A(n_8699),
.B(n_7912),
.Y(n_9039)
);

NOR2x1_ASAP7_75t_SL g9040 ( 
.A(n_8428),
.B(n_7657),
.Y(n_9040)
);

AND2x4_ASAP7_75t_L g9041 ( 
.A(n_8595),
.B(n_7938),
.Y(n_9041)
);

INVx2_ASAP7_75t_L g9042 ( 
.A(n_8594),
.Y(n_9042)
);

BUFx2_ASAP7_75t_L g9043 ( 
.A(n_8835),
.Y(n_9043)
);

OR2x2_ASAP7_75t_L g9044 ( 
.A(n_8576),
.B(n_8076),
.Y(n_9044)
);

INVx2_ASAP7_75t_L g9045 ( 
.A(n_8594),
.Y(n_9045)
);

INVx2_ASAP7_75t_L g9046 ( 
.A(n_8497),
.Y(n_9046)
);

INVx2_ASAP7_75t_L g9047 ( 
.A(n_8497),
.Y(n_9047)
);

OAI22xp5_ASAP7_75t_SL g9048 ( 
.A1(n_8779),
.A2(n_7827),
.B1(n_7835),
.B2(n_7674),
.Y(n_9048)
);

INVx1_ASAP7_75t_L g9049 ( 
.A(n_8486),
.Y(n_9049)
);

INVx2_ASAP7_75t_L g9050 ( 
.A(n_8497),
.Y(n_9050)
);

HB1xp67_ASAP7_75t_L g9051 ( 
.A(n_8735),
.Y(n_9051)
);

NAND2xp5_ASAP7_75t_L g9052 ( 
.A(n_8512),
.B(n_8840),
.Y(n_9052)
);

AND2x2_ASAP7_75t_L g9053 ( 
.A(n_8490),
.B(n_7938),
.Y(n_9053)
);

AND2x4_ASAP7_75t_L g9054 ( 
.A(n_8595),
.B(n_7938),
.Y(n_9054)
);

AND2x4_ASAP7_75t_L g9055 ( 
.A(n_8595),
.B(n_7938),
.Y(n_9055)
);

OR2x2_ASAP7_75t_L g9056 ( 
.A(n_8821),
.B(n_8248),
.Y(n_9056)
);

BUFx3_ASAP7_75t_L g9057 ( 
.A(n_8674),
.Y(n_9057)
);

NAND2x1_ASAP7_75t_L g9058 ( 
.A(n_8693),
.B(n_7657),
.Y(n_9058)
);

BUFx2_ASAP7_75t_L g9059 ( 
.A(n_8733),
.Y(n_9059)
);

NAND2xp5_ASAP7_75t_L g9060 ( 
.A(n_8890),
.B(n_7938),
.Y(n_9060)
);

AOI33xp33_ASAP7_75t_L g9061 ( 
.A1(n_8543),
.A2(n_7949),
.A3(n_7855),
.B1(n_7783),
.B2(n_8165),
.B3(n_8151),
.Y(n_9061)
);

INVx1_ASAP7_75t_L g9062 ( 
.A(n_8492),
.Y(n_9062)
);

INVx1_ASAP7_75t_L g9063 ( 
.A(n_8493),
.Y(n_9063)
);

HB1xp67_ASAP7_75t_L g9064 ( 
.A(n_8590),
.Y(n_9064)
);

INVx2_ASAP7_75t_L g9065 ( 
.A(n_8498),
.Y(n_9065)
);

INVx1_ASAP7_75t_L g9066 ( 
.A(n_8496),
.Y(n_9066)
);

INVx1_ASAP7_75t_L g9067 ( 
.A(n_8501),
.Y(n_9067)
);

INVx2_ASAP7_75t_L g9068 ( 
.A(n_8498),
.Y(n_9068)
);

INVx2_ASAP7_75t_L g9069 ( 
.A(n_8498),
.Y(n_9069)
);

AOI22xp33_ASAP7_75t_L g9070 ( 
.A1(n_8695),
.A2(n_7663),
.B1(n_7689),
.B2(n_7648),
.Y(n_9070)
);

INVx2_ASAP7_75t_L g9071 ( 
.A(n_8517),
.Y(n_9071)
);

INVx1_ASAP7_75t_L g9072 ( 
.A(n_8507),
.Y(n_9072)
);

AOI22xp33_ASAP7_75t_L g9073 ( 
.A1(n_8695),
.A2(n_8345),
.B1(n_8813),
.B2(n_8855),
.Y(n_9073)
);

BUFx3_ASAP7_75t_L g9074 ( 
.A(n_8674),
.Y(n_9074)
);

INVx2_ASAP7_75t_L g9075 ( 
.A(n_8517),
.Y(n_9075)
);

AND2x2_ASAP7_75t_L g9076 ( 
.A(n_8490),
.B(n_7722),
.Y(n_9076)
);

AND2x2_ASAP7_75t_L g9077 ( 
.A(n_8539),
.B(n_7657),
.Y(n_9077)
);

AND2x2_ASAP7_75t_L g9078 ( 
.A(n_8539),
.B(n_7657),
.Y(n_9078)
);

INVx2_ASAP7_75t_L g9079 ( 
.A(n_8517),
.Y(n_9079)
);

NOR2xp67_ASAP7_75t_L g9080 ( 
.A(n_8463),
.B(n_7950),
.Y(n_9080)
);

AO31x2_ASAP7_75t_L g9081 ( 
.A1(n_8427),
.A2(n_7882),
.A3(n_8180),
.B(n_8321),
.Y(n_9081)
);

BUFx3_ASAP7_75t_L g9082 ( 
.A(n_8612),
.Y(n_9082)
);

INVx2_ASAP7_75t_SL g9083 ( 
.A(n_8341),
.Y(n_9083)
);

INVx2_ASAP7_75t_L g9084 ( 
.A(n_8559),
.Y(n_9084)
);

AOI22xp33_ASAP7_75t_L g9085 ( 
.A1(n_8345),
.A2(n_7731),
.B1(n_7866),
.B2(n_7688),
.Y(n_9085)
);

HB1xp67_ASAP7_75t_L g9086 ( 
.A(n_8590),
.Y(n_9086)
);

INVx2_ASAP7_75t_L g9087 ( 
.A(n_8559),
.Y(n_9087)
);

AND2x2_ASAP7_75t_L g9088 ( 
.A(n_8548),
.B(n_7837),
.Y(n_9088)
);

NAND2xp5_ASAP7_75t_L g9089 ( 
.A(n_8900),
.B(n_7667),
.Y(n_9089)
);

INVx1_ASAP7_75t_L g9090 ( 
.A(n_8508),
.Y(n_9090)
);

INVx1_ASAP7_75t_L g9091 ( 
.A(n_8513),
.Y(n_9091)
);

INVx1_ASAP7_75t_L g9092 ( 
.A(n_8519),
.Y(n_9092)
);

HB1xp67_ASAP7_75t_L g9093 ( 
.A(n_8590),
.Y(n_9093)
);

NAND3xp33_ASAP7_75t_L g9094 ( 
.A(n_8725),
.B(n_8178),
.C(n_8231),
.Y(n_9094)
);

INVx1_ASAP7_75t_L g9095 ( 
.A(n_8523),
.Y(n_9095)
);

OR2x2_ASAP7_75t_L g9096 ( 
.A(n_8770),
.B(n_7996),
.Y(n_9096)
);

INVx1_ASAP7_75t_L g9097 ( 
.A(n_8524),
.Y(n_9097)
);

OR2x2_ASAP7_75t_L g9098 ( 
.A(n_8460),
.B(n_8226),
.Y(n_9098)
);

OAI21xp5_ASAP7_75t_L g9099 ( 
.A1(n_8806),
.A2(n_7710),
.B(n_7756),
.Y(n_9099)
);

INVx3_ASAP7_75t_L g9100 ( 
.A(n_8635),
.Y(n_9100)
);

AND2x2_ASAP7_75t_L g9101 ( 
.A(n_8548),
.B(n_7839),
.Y(n_9101)
);

AND2x2_ASAP7_75t_L g9102 ( 
.A(n_8389),
.B(n_8242),
.Y(n_9102)
);

CKINVDCx5p33_ASAP7_75t_R g9103 ( 
.A(n_8810),
.Y(n_9103)
);

INVx1_ASAP7_75t_L g9104 ( 
.A(n_8525),
.Y(n_9104)
);

AND2x2_ASAP7_75t_L g9105 ( 
.A(n_8389),
.B(n_7848),
.Y(n_9105)
);

OAI222xp33_ASAP7_75t_L g9106 ( 
.A1(n_8729),
.A2(n_7686),
.B1(n_8234),
.B2(n_7903),
.C1(n_7939),
.C2(n_7935),
.Y(n_9106)
);

INVx2_ASAP7_75t_L g9107 ( 
.A(n_8559),
.Y(n_9107)
);

OR2x2_ASAP7_75t_L g9108 ( 
.A(n_8460),
.B(n_8023),
.Y(n_9108)
);

INVx1_ASAP7_75t_L g9109 ( 
.A(n_8528),
.Y(n_9109)
);

INVx1_ASAP7_75t_L g9110 ( 
.A(n_8529),
.Y(n_9110)
);

INVx2_ASAP7_75t_L g9111 ( 
.A(n_8613),
.Y(n_9111)
);

INVx1_ASAP7_75t_L g9112 ( 
.A(n_8530),
.Y(n_9112)
);

BUFx2_ASAP7_75t_L g9113 ( 
.A(n_8733),
.Y(n_9113)
);

INVx1_ASAP7_75t_L g9114 ( 
.A(n_8531),
.Y(n_9114)
);

OR2x2_ASAP7_75t_L g9115 ( 
.A(n_8465),
.B(n_7927),
.Y(n_9115)
);

INVx1_ASAP7_75t_L g9116 ( 
.A(n_8533),
.Y(n_9116)
);

INVx2_ASAP7_75t_L g9117 ( 
.A(n_8613),
.Y(n_9117)
);

INVx1_ASAP7_75t_L g9118 ( 
.A(n_8542),
.Y(n_9118)
);

INVx2_ASAP7_75t_L g9119 ( 
.A(n_8613),
.Y(n_9119)
);

HB1xp67_ASAP7_75t_L g9120 ( 
.A(n_8465),
.Y(n_9120)
);

NOR2xp33_ASAP7_75t_L g9121 ( 
.A(n_8357),
.B(n_8706),
.Y(n_9121)
);

HB1xp67_ASAP7_75t_L g9122 ( 
.A(n_8468),
.Y(n_9122)
);

INVx3_ASAP7_75t_L g9123 ( 
.A(n_8635),
.Y(n_9123)
);

NOR2x1p5_ASAP7_75t_L g9124 ( 
.A(n_8463),
.B(n_7674),
.Y(n_9124)
);

BUFx3_ASAP7_75t_L g9125 ( 
.A(n_8612),
.Y(n_9125)
);

AND2x2_ASAP7_75t_L g9126 ( 
.A(n_8392),
.B(n_8408),
.Y(n_9126)
);

AND2x2_ASAP7_75t_L g9127 ( 
.A(n_8392),
.B(n_7679),
.Y(n_9127)
);

BUFx3_ASAP7_75t_L g9128 ( 
.A(n_8624),
.Y(n_9128)
);

OR2x2_ASAP7_75t_L g9129 ( 
.A(n_8468),
.B(n_8475),
.Y(n_9129)
);

AND2x2_ASAP7_75t_L g9130 ( 
.A(n_8408),
.B(n_7844),
.Y(n_9130)
);

AND2x2_ASAP7_75t_L g9131 ( 
.A(n_8411),
.B(n_8416),
.Y(n_9131)
);

AOI22xp33_ASAP7_75t_L g9132 ( 
.A1(n_8345),
.A2(n_7685),
.B1(n_7992),
.B2(n_7691),
.Y(n_9132)
);

INVxp67_ASAP7_75t_L g9133 ( 
.A(n_8886),
.Y(n_9133)
);

AND2x4_ASAP7_75t_L g9134 ( 
.A(n_8755),
.B(n_8260),
.Y(n_9134)
);

OAI33xp33_ASAP7_75t_L g9135 ( 
.A1(n_8726),
.A2(n_8228),
.A3(n_7732),
.B1(n_7989),
.B2(n_7943),
.B3(n_7811),
.Y(n_9135)
);

INVx1_ASAP7_75t_L g9136 ( 
.A(n_8544),
.Y(n_9136)
);

AND2x2_ASAP7_75t_L g9137 ( 
.A(n_8411),
.B(n_8175),
.Y(n_9137)
);

NOR4xp25_ASAP7_75t_SL g9138 ( 
.A(n_8844),
.B(n_7859),
.C(n_7929),
.D(n_8203),
.Y(n_9138)
);

BUFx2_ASAP7_75t_L g9139 ( 
.A(n_8733),
.Y(n_9139)
);

AND2x2_ASAP7_75t_L g9140 ( 
.A(n_8416),
.B(n_8191),
.Y(n_9140)
);

AND2x2_ASAP7_75t_L g9141 ( 
.A(n_8430),
.B(n_8088),
.Y(n_9141)
);

AOI22xp33_ASAP7_75t_L g9142 ( 
.A1(n_8855),
.A2(n_7715),
.B1(n_7696),
.B2(n_7718),
.Y(n_9142)
);

AND2x2_ASAP7_75t_L g9143 ( 
.A(n_8430),
.B(n_8088),
.Y(n_9143)
);

INVx2_ASAP7_75t_L g9144 ( 
.A(n_8652),
.Y(n_9144)
);

AND2x2_ASAP7_75t_L g9145 ( 
.A(n_8432),
.B(n_8168),
.Y(n_9145)
);

CKINVDCx5p33_ASAP7_75t_R g9146 ( 
.A(n_8810),
.Y(n_9146)
);

AND2x6_ASAP7_75t_L g9147 ( 
.A(n_8413),
.B(n_8106),
.Y(n_9147)
);

BUFx6f_ASAP7_75t_L g9148 ( 
.A(n_8624),
.Y(n_9148)
);

AND2x2_ASAP7_75t_L g9149 ( 
.A(n_8432),
.B(n_8174),
.Y(n_9149)
);

BUFx3_ASAP7_75t_L g9150 ( 
.A(n_8550),
.Y(n_9150)
);

NAND2xp5_ASAP7_75t_L g9151 ( 
.A(n_8725),
.B(n_8046),
.Y(n_9151)
);

AND2x4_ASAP7_75t_SL g9152 ( 
.A(n_8341),
.B(n_8115),
.Y(n_9152)
);

INVx3_ASAP7_75t_L g9153 ( 
.A(n_8635),
.Y(n_9153)
);

HB1xp67_ASAP7_75t_L g9154 ( 
.A(n_8475),
.Y(n_9154)
);

INVx1_ASAP7_75t_L g9155 ( 
.A(n_8547),
.Y(n_9155)
);

INVx1_ASAP7_75t_L g9156 ( 
.A(n_8549),
.Y(n_9156)
);

INVx2_ASAP7_75t_L g9157 ( 
.A(n_8652),
.Y(n_9157)
);

NAND3xp33_ASAP7_75t_L g9158 ( 
.A(n_8543),
.B(n_8121),
.C(n_8192),
.Y(n_9158)
);

INVxp67_ASAP7_75t_L g9159 ( 
.A(n_8785),
.Y(n_9159)
);

AND2x2_ASAP7_75t_L g9160 ( 
.A(n_8434),
.B(n_8707),
.Y(n_9160)
);

HB1xp67_ASAP7_75t_L g9161 ( 
.A(n_8483),
.Y(n_9161)
);

INVx2_ASAP7_75t_SL g9162 ( 
.A(n_8479),
.Y(n_9162)
);

INVx2_ASAP7_75t_L g9163 ( 
.A(n_8713),
.Y(n_9163)
);

AND2x2_ASAP7_75t_L g9164 ( 
.A(n_8434),
.B(n_8021),
.Y(n_9164)
);

INVx2_ASAP7_75t_L g9165 ( 
.A(n_8713),
.Y(n_9165)
);

INVx2_ASAP7_75t_L g9166 ( 
.A(n_8713),
.Y(n_9166)
);

AOI22xp33_ASAP7_75t_SL g9167 ( 
.A1(n_8745),
.A2(n_8115),
.B1(n_7886),
.B2(n_8133),
.Y(n_9167)
);

INVx2_ASAP7_75t_L g9168 ( 
.A(n_8713),
.Y(n_9168)
);

AND2x4_ASAP7_75t_L g9169 ( 
.A(n_8755),
.B(n_8260),
.Y(n_9169)
);

INVx2_ASAP7_75t_L g9170 ( 
.A(n_8762),
.Y(n_9170)
);

HB1xp67_ASAP7_75t_L g9171 ( 
.A(n_8483),
.Y(n_9171)
);

OR2x2_ASAP7_75t_L g9172 ( 
.A(n_8500),
.B(n_8751),
.Y(n_9172)
);

AND2x2_ASAP7_75t_L g9173 ( 
.A(n_8720),
.B(n_8167),
.Y(n_9173)
);

AND2x2_ASAP7_75t_L g9174 ( 
.A(n_8426),
.B(n_7933),
.Y(n_9174)
);

AND2x2_ASAP7_75t_L g9175 ( 
.A(n_8440),
.B(n_8318),
.Y(n_9175)
);

AND2x4_ASAP7_75t_SL g9176 ( 
.A(n_8733),
.B(n_8393),
.Y(n_9176)
);

NAND2x1_ASAP7_75t_L g9177 ( 
.A(n_8693),
.B(n_8290),
.Y(n_9177)
);

AND2x2_ASAP7_75t_L g9178 ( 
.A(n_8487),
.B(n_8225),
.Y(n_9178)
);

INVxp67_ASAP7_75t_L g9179 ( 
.A(n_8789),
.Y(n_9179)
);

AND2x4_ASAP7_75t_SL g9180 ( 
.A(n_8393),
.B(n_7785),
.Y(n_9180)
);

NAND2xp5_ASAP7_75t_L g9181 ( 
.A(n_8879),
.B(n_8281),
.Y(n_9181)
);

INVx1_ASAP7_75t_L g9182 ( 
.A(n_8554),
.Y(n_9182)
);

INVx4_ASAP7_75t_L g9183 ( 
.A(n_8479),
.Y(n_9183)
);

OR2x2_ASAP7_75t_L g9184 ( 
.A(n_8500),
.B(n_6826),
.Y(n_9184)
);

INVx2_ASAP7_75t_L g9185 ( 
.A(n_8762),
.Y(n_9185)
);

HB1xp67_ASAP7_75t_L g9186 ( 
.A(n_8754),
.Y(n_9186)
);

INVx1_ASAP7_75t_L g9187 ( 
.A(n_8557),
.Y(n_9187)
);

NAND2xp5_ASAP7_75t_L g9188 ( 
.A(n_8879),
.B(n_7819),
.Y(n_9188)
);

INVx1_ASAP7_75t_L g9189 ( 
.A(n_8567),
.Y(n_9189)
);

AND2x2_ASAP7_75t_L g9190 ( 
.A(n_8504),
.B(n_8225),
.Y(n_9190)
);

AND2x2_ASAP7_75t_L g9191 ( 
.A(n_8335),
.B(n_8132),
.Y(n_9191)
);

AND2x2_ASAP7_75t_L g9192 ( 
.A(n_8335),
.B(n_8135),
.Y(n_9192)
);

NAND2xp5_ASAP7_75t_L g9193 ( 
.A(n_8336),
.B(n_7959),
.Y(n_9193)
);

INVx2_ASAP7_75t_L g9194 ( 
.A(n_8762),
.Y(n_9194)
);

INVx1_ASAP7_75t_L g9195 ( 
.A(n_8569),
.Y(n_9195)
);

INVx1_ASAP7_75t_L g9196 ( 
.A(n_8581),
.Y(n_9196)
);

NAND2xp5_ASAP7_75t_L g9197 ( 
.A(n_8336),
.B(n_7806),
.Y(n_9197)
);

INVx3_ASAP7_75t_L g9198 ( 
.A(n_8393),
.Y(n_9198)
);

AND2x2_ASAP7_75t_L g9199 ( 
.A(n_8727),
.B(n_8145),
.Y(n_9199)
);

BUFx6f_ASAP7_75t_L g9200 ( 
.A(n_8479),
.Y(n_9200)
);

AND2x2_ASAP7_75t_L g9201 ( 
.A(n_8727),
.B(n_8738),
.Y(n_9201)
);

OR2x2_ASAP7_75t_L g9202 ( 
.A(n_8363),
.B(n_6826),
.Y(n_9202)
);

INVx1_ASAP7_75t_L g9203 ( 
.A(n_8584),
.Y(n_9203)
);

AND2x2_ASAP7_75t_L g9204 ( 
.A(n_8738),
.B(n_7830),
.Y(n_9204)
);

INVx2_ASAP7_75t_L g9205 ( 
.A(n_8762),
.Y(n_9205)
);

INVx3_ASAP7_75t_L g9206 ( 
.A(n_8403),
.Y(n_9206)
);

BUFx4f_ASAP7_75t_SL g9207 ( 
.A(n_8463),
.Y(n_9207)
);

AND2x2_ASAP7_75t_L g9208 ( 
.A(n_8553),
.B(n_7831),
.Y(n_9208)
);

OAI22xp33_ASAP7_75t_L g9209 ( 
.A1(n_8649),
.A2(n_7749),
.B1(n_8003),
.B2(n_7978),
.Y(n_9209)
);

AOI22xp5_ASAP7_75t_L g9210 ( 
.A1(n_8514),
.A2(n_8057),
.B1(n_8054),
.B2(n_8050),
.Y(n_9210)
);

INVxp67_ASAP7_75t_SL g9211 ( 
.A(n_8744),
.Y(n_9211)
);

INVx2_ASAP7_75t_L g9212 ( 
.A(n_8798),
.Y(n_9212)
);

INVx2_ASAP7_75t_L g9213 ( 
.A(n_8798),
.Y(n_9213)
);

NOR2xp33_ASAP7_75t_L g9214 ( 
.A(n_8706),
.B(n_8091),
.Y(n_9214)
);

AND2x2_ASAP7_75t_L g9215 ( 
.A(n_8578),
.B(n_7984),
.Y(n_9215)
);

OR2x2_ASAP7_75t_L g9216 ( 
.A(n_8758),
.B(n_6826),
.Y(n_9216)
);

AND2x2_ASAP7_75t_L g9217 ( 
.A(n_8601),
.B(n_7988),
.Y(n_9217)
);

INVx1_ASAP7_75t_L g9218 ( 
.A(n_8587),
.Y(n_9218)
);

AND2x2_ASAP7_75t_L g9219 ( 
.A(n_8746),
.B(n_7986),
.Y(n_9219)
);

HB1xp67_ASAP7_75t_L g9220 ( 
.A(n_8763),
.Y(n_9220)
);

INVx1_ASAP7_75t_L g9221 ( 
.A(n_8593),
.Y(n_9221)
);

INVx2_ASAP7_75t_L g9222 ( 
.A(n_8798),
.Y(n_9222)
);

AND2x2_ASAP7_75t_L g9223 ( 
.A(n_8795),
.B(n_7983),
.Y(n_9223)
);

INVx1_ASAP7_75t_L g9224 ( 
.A(n_8598),
.Y(n_9224)
);

HB1xp67_ASAP7_75t_L g9225 ( 
.A(n_8781),
.Y(n_9225)
);

INVx2_ASAP7_75t_L g9226 ( 
.A(n_8798),
.Y(n_9226)
);

BUFx3_ASAP7_75t_L g9227 ( 
.A(n_8485),
.Y(n_9227)
);

INVx1_ASAP7_75t_L g9228 ( 
.A(n_8599),
.Y(n_9228)
);

INVx1_ASAP7_75t_SL g9229 ( 
.A(n_8374),
.Y(n_9229)
);

INVx2_ASAP7_75t_L g9230 ( 
.A(n_8830),
.Y(n_9230)
);

INVx2_ASAP7_75t_L g9231 ( 
.A(n_8830),
.Y(n_9231)
);

NAND2xp5_ASAP7_75t_L g9232 ( 
.A(n_8382),
.B(n_7917),
.Y(n_9232)
);

INVx2_ASAP7_75t_L g9233 ( 
.A(n_8830),
.Y(n_9233)
);

INVx2_ASAP7_75t_L g9234 ( 
.A(n_8830),
.Y(n_9234)
);

OR2x2_ASAP7_75t_SL g9235 ( 
.A(n_8479),
.B(n_6829),
.Y(n_9235)
);

INVx1_ASAP7_75t_L g9236 ( 
.A(n_8604),
.Y(n_9236)
);

BUFx2_ASAP7_75t_L g9237 ( 
.A(n_8403),
.Y(n_9237)
);

INVx1_ASAP7_75t_L g9238 ( 
.A(n_8608),
.Y(n_9238)
);

INVx1_ASAP7_75t_L g9239 ( 
.A(n_8610),
.Y(n_9239)
);

INVx2_ASAP7_75t_L g9240 ( 
.A(n_8650),
.Y(n_9240)
);

HB1xp67_ASAP7_75t_L g9241 ( 
.A(n_8812),
.Y(n_9241)
);

INVx2_ASAP7_75t_L g9242 ( 
.A(n_8650),
.Y(n_9242)
);

AND2x2_ASAP7_75t_L g9243 ( 
.A(n_8795),
.B(n_8266),
.Y(n_9243)
);

INVx1_ASAP7_75t_L g9244 ( 
.A(n_8617),
.Y(n_9244)
);

AND2x2_ASAP7_75t_L g9245 ( 
.A(n_8803),
.B(n_8266),
.Y(n_9245)
);

INVx2_ASAP7_75t_L g9246 ( 
.A(n_8650),
.Y(n_9246)
);

INVx1_ASAP7_75t_L g9247 ( 
.A(n_8619),
.Y(n_9247)
);

INVx1_ASAP7_75t_L g9248 ( 
.A(n_8621),
.Y(n_9248)
);

INVx1_ASAP7_75t_L g9249 ( 
.A(n_8622),
.Y(n_9249)
);

INVx1_ASAP7_75t_L g9250 ( 
.A(n_8627),
.Y(n_9250)
);

INVx1_ASAP7_75t_L g9251 ( 
.A(n_8630),
.Y(n_9251)
);

HB1xp67_ASAP7_75t_L g9252 ( 
.A(n_8818),
.Y(n_9252)
);

BUFx2_ASAP7_75t_L g9253 ( 
.A(n_8403),
.Y(n_9253)
);

INVx2_ASAP7_75t_L g9254 ( 
.A(n_8660),
.Y(n_9254)
);

INVx2_ASAP7_75t_L g9255 ( 
.A(n_8660),
.Y(n_9255)
);

HB1xp67_ASAP7_75t_L g9256 ( 
.A(n_8828),
.Y(n_9256)
);

NAND2xp5_ASAP7_75t_SL g9257 ( 
.A(n_8561),
.B(n_8195),
.Y(n_9257)
);

BUFx2_ASAP7_75t_L g9258 ( 
.A(n_8347),
.Y(n_9258)
);

OAI21x1_ASAP7_75t_L g9259 ( 
.A1(n_8753),
.A2(n_7142),
.B(n_6979),
.Y(n_9259)
);

OAI211xp5_ASAP7_75t_L g9260 ( 
.A1(n_8482),
.A2(n_8140),
.B(n_7843),
.C(n_7842),
.Y(n_9260)
);

INVx1_ASAP7_75t_L g9261 ( 
.A(n_8634),
.Y(n_9261)
);

AND2x2_ASAP7_75t_L g9262 ( 
.A(n_8803),
.B(n_8293),
.Y(n_9262)
);

INVx1_ASAP7_75t_L g9263 ( 
.A(n_8642),
.Y(n_9263)
);

AND2x2_ASAP7_75t_L g9264 ( 
.A(n_8540),
.B(n_8293),
.Y(n_9264)
);

INVx2_ASAP7_75t_L g9265 ( 
.A(n_8660),
.Y(n_9265)
);

INVx2_ASAP7_75t_L g9266 ( 
.A(n_8675),
.Y(n_9266)
);

OAI22xp33_ASAP7_75t_L g9267 ( 
.A1(n_8867),
.A2(n_8185),
.B1(n_8188),
.B2(n_8111),
.Y(n_9267)
);

INVx1_ASAP7_75t_L g9268 ( 
.A(n_8643),
.Y(n_9268)
);

AND2x2_ASAP7_75t_L g9269 ( 
.A(n_8540),
.B(n_8295),
.Y(n_9269)
);

NAND2xp5_ASAP7_75t_L g9270 ( 
.A(n_8382),
.B(n_8090),
.Y(n_9270)
);

INVx2_ASAP7_75t_L g9271 ( 
.A(n_8675),
.Y(n_9271)
);

INVx2_ASAP7_75t_L g9272 ( 
.A(n_8675),
.Y(n_9272)
);

AOI22xp33_ASAP7_75t_L g9273 ( 
.A1(n_8855),
.A2(n_8072),
.B1(n_7860),
.B2(n_7861),
.Y(n_9273)
);

AND2x2_ASAP7_75t_L g9274 ( 
.A(n_8792),
.B(n_8295),
.Y(n_9274)
);

INVx1_ASAP7_75t_L g9275 ( 
.A(n_8658),
.Y(n_9275)
);

AND2x2_ASAP7_75t_L g9276 ( 
.A(n_8792),
.B(n_8309),
.Y(n_9276)
);

INVx2_ASAP7_75t_L g9277 ( 
.A(n_8702),
.Y(n_9277)
);

BUFx2_ASAP7_75t_SL g9278 ( 
.A(n_8505),
.Y(n_9278)
);

INVx1_ASAP7_75t_L g9279 ( 
.A(n_8664),
.Y(n_9279)
);

NAND2x1_ASAP7_75t_L g9280 ( 
.A(n_8823),
.B(n_8309),
.Y(n_9280)
);

AND2x4_ASAP7_75t_L g9281 ( 
.A(n_8755),
.B(n_8347),
.Y(n_9281)
);

AND2x2_ASAP7_75t_L g9282 ( 
.A(n_8807),
.B(n_8150),
.Y(n_9282)
);

INVx2_ASAP7_75t_L g9283 ( 
.A(n_8702),
.Y(n_9283)
);

INVx1_ASAP7_75t_L g9284 ( 
.A(n_8665),
.Y(n_9284)
);

OR2x2_ASAP7_75t_L g9285 ( 
.A(n_8423),
.B(n_6826),
.Y(n_9285)
);

INVx1_ASAP7_75t_L g9286 ( 
.A(n_8667),
.Y(n_9286)
);

AND2x4_ASAP7_75t_L g9287 ( 
.A(n_8347),
.B(n_7142),
.Y(n_9287)
);

NAND2xp5_ASAP7_75t_L g9288 ( 
.A(n_8396),
.B(n_8217),
.Y(n_9288)
);

INVx2_ASAP7_75t_L g9289 ( 
.A(n_8702),
.Y(n_9289)
);

INVx1_ASAP7_75t_L g9290 ( 
.A(n_8671),
.Y(n_9290)
);

BUFx2_ASAP7_75t_L g9291 ( 
.A(n_8485),
.Y(n_9291)
);

INVx1_ASAP7_75t_L g9292 ( 
.A(n_8673),
.Y(n_9292)
);

AND2x2_ASAP7_75t_L g9293 ( 
.A(n_8807),
.B(n_8153),
.Y(n_9293)
);

INVx1_ASAP7_75t_L g9294 ( 
.A(n_8677),
.Y(n_9294)
);

INVx1_ASAP7_75t_L g9295 ( 
.A(n_8681),
.Y(n_9295)
);

BUFx3_ASAP7_75t_L g9296 ( 
.A(n_8511),
.Y(n_9296)
);

INVx1_ASAP7_75t_L g9297 ( 
.A(n_8690),
.Y(n_9297)
);

NAND2xp5_ASAP7_75t_L g9298 ( 
.A(n_8396),
.B(n_7025),
.Y(n_9298)
);

INVx1_ASAP7_75t_SL g9299 ( 
.A(n_8469),
.Y(n_9299)
);

INVx1_ASAP7_75t_L g9300 ( 
.A(n_8698),
.Y(n_9300)
);

INVx1_ASAP7_75t_L g9301 ( 
.A(n_8700),
.Y(n_9301)
);

INVx2_ASAP7_75t_L g9302 ( 
.A(n_8823),
.Y(n_9302)
);

BUFx2_ASAP7_75t_L g9303 ( 
.A(n_8511),
.Y(n_9303)
);

INVx2_ASAP7_75t_L g9304 ( 
.A(n_8823),
.Y(n_9304)
);

AND2x2_ASAP7_75t_L g9305 ( 
.A(n_8522),
.B(n_8625),
.Y(n_9305)
);

AND2x2_ASAP7_75t_L g9306 ( 
.A(n_8714),
.B(n_8154),
.Y(n_9306)
);

HB1xp67_ASAP7_75t_L g9307 ( 
.A(n_8832),
.Y(n_9307)
);

AND2x2_ASAP7_75t_L g9308 ( 
.A(n_8836),
.B(n_8880),
.Y(n_9308)
);

HB1xp67_ASAP7_75t_L g9309 ( 
.A(n_8639),
.Y(n_9309)
);

INVx1_ASAP7_75t_L g9310 ( 
.A(n_8704),
.Y(n_9310)
);

HB1xp67_ASAP7_75t_L g9311 ( 
.A(n_8639),
.Y(n_9311)
);

INVx1_ASAP7_75t_L g9312 ( 
.A(n_8708),
.Y(n_9312)
);

INVx1_ASAP7_75t_L g9313 ( 
.A(n_8710),
.Y(n_9313)
);

INVx1_ASAP7_75t_SL g9314 ( 
.A(n_8552),
.Y(n_9314)
);

OAI221xp5_ASAP7_75t_L g9315 ( 
.A1(n_8417),
.A2(n_8123),
.B1(n_8220),
.B2(n_8218),
.C(n_7716),
.Y(n_9315)
);

INVx2_ASAP7_75t_L g9316 ( 
.A(n_8823),
.Y(n_9316)
);

AND2x2_ASAP7_75t_L g9317 ( 
.A(n_8427),
.B(n_8162),
.Y(n_9317)
);

INVx1_ASAP7_75t_L g9318 ( 
.A(n_8711),
.Y(n_9318)
);

OAI21xp5_ASAP7_75t_L g9319 ( 
.A1(n_8470),
.A2(n_7793),
.B(n_7796),
.Y(n_9319)
);

INVx2_ASAP7_75t_L g9320 ( 
.A(n_8546),
.Y(n_9320)
);

INVx1_ASAP7_75t_L g9321 ( 
.A(n_8712),
.Y(n_9321)
);

INVx1_ASAP7_75t_L g9322 ( 
.A(n_8715),
.Y(n_9322)
);

BUFx3_ASAP7_75t_L g9323 ( 
.A(n_8552),
.Y(n_9323)
);

INVx1_ASAP7_75t_L g9324 ( 
.A(n_8728),
.Y(n_9324)
);

AND2x2_ASAP7_75t_L g9325 ( 
.A(n_8670),
.B(n_7771),
.Y(n_9325)
);

INVx2_ASAP7_75t_L g9326 ( 
.A(n_8546),
.Y(n_9326)
);

INVx1_ASAP7_75t_L g9327 ( 
.A(n_8732),
.Y(n_9327)
);

AND2x2_ASAP7_75t_L g9328 ( 
.A(n_8670),
.B(n_7870),
.Y(n_9328)
);

BUFx2_ASAP7_75t_L g9329 ( 
.A(n_8558),
.Y(n_9329)
);

NAND2xp5_ASAP7_75t_L g9330 ( 
.A(n_8526),
.B(n_7961),
.Y(n_9330)
);

INVx2_ASAP7_75t_L g9331 ( 
.A(n_8546),
.Y(n_9331)
);

AND2x4_ASAP7_75t_L g9332 ( 
.A(n_8370),
.B(n_7178),
.Y(n_9332)
);

AND2x2_ASAP7_75t_L g9333 ( 
.A(n_8739),
.B(n_7954),
.Y(n_9333)
);

BUFx8_ASAP7_75t_L g9334 ( 
.A(n_8489),
.Y(n_9334)
);

INVx1_ASAP7_75t_L g9335 ( 
.A(n_8736),
.Y(n_9335)
);

BUFx2_ASAP7_75t_L g9336 ( 
.A(n_8558),
.Y(n_9336)
);

INVx3_ASAP7_75t_L g9337 ( 
.A(n_8489),
.Y(n_9337)
);

INVx1_ASAP7_75t_L g9338 ( 
.A(n_8805),
.Y(n_9338)
);

AND2x2_ASAP7_75t_L g9339 ( 
.A(n_8739),
.B(n_8128),
.Y(n_9339)
);

INVx4_ASAP7_75t_L g9340 ( 
.A(n_8489),
.Y(n_9340)
);

OR2x2_ASAP7_75t_L g9341 ( 
.A(n_8566),
.B(n_8250),
.Y(n_9341)
);

AND2x2_ASAP7_75t_L g9342 ( 
.A(n_8825),
.B(n_7824),
.Y(n_9342)
);

HB1xp67_ASAP7_75t_L g9343 ( 
.A(n_8639),
.Y(n_9343)
);

INVx3_ASAP7_75t_L g9344 ( 
.A(n_8489),
.Y(n_9344)
);

INVx2_ASAP7_75t_L g9345 ( 
.A(n_8546),
.Y(n_9345)
);

HB1xp67_ASAP7_75t_L g9346 ( 
.A(n_8669),
.Y(n_9346)
);

AND2x2_ASAP7_75t_L g9347 ( 
.A(n_8592),
.B(n_8106),
.Y(n_9347)
);

INVx1_ASAP7_75t_L g9348 ( 
.A(n_8805),
.Y(n_9348)
);

AND2x4_ASAP7_75t_L g9349 ( 
.A(n_8370),
.B(n_7178),
.Y(n_9349)
);

INVx2_ASAP7_75t_SL g9350 ( 
.A(n_8644),
.Y(n_9350)
);

AND2x4_ASAP7_75t_SL g9351 ( 
.A(n_8814),
.B(n_7873),
.Y(n_9351)
);

HB1xp67_ASAP7_75t_L g9352 ( 
.A(n_8669),
.Y(n_9352)
);

AND2x2_ASAP7_75t_L g9353 ( 
.A(n_8592),
.B(n_8106),
.Y(n_9353)
);

BUFx3_ASAP7_75t_L g9354 ( 
.A(n_8494),
.Y(n_9354)
);

INVx1_ASAP7_75t_L g9355 ( 
.A(n_8815),
.Y(n_9355)
);

INVx1_ASAP7_75t_L g9356 ( 
.A(n_8815),
.Y(n_9356)
);

INVx1_ASAP7_75t_L g9357 ( 
.A(n_8822),
.Y(n_9357)
);

OAI221xp5_ASAP7_75t_L g9358 ( 
.A1(n_8816),
.A2(n_8190),
.B1(n_8012),
.B2(n_8127),
.C(n_7852),
.Y(n_9358)
);

OR2x2_ASAP7_75t_L g9359 ( 
.A(n_8566),
.B(n_8258),
.Y(n_9359)
);

INVx1_ASAP7_75t_SL g9360 ( 
.A(n_8413),
.Y(n_9360)
);

AND2x2_ASAP7_75t_L g9361 ( 
.A(n_8387),
.B(n_8106),
.Y(n_9361)
);

INVx2_ASAP7_75t_R g9362 ( 
.A(n_8791),
.Y(n_9362)
);

INVx2_ASAP7_75t_L g9363 ( 
.A(n_8644),
.Y(n_9363)
);

AND2x2_ASAP7_75t_L g9364 ( 
.A(n_8387),
.B(n_7318),
.Y(n_9364)
);

AOI22xp33_ASAP7_75t_L g9365 ( 
.A1(n_8538),
.A2(n_7851),
.B1(n_7849),
.B2(n_8018),
.Y(n_9365)
);

INVx2_ASAP7_75t_L g9366 ( 
.A(n_8644),
.Y(n_9366)
);

BUFx2_ASAP7_75t_L g9367 ( 
.A(n_8457),
.Y(n_9367)
);

INVx1_ASAP7_75t_L g9368 ( 
.A(n_8822),
.Y(n_9368)
);

NAND2xp5_ASAP7_75t_L g9369 ( 
.A(n_8526),
.B(n_7966),
.Y(n_9369)
);

INVx1_ASAP7_75t_L g9370 ( 
.A(n_8849),
.Y(n_9370)
);

INVx1_ASAP7_75t_L g9371 ( 
.A(n_8849),
.Y(n_9371)
);

AND2x2_ASAP7_75t_L g9372 ( 
.A(n_8757),
.B(n_7318),
.Y(n_9372)
);

INVx2_ASAP7_75t_L g9373 ( 
.A(n_8644),
.Y(n_9373)
);

INVx2_ASAP7_75t_L g9374 ( 
.A(n_8342),
.Y(n_9374)
);

INVx2_ASAP7_75t_L g9375 ( 
.A(n_8342),
.Y(n_9375)
);

NAND2xp5_ASAP7_75t_L g9376 ( 
.A(n_8532),
.B(n_7985),
.Y(n_9376)
);

OR2x2_ASAP7_75t_L g9377 ( 
.A(n_8568),
.B(n_8271),
.Y(n_9377)
);

OR2x2_ASAP7_75t_L g9378 ( 
.A(n_8568),
.B(n_8277),
.Y(n_9378)
);

INVx3_ASAP7_75t_L g9379 ( 
.A(n_8494),
.Y(n_9379)
);

AND2x2_ASAP7_75t_L g9380 ( 
.A(n_8757),
.B(n_7370),
.Y(n_9380)
);

INVx1_ASAP7_75t_L g9381 ( 
.A(n_8851),
.Y(n_9381)
);

OR2x2_ASAP7_75t_L g9382 ( 
.A(n_8898),
.B(n_7486),
.Y(n_9382)
);

HB1xp67_ASAP7_75t_L g9383 ( 
.A(n_8669),
.Y(n_9383)
);

AOI21xp5_ASAP7_75t_L g9384 ( 
.A1(n_8883),
.A2(n_8272),
.B(n_8246),
.Y(n_9384)
);

INVx2_ASAP7_75t_L g9385 ( 
.A(n_8360),
.Y(n_9385)
);

INVx1_ASAP7_75t_L g9386 ( 
.A(n_8851),
.Y(n_9386)
);

AND2x4_ASAP7_75t_L g9387 ( 
.A(n_8370),
.B(n_7178),
.Y(n_9387)
);

NAND2x1_ASAP7_75t_L g9388 ( 
.A(n_8457),
.B(n_6979),
.Y(n_9388)
);

BUFx2_ASAP7_75t_L g9389 ( 
.A(n_8457),
.Y(n_9389)
);

INVx2_ASAP7_75t_L g9390 ( 
.A(n_8360),
.Y(n_9390)
);

INVx3_ASAP7_75t_L g9391 ( 
.A(n_8494),
.Y(n_9391)
);

OAI21xp5_ASAP7_75t_L g9392 ( 
.A1(n_8482),
.A2(n_7967),
.B(n_7999),
.Y(n_9392)
);

INVx1_ASAP7_75t_L g9393 ( 
.A(n_8858),
.Y(n_9393)
);

INVx2_ASAP7_75t_L g9394 ( 
.A(n_8656),
.Y(n_9394)
);

INVx2_ASAP7_75t_L g9395 ( 
.A(n_8656),
.Y(n_9395)
);

AND2x2_ASAP7_75t_L g9396 ( 
.A(n_8775),
.B(n_8784),
.Y(n_9396)
);

INVx2_ASAP7_75t_L g9397 ( 
.A(n_8662),
.Y(n_9397)
);

NOR2x1_ASAP7_75t_SL g9398 ( 
.A(n_8790),
.B(n_7899),
.Y(n_9398)
);

AO31x2_ASAP7_75t_L g9399 ( 
.A1(n_8520),
.A2(n_8296),
.A3(n_8316),
.B(n_8078),
.Y(n_9399)
);

AND2x2_ASAP7_75t_L g9400 ( 
.A(n_8775),
.B(n_7370),
.Y(n_9400)
);

INVx1_ASAP7_75t_L g9401 ( 
.A(n_8858),
.Y(n_9401)
);

AND2x2_ASAP7_75t_L g9402 ( 
.A(n_8784),
.B(n_7423),
.Y(n_9402)
);

AND2x2_ASAP7_75t_L g9403 ( 
.A(n_8866),
.B(n_7423),
.Y(n_9403)
);

NOR2x1_ASAP7_75t_SL g9404 ( 
.A(n_8790),
.B(n_7928),
.Y(n_9404)
);

INVxp67_ASAP7_75t_L g9405 ( 
.A(n_8442),
.Y(n_9405)
);

HB1xp67_ASAP7_75t_L g9406 ( 
.A(n_8506),
.Y(n_9406)
);

INVx3_ASAP7_75t_L g9407 ( 
.A(n_8494),
.Y(n_9407)
);

NAND2xp5_ASAP7_75t_L g9408 ( 
.A(n_8532),
.B(n_8274),
.Y(n_9408)
);

INVx2_ASAP7_75t_L g9409 ( 
.A(n_8662),
.Y(n_9409)
);

NAND2xp5_ASAP7_75t_L g9410 ( 
.A(n_8534),
.B(n_8286),
.Y(n_9410)
);

OR2x2_ASAP7_75t_L g9411 ( 
.A(n_8780),
.B(n_7486),
.Y(n_9411)
);

OR2x2_ASAP7_75t_L g9412 ( 
.A(n_8368),
.B(n_7601),
.Y(n_9412)
);

INVx1_ASAP7_75t_L g9413 ( 
.A(n_8860),
.Y(n_9413)
);

AND2x2_ASAP7_75t_L g9414 ( 
.A(n_8866),
.B(n_7459),
.Y(n_9414)
);

INVx1_ASAP7_75t_L g9415 ( 
.A(n_8860),
.Y(n_9415)
);

NAND2xp5_ASAP7_75t_L g9416 ( 
.A(n_8534),
.B(n_7990),
.Y(n_9416)
);

INVx1_ASAP7_75t_L g9417 ( 
.A(n_8869),
.Y(n_9417)
);

AND2x2_ASAP7_75t_L g9418 ( 
.A(n_8866),
.B(n_7459),
.Y(n_9418)
);

AND2x2_ASAP7_75t_L g9419 ( 
.A(n_8747),
.B(n_7173),
.Y(n_9419)
);

INVx2_ASAP7_75t_L g9420 ( 
.A(n_8871),
.Y(n_9420)
);

HB1xp67_ASAP7_75t_L g9421 ( 
.A(n_8506),
.Y(n_9421)
);

OAI22xp33_ASAP7_75t_L g9422 ( 
.A1(n_8843),
.A2(n_8244),
.B1(n_8330),
.B2(n_8314),
.Y(n_9422)
);

INVx1_ASAP7_75t_L g9423 ( 
.A(n_8869),
.Y(n_9423)
);

NAND2xp5_ASAP7_75t_L g9424 ( 
.A(n_8551),
.B(n_8560),
.Y(n_9424)
);

NOR2xp33_ASAP7_75t_L g9425 ( 
.A(n_8505),
.B(n_7960),
.Y(n_9425)
);

INVx3_ASAP7_75t_L g9426 ( 
.A(n_8871),
.Y(n_9426)
);

OR2x2_ASAP7_75t_L g9427 ( 
.A(n_8397),
.B(n_7601),
.Y(n_9427)
);

NOR2x1p5_ASAP7_75t_L g9428 ( 
.A(n_8505),
.B(n_7960),
.Y(n_9428)
);

AND2x2_ASAP7_75t_L g9429 ( 
.A(n_8747),
.B(n_7173),
.Y(n_9429)
);

OR2x2_ASAP7_75t_L g9430 ( 
.A(n_8394),
.B(n_8317),
.Y(n_9430)
);

HB1xp67_ASAP7_75t_L g9431 ( 
.A(n_8786),
.Y(n_9431)
);

HB1xp67_ASAP7_75t_L g9432 ( 
.A(n_8786),
.Y(n_9432)
);

NAND2xp5_ASAP7_75t_L g9433 ( 
.A(n_8551),
.B(n_8130),
.Y(n_9433)
);

NAND2xp5_ASAP7_75t_L g9434 ( 
.A(n_8560),
.B(n_8166),
.Y(n_9434)
);

INVx1_ASAP7_75t_L g9435 ( 
.A(n_8870),
.Y(n_9435)
);

INVx1_ASAP7_75t_L g9436 ( 
.A(n_8870),
.Y(n_9436)
);

INVx1_ASAP7_75t_L g9437 ( 
.A(n_8872),
.Y(n_9437)
);

INVx2_ASAP7_75t_L g9438 ( 
.A(n_8871),
.Y(n_9438)
);

INVx1_ASAP7_75t_L g9439 ( 
.A(n_8872),
.Y(n_9439)
);

OAI221xp5_ASAP7_75t_L g9440 ( 
.A1(n_8914),
.A2(n_7781),
.B1(n_7774),
.B2(n_7763),
.C(n_7995),
.Y(n_9440)
);

INVx1_ASAP7_75t_L g9441 ( 
.A(n_8875),
.Y(n_9441)
);

AND2x2_ASAP7_75t_L g9442 ( 
.A(n_8748),
.B(n_7207),
.Y(n_9442)
);

HB1xp67_ASAP7_75t_L g9443 ( 
.A(n_8787),
.Y(n_9443)
);

NAND2xp5_ASAP7_75t_L g9444 ( 
.A(n_8563),
.B(n_7993),
.Y(n_9444)
);

INVx1_ASAP7_75t_L g9445 ( 
.A(n_8875),
.Y(n_9445)
);

INVx2_ASAP7_75t_L g9446 ( 
.A(n_8915),
.Y(n_9446)
);

BUFx6f_ASAP7_75t_L g9447 ( 
.A(n_8459),
.Y(n_9447)
);

AND2x2_ASAP7_75t_L g9448 ( 
.A(n_8748),
.B(n_7207),
.Y(n_9448)
);

INVx1_ASAP7_75t_L g9449 ( 
.A(n_8878),
.Y(n_9449)
);

INVx2_ASAP7_75t_SL g9450 ( 
.A(n_8573),
.Y(n_9450)
);

AND2x2_ASAP7_75t_L g9451 ( 
.A(n_8814),
.B(n_7982),
.Y(n_9451)
);

INVx1_ASAP7_75t_L g9452 ( 
.A(n_8878),
.Y(n_9452)
);

NAND2x1_ASAP7_75t_L g9453 ( 
.A(n_8457),
.B(n_7142),
.Y(n_9453)
);

INVx2_ASAP7_75t_L g9454 ( 
.A(n_8915),
.Y(n_9454)
);

OR2x2_ASAP7_75t_L g9455 ( 
.A(n_8572),
.B(n_8141),
.Y(n_9455)
);

NAND2xp5_ASAP7_75t_L g9456 ( 
.A(n_8563),
.B(n_8186),
.Y(n_9456)
);

NAND2xp5_ASAP7_75t_L g9457 ( 
.A(n_8442),
.B(n_8007),
.Y(n_9457)
);

INVx2_ASAP7_75t_SL g9458 ( 
.A(n_8573),
.Y(n_9458)
);

HB1xp67_ASAP7_75t_L g9459 ( 
.A(n_8787),
.Y(n_9459)
);

NAND2xp5_ASAP7_75t_L g9460 ( 
.A(n_8491),
.B(n_7029),
.Y(n_9460)
);

INVx2_ASAP7_75t_L g9461 ( 
.A(n_8915),
.Y(n_9461)
);

INVx1_ASAP7_75t_L g9462 ( 
.A(n_8910),
.Y(n_9462)
);

INVx2_ASAP7_75t_L g9463 ( 
.A(n_8915),
.Y(n_9463)
);

NAND2xp5_ASAP7_75t_L g9464 ( 
.A(n_8491),
.B(n_7035),
.Y(n_9464)
);

INVx1_ASAP7_75t_L g9465 ( 
.A(n_8910),
.Y(n_9465)
);

INVx2_ASAP7_75t_L g9466 ( 
.A(n_8647),
.Y(n_9466)
);

INVx2_ASAP7_75t_L g9467 ( 
.A(n_8647),
.Y(n_9467)
);

AND2x2_ASAP7_75t_L g9468 ( 
.A(n_8814),
.B(n_8105),
.Y(n_9468)
);

INVx1_ASAP7_75t_L g9469 ( 
.A(n_8912),
.Y(n_9469)
);

INVx1_ASAP7_75t_L g9470 ( 
.A(n_8912),
.Y(n_9470)
);

INVxp67_ASAP7_75t_L g9471 ( 
.A(n_8521),
.Y(n_9471)
);

INVxp67_ASAP7_75t_L g9472 ( 
.A(n_8521),
.Y(n_9472)
);

INVx2_ASAP7_75t_L g9473 ( 
.A(n_8774),
.Y(n_9473)
);

NAND2xp5_ASAP7_75t_L g9474 ( 
.A(n_8577),
.B(n_7035),
.Y(n_9474)
);

INVx2_ASAP7_75t_SL g9475 ( 
.A(n_8574),
.Y(n_9475)
);

NAND2xp5_ASAP7_75t_L g9476 ( 
.A(n_8577),
.B(n_8793),
.Y(n_9476)
);

INVx1_ASAP7_75t_L g9477 ( 
.A(n_8765),
.Y(n_9477)
);

AND2x2_ASAP7_75t_L g9478 ( 
.A(n_8819),
.B(n_8574),
.Y(n_9478)
);

HB1xp67_ASAP7_75t_L g9479 ( 
.A(n_8788),
.Y(n_9479)
);

INVx1_ASAP7_75t_L g9480 ( 
.A(n_8767),
.Y(n_9480)
);

AND2x2_ASAP7_75t_L g9481 ( 
.A(n_8819),
.B(n_8122),
.Y(n_9481)
);

AND2x2_ASAP7_75t_L g9482 ( 
.A(n_8819),
.B(n_8001),
.Y(n_9482)
);

INVx2_ASAP7_75t_L g9483 ( 
.A(n_9057),
.Y(n_9483)
);

INVx2_ASAP7_75t_L g9484 ( 
.A(n_9057),
.Y(n_9484)
);

NAND2xp5_ASAP7_75t_L g9485 ( 
.A(n_9151),
.B(n_8888),
.Y(n_9485)
);

INVx2_ASAP7_75t_L g9486 ( 
.A(n_9074),
.Y(n_9486)
);

OR2x2_ASAP7_75t_L g9487 ( 
.A(n_8940),
.B(n_8572),
.Y(n_9487)
);

AND2x2_ASAP7_75t_L g9488 ( 
.A(n_9074),
.B(n_8459),
.Y(n_9488)
);

INVx2_ASAP7_75t_SL g9489 ( 
.A(n_9037),
.Y(n_9489)
);

AOI22xp33_ASAP7_75t_L g9490 ( 
.A1(n_9135),
.A2(n_8811),
.B1(n_8809),
.B2(n_8609),
.Y(n_9490)
);

INVx1_ASAP7_75t_L g9491 ( 
.A(n_9186),
.Y(n_9491)
);

BUFx3_ASAP7_75t_L g9492 ( 
.A(n_8929),
.Y(n_9492)
);

AND2x2_ASAP7_75t_L g9493 ( 
.A(n_9152),
.B(n_8476),
.Y(n_9493)
);

AND2x4_ASAP7_75t_L g9494 ( 
.A(n_9152),
.B(n_8476),
.Y(n_9494)
);

AND2x2_ASAP7_75t_L g9495 ( 
.A(n_9032),
.B(n_8648),
.Y(n_9495)
);

INVx1_ASAP7_75t_L g9496 ( 
.A(n_9186),
.Y(n_9496)
);

INVx1_ASAP7_75t_L g9497 ( 
.A(n_9220),
.Y(n_9497)
);

BUFx3_ASAP7_75t_L g9498 ( 
.A(n_8929),
.Y(n_9498)
);

INVx3_ASAP7_75t_L g9499 ( 
.A(n_8929),
.Y(n_9499)
);

NAND2x1_ASAP7_75t_L g9500 ( 
.A(n_9134),
.B(n_8480),
.Y(n_9500)
);

BUFx2_ASAP7_75t_L g9501 ( 
.A(n_8949),
.Y(n_9501)
);

INVx3_ASAP7_75t_L g9502 ( 
.A(n_8929),
.Y(n_9502)
);

BUFx2_ASAP7_75t_L g9503 ( 
.A(n_8949),
.Y(n_9503)
);

INVx5_ASAP7_75t_L g9504 ( 
.A(n_9037),
.Y(n_9504)
);

INVx3_ASAP7_75t_L g9505 ( 
.A(n_9200),
.Y(n_9505)
);

INVx1_ASAP7_75t_L g9506 ( 
.A(n_9220),
.Y(n_9506)
);

INVx2_ASAP7_75t_SL g9507 ( 
.A(n_9037),
.Y(n_9507)
);

AND2x2_ASAP7_75t_L g9508 ( 
.A(n_8934),
.B(n_8648),
.Y(n_9508)
);

OR2x2_ASAP7_75t_L g9509 ( 
.A(n_9229),
.B(n_8575),
.Y(n_9509)
);

INVx1_ASAP7_75t_L g9510 ( 
.A(n_9225),
.Y(n_9510)
);

AND2x2_ASAP7_75t_L g9511 ( 
.A(n_8948),
.B(n_8648),
.Y(n_9511)
);

AND2x2_ASAP7_75t_L g9512 ( 
.A(n_8951),
.B(n_8663),
.Y(n_9512)
);

HB1xp67_ASAP7_75t_L g9513 ( 
.A(n_9064),
.Y(n_9513)
);

NAND2xp5_ASAP7_75t_L g9514 ( 
.A(n_8924),
.B(n_8888),
.Y(n_9514)
);

INVx2_ASAP7_75t_L g9515 ( 
.A(n_8996),
.Y(n_9515)
);

INVx1_ASAP7_75t_L g9516 ( 
.A(n_9225),
.Y(n_9516)
);

INVx2_ASAP7_75t_L g9517 ( 
.A(n_8996),
.Y(n_9517)
);

INVx2_ASAP7_75t_L g9518 ( 
.A(n_9008),
.Y(n_9518)
);

INVx2_ASAP7_75t_L g9519 ( 
.A(n_9008),
.Y(n_9519)
);

AO21x2_ASAP7_75t_L g9520 ( 
.A1(n_9064),
.A2(n_8618),
.B(n_8723),
.Y(n_9520)
);

INVx2_ASAP7_75t_L g9521 ( 
.A(n_9022),
.Y(n_9521)
);

INVx2_ASAP7_75t_L g9522 ( 
.A(n_9022),
.Y(n_9522)
);

INVx2_ASAP7_75t_SL g9523 ( 
.A(n_9037),
.Y(n_9523)
);

INVx1_ASAP7_75t_L g9524 ( 
.A(n_9241),
.Y(n_9524)
);

INVx2_ASAP7_75t_L g9525 ( 
.A(n_9148),
.Y(n_9525)
);

BUFx3_ASAP7_75t_L g9526 ( 
.A(n_9334),
.Y(n_9526)
);

BUFx2_ASAP7_75t_L g9527 ( 
.A(n_9334),
.Y(n_9527)
);

HB1xp67_ASAP7_75t_L g9528 ( 
.A(n_9086),
.Y(n_9528)
);

NAND2xp5_ASAP7_75t_L g9529 ( 
.A(n_8924),
.B(n_8555),
.Y(n_9529)
);

BUFx3_ASAP7_75t_L g9530 ( 
.A(n_9334),
.Y(n_9530)
);

BUFx6f_ASAP7_75t_L g9531 ( 
.A(n_9148),
.Y(n_9531)
);

INVx1_ASAP7_75t_L g9532 ( 
.A(n_9241),
.Y(n_9532)
);

AND2x2_ASAP7_75t_L g9533 ( 
.A(n_9180),
.B(n_8663),
.Y(n_9533)
);

AND2x2_ASAP7_75t_L g9534 ( 
.A(n_9180),
.B(n_8663),
.Y(n_9534)
);

INVx2_ASAP7_75t_L g9535 ( 
.A(n_9148),
.Y(n_9535)
);

HB1xp67_ASAP7_75t_L g9536 ( 
.A(n_9086),
.Y(n_9536)
);

HB1xp67_ASAP7_75t_L g9537 ( 
.A(n_9093),
.Y(n_9537)
);

AND2x2_ASAP7_75t_L g9538 ( 
.A(n_8954),
.B(n_8881),
.Y(n_9538)
);

INVx1_ASAP7_75t_L g9539 ( 
.A(n_9252),
.Y(n_9539)
);

BUFx6f_ASAP7_75t_L g9540 ( 
.A(n_9148),
.Y(n_9540)
);

INVx2_ASAP7_75t_L g9541 ( 
.A(n_9100),
.Y(n_9541)
);

AND2x2_ASAP7_75t_L g9542 ( 
.A(n_9000),
.B(n_8881),
.Y(n_9542)
);

INVx2_ASAP7_75t_L g9543 ( 
.A(n_9100),
.Y(n_9543)
);

AND2x2_ASAP7_75t_L g9544 ( 
.A(n_9009),
.B(n_8881),
.Y(n_9544)
);

INVx1_ASAP7_75t_L g9545 ( 
.A(n_9252),
.Y(n_9545)
);

NOR2xp33_ASAP7_75t_L g9546 ( 
.A(n_9299),
.B(n_8752),
.Y(n_9546)
);

INVx2_ASAP7_75t_L g9547 ( 
.A(n_9082),
.Y(n_9547)
);

AND2x2_ASAP7_75t_L g9548 ( 
.A(n_8927),
.B(n_8616),
.Y(n_9548)
);

NAND2xp5_ASAP7_75t_L g9549 ( 
.A(n_9256),
.B(n_8555),
.Y(n_9549)
);

INVx2_ASAP7_75t_L g9550 ( 
.A(n_9082),
.Y(n_9550)
);

BUFx3_ASAP7_75t_L g9551 ( 
.A(n_9125),
.Y(n_9551)
);

INVx1_ASAP7_75t_L g9552 ( 
.A(n_9256),
.Y(n_9552)
);

INVx2_ASAP7_75t_SL g9553 ( 
.A(n_9176),
.Y(n_9553)
);

AND2x2_ASAP7_75t_L g9554 ( 
.A(n_9201),
.B(n_8616),
.Y(n_9554)
);

HB1xp67_ASAP7_75t_L g9555 ( 
.A(n_9093),
.Y(n_9555)
);

AND2x2_ASAP7_75t_L g9556 ( 
.A(n_9291),
.B(n_8629),
.Y(n_9556)
);

INVx1_ASAP7_75t_L g9557 ( 
.A(n_9307),
.Y(n_9557)
);

HB1xp67_ASAP7_75t_L g9558 ( 
.A(n_9035),
.Y(n_9558)
);

INVx1_ASAP7_75t_L g9559 ( 
.A(n_9307),
.Y(n_9559)
);

AND2x4_ASAP7_75t_L g9560 ( 
.A(n_9176),
.B(n_8381),
.Y(n_9560)
);

INVx2_ASAP7_75t_L g9561 ( 
.A(n_9125),
.Y(n_9561)
);

INVx4_ASAP7_75t_L g9562 ( 
.A(n_9207),
.Y(n_9562)
);

AND2x2_ASAP7_75t_L g9563 ( 
.A(n_9303),
.B(n_8629),
.Y(n_9563)
);

INVx1_ASAP7_75t_L g9564 ( 
.A(n_9035),
.Y(n_9564)
);

OR2x2_ASAP7_75t_L g9565 ( 
.A(n_9052),
.B(n_8575),
.Y(n_9565)
);

AND2x2_ASAP7_75t_L g9566 ( 
.A(n_9329),
.B(n_8633),
.Y(n_9566)
);

AND2x4_ASAP7_75t_L g9567 ( 
.A(n_9237),
.B(n_8381),
.Y(n_9567)
);

INVx1_ASAP7_75t_L g9568 ( 
.A(n_9051),
.Y(n_9568)
);

HB1xp67_ASAP7_75t_L g9569 ( 
.A(n_9051),
.Y(n_9569)
);

INVx1_ASAP7_75t_L g9570 ( 
.A(n_8962),
.Y(n_9570)
);

INVx1_ASAP7_75t_L g9571 ( 
.A(n_8962),
.Y(n_9571)
);

AND2x2_ASAP7_75t_L g9572 ( 
.A(n_9336),
.B(n_8633),
.Y(n_9572)
);

INVx2_ASAP7_75t_SL g9573 ( 
.A(n_9200),
.Y(n_9573)
);

INVx1_ASAP7_75t_L g9574 ( 
.A(n_8968),
.Y(n_9574)
);

INVx1_ASAP7_75t_L g9575 ( 
.A(n_8968),
.Y(n_9575)
);

BUFx2_ASAP7_75t_L g9576 ( 
.A(n_9123),
.Y(n_9576)
);

AND2x4_ASAP7_75t_L g9577 ( 
.A(n_9253),
.B(n_8381),
.Y(n_9577)
);

AND2x2_ASAP7_75t_L g9578 ( 
.A(n_9305),
.B(n_8637),
.Y(n_9578)
);

AND2x2_ASAP7_75t_L g9579 ( 
.A(n_9126),
.B(n_8637),
.Y(n_9579)
);

INVx2_ASAP7_75t_L g9580 ( 
.A(n_9123),
.Y(n_9580)
);

BUFx2_ASAP7_75t_L g9581 ( 
.A(n_9153),
.Y(n_9581)
);

HB1xp67_ASAP7_75t_L g9582 ( 
.A(n_9007),
.Y(n_9582)
);

AND2x2_ASAP7_75t_L g9583 ( 
.A(n_9131),
.B(n_8414),
.Y(n_9583)
);

NAND2xp5_ASAP7_75t_L g9584 ( 
.A(n_9211),
.B(n_8369),
.Y(n_9584)
);

NAND2xp5_ASAP7_75t_L g9585 ( 
.A(n_9211),
.B(n_8369),
.Y(n_9585)
);

INVx1_ASAP7_75t_L g9586 ( 
.A(n_8973),
.Y(n_9586)
);

INVx2_ASAP7_75t_L g9587 ( 
.A(n_9153),
.Y(n_9587)
);

HB1xp67_ASAP7_75t_L g9588 ( 
.A(n_9007),
.Y(n_9588)
);

INVx2_ASAP7_75t_L g9589 ( 
.A(n_9198),
.Y(n_9589)
);

OR2x2_ASAP7_75t_L g9590 ( 
.A(n_9298),
.B(n_8579),
.Y(n_9590)
);

OR2x2_ASAP7_75t_L g9591 ( 
.A(n_9330),
.B(n_8579),
.Y(n_9591)
);

BUFx2_ASAP7_75t_L g9592 ( 
.A(n_9183),
.Y(n_9592)
);

INVx1_ASAP7_75t_L g9593 ( 
.A(n_8973),
.Y(n_9593)
);

INVx2_ASAP7_75t_L g9594 ( 
.A(n_9198),
.Y(n_9594)
);

AND2x2_ASAP7_75t_L g9595 ( 
.A(n_9141),
.B(n_8414),
.Y(n_9595)
);

AND2x2_ASAP7_75t_L g9596 ( 
.A(n_9143),
.B(n_8414),
.Y(n_9596)
);

NOR2xp33_ASAP7_75t_L g9597 ( 
.A(n_9207),
.B(n_8752),
.Y(n_9597)
);

AND2x2_ASAP7_75t_L g9598 ( 
.A(n_9396),
.B(n_8717),
.Y(n_9598)
);

AOI22xp33_ASAP7_75t_SL g9599 ( 
.A1(n_9094),
.A2(n_8811),
.B1(n_8824),
.B2(n_8853),
.Y(n_9599)
);

NOR2xp67_ASAP7_75t_L g9600 ( 
.A(n_9183),
.B(n_8917),
.Y(n_9600)
);

NAND2xp5_ASAP7_75t_L g9601 ( 
.A(n_8993),
.B(n_8375),
.Y(n_9601)
);

AOI221xp5_ASAP7_75t_L g9602 ( 
.A1(n_8981),
.A2(n_8709),
.B1(n_8876),
.B2(n_8894),
.C(n_8773),
.Y(n_9602)
);

NAND2xp5_ASAP7_75t_L g9603 ( 
.A(n_8993),
.B(n_8375),
.Y(n_9603)
);

INVx2_ASAP7_75t_L g9604 ( 
.A(n_9206),
.Y(n_9604)
);

BUFx2_ASAP7_75t_L g9605 ( 
.A(n_9340),
.Y(n_9605)
);

INVxp67_ASAP7_75t_L g9606 ( 
.A(n_9002),
.Y(n_9606)
);

INVx2_ASAP7_75t_L g9607 ( 
.A(n_9206),
.Y(n_9607)
);

INVx1_ASAP7_75t_L g9608 ( 
.A(n_9002),
.Y(n_9608)
);

INVx1_ASAP7_75t_SL g9609 ( 
.A(n_8983),
.Y(n_9609)
);

INVx2_ASAP7_75t_SL g9610 ( 
.A(n_9200),
.Y(n_9610)
);

AND2x2_ASAP7_75t_L g9611 ( 
.A(n_8925),
.B(n_8717),
.Y(n_9611)
);

AND2x2_ASAP7_75t_L g9612 ( 
.A(n_8966),
.B(n_8520),
.Y(n_9612)
);

NAND2xp5_ASAP7_75t_L g9613 ( 
.A(n_8981),
.B(n_8380),
.Y(n_9613)
);

OR2x2_ASAP7_75t_L g9614 ( 
.A(n_9369),
.B(n_9376),
.Y(n_9614)
);

INVx2_ASAP7_75t_L g9615 ( 
.A(n_9128),
.Y(n_9615)
);

INVx2_ASAP7_75t_L g9616 ( 
.A(n_9128),
.Y(n_9616)
);

AND2x2_ASAP7_75t_L g9617 ( 
.A(n_8966),
.B(n_8976),
.Y(n_9617)
);

INVx1_ASAP7_75t_L g9618 ( 
.A(n_9120),
.Y(n_9618)
);

NOR2xp33_ASAP7_75t_L g9619 ( 
.A(n_9121),
.B(n_7998),
.Y(n_9619)
);

INVx2_ASAP7_75t_L g9620 ( 
.A(n_9200),
.Y(n_9620)
);

INVx1_ASAP7_75t_L g9621 ( 
.A(n_9120),
.Y(n_9621)
);

OR2x2_ASAP7_75t_L g9622 ( 
.A(n_9089),
.B(n_9028),
.Y(n_9622)
);

INVx1_ASAP7_75t_L g9623 ( 
.A(n_9122),
.Y(n_9623)
);

NAND2xp5_ASAP7_75t_SL g9624 ( 
.A(n_9073),
.B(n_8709),
.Y(n_9624)
);

BUFx2_ASAP7_75t_L g9625 ( 
.A(n_9340),
.Y(n_9625)
);

INVx1_ASAP7_75t_L g9626 ( 
.A(n_9122),
.Y(n_9626)
);

INVx1_ASAP7_75t_L g9627 ( 
.A(n_9154),
.Y(n_9627)
);

INVx1_ASAP7_75t_L g9628 ( 
.A(n_9154),
.Y(n_9628)
);

INVx2_ASAP7_75t_L g9629 ( 
.A(n_9150),
.Y(n_9629)
);

AND2x2_ASAP7_75t_L g9630 ( 
.A(n_8976),
.B(n_8480),
.Y(n_9630)
);

NAND2xp5_ASAP7_75t_L g9631 ( 
.A(n_9133),
.B(n_8380),
.Y(n_9631)
);

INVx2_ASAP7_75t_L g9632 ( 
.A(n_9150),
.Y(n_9632)
);

NOR2xp33_ASAP7_75t_L g9633 ( 
.A(n_9121),
.B(n_7998),
.Y(n_9633)
);

OAI211xp5_ASAP7_75t_L g9634 ( 
.A1(n_9073),
.A2(n_8694),
.B(n_8913),
.C(n_8906),
.Y(n_9634)
);

AND2x4_ASAP7_75t_L g9635 ( 
.A(n_9354),
.B(n_8356),
.Y(n_9635)
);

INVx1_ASAP7_75t_L g9636 ( 
.A(n_9161),
.Y(n_9636)
);

INVx2_ASAP7_75t_L g9637 ( 
.A(n_9227),
.Y(n_9637)
);

INVx2_ASAP7_75t_L g9638 ( 
.A(n_9227),
.Y(n_9638)
);

INVx1_ASAP7_75t_L g9639 ( 
.A(n_9161),
.Y(n_9639)
);

INVx2_ASAP7_75t_L g9640 ( 
.A(n_9296),
.Y(n_9640)
);

NOR2x1_ASAP7_75t_L g9641 ( 
.A(n_9354),
.B(n_9214),
.Y(n_9641)
);

INVx3_ASAP7_75t_L g9642 ( 
.A(n_9388),
.Y(n_9642)
);

INVx1_ASAP7_75t_L g9643 ( 
.A(n_9171),
.Y(n_9643)
);

INVx1_ASAP7_75t_L g9644 ( 
.A(n_9171),
.Y(n_9644)
);

INVxp67_ASAP7_75t_L g9645 ( 
.A(n_9023),
.Y(n_9645)
);

INVx1_ASAP7_75t_L g9646 ( 
.A(n_9431),
.Y(n_9646)
);

AND2x2_ASAP7_75t_L g9647 ( 
.A(n_9160),
.B(n_8480),
.Y(n_9647)
);

INVx1_ASAP7_75t_L g9648 ( 
.A(n_9431),
.Y(n_9648)
);

AND2x2_ASAP7_75t_L g9649 ( 
.A(n_9076),
.B(n_8480),
.Y(n_9649)
);

NAND2xp5_ASAP7_75t_L g9650 ( 
.A(n_9133),
.B(n_8384),
.Y(n_9650)
);

AND2x2_ASAP7_75t_L g9651 ( 
.A(n_8953),
.B(n_8901),
.Y(n_9651)
);

AND2x2_ASAP7_75t_L g9652 ( 
.A(n_8956),
.B(n_8901),
.Y(n_9652)
);

BUFx12f_ASAP7_75t_L g9653 ( 
.A(n_9103),
.Y(n_9653)
);

INVx2_ASAP7_75t_L g9654 ( 
.A(n_9296),
.Y(n_9654)
);

NOR2x1_ASAP7_75t_SL g9655 ( 
.A(n_9350),
.B(n_8790),
.Y(n_9655)
);

NAND2x1_ASAP7_75t_L g9656 ( 
.A(n_9134),
.B(n_8742),
.Y(n_9656)
);

OR2x2_ASAP7_75t_L g9657 ( 
.A(n_9030),
.B(n_8580),
.Y(n_9657)
);

INVxp67_ASAP7_75t_SL g9658 ( 
.A(n_9033),
.Y(n_9658)
);

AND2x2_ASAP7_75t_L g9659 ( 
.A(n_9031),
.B(n_8901),
.Y(n_9659)
);

NOR2xp67_ASAP7_75t_L g9660 ( 
.A(n_9103),
.B(n_8917),
.Y(n_9660)
);

OR2x2_ASAP7_75t_L g9661 ( 
.A(n_9424),
.B(n_8580),
.Y(n_9661)
);

AND2x4_ASAP7_75t_L g9662 ( 
.A(n_9281),
.B(n_8356),
.Y(n_9662)
);

INVx1_ASAP7_75t_L g9663 ( 
.A(n_9432),
.Y(n_9663)
);

AND2x2_ASAP7_75t_L g9664 ( 
.A(n_9043),
.B(n_8743),
.Y(n_9664)
);

INVx1_ASAP7_75t_L g9665 ( 
.A(n_9432),
.Y(n_9665)
);

INVx1_ASAP7_75t_L g9666 ( 
.A(n_9443),
.Y(n_9666)
);

AND2x2_ASAP7_75t_SL g9667 ( 
.A(n_9214),
.B(n_8743),
.Y(n_9667)
);

INVx1_ASAP7_75t_L g9668 ( 
.A(n_9443),
.Y(n_9668)
);

INVx2_ASAP7_75t_L g9669 ( 
.A(n_9323),
.Y(n_9669)
);

INVx2_ASAP7_75t_L g9670 ( 
.A(n_9323),
.Y(n_9670)
);

OR2x2_ASAP7_75t_L g9671 ( 
.A(n_9172),
.B(n_8583),
.Y(n_9671)
);

INVx1_ASAP7_75t_SL g9672 ( 
.A(n_8983),
.Y(n_9672)
);

INVx1_ASAP7_75t_L g9673 ( 
.A(n_9459),
.Y(n_9673)
);

INVx2_ASAP7_75t_L g9674 ( 
.A(n_9447),
.Y(n_9674)
);

OAI22xp33_ASAP7_75t_L g9675 ( 
.A1(n_9158),
.A2(n_8756),
.B1(n_8516),
.B2(n_8527),
.Y(n_9675)
);

INVx2_ASAP7_75t_L g9676 ( 
.A(n_9447),
.Y(n_9676)
);

AND2x2_ASAP7_75t_L g9677 ( 
.A(n_9314),
.B(n_8743),
.Y(n_9677)
);

INVx2_ASAP7_75t_L g9678 ( 
.A(n_9019),
.Y(n_9678)
);

NAND2xp5_ASAP7_75t_L g9679 ( 
.A(n_9033),
.B(n_9159),
.Y(n_9679)
);

INVx2_ASAP7_75t_L g9680 ( 
.A(n_9019),
.Y(n_9680)
);

INVxp67_ASAP7_75t_SL g9681 ( 
.A(n_9019),
.Y(n_9681)
);

NAND2x1p5_ASAP7_75t_L g9682 ( 
.A(n_9281),
.B(n_8917),
.Y(n_9682)
);

INVx2_ASAP7_75t_L g9683 ( 
.A(n_9041),
.Y(n_9683)
);

INVxp67_ASAP7_75t_SL g9684 ( 
.A(n_9459),
.Y(n_9684)
);

INVx2_ASAP7_75t_L g9685 ( 
.A(n_9041),
.Y(n_9685)
);

INVx3_ASAP7_75t_L g9686 ( 
.A(n_9453),
.Y(n_9686)
);

HB1xp67_ASAP7_75t_L g9687 ( 
.A(n_9346),
.Y(n_9687)
);

AND2x2_ASAP7_75t_L g9688 ( 
.A(n_8980),
.B(n_8760),
.Y(n_9688)
);

INVx2_ASAP7_75t_L g9689 ( 
.A(n_9041),
.Y(n_9689)
);

AND2x2_ASAP7_75t_L g9690 ( 
.A(n_8986),
.B(n_8760),
.Y(n_9690)
);

AND2x2_ASAP7_75t_L g9691 ( 
.A(n_8987),
.B(n_8760),
.Y(n_9691)
);

INVx1_ASAP7_75t_L g9692 ( 
.A(n_9479),
.Y(n_9692)
);

INVx2_ASAP7_75t_L g9693 ( 
.A(n_9054),
.Y(n_9693)
);

AND2x2_ASAP7_75t_L g9694 ( 
.A(n_8989),
.B(n_8778),
.Y(n_9694)
);

AO21x2_ASAP7_75t_L g9695 ( 
.A1(n_9106),
.A2(n_8853),
.B(n_8661),
.Y(n_9695)
);

INVx1_ASAP7_75t_L g9696 ( 
.A(n_9479),
.Y(n_9696)
);

INVx1_ASAP7_75t_L g9697 ( 
.A(n_9406),
.Y(n_9697)
);

AND2x2_ASAP7_75t_L g9698 ( 
.A(n_8990),
.B(n_8778),
.Y(n_9698)
);

INVx1_ASAP7_75t_L g9699 ( 
.A(n_9406),
.Y(n_9699)
);

AND2x4_ASAP7_75t_L g9700 ( 
.A(n_9281),
.B(n_8356),
.Y(n_9700)
);

AND2x2_ASAP7_75t_L g9701 ( 
.A(n_8998),
.B(n_8778),
.Y(n_9701)
);

INVx1_ASAP7_75t_L g9702 ( 
.A(n_9421),
.Y(n_9702)
);

AND2x2_ASAP7_75t_L g9703 ( 
.A(n_9016),
.B(n_8865),
.Y(n_9703)
);

NAND2xp5_ASAP7_75t_L g9704 ( 
.A(n_9159),
.B(n_8384),
.Y(n_9704)
);

OR2x2_ASAP7_75t_L g9705 ( 
.A(n_8936),
.B(n_8583),
.Y(n_9705)
);

AND2x2_ASAP7_75t_L g9706 ( 
.A(n_9034),
.B(n_8865),
.Y(n_9706)
);

INVx1_ASAP7_75t_L g9707 ( 
.A(n_9421),
.Y(n_9707)
);

AND2x2_ASAP7_75t_L g9708 ( 
.A(n_9053),
.B(n_8605),
.Y(n_9708)
);

INVx2_ASAP7_75t_L g9709 ( 
.A(n_9447),
.Y(n_9709)
);

INVx1_ASAP7_75t_L g9710 ( 
.A(n_9346),
.Y(n_9710)
);

HB1xp67_ASAP7_75t_L g9711 ( 
.A(n_9352),
.Y(n_9711)
);

INVx3_ASAP7_75t_L g9712 ( 
.A(n_9054),
.Y(n_9712)
);

INVx1_ASAP7_75t_L g9713 ( 
.A(n_9352),
.Y(n_9713)
);

INVx1_ASAP7_75t_L g9714 ( 
.A(n_9383),
.Y(n_9714)
);

INVx1_ASAP7_75t_L g9715 ( 
.A(n_9383),
.Y(n_9715)
);

OR2x2_ASAP7_75t_L g9716 ( 
.A(n_8937),
.B(n_8935),
.Y(n_9716)
);

INVx2_ASAP7_75t_L g9717 ( 
.A(n_9447),
.Y(n_9717)
);

HB1xp67_ASAP7_75t_L g9718 ( 
.A(n_9309),
.Y(n_9718)
);

INVx2_ASAP7_75t_L g9719 ( 
.A(n_9146),
.Y(n_9719)
);

INVx1_ASAP7_75t_L g9720 ( 
.A(n_9309),
.Y(n_9720)
);

INVx1_ASAP7_75t_L g9721 ( 
.A(n_9311),
.Y(n_9721)
);

BUFx2_ASAP7_75t_L g9722 ( 
.A(n_9146),
.Y(n_9722)
);

INVx2_ASAP7_75t_L g9723 ( 
.A(n_9054),
.Y(n_9723)
);

INVx1_ASAP7_75t_L g9724 ( 
.A(n_9311),
.Y(n_9724)
);

NAND2x1_ASAP7_75t_L g9725 ( 
.A(n_9134),
.B(n_8742),
.Y(n_9725)
);

INVx1_ASAP7_75t_L g9726 ( 
.A(n_9343),
.Y(n_9726)
);

INVx1_ASAP7_75t_L g9727 ( 
.A(n_9343),
.Y(n_9727)
);

AND2x2_ASAP7_75t_L g9728 ( 
.A(n_9360),
.B(n_8605),
.Y(n_9728)
);

NAND2xp5_ASAP7_75t_L g9729 ( 
.A(n_9179),
.B(n_8395),
.Y(n_9729)
);

BUFx6f_ASAP7_75t_L g9730 ( 
.A(n_9258),
.Y(n_9730)
);

INVx3_ASAP7_75t_L g9731 ( 
.A(n_9055),
.Y(n_9731)
);

BUFx2_ASAP7_75t_L g9732 ( 
.A(n_9337),
.Y(n_9732)
);

INVx2_ASAP7_75t_SL g9733 ( 
.A(n_9124),
.Y(n_9733)
);

AND2x4_ASAP7_75t_L g9734 ( 
.A(n_9337),
.B(n_9344),
.Y(n_9734)
);

INVx2_ASAP7_75t_L g9735 ( 
.A(n_9055),
.Y(n_9735)
);

INVx2_ASAP7_75t_L g9736 ( 
.A(n_9055),
.Y(n_9736)
);

INVx1_ASAP7_75t_L g9737 ( 
.A(n_9338),
.Y(n_9737)
);

AND2x4_ASAP7_75t_L g9738 ( 
.A(n_9344),
.B(n_8607),
.Y(n_9738)
);

AND2x2_ASAP7_75t_L g9739 ( 
.A(n_9088),
.B(n_8607),
.Y(n_9739)
);

INVx2_ASAP7_75t_SL g9740 ( 
.A(n_9428),
.Y(n_9740)
);

BUFx3_ASAP7_75t_L g9741 ( 
.A(n_9379),
.Y(n_9741)
);

AND2x2_ASAP7_75t_L g9742 ( 
.A(n_9101),
.B(n_8614),
.Y(n_9742)
);

INVx2_ASAP7_75t_L g9743 ( 
.A(n_9379),
.Y(n_9743)
);

INVx1_ASAP7_75t_L g9744 ( 
.A(n_9348),
.Y(n_9744)
);

AND2x2_ASAP7_75t_L g9745 ( 
.A(n_9478),
.B(n_8614),
.Y(n_9745)
);

INVx2_ASAP7_75t_L g9746 ( 
.A(n_9391),
.Y(n_9746)
);

OR2x2_ASAP7_75t_L g9747 ( 
.A(n_9098),
.B(n_8585),
.Y(n_9747)
);

AND2x2_ASAP7_75t_L g9748 ( 
.A(n_9127),
.B(n_8863),
.Y(n_9748)
);

INVx2_ASAP7_75t_L g9749 ( 
.A(n_9391),
.Y(n_9749)
);

INVx2_ASAP7_75t_L g9750 ( 
.A(n_9407),
.Y(n_9750)
);

INVx1_ASAP7_75t_L g9751 ( 
.A(n_9355),
.Y(n_9751)
);

INVx2_ASAP7_75t_L g9752 ( 
.A(n_9407),
.Y(n_9752)
);

HB1xp67_ASAP7_75t_L g9753 ( 
.A(n_9179),
.Y(n_9753)
);

AND2x2_ASAP7_75t_L g9754 ( 
.A(n_9173),
.B(n_8863),
.Y(n_9754)
);

OR2x2_ASAP7_75t_L g9755 ( 
.A(n_9394),
.B(n_8585),
.Y(n_9755)
);

INVx2_ASAP7_75t_L g9756 ( 
.A(n_9450),
.Y(n_9756)
);

INVx2_ASAP7_75t_L g9757 ( 
.A(n_9450),
.Y(n_9757)
);

AOI22xp33_ASAP7_75t_L g9758 ( 
.A1(n_9135),
.A2(n_8811),
.B1(n_8853),
.B2(n_8406),
.Y(n_9758)
);

INVx2_ASAP7_75t_L g9759 ( 
.A(n_9458),
.Y(n_9759)
);

AND2x2_ASAP7_75t_L g9760 ( 
.A(n_9425),
.B(n_8877),
.Y(n_9760)
);

AND2x4_ASAP7_75t_L g9761 ( 
.A(n_9162),
.B(n_8788),
.Y(n_9761)
);

INVx2_ASAP7_75t_L g9762 ( 
.A(n_9458),
.Y(n_9762)
);

AND2x2_ASAP7_75t_L g9763 ( 
.A(n_9425),
.B(n_8877),
.Y(n_9763)
);

INVx1_ASAP7_75t_L g9764 ( 
.A(n_9356),
.Y(n_9764)
);

INVx1_ASAP7_75t_L g9765 ( 
.A(n_9357),
.Y(n_9765)
);

AND2x2_ASAP7_75t_L g9766 ( 
.A(n_9178),
.B(n_8834),
.Y(n_9766)
);

INVx2_ASAP7_75t_SL g9767 ( 
.A(n_9169),
.Y(n_9767)
);

AND2x2_ASAP7_75t_L g9768 ( 
.A(n_9190),
.B(n_8834),
.Y(n_9768)
);

OR2x2_ASAP7_75t_L g9769 ( 
.A(n_9394),
.B(n_8586),
.Y(n_9769)
);

INVx1_ASAP7_75t_L g9770 ( 
.A(n_9368),
.Y(n_9770)
);

INVx2_ASAP7_75t_L g9771 ( 
.A(n_9475),
.Y(n_9771)
);

AND2x4_ASAP7_75t_SL g9772 ( 
.A(n_9169),
.B(n_8790),
.Y(n_9772)
);

INVxp67_ASAP7_75t_L g9773 ( 
.A(n_8922),
.Y(n_9773)
);

INVx1_ASAP7_75t_L g9774 ( 
.A(n_9370),
.Y(n_9774)
);

INVx2_ASAP7_75t_SL g9775 ( 
.A(n_9169),
.Y(n_9775)
);

AND2x4_ASAP7_75t_L g9776 ( 
.A(n_8926),
.B(n_8794),
.Y(n_9776)
);

INVx1_ASAP7_75t_L g9777 ( 
.A(n_9371),
.Y(n_9777)
);

AND2x2_ASAP7_75t_L g9778 ( 
.A(n_9208),
.B(n_8834),
.Y(n_9778)
);

AND2x2_ASAP7_75t_L g9779 ( 
.A(n_9137),
.B(n_8679),
.Y(n_9779)
);

AND2x2_ASAP7_75t_L g9780 ( 
.A(n_9102),
.B(n_8679),
.Y(n_9780)
);

HB1xp67_ASAP7_75t_L g9781 ( 
.A(n_9395),
.Y(n_9781)
);

BUFx3_ASAP7_75t_L g9782 ( 
.A(n_9059),
.Y(n_9782)
);

AND2x2_ASAP7_75t_L g9783 ( 
.A(n_9145),
.B(n_8685),
.Y(n_9783)
);

OR2x2_ASAP7_75t_L g9784 ( 
.A(n_9395),
.B(n_8586),
.Y(n_9784)
);

NAND2xp5_ASAP7_75t_L g9785 ( 
.A(n_8923),
.B(n_8395),
.Y(n_9785)
);

AND2x2_ASAP7_75t_L g9786 ( 
.A(n_9149),
.B(n_8685),
.Y(n_9786)
);

NAND2xp5_ASAP7_75t_L g9787 ( 
.A(n_8930),
.B(n_8400),
.Y(n_9787)
);

INVx4_ASAP7_75t_L g9788 ( 
.A(n_9426),
.Y(n_9788)
);

HB1xp67_ASAP7_75t_L g9789 ( 
.A(n_9397),
.Y(n_9789)
);

INVx3_ASAP7_75t_L g9790 ( 
.A(n_9287),
.Y(n_9790)
);

NAND2xp5_ASAP7_75t_L g9791 ( 
.A(n_9270),
.B(n_8400),
.Y(n_9791)
);

OR2x2_ASAP7_75t_L g9792 ( 
.A(n_9397),
.B(n_8588),
.Y(n_9792)
);

AND2x2_ASAP7_75t_L g9793 ( 
.A(n_9204),
.B(n_8688),
.Y(n_9793)
);

AND2x2_ASAP7_75t_L g9794 ( 
.A(n_9199),
.B(n_8688),
.Y(n_9794)
);

HB1xp67_ASAP7_75t_L g9795 ( 
.A(n_9409),
.Y(n_9795)
);

NAND2xp5_ASAP7_75t_L g9796 ( 
.A(n_9061),
.B(n_8402),
.Y(n_9796)
);

INVx2_ASAP7_75t_L g9797 ( 
.A(n_8975),
.Y(n_9797)
);

BUFx2_ASAP7_75t_L g9798 ( 
.A(n_9113),
.Y(n_9798)
);

HB1xp67_ASAP7_75t_L g9799 ( 
.A(n_9409),
.Y(n_9799)
);

AO21x2_ASAP7_75t_L g9800 ( 
.A1(n_9106),
.A2(n_8661),
.B(n_8659),
.Y(n_9800)
);

INVx2_ASAP7_75t_L g9801 ( 
.A(n_8975),
.Y(n_9801)
);

AND2x2_ASAP7_75t_L g9802 ( 
.A(n_9308),
.B(n_8588),
.Y(n_9802)
);

INVx2_ASAP7_75t_L g9803 ( 
.A(n_9029),
.Y(n_9803)
);

BUFx2_ASAP7_75t_L g9804 ( 
.A(n_9139),
.Y(n_9804)
);

INVx1_ASAP7_75t_L g9805 ( 
.A(n_9381),
.Y(n_9805)
);

AND2x2_ASAP7_75t_SL g9806 ( 
.A(n_9061),
.B(n_8424),
.Y(n_9806)
);

INVx1_ASAP7_75t_L g9807 ( 
.A(n_9386),
.Y(n_9807)
);

INVx1_ASAP7_75t_L g9808 ( 
.A(n_9393),
.Y(n_9808)
);

INVx1_ASAP7_75t_L g9809 ( 
.A(n_9401),
.Y(n_9809)
);

INVx1_ASAP7_75t_L g9810 ( 
.A(n_9413),
.Y(n_9810)
);

HB1xp67_ASAP7_75t_L g9811 ( 
.A(n_9405),
.Y(n_9811)
);

AND2x2_ASAP7_75t_L g9812 ( 
.A(n_9140),
.B(n_8589),
.Y(n_9812)
);

INVx2_ASAP7_75t_L g9813 ( 
.A(n_9029),
.Y(n_9813)
);

AND2x2_ASAP7_75t_L g9814 ( 
.A(n_9130),
.B(n_9215),
.Y(n_9814)
);

INVx2_ASAP7_75t_L g9815 ( 
.A(n_9475),
.Y(n_9815)
);

AND2x2_ASAP7_75t_L g9816 ( 
.A(n_9217),
.B(n_8589),
.Y(n_9816)
);

AND2x2_ASAP7_75t_L g9817 ( 
.A(n_9105),
.B(n_9347),
.Y(n_9817)
);

HB1xp67_ASAP7_75t_L g9818 ( 
.A(n_9405),
.Y(n_9818)
);

INVx1_ASAP7_75t_L g9819 ( 
.A(n_9415),
.Y(n_9819)
);

INVx3_ASAP7_75t_L g9820 ( 
.A(n_9287),
.Y(n_9820)
);

INVx1_ASAP7_75t_L g9821 ( 
.A(n_9417),
.Y(n_9821)
);

INVx1_ASAP7_75t_L g9822 ( 
.A(n_9423),
.Y(n_9822)
);

BUFx4f_ASAP7_75t_L g9823 ( 
.A(n_9021),
.Y(n_9823)
);

INVx1_ASAP7_75t_L g9824 ( 
.A(n_9435),
.Y(n_9824)
);

INVx1_ASAP7_75t_L g9825 ( 
.A(n_9436),
.Y(n_9825)
);

AND2x2_ASAP7_75t_L g9826 ( 
.A(n_9353),
.B(n_8597),
.Y(n_9826)
);

INVx1_ASAP7_75t_L g9827 ( 
.A(n_9437),
.Y(n_9827)
);

NAND2xp5_ASAP7_75t_L g9828 ( 
.A(n_8933),
.B(n_8402),
.Y(n_9828)
);

INVx1_ASAP7_75t_L g9829 ( 
.A(n_9439),
.Y(n_9829)
);

INVx1_ASAP7_75t_L g9830 ( 
.A(n_9441),
.Y(n_9830)
);

AND2x2_ASAP7_75t_L g9831 ( 
.A(n_8961),
.B(n_8597),
.Y(n_9831)
);

INVx1_ASAP7_75t_L g9832 ( 
.A(n_9445),
.Y(n_9832)
);

OR2x2_ASAP7_75t_L g9833 ( 
.A(n_9129),
.B(n_8600),
.Y(n_9833)
);

AND2x2_ASAP7_75t_L g9834 ( 
.A(n_8971),
.B(n_8600),
.Y(n_9834)
);

OR2x2_ASAP7_75t_L g9835 ( 
.A(n_8958),
.B(n_8602),
.Y(n_9835)
);

INVx2_ASAP7_75t_L g9836 ( 
.A(n_9235),
.Y(n_9836)
);

OR2x2_ASAP7_75t_L g9837 ( 
.A(n_8999),
.B(n_8602),
.Y(n_9837)
);

INVx3_ASAP7_75t_L g9838 ( 
.A(n_9287),
.Y(n_9838)
);

BUFx2_ASAP7_75t_L g9839 ( 
.A(n_9147),
.Y(n_9839)
);

CKINVDCx5p33_ASAP7_75t_R g9840 ( 
.A(n_9278),
.Y(n_9840)
);

OR2x2_ASAP7_75t_L g9841 ( 
.A(n_9193),
.B(n_8847),
.Y(n_9841)
);

AO21x2_ASAP7_75t_L g9842 ( 
.A1(n_9209),
.A2(n_8666),
.B(n_8659),
.Y(n_9842)
);

INVx2_ASAP7_75t_L g9843 ( 
.A(n_9426),
.Y(n_9843)
);

INVx2_ASAP7_75t_SL g9844 ( 
.A(n_9350),
.Y(n_9844)
);

INVx2_ASAP7_75t_L g9845 ( 
.A(n_9259),
.Y(n_9845)
);

INVx2_ASAP7_75t_SL g9846 ( 
.A(n_8926),
.Y(n_9846)
);

OR2x2_ASAP7_75t_L g9847 ( 
.A(n_8957),
.B(n_9410),
.Y(n_9847)
);

NAND2xp5_ASAP7_75t_L g9848 ( 
.A(n_8933),
.B(n_8404),
.Y(n_9848)
);

INVx1_ASAP7_75t_L g9849 ( 
.A(n_9449),
.Y(n_9849)
);

AND2x2_ASAP7_75t_L g9850 ( 
.A(n_9219),
.B(n_8796),
.Y(n_9850)
);

INVx1_ASAP7_75t_L g9851 ( 
.A(n_9452),
.Y(n_9851)
);

INVx1_ASAP7_75t_L g9852 ( 
.A(n_9462),
.Y(n_9852)
);

AND2x2_ASAP7_75t_L g9853 ( 
.A(n_9468),
.B(n_9481),
.Y(n_9853)
);

AND2x2_ASAP7_75t_L g9854 ( 
.A(n_8932),
.B(n_8797),
.Y(n_9854)
);

INVx2_ASAP7_75t_L g9855 ( 
.A(n_9259),
.Y(n_9855)
);

OAI33xp33_ASAP7_75t_L g9856 ( 
.A1(n_8991),
.A2(n_8631),
.A3(n_8509),
.B1(n_8749),
.B2(n_8800),
.B3(n_8799),
.Y(n_9856)
);

INVx1_ASAP7_75t_L g9857 ( 
.A(n_9465),
.Y(n_9857)
);

AOI22xp33_ASAP7_75t_SL g9858 ( 
.A1(n_9260),
.A2(n_8894),
.B1(n_8406),
.B2(n_8424),
.Y(n_9858)
);

INVx1_ASAP7_75t_L g9859 ( 
.A(n_9469),
.Y(n_9859)
);

INVx2_ASAP7_75t_L g9860 ( 
.A(n_9280),
.Y(n_9860)
);

AND2x2_ASAP7_75t_L g9861 ( 
.A(n_9342),
.B(n_8794),
.Y(n_9861)
);

INVx3_ASAP7_75t_L g9862 ( 
.A(n_9332),
.Y(n_9862)
);

NAND2xp5_ASAP7_75t_L g9863 ( 
.A(n_9471),
.B(n_8404),
.Y(n_9863)
);

NAND2xp5_ASAP7_75t_L g9864 ( 
.A(n_9471),
.B(n_8418),
.Y(n_9864)
);

INVx1_ASAP7_75t_L g9865 ( 
.A(n_9470),
.Y(n_9865)
);

INVx4_ASAP7_75t_L g9866 ( 
.A(n_9083),
.Y(n_9866)
);

OR2x6_ASAP7_75t_L g9867 ( 
.A(n_9083),
.B(n_8774),
.Y(n_9867)
);

INVx3_ASAP7_75t_L g9868 ( 
.A(n_9332),
.Y(n_9868)
);

NAND2xp5_ASAP7_75t_L g9869 ( 
.A(n_9472),
.B(n_8418),
.Y(n_9869)
);

INVx2_ASAP7_75t_SL g9870 ( 
.A(n_8938),
.Y(n_9870)
);

AND2x2_ASAP7_75t_L g9871 ( 
.A(n_9164),
.B(n_8691),
.Y(n_9871)
);

OR2x2_ASAP7_75t_L g9872 ( 
.A(n_9374),
.B(n_8582),
.Y(n_9872)
);

NOR2xp33_ASAP7_75t_R g9873 ( 
.A(n_9147),
.B(n_8008),
.Y(n_9873)
);

INVx2_ASAP7_75t_SL g9874 ( 
.A(n_8938),
.Y(n_9874)
);

AND2x2_ASAP7_75t_L g9875 ( 
.A(n_9175),
.B(n_8691),
.Y(n_9875)
);

AND2x2_ASAP7_75t_L g9876 ( 
.A(n_9328),
.B(n_8697),
.Y(n_9876)
);

AND2x2_ASAP7_75t_L g9877 ( 
.A(n_9174),
.B(n_8697),
.Y(n_9877)
);

INVx1_ASAP7_75t_L g9878 ( 
.A(n_9477),
.Y(n_9878)
);

OAI31xp33_ASAP7_75t_SL g9879 ( 
.A1(n_9209),
.A2(n_8903),
.A3(n_8916),
.B(n_8896),
.Y(n_9879)
);

INVx2_ASAP7_75t_L g9880 ( 
.A(n_9036),
.Y(n_9880)
);

INVx3_ASAP7_75t_L g9881 ( 
.A(n_9332),
.Y(n_9881)
);

BUFx2_ASAP7_75t_L g9882 ( 
.A(n_9147),
.Y(n_9882)
);

INVx2_ASAP7_75t_L g9883 ( 
.A(n_9036),
.Y(n_9883)
);

AOI22xp33_ASAP7_75t_L g9884 ( 
.A1(n_9085),
.A2(n_8406),
.B1(n_8409),
.B2(n_8424),
.Y(n_9884)
);

INVx1_ASAP7_75t_L g9885 ( 
.A(n_9480),
.Y(n_9885)
);

INVx2_ASAP7_75t_L g9886 ( 
.A(n_9038),
.Y(n_9886)
);

INVx2_ASAP7_75t_L g9887 ( 
.A(n_9038),
.Y(n_9887)
);

INVx1_ASAP7_75t_L g9888 ( 
.A(n_8939),
.Y(n_9888)
);

INVx1_ASAP7_75t_L g9889 ( 
.A(n_8942),
.Y(n_9889)
);

INVx2_ASAP7_75t_L g9890 ( 
.A(n_9042),
.Y(n_9890)
);

AND2x2_ASAP7_75t_L g9891 ( 
.A(n_9361),
.B(n_8928),
.Y(n_9891)
);

INVx1_ASAP7_75t_L g9892 ( 
.A(n_8946),
.Y(n_9892)
);

NAND2xp5_ASAP7_75t_L g9893 ( 
.A(n_9472),
.B(n_8422),
.Y(n_9893)
);

INVx1_ASAP7_75t_L g9894 ( 
.A(n_8952),
.Y(n_9894)
);

AO21x2_ASAP7_75t_L g9895 ( 
.A1(n_9080),
.A2(n_8678),
.B(n_8666),
.Y(n_9895)
);

HB1xp67_ASAP7_75t_L g9896 ( 
.A(n_9042),
.Y(n_9896)
);

AND2x2_ASAP7_75t_L g9897 ( 
.A(n_9306),
.B(n_8678),
.Y(n_9897)
);

AND2x2_ASAP7_75t_L g9898 ( 
.A(n_9282),
.B(n_8680),
.Y(n_9898)
);

AND2x2_ASAP7_75t_L g9899 ( 
.A(n_9293),
.B(n_8680),
.Y(n_9899)
);

AND2x4_ASAP7_75t_L g9900 ( 
.A(n_8943),
.B(n_8683),
.Y(n_9900)
);

AND2x2_ASAP7_75t_L g9901 ( 
.A(n_8931),
.B(n_9351),
.Y(n_9901)
);

AOI22xp5_ASAP7_75t_L g9902 ( 
.A1(n_9167),
.A2(n_8409),
.B1(n_8771),
.B2(n_8907),
.Y(n_9902)
);

AND2x4_ASAP7_75t_L g9903 ( 
.A(n_8943),
.B(n_8683),
.Y(n_9903)
);

INVx1_ASAP7_75t_L g9904 ( 
.A(n_8955),
.Y(n_9904)
);

INVx2_ASAP7_75t_L g9905 ( 
.A(n_9045),
.Y(n_9905)
);

INVx1_ASAP7_75t_L g9906 ( 
.A(n_8959),
.Y(n_9906)
);

INVx1_ASAP7_75t_L g9907 ( 
.A(n_8963),
.Y(n_9907)
);

BUFx2_ASAP7_75t_L g9908 ( 
.A(n_9147),
.Y(n_9908)
);

BUFx5_ASAP7_75t_L g9909 ( 
.A(n_9147),
.Y(n_9909)
);

AND2x2_ASAP7_75t_L g9910 ( 
.A(n_9351),
.B(n_8684),
.Y(n_9910)
);

AND2x2_ASAP7_75t_L g9911 ( 
.A(n_9325),
.B(n_8684),
.Y(n_9911)
);

INVx1_ASAP7_75t_L g9912 ( 
.A(n_8965),
.Y(n_9912)
);

AND2x2_ASAP7_75t_L g9913 ( 
.A(n_9451),
.B(n_8687),
.Y(n_9913)
);

AND2x2_ASAP7_75t_L g9914 ( 
.A(n_9077),
.B(n_8687),
.Y(n_9914)
);

OR2x2_ASAP7_75t_L g9915 ( 
.A(n_9374),
.B(n_8422),
.Y(n_9915)
);

AND2x2_ASAP7_75t_L g9916 ( 
.A(n_9078),
.B(n_8692),
.Y(n_9916)
);

OR2x2_ASAP7_75t_L g9917 ( 
.A(n_9375),
.B(n_8425),
.Y(n_9917)
);

AND2x4_ASAP7_75t_L g9918 ( 
.A(n_8944),
.B(n_8692),
.Y(n_9918)
);

AOI22xp33_ASAP7_75t_L g9919 ( 
.A1(n_9085),
.A2(n_8409),
.B1(n_8907),
.B2(n_8771),
.Y(n_9919)
);

NAND2xp5_ASAP7_75t_L g9920 ( 
.A(n_9466),
.B(n_8425),
.Y(n_9920)
);

OR2x2_ASAP7_75t_L g9921 ( 
.A(n_9375),
.B(n_8429),
.Y(n_9921)
);

AND2x2_ASAP7_75t_L g9922 ( 
.A(n_9482),
.B(n_8718),
.Y(n_9922)
);

BUFx3_ASAP7_75t_L g9923 ( 
.A(n_9367),
.Y(n_9923)
);

AND2x2_ASAP7_75t_L g9924 ( 
.A(n_9403),
.B(n_8718),
.Y(n_9924)
);

INVx1_ASAP7_75t_L g9925 ( 
.A(n_8967),
.Y(n_9925)
);

INVx2_ASAP7_75t_SL g9926 ( 
.A(n_8944),
.Y(n_9926)
);

AND2x2_ASAP7_75t_L g9927 ( 
.A(n_9414),
.B(n_8719),
.Y(n_9927)
);

INVx2_ASAP7_75t_L g9928 ( 
.A(n_9045),
.Y(n_9928)
);

INVx2_ASAP7_75t_L g9929 ( 
.A(n_9385),
.Y(n_9929)
);

AND2x2_ASAP7_75t_L g9930 ( 
.A(n_9418),
.B(n_8719),
.Y(n_9930)
);

INVx1_ASAP7_75t_L g9931 ( 
.A(n_8972),
.Y(n_9931)
);

AND2x2_ASAP7_75t_L g9932 ( 
.A(n_9191),
.B(n_8730),
.Y(n_9932)
);

INVx2_ASAP7_75t_L g9933 ( 
.A(n_9385),
.Y(n_9933)
);

INVx2_ASAP7_75t_L g9934 ( 
.A(n_9390),
.Y(n_9934)
);

INVx2_ASAP7_75t_L g9935 ( 
.A(n_9390),
.Y(n_9935)
);

BUFx2_ASAP7_75t_L g9936 ( 
.A(n_9389),
.Y(n_9936)
);

BUFx2_ASAP7_75t_L g9937 ( 
.A(n_9144),
.Y(n_9937)
);

INVx1_ASAP7_75t_L g9938 ( 
.A(n_8974),
.Y(n_9938)
);

INVx2_ASAP7_75t_L g9939 ( 
.A(n_9349),
.Y(n_9939)
);

NOR2x1_ASAP7_75t_L g9940 ( 
.A(n_9046),
.B(n_8730),
.Y(n_9940)
);

OR2x2_ASAP7_75t_L g9941 ( 
.A(n_8992),
.B(n_8429),
.Y(n_9941)
);

OR2x2_ASAP7_75t_L g9942 ( 
.A(n_9027),
.B(n_8438),
.Y(n_9942)
);

INVx1_ASAP7_75t_L g9943 ( 
.A(n_8977),
.Y(n_9943)
);

AND2x2_ASAP7_75t_L g9944 ( 
.A(n_9192),
.B(n_8734),
.Y(n_9944)
);

HB1xp67_ASAP7_75t_L g9945 ( 
.A(n_9466),
.Y(n_9945)
);

AOI22xp33_ASAP7_75t_L g9946 ( 
.A1(n_9070),
.A2(n_8907),
.B1(n_8771),
.B2(n_8448),
.Y(n_9946)
);

INVx1_ASAP7_75t_L g9947 ( 
.A(n_8978),
.Y(n_9947)
);

AND2x2_ASAP7_75t_L g9948 ( 
.A(n_9398),
.B(n_8734),
.Y(n_9948)
);

INVx1_ASAP7_75t_L g9949 ( 
.A(n_8979),
.Y(n_9949)
);

AND2x2_ASAP7_75t_L g9950 ( 
.A(n_9404),
.B(n_8740),
.Y(n_9950)
);

AND2x2_ASAP7_75t_L g9951 ( 
.A(n_9362),
.B(n_8740),
.Y(n_9951)
);

BUFx3_ASAP7_75t_L g9952 ( 
.A(n_9144),
.Y(n_9952)
);

NAND2xp5_ASAP7_75t_L g9953 ( 
.A(n_9467),
.B(n_8438),
.Y(n_9953)
);

INVx1_ASAP7_75t_L g9954 ( 
.A(n_8984),
.Y(n_9954)
);

INVx2_ASAP7_75t_L g9955 ( 
.A(n_9349),
.Y(n_9955)
);

OAI22xp5_ASAP7_75t_L g9956 ( 
.A1(n_9070),
.A2(n_8005),
.B1(n_7970),
.B2(n_7972),
.Y(n_9956)
);

INVx2_ASAP7_75t_L g9957 ( 
.A(n_9349),
.Y(n_9957)
);

INVx2_ASAP7_75t_L g9958 ( 
.A(n_9504),
.Y(n_9958)
);

INVxp67_ASAP7_75t_L g9959 ( 
.A(n_9619),
.Y(n_9959)
);

AND2x2_ASAP7_75t_L g9960 ( 
.A(n_9501),
.B(n_9362),
.Y(n_9960)
);

AND2x2_ASAP7_75t_L g9961 ( 
.A(n_9503),
.B(n_9333),
.Y(n_9961)
);

INVx1_ASAP7_75t_L g9962 ( 
.A(n_9582),
.Y(n_9962)
);

NAND2x1p5_ASAP7_75t_L g9963 ( 
.A(n_9494),
.B(n_9058),
.Y(n_9963)
);

INVx1_ASAP7_75t_L g9964 ( 
.A(n_9582),
.Y(n_9964)
);

NAND2xp5_ASAP7_75t_L g9965 ( 
.A(n_9483),
.B(n_9157),
.Y(n_9965)
);

NAND4xp25_ASAP7_75t_SL g9966 ( 
.A(n_9858),
.B(n_8997),
.C(n_8941),
.D(n_9132),
.Y(n_9966)
);

AND2x2_ASAP7_75t_L g9967 ( 
.A(n_9488),
.B(n_9493),
.Y(n_9967)
);

AND2x2_ASAP7_75t_L g9968 ( 
.A(n_9556),
.B(n_9317),
.Y(n_9968)
);

AND2x4_ASAP7_75t_SL g9969 ( 
.A(n_9494),
.B(n_9157),
.Y(n_9969)
);

INVx1_ASAP7_75t_L g9970 ( 
.A(n_9588),
.Y(n_9970)
);

INVx2_ASAP7_75t_L g9971 ( 
.A(n_9504),
.Y(n_9971)
);

AND2x4_ASAP7_75t_L g9972 ( 
.A(n_9504),
.B(n_9467),
.Y(n_9972)
);

INVx1_ASAP7_75t_L g9973 ( 
.A(n_9588),
.Y(n_9973)
);

AND2x2_ASAP7_75t_SL g9974 ( 
.A(n_9667),
.B(n_9806),
.Y(n_9974)
);

INVx1_ASAP7_75t_L g9975 ( 
.A(n_9658),
.Y(n_9975)
);

NAND2xp5_ASAP7_75t_L g9976 ( 
.A(n_9483),
.B(n_9473),
.Y(n_9976)
);

AND2x4_ASAP7_75t_SL g9977 ( 
.A(n_9562),
.B(n_9420),
.Y(n_9977)
);

AND2x4_ASAP7_75t_L g9978 ( 
.A(n_9504),
.B(n_9473),
.Y(n_9978)
);

INVx1_ASAP7_75t_L g9979 ( 
.A(n_9658),
.Y(n_9979)
);

HB1xp67_ASAP7_75t_L g9980 ( 
.A(n_9558),
.Y(n_9980)
);

INVx1_ASAP7_75t_L g9981 ( 
.A(n_9684),
.Y(n_9981)
);

AND2x2_ASAP7_75t_L g9982 ( 
.A(n_9563),
.B(n_9223),
.Y(n_9982)
);

OR2x2_ASAP7_75t_L g9983 ( 
.A(n_9484),
.B(n_9003),
.Y(n_9983)
);

AND2x2_ASAP7_75t_L g9984 ( 
.A(n_9566),
.B(n_9339),
.Y(n_9984)
);

INVx1_ASAP7_75t_L g9985 ( 
.A(n_9684),
.Y(n_9985)
);

INVx2_ASAP7_75t_L g9986 ( 
.A(n_9682),
.Y(n_9986)
);

NOR3xp33_ASAP7_75t_L g9987 ( 
.A(n_9624),
.B(n_9048),
.C(n_9167),
.Y(n_9987)
);

AND2x2_ASAP7_75t_L g9988 ( 
.A(n_9572),
.B(n_9419),
.Y(n_9988)
);

INVxp67_ASAP7_75t_SL g9989 ( 
.A(n_9558),
.Y(n_9989)
);

HB1xp67_ASAP7_75t_L g9990 ( 
.A(n_9569),
.Y(n_9990)
);

NAND3xp33_ASAP7_75t_L g9991 ( 
.A(n_9858),
.B(n_9132),
.C(n_9392),
.Y(n_9991)
);

AND2x2_ASAP7_75t_L g9992 ( 
.A(n_9853),
.B(n_9429),
.Y(n_9992)
);

HB1xp67_ASAP7_75t_L g9993 ( 
.A(n_9569),
.Y(n_9993)
);

INVx2_ASAP7_75t_L g9994 ( 
.A(n_9682),
.Y(n_9994)
);

BUFx2_ASAP7_75t_L g9995 ( 
.A(n_9653),
.Y(n_9995)
);

INVx3_ASAP7_75t_L g9996 ( 
.A(n_9531),
.Y(n_9996)
);

NAND2xp5_ASAP7_75t_L g9997 ( 
.A(n_9484),
.B(n_9060),
.Y(n_9997)
);

AND2x2_ASAP7_75t_L g9998 ( 
.A(n_9527),
.B(n_9442),
.Y(n_9998)
);

AND2x4_ASAP7_75t_L g9999 ( 
.A(n_9712),
.B(n_9420),
.Y(n_9999)
);

HB1xp67_ASAP7_75t_L g10000 ( 
.A(n_9895),
.Y(n_10000)
);

INVx3_ASAP7_75t_R g10001 ( 
.A(n_9592),
.Y(n_10001)
);

NAND2xp5_ASAP7_75t_L g10002 ( 
.A(n_9486),
.B(n_9039),
.Y(n_10002)
);

NAND2xp5_ASAP7_75t_L g10003 ( 
.A(n_9486),
.B(n_9476),
.Y(n_10003)
);

NAND2xp5_ASAP7_75t_L g10004 ( 
.A(n_9767),
.B(n_9438),
.Y(n_10004)
);

AND2x2_ASAP7_75t_L g10005 ( 
.A(n_9578),
.B(n_9448),
.Y(n_10005)
);

AND2x2_ASAP7_75t_L g10006 ( 
.A(n_9611),
.B(n_9243),
.Y(n_10006)
);

NAND2xp5_ASAP7_75t_L g10007 ( 
.A(n_9775),
.B(n_9438),
.Y(n_10007)
);

INVx1_ASAP7_75t_L g10008 ( 
.A(n_9687),
.Y(n_10008)
);

OR2x2_ASAP7_75t_L g10009 ( 
.A(n_9613),
.B(n_9181),
.Y(n_10009)
);

NAND2xp5_ASAP7_75t_L g10010 ( 
.A(n_9814),
.B(n_8945),
.Y(n_10010)
);

NOR3xp33_ASAP7_75t_L g10011 ( 
.A(n_9624),
.B(n_9422),
.C(n_9319),
.Y(n_10011)
);

OR2x2_ASAP7_75t_L g10012 ( 
.A(n_9613),
.B(n_8947),
.Y(n_10012)
);

INVx2_ASAP7_75t_L g10013 ( 
.A(n_9531),
.Y(n_10013)
);

INVx2_ASAP7_75t_L g10014 ( 
.A(n_9531),
.Y(n_10014)
);

OR2x2_ASAP7_75t_L g10015 ( 
.A(n_9509),
.B(n_9416),
.Y(n_10015)
);

NAND2xp5_ASAP7_75t_L g10016 ( 
.A(n_9730),
.B(n_8945),
.Y(n_10016)
);

HB1xp67_ASAP7_75t_L g10017 ( 
.A(n_9895),
.Y(n_10017)
);

OR2x6_ASAP7_75t_L g10018 ( 
.A(n_9562),
.B(n_9722),
.Y(n_10018)
);

OR2x2_ASAP7_75t_L g10019 ( 
.A(n_9835),
.B(n_9444),
.Y(n_10019)
);

AND2x4_ASAP7_75t_L g10020 ( 
.A(n_9712),
.B(n_9046),
.Y(n_10020)
);

INVxp67_ASAP7_75t_SL g10021 ( 
.A(n_9773),
.Y(n_10021)
);

NAND2xp5_ASAP7_75t_L g10022 ( 
.A(n_9730),
.B(n_8950),
.Y(n_10022)
);

INVx1_ASAP7_75t_L g10023 ( 
.A(n_9687),
.Y(n_10023)
);

OR2x2_ASAP7_75t_L g10024 ( 
.A(n_9837),
.B(n_9232),
.Y(n_10024)
);

AND2x2_ASAP7_75t_L g10025 ( 
.A(n_9609),
.B(n_9245),
.Y(n_10025)
);

NAND2xp5_ASAP7_75t_L g10026 ( 
.A(n_9730),
.B(n_8950),
.Y(n_10026)
);

NAND2xp5_ASAP7_75t_L g10027 ( 
.A(n_9936),
.B(n_8960),
.Y(n_10027)
);

INVx1_ASAP7_75t_L g10028 ( 
.A(n_9711),
.Y(n_10028)
);

NAND2xp5_ASAP7_75t_L g10029 ( 
.A(n_9732),
.B(n_8960),
.Y(n_10029)
);

AND2x4_ASAP7_75t_L g10030 ( 
.A(n_9731),
.B(n_9662),
.Y(n_10030)
);

INVx2_ASAP7_75t_L g10031 ( 
.A(n_9540),
.Y(n_10031)
);

AND2x2_ASAP7_75t_L g10032 ( 
.A(n_9609),
.B(n_9262),
.Y(n_10032)
);

AND2x2_ASAP7_75t_L g10033 ( 
.A(n_9672),
.B(n_9274),
.Y(n_10033)
);

NAND2xp5_ASAP7_75t_L g10034 ( 
.A(n_9525),
.B(n_8964),
.Y(n_10034)
);

INVx1_ASAP7_75t_L g10035 ( 
.A(n_9711),
.Y(n_10035)
);

NAND2xp5_ASAP7_75t_L g10036 ( 
.A(n_9535),
.B(n_8964),
.Y(n_10036)
);

OR2x2_ASAP7_75t_L g10037 ( 
.A(n_9798),
.B(n_9197),
.Y(n_10037)
);

NOR2xp33_ASAP7_75t_L g10038 ( 
.A(n_9672),
.B(n_8008),
.Y(n_10038)
);

NAND2xp5_ASAP7_75t_L g10039 ( 
.A(n_9629),
.B(n_8969),
.Y(n_10039)
);

INVx2_ASAP7_75t_L g10040 ( 
.A(n_9540),
.Y(n_10040)
);

NAND3xp33_ASAP7_75t_L g10041 ( 
.A(n_9879),
.B(n_9365),
.C(n_9138),
.Y(n_10041)
);

INVx1_ASAP7_75t_L g10042 ( 
.A(n_9718),
.Y(n_10042)
);

AND2x2_ASAP7_75t_L g10043 ( 
.A(n_9598),
.B(n_9276),
.Y(n_10043)
);

INVx1_ASAP7_75t_L g10044 ( 
.A(n_9718),
.Y(n_10044)
);

INVx1_ASAP7_75t_L g10045 ( 
.A(n_9811),
.Y(n_10045)
);

INVx1_ASAP7_75t_L g10046 ( 
.A(n_9811),
.Y(n_10046)
);

AND2x2_ASAP7_75t_L g10047 ( 
.A(n_9554),
.B(n_9372),
.Y(n_10047)
);

INVx1_ASAP7_75t_L g10048 ( 
.A(n_9818),
.Y(n_10048)
);

AND2x2_ASAP7_75t_L g10049 ( 
.A(n_9508),
.B(n_9380),
.Y(n_10049)
);

INVx1_ASAP7_75t_L g10050 ( 
.A(n_9818),
.Y(n_10050)
);

AND2x2_ASAP7_75t_L g10051 ( 
.A(n_9901),
.B(n_9400),
.Y(n_10051)
);

AND2x4_ASAP7_75t_L g10052 ( 
.A(n_9731),
.B(n_9047),
.Y(n_10052)
);

INVx1_ASAP7_75t_L g10053 ( 
.A(n_9896),
.Y(n_10053)
);

INVx1_ASAP7_75t_L g10054 ( 
.A(n_9896),
.Y(n_10054)
);

INVx2_ASAP7_75t_L g10055 ( 
.A(n_9540),
.Y(n_10055)
);

INVx2_ASAP7_75t_L g10056 ( 
.A(n_9642),
.Y(n_10056)
);

INVx1_ASAP7_75t_L g10057 ( 
.A(n_9945),
.Y(n_10057)
);

AND2x2_ASAP7_75t_L g10058 ( 
.A(n_9495),
.B(n_9402),
.Y(n_10058)
);

INVx2_ASAP7_75t_L g10059 ( 
.A(n_9642),
.Y(n_10059)
);

AND2x2_ASAP7_75t_L g10060 ( 
.A(n_9677),
.B(n_9548),
.Y(n_10060)
);

INVx1_ASAP7_75t_L g10061 ( 
.A(n_9945),
.Y(n_10061)
);

AND2x2_ASAP7_75t_L g10062 ( 
.A(n_9533),
.B(n_9320),
.Y(n_10062)
);

INVx2_ASAP7_75t_L g10063 ( 
.A(n_9686),
.Y(n_10063)
);

AND2x2_ASAP7_75t_L g10064 ( 
.A(n_9534),
.B(n_9320),
.Y(n_10064)
);

INVx1_ASAP7_75t_L g10065 ( 
.A(n_9781),
.Y(n_10065)
);

INVx1_ASAP7_75t_L g10066 ( 
.A(n_9781),
.Y(n_10066)
);

AND2x2_ASAP7_75t_L g10067 ( 
.A(n_9688),
.B(n_9326),
.Y(n_10067)
);

NOR2xp33_ASAP7_75t_L g10068 ( 
.A(n_9619),
.B(n_8017),
.Y(n_10068)
);

NAND2xp5_ASAP7_75t_SL g10069 ( 
.A(n_9806),
.B(n_9210),
.Y(n_10069)
);

AND2x4_ASAP7_75t_L g10070 ( 
.A(n_9662),
.B(n_9047),
.Y(n_10070)
);

INVx2_ASAP7_75t_L g10071 ( 
.A(n_9686),
.Y(n_10071)
);

INVx2_ASAP7_75t_L g10072 ( 
.A(n_9576),
.Y(n_10072)
);

INVx1_ASAP7_75t_L g10073 ( 
.A(n_9789),
.Y(n_10073)
);

AND2x2_ASAP7_75t_L g10074 ( 
.A(n_9690),
.B(n_9691),
.Y(n_10074)
);

AND2x2_ASAP7_75t_L g10075 ( 
.A(n_9694),
.B(n_9326),
.Y(n_10075)
);

AND2x2_ASAP7_75t_L g10076 ( 
.A(n_9698),
.B(n_9701),
.Y(n_10076)
);

INVx1_ASAP7_75t_L g10077 ( 
.A(n_9789),
.Y(n_10077)
);

AND2x4_ASAP7_75t_L g10078 ( 
.A(n_9700),
.B(n_9050),
.Y(n_10078)
);

AND2x2_ASAP7_75t_SL g10079 ( 
.A(n_9667),
.B(n_9188),
.Y(n_10079)
);

AND2x2_ASAP7_75t_L g10080 ( 
.A(n_9526),
.B(n_9331),
.Y(n_10080)
);

OR2x2_ASAP7_75t_L g10081 ( 
.A(n_9804),
.B(n_9456),
.Y(n_10081)
);

INVx1_ASAP7_75t_L g10082 ( 
.A(n_9795),
.Y(n_10082)
);

INVx2_ASAP7_75t_SL g10083 ( 
.A(n_9772),
.Y(n_10083)
);

INVx1_ASAP7_75t_L g10084 ( 
.A(n_9795),
.Y(n_10084)
);

AND2x4_ASAP7_75t_L g10085 ( 
.A(n_9700),
.B(n_9050),
.Y(n_10085)
);

AND2x2_ASAP7_75t_L g10086 ( 
.A(n_9526),
.B(n_9331),
.Y(n_10086)
);

NOR2xp33_ASAP7_75t_L g10087 ( 
.A(n_9633),
.B(n_8017),
.Y(n_10087)
);

INVx2_ASAP7_75t_L g10088 ( 
.A(n_9581),
.Y(n_10088)
);

INVx1_ASAP7_75t_L g10089 ( 
.A(n_9799),
.Y(n_10089)
);

INVx2_ASAP7_75t_L g10090 ( 
.A(n_9551),
.Y(n_10090)
);

INVx2_ASAP7_75t_L g10091 ( 
.A(n_9551),
.Y(n_10091)
);

INVx1_ASAP7_75t_L g10092 ( 
.A(n_9799),
.Y(n_10092)
);

NAND2xp5_ASAP7_75t_L g10093 ( 
.A(n_9632),
.B(n_8969),
.Y(n_10093)
);

INVx1_ASAP7_75t_L g10094 ( 
.A(n_9513),
.Y(n_10094)
);

INVx1_ASAP7_75t_L g10095 ( 
.A(n_9513),
.Y(n_10095)
);

INVx1_ASAP7_75t_L g10096 ( 
.A(n_9528),
.Y(n_10096)
);

NAND2x1p5_ASAP7_75t_L g10097 ( 
.A(n_9500),
.B(n_9660),
.Y(n_10097)
);

NAND2xp33_ASAP7_75t_SL g10098 ( 
.A(n_9873),
.B(n_9026),
.Y(n_10098)
);

OR2x2_ASAP7_75t_L g10099 ( 
.A(n_9645),
.B(n_9457),
.Y(n_10099)
);

AND2x2_ASAP7_75t_L g10100 ( 
.A(n_9530),
.B(n_9345),
.Y(n_10100)
);

NAND2xp5_ASAP7_75t_L g10101 ( 
.A(n_9844),
.B(n_8970),
.Y(n_10101)
);

HB1xp67_ASAP7_75t_L g10102 ( 
.A(n_9940),
.Y(n_10102)
);

AND2x4_ASAP7_75t_L g10103 ( 
.A(n_9492),
.B(n_9065),
.Y(n_10103)
);

INVx1_ASAP7_75t_L g10104 ( 
.A(n_9528),
.Y(n_10104)
);

AND2x2_ASAP7_75t_L g10105 ( 
.A(n_9530),
.B(n_9345),
.Y(n_10105)
);

AND2x2_ASAP7_75t_L g10106 ( 
.A(n_9583),
.B(n_9363),
.Y(n_10106)
);

NAND2xp5_ASAP7_75t_SL g10107 ( 
.A(n_9902),
.B(n_9422),
.Y(n_10107)
);

INVx2_ASAP7_75t_L g10108 ( 
.A(n_9867),
.Y(n_10108)
);

AND2x2_ASAP7_75t_L g10109 ( 
.A(n_9617),
.B(n_9363),
.Y(n_10109)
);

INVx1_ASAP7_75t_L g10110 ( 
.A(n_9536),
.Y(n_10110)
);

NAND2xp5_ASAP7_75t_L g10111 ( 
.A(n_9674),
.B(n_8970),
.Y(n_10111)
);

HB1xp67_ASAP7_75t_L g10112 ( 
.A(n_9867),
.Y(n_10112)
);

OR2x2_ASAP7_75t_L g10113 ( 
.A(n_9645),
.B(n_9408),
.Y(n_10113)
);

AND2x2_ASAP7_75t_L g10114 ( 
.A(n_9659),
.B(n_9366),
.Y(n_10114)
);

AND2x2_ASAP7_75t_L g10115 ( 
.A(n_9538),
.B(n_9366),
.Y(n_10115)
);

INVx1_ASAP7_75t_L g10116 ( 
.A(n_9536),
.Y(n_10116)
);

INVx3_ASAP7_75t_L g10117 ( 
.A(n_9560),
.Y(n_10117)
);

BUFx6f_ASAP7_75t_L g10118 ( 
.A(n_9492),
.Y(n_10118)
);

INVx1_ASAP7_75t_L g10119 ( 
.A(n_9537),
.Y(n_10119)
);

INVx1_ASAP7_75t_L g10120 ( 
.A(n_9537),
.Y(n_10120)
);

INVx1_ASAP7_75t_L g10121 ( 
.A(n_9555),
.Y(n_10121)
);

INVx1_ASAP7_75t_L g10122 ( 
.A(n_9555),
.Y(n_10122)
);

AOI22xp33_ASAP7_75t_L g10123 ( 
.A1(n_9842),
.A2(n_9099),
.B1(n_9257),
.B2(n_9358),
.Y(n_10123)
);

AND2x2_ASAP7_75t_L g10124 ( 
.A(n_9542),
.B(n_9373),
.Y(n_10124)
);

INVx2_ASAP7_75t_L g10125 ( 
.A(n_9867),
.Y(n_10125)
);

AND2x2_ASAP7_75t_L g10126 ( 
.A(n_9544),
.B(n_9373),
.Y(n_10126)
);

NAND2xp5_ASAP7_75t_L g10127 ( 
.A(n_9676),
.B(n_8982),
.Y(n_10127)
);

NOR2xp67_ASAP7_75t_L g10128 ( 
.A(n_9606),
.B(n_9302),
.Y(n_10128)
);

INVx1_ASAP7_75t_L g10129 ( 
.A(n_9753),
.Y(n_10129)
);

AND2x2_ASAP7_75t_L g10130 ( 
.A(n_9754),
.B(n_9364),
.Y(n_10130)
);

OR2x2_ASAP7_75t_L g10131 ( 
.A(n_9485),
.B(n_9108),
.Y(n_10131)
);

AND2x2_ASAP7_75t_L g10132 ( 
.A(n_9891),
.B(n_9040),
.Y(n_10132)
);

INVx2_ASAP7_75t_SL g10133 ( 
.A(n_9772),
.Y(n_10133)
);

NAND2xp5_ASAP7_75t_L g10134 ( 
.A(n_9709),
.B(n_8982),
.Y(n_10134)
);

INVx2_ASAP7_75t_L g10135 ( 
.A(n_9498),
.Y(n_10135)
);

INVx1_ASAP7_75t_L g10136 ( 
.A(n_9753),
.Y(n_10136)
);

AND2x2_ASAP7_75t_L g10137 ( 
.A(n_9922),
.B(n_9264),
.Y(n_10137)
);

NAND2xp5_ASAP7_75t_L g10138 ( 
.A(n_9717),
.B(n_8988),
.Y(n_10138)
);

AND2x2_ASAP7_75t_L g10139 ( 
.A(n_9664),
.B(n_9269),
.Y(n_10139)
);

AND2x4_ASAP7_75t_L g10140 ( 
.A(n_9498),
.B(n_9065),
.Y(n_10140)
);

INVx2_ASAP7_75t_L g10141 ( 
.A(n_9790),
.Y(n_10141)
);

NOR3xp33_ASAP7_75t_L g10142 ( 
.A(n_9733),
.B(n_9267),
.C(n_9440),
.Y(n_10142)
);

INVx1_ASAP7_75t_L g10143 ( 
.A(n_9681),
.Y(n_10143)
);

HB1xp67_ASAP7_75t_L g10144 ( 
.A(n_9951),
.Y(n_10144)
);

NOR2x1_ASAP7_75t_SL g10145 ( 
.A(n_9842),
.B(n_9302),
.Y(n_10145)
);

NAND2xp5_ASAP7_75t_L g10146 ( 
.A(n_9932),
.B(n_8988),
.Y(n_10146)
);

INVx1_ASAP7_75t_L g10147 ( 
.A(n_9681),
.Y(n_10147)
);

AND2x2_ASAP7_75t_L g10148 ( 
.A(n_9817),
.B(n_9068),
.Y(n_10148)
);

AND2x2_ASAP7_75t_L g10149 ( 
.A(n_9595),
.B(n_9068),
.Y(n_10149)
);

INVx3_ASAP7_75t_L g10150 ( 
.A(n_9560),
.Y(n_10150)
);

AND2x4_ASAP7_75t_L g10151 ( 
.A(n_9600),
.B(n_9069),
.Y(n_10151)
);

AND2x2_ASAP7_75t_L g10152 ( 
.A(n_9596),
.B(n_9069),
.Y(n_10152)
);

INVxp67_ASAP7_75t_L g10153 ( 
.A(n_9633),
.Y(n_10153)
);

AND2x2_ASAP7_75t_L g10154 ( 
.A(n_9778),
.B(n_9071),
.Y(n_10154)
);

AOI22xp5_ASAP7_75t_L g10155 ( 
.A1(n_9956),
.A2(n_9257),
.B1(n_9365),
.B2(n_9273),
.Y(n_10155)
);

AND2x2_ASAP7_75t_L g10156 ( 
.A(n_9703),
.B(n_9071),
.Y(n_10156)
);

OR2x2_ASAP7_75t_L g10157 ( 
.A(n_9485),
.B(n_9096),
.Y(n_10157)
);

AND2x2_ASAP7_75t_L g10158 ( 
.A(n_9706),
.B(n_9075),
.Y(n_10158)
);

AND2x4_ASAP7_75t_L g10159 ( 
.A(n_9567),
.B(n_9075),
.Y(n_10159)
);

OAI21xp5_ASAP7_75t_SL g10160 ( 
.A1(n_9879),
.A2(n_9142),
.B(n_9273),
.Y(n_10160)
);

NAND2xp5_ASAP7_75t_L g10161 ( 
.A(n_9944),
.B(n_9012),
.Y(n_10161)
);

AND2x4_ASAP7_75t_L g10162 ( 
.A(n_9567),
.B(n_9577),
.Y(n_10162)
);

INVx2_ASAP7_75t_L g10163 ( 
.A(n_9790),
.Y(n_10163)
);

NAND2xp5_ASAP7_75t_L g10164 ( 
.A(n_9547),
.B(n_9012),
.Y(n_10164)
);

AND2x2_ASAP7_75t_L g10165 ( 
.A(n_9651),
.B(n_9079),
.Y(n_10165)
);

NAND2xp5_ASAP7_75t_L g10166 ( 
.A(n_9550),
.B(n_9013),
.Y(n_10166)
);

AND2x2_ASAP7_75t_L g10167 ( 
.A(n_9652),
.B(n_9079),
.Y(n_10167)
);

AND2x2_ASAP7_75t_L g10168 ( 
.A(n_9748),
.B(n_9084),
.Y(n_10168)
);

OR2x2_ASAP7_75t_L g10169 ( 
.A(n_9747),
.B(n_9411),
.Y(n_10169)
);

AND2x2_ASAP7_75t_L g10170 ( 
.A(n_9766),
.B(n_9084),
.Y(n_10170)
);

NAND2x1_ASAP7_75t_SL g10171 ( 
.A(n_9499),
.B(n_9387),
.Y(n_10171)
);

INVx2_ASAP7_75t_L g10172 ( 
.A(n_9820),
.Y(n_10172)
);

INVx3_ASAP7_75t_L g10173 ( 
.A(n_9577),
.Y(n_10173)
);

OR2x2_ASAP7_75t_L g10174 ( 
.A(n_9622),
.B(n_9382),
.Y(n_10174)
);

INVx1_ASAP7_75t_SL g10175 ( 
.A(n_9840),
.Y(n_10175)
);

INVx1_ASAP7_75t_L g10176 ( 
.A(n_9697),
.Y(n_10176)
);

NAND2xp5_ASAP7_75t_L g10177 ( 
.A(n_9561),
.B(n_9615),
.Y(n_10177)
);

AND2x2_ASAP7_75t_L g10178 ( 
.A(n_9768),
.B(n_9087),
.Y(n_10178)
);

INVx3_ASAP7_75t_L g10179 ( 
.A(n_9635),
.Y(n_10179)
);

INVx1_ASAP7_75t_L g10180 ( 
.A(n_9699),
.Y(n_10180)
);

INVx1_ASAP7_75t_L g10181 ( 
.A(n_9702),
.Y(n_10181)
);

AND2x2_ASAP7_75t_L g10182 ( 
.A(n_9511),
.B(n_9087),
.Y(n_10182)
);

AND2x2_ASAP7_75t_L g10183 ( 
.A(n_9512),
.B(n_9647),
.Y(n_10183)
);

INVx1_ASAP7_75t_L g10184 ( 
.A(n_9707),
.Y(n_10184)
);

NAND2xp5_ASAP7_75t_L g10185 ( 
.A(n_9616),
.B(n_9013),
.Y(n_10185)
);

INVx1_ASAP7_75t_L g10186 ( 
.A(n_9646),
.Y(n_10186)
);

INVx2_ASAP7_75t_SL g10187 ( 
.A(n_9823),
.Y(n_10187)
);

OR2x2_ASAP7_75t_L g10188 ( 
.A(n_9716),
.B(n_9216),
.Y(n_10188)
);

AND2x4_ASAP7_75t_L g10189 ( 
.A(n_9635),
.B(n_9107),
.Y(n_10189)
);

AND2x2_ASAP7_75t_L g10190 ( 
.A(n_9553),
.B(n_9107),
.Y(n_10190)
);

INVx2_ASAP7_75t_L g10191 ( 
.A(n_9820),
.Y(n_10191)
);

AND2x2_ASAP7_75t_L g10192 ( 
.A(n_9910),
.B(n_9111),
.Y(n_10192)
);

NAND2xp5_ASAP7_75t_L g10193 ( 
.A(n_9923),
.B(n_9018),
.Y(n_10193)
);

AND2x2_ASAP7_75t_L g10194 ( 
.A(n_9898),
.B(n_9111),
.Y(n_10194)
);

INVxp67_ASAP7_75t_L g10195 ( 
.A(n_9605),
.Y(n_10195)
);

NAND2xp5_ASAP7_75t_L g10196 ( 
.A(n_9923),
.B(n_9018),
.Y(n_10196)
);

INVx1_ASAP7_75t_L g10197 ( 
.A(n_9648),
.Y(n_10197)
);

INVx1_ASAP7_75t_L g10198 ( 
.A(n_9663),
.Y(n_10198)
);

NAND2xp5_ASAP7_75t_L g10199 ( 
.A(n_9952),
.B(n_9637),
.Y(n_10199)
);

HB1xp67_ASAP7_75t_L g10200 ( 
.A(n_9606),
.Y(n_10200)
);

AND2x2_ASAP7_75t_L g10201 ( 
.A(n_9899),
.B(n_9117),
.Y(n_10201)
);

AND2x2_ASAP7_75t_L g10202 ( 
.A(n_9913),
.B(n_9117),
.Y(n_10202)
);

INVx2_ASAP7_75t_SL g10203 ( 
.A(n_9823),
.Y(n_10203)
);

INVx1_ASAP7_75t_L g10204 ( 
.A(n_9665),
.Y(n_10204)
);

OR2x2_ASAP7_75t_L g10205 ( 
.A(n_9846),
.B(n_9870),
.Y(n_10205)
);

INVx2_ASAP7_75t_L g10206 ( 
.A(n_9838),
.Y(n_10206)
);

INVx2_ASAP7_75t_L g10207 ( 
.A(n_9838),
.Y(n_10207)
);

AND2x2_ASAP7_75t_L g10208 ( 
.A(n_9579),
.B(n_9119),
.Y(n_10208)
);

HB1xp67_ASAP7_75t_L g10209 ( 
.A(n_9625),
.Y(n_10209)
);

INVx2_ASAP7_75t_SL g10210 ( 
.A(n_9840),
.Y(n_10210)
);

OR2x2_ASAP7_75t_L g10211 ( 
.A(n_9874),
.B(n_9288),
.Y(n_10211)
);

BUFx2_ASAP7_75t_L g10212 ( 
.A(n_9873),
.Y(n_10212)
);

INVx1_ASAP7_75t_L g10213 ( 
.A(n_9666),
.Y(n_10213)
);

INVx1_ASAP7_75t_L g10214 ( 
.A(n_9668),
.Y(n_10214)
);

INVx2_ASAP7_75t_L g10215 ( 
.A(n_9862),
.Y(n_10215)
);

AND2x2_ASAP7_75t_L g10216 ( 
.A(n_9760),
.B(n_9119),
.Y(n_10216)
);

INVx1_ASAP7_75t_L g10217 ( 
.A(n_9710),
.Y(n_10217)
);

INVx1_ASAP7_75t_L g10218 ( 
.A(n_9713),
.Y(n_10218)
);

AND2x2_ASAP7_75t_L g10219 ( 
.A(n_9763),
.B(n_9024),
.Y(n_10219)
);

OR2x2_ASAP7_75t_L g10220 ( 
.A(n_9926),
.B(n_9460),
.Y(n_10220)
);

INVx1_ASAP7_75t_L g10221 ( 
.A(n_9714),
.Y(n_10221)
);

INVx1_ASAP7_75t_L g10222 ( 
.A(n_9715),
.Y(n_10222)
);

AOI211xp5_ASAP7_75t_L g10223 ( 
.A1(n_9602),
.A2(n_9267),
.B(n_9315),
.C(n_9011),
.Y(n_10223)
);

NAND2xp5_ASAP7_75t_L g10224 ( 
.A(n_9952),
.B(n_9024),
.Y(n_10224)
);

INVx1_ASAP7_75t_L g10225 ( 
.A(n_9720),
.Y(n_10225)
);

INVx1_ASAP7_75t_L g10226 ( 
.A(n_9721),
.Y(n_10226)
);

INVx2_ASAP7_75t_L g10227 ( 
.A(n_9862),
.Y(n_10227)
);

AND2x2_ASAP7_75t_L g10228 ( 
.A(n_9897),
.B(n_9728),
.Y(n_10228)
);

INVx2_ASAP7_75t_L g10229 ( 
.A(n_9868),
.Y(n_10229)
);

AOI22xp5_ASAP7_75t_L g10230 ( 
.A1(n_9956),
.A2(n_9142),
.B1(n_9177),
.B2(n_9384),
.Y(n_10230)
);

INVx1_ASAP7_75t_L g10231 ( 
.A(n_9724),
.Y(n_10231)
);

AND2x2_ASAP7_75t_L g10232 ( 
.A(n_9911),
.B(n_9163),
.Y(n_10232)
);

INVx1_ASAP7_75t_L g10233 ( 
.A(n_9726),
.Y(n_10233)
);

AND2x4_ASAP7_75t_L g10234 ( 
.A(n_9489),
.B(n_9507),
.Y(n_10234)
);

INVx3_ASAP7_75t_L g10235 ( 
.A(n_9788),
.Y(n_10235)
);

INVx1_ASAP7_75t_L g10236 ( 
.A(n_9727),
.Y(n_10236)
);

AND2x2_ASAP7_75t_L g10237 ( 
.A(n_9861),
.B(n_9163),
.Y(n_10237)
);

NAND2x1p5_ASAP7_75t_L g10238 ( 
.A(n_9839),
.B(n_9446),
.Y(n_10238)
);

NAND2xp5_ASAP7_75t_L g10239 ( 
.A(n_9638),
.B(n_9165),
.Y(n_10239)
);

AND2x4_ASAP7_75t_L g10240 ( 
.A(n_9523),
.B(n_9165),
.Y(n_10240)
);

INVx1_ASAP7_75t_L g10241 ( 
.A(n_9673),
.Y(n_10241)
);

INVxp67_ASAP7_75t_L g10242 ( 
.A(n_9655),
.Y(n_10242)
);

AND2x2_ASAP7_75t_L g10243 ( 
.A(n_9854),
.B(n_9739),
.Y(n_10243)
);

NAND2xp5_ASAP7_75t_L g10244 ( 
.A(n_9640),
.B(n_9166),
.Y(n_10244)
);

AND2x2_ASAP7_75t_L g10245 ( 
.A(n_9742),
.B(n_9166),
.Y(n_10245)
);

AND2x2_ASAP7_75t_L g10246 ( 
.A(n_9850),
.B(n_9168),
.Y(n_10246)
);

OR2x2_ASAP7_75t_L g10247 ( 
.A(n_9591),
.B(n_9464),
.Y(n_10247)
);

INVx1_ASAP7_75t_L g10248 ( 
.A(n_9692),
.Y(n_10248)
);

OAI22xp5_ASAP7_75t_L g10249 ( 
.A1(n_9758),
.A2(n_7904),
.B1(n_7925),
.B2(n_7921),
.Y(n_10249)
);

INVx1_ASAP7_75t_L g10250 ( 
.A(n_9696),
.Y(n_10250)
);

AND2x2_ASAP7_75t_L g10251 ( 
.A(n_9649),
.B(n_9168),
.Y(n_10251)
);

OAI221xp5_ASAP7_75t_SL g10252 ( 
.A1(n_9490),
.A2(n_9044),
.B1(n_9115),
.B2(n_9455),
.C(n_9202),
.Y(n_10252)
);

AND2x2_ASAP7_75t_L g10253 ( 
.A(n_9654),
.B(n_9170),
.Y(n_10253)
);

AND2x4_ASAP7_75t_L g10254 ( 
.A(n_9499),
.B(n_9170),
.Y(n_10254)
);

INVx1_ASAP7_75t_SL g10255 ( 
.A(n_9948),
.Y(n_10255)
);

AND2x2_ASAP7_75t_L g10256 ( 
.A(n_9669),
.B(n_9670),
.Y(n_10256)
);

OR2x2_ASAP7_75t_L g10257 ( 
.A(n_9847),
.B(n_9474),
.Y(n_10257)
);

NAND3xp33_ASAP7_75t_L g10258 ( 
.A(n_9884),
.B(n_9316),
.C(n_9304),
.Y(n_10258)
);

AND2x2_ASAP7_75t_L g10259 ( 
.A(n_9708),
.B(n_9185),
.Y(n_10259)
);

AND2x2_ASAP7_75t_L g10260 ( 
.A(n_9745),
.B(n_9185),
.Y(n_10260)
);

INVx1_ASAP7_75t_L g10261 ( 
.A(n_9618),
.Y(n_10261)
);

INVx2_ASAP7_75t_L g10262 ( 
.A(n_9868),
.Y(n_10262)
);

INVx1_ASAP7_75t_L g10263 ( 
.A(n_9621),
.Y(n_10263)
);

INVx1_ASAP7_75t_L g10264 ( 
.A(n_9623),
.Y(n_10264)
);

AND2x4_ASAP7_75t_SL g10265 ( 
.A(n_9719),
.B(n_9446),
.Y(n_10265)
);

NAND2xp5_ASAP7_75t_SL g10266 ( 
.A(n_9902),
.B(n_9304),
.Y(n_10266)
);

NOR2xp33_ASAP7_75t_L g10267 ( 
.A(n_9773),
.B(n_7825),
.Y(n_10267)
);

NAND2x1p5_ASAP7_75t_L g10268 ( 
.A(n_9882),
.B(n_9454),
.Y(n_10268)
);

NAND2xp5_ASAP7_75t_L g10269 ( 
.A(n_9782),
.B(n_9194),
.Y(n_10269)
);

AND2x4_ASAP7_75t_L g10270 ( 
.A(n_9502),
.B(n_9194),
.Y(n_10270)
);

AND2x2_ASAP7_75t_L g10271 ( 
.A(n_9546),
.B(n_9205),
.Y(n_10271)
);

INVx1_ASAP7_75t_L g10272 ( 
.A(n_9626),
.Y(n_10272)
);

INVx2_ASAP7_75t_L g10273 ( 
.A(n_9881),
.Y(n_10273)
);

OR2x2_ASAP7_75t_L g10274 ( 
.A(n_9828),
.B(n_9848),
.Y(n_10274)
);

AND2x2_ASAP7_75t_L g10275 ( 
.A(n_9546),
.B(n_9205),
.Y(n_10275)
);

OR2x2_ASAP7_75t_L g10276 ( 
.A(n_9828),
.B(n_9056),
.Y(n_10276)
);

AND2x4_ASAP7_75t_L g10277 ( 
.A(n_9502),
.B(n_9212),
.Y(n_10277)
);

NOR2x1_ASAP7_75t_L g10278 ( 
.A(n_9788),
.B(n_9212),
.Y(n_10278)
);

NAND2xp5_ASAP7_75t_L g10279 ( 
.A(n_9782),
.B(n_9213),
.Y(n_10279)
);

INVx1_ASAP7_75t_L g10280 ( 
.A(n_9627),
.Y(n_10280)
);

HB1xp67_ASAP7_75t_L g10281 ( 
.A(n_9741),
.Y(n_10281)
);

OR2x2_ASAP7_75t_L g10282 ( 
.A(n_9848),
.B(n_9433),
.Y(n_10282)
);

INVx1_ASAP7_75t_L g10283 ( 
.A(n_9628),
.Y(n_10283)
);

NAND2xp5_ASAP7_75t_L g10284 ( 
.A(n_9937),
.B(n_9213),
.Y(n_10284)
);

AND2x4_ASAP7_75t_L g10285 ( 
.A(n_9741),
.B(n_9222),
.Y(n_10285)
);

AND2x4_ASAP7_75t_L g10286 ( 
.A(n_9515),
.B(n_9222),
.Y(n_10286)
);

AND2x2_ASAP7_75t_L g10287 ( 
.A(n_9802),
.B(n_9226),
.Y(n_10287)
);

INVx1_ASAP7_75t_L g10288 ( 
.A(n_9636),
.Y(n_10288)
);

HB1xp67_ASAP7_75t_L g10289 ( 
.A(n_9641),
.Y(n_10289)
);

INVx1_ASAP7_75t_L g10290 ( 
.A(n_9639),
.Y(n_10290)
);

AND2x2_ASAP7_75t_L g10291 ( 
.A(n_9612),
.B(n_9226),
.Y(n_10291)
);

AND2x2_ASAP7_75t_L g10292 ( 
.A(n_9816),
.B(n_9230),
.Y(n_10292)
);

AND2x2_ASAP7_75t_L g10293 ( 
.A(n_9914),
.B(n_9230),
.Y(n_10293)
);

NAND2xp5_ASAP7_75t_L g10294 ( 
.A(n_9761),
.B(n_9573),
.Y(n_10294)
);

AND2x2_ASAP7_75t_SL g10295 ( 
.A(n_9908),
.B(n_9316),
.Y(n_10295)
);

AND2x2_ASAP7_75t_L g10296 ( 
.A(n_9916),
.B(n_9231),
.Y(n_10296)
);

AND2x2_ASAP7_75t_L g10297 ( 
.A(n_9812),
.B(n_9231),
.Y(n_10297)
);

OR2x2_ASAP7_75t_L g10298 ( 
.A(n_9565),
.B(n_9434),
.Y(n_10298)
);

INVx2_ASAP7_75t_L g10299 ( 
.A(n_9881),
.Y(n_10299)
);

AND2x2_ASAP7_75t_L g10300 ( 
.A(n_9740),
.B(n_9831),
.Y(n_10300)
);

INVx1_ASAP7_75t_L g10301 ( 
.A(n_9643),
.Y(n_10301)
);

OR2x2_ASAP7_75t_L g10302 ( 
.A(n_9791),
.B(n_9233),
.Y(n_10302)
);

OR2x2_ASAP7_75t_L g10303 ( 
.A(n_9791),
.B(n_9233),
.Y(n_10303)
);

NAND3xp33_ASAP7_75t_L g10304 ( 
.A(n_9884),
.B(n_9461),
.C(n_9454),
.Y(n_10304)
);

INVx2_ASAP7_75t_L g10305 ( 
.A(n_9515),
.Y(n_10305)
);

AND2x2_ASAP7_75t_L g10306 ( 
.A(n_9834),
.B(n_9234),
.Y(n_10306)
);

INVx2_ASAP7_75t_SL g10307 ( 
.A(n_9734),
.Y(n_10307)
);

NAND2xp5_ASAP7_75t_L g10308 ( 
.A(n_9761),
.B(n_9234),
.Y(n_10308)
);

INVx1_ASAP7_75t_L g10309 ( 
.A(n_9644),
.Y(n_10309)
);

NAND4xp25_ASAP7_75t_SL g10310 ( 
.A(n_9602),
.B(n_8826),
.C(n_8110),
.D(n_8280),
.Y(n_10310)
);

INVx1_ASAP7_75t_L g10311 ( 
.A(n_9584),
.Y(n_10311)
);

OR2x2_ASAP7_75t_L g10312 ( 
.A(n_9487),
.B(n_9049),
.Y(n_10312)
);

INVx2_ASAP7_75t_L g10313 ( 
.A(n_9517),
.Y(n_10313)
);

AND2x2_ASAP7_75t_L g10314 ( 
.A(n_9924),
.B(n_9461),
.Y(n_10314)
);

AND2x2_ASAP7_75t_L g10315 ( 
.A(n_9927),
.B(n_9463),
.Y(n_10315)
);

AND2x2_ASAP7_75t_L g10316 ( 
.A(n_9930),
.B(n_9463),
.Y(n_10316)
);

HB1xp67_ASAP7_75t_L g10317 ( 
.A(n_9656),
.Y(n_10317)
);

INVx1_ASAP7_75t_L g10318 ( 
.A(n_9584),
.Y(n_10318)
);

NAND2xp5_ASAP7_75t_L g10319 ( 
.A(n_9610),
.B(n_9062),
.Y(n_10319)
);

NAND2xp5_ASAP7_75t_L g10320 ( 
.A(n_9589),
.B(n_9594),
.Y(n_10320)
);

INVx2_ASAP7_75t_L g10321 ( 
.A(n_9517),
.Y(n_10321)
);

INVx2_ASAP7_75t_L g10322 ( 
.A(n_9518),
.Y(n_10322)
);

AND2x2_ASAP7_75t_L g10323 ( 
.A(n_9597),
.B(n_9240),
.Y(n_10323)
);

INVx2_ASAP7_75t_L g10324 ( 
.A(n_9518),
.Y(n_10324)
);

INVx2_ASAP7_75t_L g10325 ( 
.A(n_9519),
.Y(n_10325)
);

INVx2_ASAP7_75t_L g10326 ( 
.A(n_9519),
.Y(n_10326)
);

HB1xp67_ASAP7_75t_L g10327 ( 
.A(n_9725),
.Y(n_10327)
);

INVx1_ASAP7_75t_L g10328 ( 
.A(n_9585),
.Y(n_10328)
);

INVx1_ASAP7_75t_L g10329 ( 
.A(n_9585),
.Y(n_10329)
);

NAND2xp5_ASAP7_75t_L g10330 ( 
.A(n_9589),
.B(n_9063),
.Y(n_10330)
);

INVx1_ASAP7_75t_L g10331 ( 
.A(n_9491),
.Y(n_10331)
);

BUFx2_ASAP7_75t_L g10332 ( 
.A(n_9734),
.Y(n_10332)
);

INVx2_ASAP7_75t_L g10333 ( 
.A(n_9521),
.Y(n_10333)
);

OR2x2_ASAP7_75t_L g10334 ( 
.A(n_9941),
.B(n_9066),
.Y(n_10334)
);

NAND2xp5_ASAP7_75t_L g10335 ( 
.A(n_9594),
.B(n_9067),
.Y(n_10335)
);

AND2x2_ASAP7_75t_L g10336 ( 
.A(n_9597),
.B(n_9240),
.Y(n_10336)
);

NAND2xp5_ASAP7_75t_L g10337 ( 
.A(n_9604),
.B(n_9072),
.Y(n_10337)
);

NAND2xp5_ASAP7_75t_L g10338 ( 
.A(n_9604),
.B(n_9090),
.Y(n_10338)
);

NAND3xp33_ASAP7_75t_L g10339 ( 
.A(n_9758),
.B(n_9092),
.C(n_9091),
.Y(n_10339)
);

HB1xp67_ASAP7_75t_L g10340 ( 
.A(n_9521),
.Y(n_10340)
);

OAI21xp33_ASAP7_75t_L g10341 ( 
.A1(n_9490),
.A2(n_9011),
.B(n_9095),
.Y(n_10341)
);

AND2x2_ASAP7_75t_L g10342 ( 
.A(n_9826),
.B(n_9242),
.Y(n_10342)
);

AND2x2_ASAP7_75t_L g10343 ( 
.A(n_9877),
.B(n_9950),
.Y(n_10343)
);

AND2x4_ASAP7_75t_L g10344 ( 
.A(n_9522),
.B(n_9242),
.Y(n_10344)
);

AND2x4_ASAP7_75t_L g10345 ( 
.A(n_9522),
.B(n_9246),
.Y(n_10345)
);

AND2x2_ASAP7_75t_L g10346 ( 
.A(n_9630),
.B(n_9246),
.Y(n_10346)
);

INVx1_ASAP7_75t_SL g10347 ( 
.A(n_9671),
.Y(n_10347)
);

HB1xp67_ASAP7_75t_L g10348 ( 
.A(n_9541),
.Y(n_10348)
);

OR2x2_ASAP7_75t_L g10349 ( 
.A(n_9833),
.B(n_9097),
.Y(n_10349)
);

INVx1_ASAP7_75t_L g10350 ( 
.A(n_9679),
.Y(n_10350)
);

AND2x2_ASAP7_75t_L g10351 ( 
.A(n_9793),
.B(n_9254),
.Y(n_10351)
);

NAND2xp5_ASAP7_75t_L g10352 ( 
.A(n_9607),
.B(n_9104),
.Y(n_10352)
);

AND2x2_ASAP7_75t_L g10353 ( 
.A(n_9876),
.B(n_9254),
.Y(n_10353)
);

NAND2xp5_ASAP7_75t_L g10354 ( 
.A(n_9607),
.B(n_9109),
.Y(n_10354)
);

OR2x2_ASAP7_75t_L g10355 ( 
.A(n_9590),
.B(n_9110),
.Y(n_10355)
);

INVx1_ASAP7_75t_L g10356 ( 
.A(n_9679),
.Y(n_10356)
);

INVx2_ASAP7_75t_L g10357 ( 
.A(n_9541),
.Y(n_10357)
);

NAND2xp5_ASAP7_75t_L g10358 ( 
.A(n_9543),
.B(n_9112),
.Y(n_10358)
);

AND2x2_ASAP7_75t_L g10359 ( 
.A(n_9875),
.B(n_9255),
.Y(n_10359)
);

INVx1_ASAP7_75t_L g10360 ( 
.A(n_9496),
.Y(n_10360)
);

HB1xp67_ASAP7_75t_L g10361 ( 
.A(n_9543),
.Y(n_10361)
);

INVx1_ASAP7_75t_L g10362 ( 
.A(n_9497),
.Y(n_10362)
);

AND2x4_ASAP7_75t_L g10363 ( 
.A(n_9580),
.B(n_9255),
.Y(n_10363)
);

NAND2xp5_ASAP7_75t_L g10364 ( 
.A(n_9580),
.B(n_9114),
.Y(n_10364)
);

OR2x2_ASAP7_75t_L g10365 ( 
.A(n_9657),
.B(n_9116),
.Y(n_10365)
);

INVx1_ASAP7_75t_L g10366 ( 
.A(n_9506),
.Y(n_10366)
);

AND2x2_ASAP7_75t_L g10367 ( 
.A(n_9794),
.B(n_9265),
.Y(n_10367)
);

BUFx2_ASAP7_75t_L g10368 ( 
.A(n_9860),
.Y(n_10368)
);

OR2x2_ASAP7_75t_L g10369 ( 
.A(n_9705),
.B(n_9118),
.Y(n_10369)
);

OR2x2_ASAP7_75t_L g10370 ( 
.A(n_9942),
.B(n_9136),
.Y(n_10370)
);

INVx1_ASAP7_75t_L g10371 ( 
.A(n_9510),
.Y(n_10371)
);

INVx1_ASAP7_75t_L g10372 ( 
.A(n_9516),
.Y(n_10372)
);

AND2x2_ASAP7_75t_L g10373 ( 
.A(n_9967),
.B(n_9866),
.Y(n_10373)
);

INVx2_ASAP7_75t_L g10374 ( 
.A(n_10171),
.Y(n_10374)
);

AND2x2_ASAP7_75t_L g10375 ( 
.A(n_9969),
.B(n_9866),
.Y(n_10375)
);

AND2x4_ASAP7_75t_L g10376 ( 
.A(n_10030),
.B(n_9683),
.Y(n_10376)
);

INVx1_ASAP7_75t_L g10377 ( 
.A(n_10000),
.Y(n_10377)
);

INVx2_ASAP7_75t_L g10378 ( 
.A(n_10030),
.Y(n_10378)
);

AND2x2_ASAP7_75t_L g10379 ( 
.A(n_10228),
.B(n_9756),
.Y(n_10379)
);

BUFx12f_ASAP7_75t_L g10380 ( 
.A(n_9995),
.Y(n_10380)
);

INVx2_ASAP7_75t_L g10381 ( 
.A(n_10173),
.Y(n_10381)
);

AND2x4_ASAP7_75t_SL g10382 ( 
.A(n_10018),
.B(n_9723),
.Y(n_10382)
);

INVx1_ASAP7_75t_SL g10383 ( 
.A(n_9960),
.Y(n_10383)
);

AND2x2_ASAP7_75t_L g10384 ( 
.A(n_9998),
.B(n_9757),
.Y(n_10384)
);

AND2x2_ASAP7_75t_L g10385 ( 
.A(n_10074),
.B(n_9759),
.Y(n_10385)
);

INVx2_ASAP7_75t_L g10386 ( 
.A(n_10173),
.Y(n_10386)
);

OR2x2_ASAP7_75t_L g10387 ( 
.A(n_10144),
.B(n_9661),
.Y(n_10387)
);

INVx2_ASAP7_75t_L g10388 ( 
.A(n_10179),
.Y(n_10388)
);

INVx1_ASAP7_75t_L g10389 ( 
.A(n_10017),
.Y(n_10389)
);

INVx2_ASAP7_75t_L g10390 ( 
.A(n_10179),
.Y(n_10390)
);

NAND2xp5_ASAP7_75t_L g10391 ( 
.A(n_9961),
.B(n_9735),
.Y(n_10391)
);

INVx2_ASAP7_75t_L g10392 ( 
.A(n_10097),
.Y(n_10392)
);

AND2x2_ASAP7_75t_L g10393 ( 
.A(n_10076),
.B(n_9762),
.Y(n_10393)
);

AND2x2_ASAP7_75t_L g10394 ( 
.A(n_9982),
.B(n_9771),
.Y(n_10394)
);

AND2x2_ASAP7_75t_L g10395 ( 
.A(n_10243),
.B(n_9736),
.Y(n_10395)
);

INVx2_ASAP7_75t_L g10396 ( 
.A(n_10117),
.Y(n_10396)
);

INVx1_ASAP7_75t_L g10397 ( 
.A(n_10145),
.Y(n_10397)
);

INVx1_ASAP7_75t_L g10398 ( 
.A(n_10145),
.Y(n_10398)
);

NAND2xp5_ASAP7_75t_L g10399 ( 
.A(n_9974),
.B(n_9683),
.Y(n_10399)
);

INVx1_ASAP7_75t_L g10400 ( 
.A(n_9980),
.Y(n_10400)
);

INVxp67_ASAP7_75t_SL g10401 ( 
.A(n_9990),
.Y(n_10401)
);

INVx2_ASAP7_75t_L g10402 ( 
.A(n_10117),
.Y(n_10402)
);

OR2x2_ASAP7_75t_L g10403 ( 
.A(n_10205),
.B(n_9983),
.Y(n_10403)
);

AND2x2_ASAP7_75t_L g10404 ( 
.A(n_10060),
.B(n_9587),
.Y(n_10404)
);

AND2x2_ASAP7_75t_L g10405 ( 
.A(n_10343),
.B(n_9587),
.Y(n_10405)
);

AND2x2_ASAP7_75t_L g10406 ( 
.A(n_10139),
.B(n_9743),
.Y(n_10406)
);

AND2x2_ASAP7_75t_L g10407 ( 
.A(n_9984),
.B(n_9746),
.Y(n_10407)
);

HB1xp67_ASAP7_75t_L g10408 ( 
.A(n_10128),
.Y(n_10408)
);

INVx1_ASAP7_75t_L g10409 ( 
.A(n_9993),
.Y(n_10409)
);

OR2x2_ASAP7_75t_L g10410 ( 
.A(n_10010),
.B(n_9965),
.Y(n_10410)
);

NAND2xp5_ASAP7_75t_L g10411 ( 
.A(n_10021),
.B(n_9968),
.Y(n_10411)
);

HB1xp67_ASAP7_75t_L g10412 ( 
.A(n_10102),
.Y(n_10412)
);

AND2x4_ASAP7_75t_L g10413 ( 
.A(n_10162),
.B(n_9685),
.Y(n_10413)
);

AND2x4_ASAP7_75t_L g10414 ( 
.A(n_10162),
.B(n_9685),
.Y(n_10414)
);

AND2x2_ASAP7_75t_L g10415 ( 
.A(n_10006),
.B(n_9749),
.Y(n_10415)
);

AND2x2_ASAP7_75t_L g10416 ( 
.A(n_9992),
.B(n_9750),
.Y(n_10416)
);

OR2x2_ASAP7_75t_L g10417 ( 
.A(n_9976),
.B(n_10027),
.Y(n_10417)
);

NAND2xp5_ASAP7_75t_L g10418 ( 
.A(n_10295),
.B(n_10255),
.Y(n_10418)
);

INVx2_ASAP7_75t_L g10419 ( 
.A(n_10150),
.Y(n_10419)
);

NAND2xp5_ASAP7_75t_L g10420 ( 
.A(n_10332),
.B(n_9689),
.Y(n_10420)
);

AND2x2_ASAP7_75t_L g10421 ( 
.A(n_9988),
.B(n_9752),
.Y(n_10421)
);

AND2x2_ASAP7_75t_L g10422 ( 
.A(n_10051),
.B(n_9689),
.Y(n_10422)
);

AND2x2_ASAP7_75t_L g10423 ( 
.A(n_10137),
.B(n_9693),
.Y(n_10423)
);

OR2x2_ASAP7_75t_L g10424 ( 
.A(n_10113),
.B(n_10211),
.Y(n_10424)
);

AND2x2_ASAP7_75t_L g10425 ( 
.A(n_10114),
.B(n_9693),
.Y(n_10425)
);

INVx1_ASAP7_75t_L g10426 ( 
.A(n_10143),
.Y(n_10426)
);

INVx1_ASAP7_75t_L g10427 ( 
.A(n_10143),
.Y(n_10427)
);

OR2x2_ASAP7_75t_L g10428 ( 
.A(n_10072),
.B(n_9755),
.Y(n_10428)
);

AND2x2_ASAP7_75t_L g10429 ( 
.A(n_10271),
.B(n_9815),
.Y(n_10429)
);

AND2x2_ASAP7_75t_L g10430 ( 
.A(n_10275),
.B(n_9815),
.Y(n_10430)
);

AND2x2_ASAP7_75t_L g10431 ( 
.A(n_10183),
.B(n_9871),
.Y(n_10431)
);

AND2x2_ASAP7_75t_L g10432 ( 
.A(n_10080),
.B(n_9779),
.Y(n_10432)
);

INVxp67_ASAP7_75t_SL g10433 ( 
.A(n_10289),
.Y(n_10433)
);

INVx1_ASAP7_75t_L g10434 ( 
.A(n_9962),
.Y(n_10434)
);

OR2x2_ASAP7_75t_L g10435 ( 
.A(n_10088),
.B(n_9769),
.Y(n_10435)
);

HB1xp67_ASAP7_75t_L g10436 ( 
.A(n_10317),
.Y(n_10436)
);

INVx1_ASAP7_75t_L g10437 ( 
.A(n_9962),
.Y(n_10437)
);

OR2x2_ASAP7_75t_L g10438 ( 
.A(n_10209),
.B(n_9784),
.Y(n_10438)
);

INVx1_ASAP7_75t_L g10439 ( 
.A(n_10147),
.Y(n_10439)
);

AND2x4_ASAP7_75t_L g10440 ( 
.A(n_10150),
.B(n_9505),
.Y(n_10440)
);

OR2x2_ASAP7_75t_L g10441 ( 
.A(n_10003),
.B(n_9792),
.Y(n_10441)
);

NOR2xp33_ASAP7_75t_L g10442 ( 
.A(n_10175),
.B(n_9614),
.Y(n_10442)
);

INVx1_ASAP7_75t_L g10443 ( 
.A(n_10147),
.Y(n_10443)
);

OR2x2_ASAP7_75t_L g10444 ( 
.A(n_10081),
.B(n_9564),
.Y(n_10444)
);

AND2x2_ASAP7_75t_L g10445 ( 
.A(n_10086),
.B(n_10100),
.Y(n_10445)
);

AND2x2_ASAP7_75t_L g10446 ( 
.A(n_10105),
.B(n_10025),
.Y(n_10446)
);

NOR2xp33_ASAP7_75t_L g10447 ( 
.A(n_10187),
.B(n_9620),
.Y(n_10447)
);

AND2x4_ASAP7_75t_L g10448 ( 
.A(n_10020),
.B(n_9505),
.Y(n_10448)
);

AND2x2_ASAP7_75t_L g10449 ( 
.A(n_10032),
.B(n_9738),
.Y(n_10449)
);

NOR2xp33_ASAP7_75t_SL g10450 ( 
.A(n_10203),
.B(n_9568),
.Y(n_10450)
);

AND2x2_ASAP7_75t_L g10451 ( 
.A(n_10246),
.B(n_9738),
.Y(n_10451)
);

NAND2xp5_ASAP7_75t_L g10452 ( 
.A(n_10112),
.B(n_10079),
.Y(n_10452)
);

INVx4_ASAP7_75t_L g10453 ( 
.A(n_10118),
.Y(n_10453)
);

HB1xp67_ASAP7_75t_L g10454 ( 
.A(n_10327),
.Y(n_10454)
);

AND2x2_ASAP7_75t_L g10455 ( 
.A(n_10058),
.B(n_9780),
.Y(n_10455)
);

AND2x4_ASAP7_75t_L g10456 ( 
.A(n_10020),
.B(n_9797),
.Y(n_10456)
);

NAND2xp5_ASAP7_75t_L g10457 ( 
.A(n_10281),
.B(n_9900),
.Y(n_10457)
);

HB1xp67_ASAP7_75t_L g10458 ( 
.A(n_10001),
.Y(n_10458)
);

AND2x4_ASAP7_75t_L g10459 ( 
.A(n_10052),
.B(n_9797),
.Y(n_10459)
);

AND2x2_ASAP7_75t_L g10460 ( 
.A(n_10148),
.B(n_9783),
.Y(n_10460)
);

AND2x2_ASAP7_75t_L g10461 ( 
.A(n_10067),
.B(n_9786),
.Y(n_10461)
);

INVx1_ASAP7_75t_L g10462 ( 
.A(n_9964),
.Y(n_10462)
);

NAND2xp5_ASAP7_75t_L g10463 ( 
.A(n_10189),
.B(n_9900),
.Y(n_10463)
);

NAND2xp5_ASAP7_75t_L g10464 ( 
.A(n_10189),
.B(n_9903),
.Y(n_10464)
);

INVx1_ASAP7_75t_L g10465 ( 
.A(n_9964),
.Y(n_10465)
);

AND2x2_ASAP7_75t_L g10466 ( 
.A(n_10075),
.B(n_9776),
.Y(n_10466)
);

INVx2_ASAP7_75t_L g10467 ( 
.A(n_9972),
.Y(n_10467)
);

NAND2xp5_ASAP7_75t_L g10468 ( 
.A(n_10307),
.B(n_9903),
.Y(n_10468)
);

OR2x2_ASAP7_75t_L g10469 ( 
.A(n_10220),
.B(n_9785),
.Y(n_10469)
);

AND2x2_ASAP7_75t_L g10470 ( 
.A(n_10049),
.B(n_9776),
.Y(n_10470)
);

OR2x2_ASAP7_75t_L g10471 ( 
.A(n_10193),
.B(n_9785),
.Y(n_10471)
);

INVx1_ASAP7_75t_L g10472 ( 
.A(n_9970),
.Y(n_10472)
);

OR2x2_ASAP7_75t_L g10473 ( 
.A(n_10196),
.B(n_9787),
.Y(n_10473)
);

INVx1_ASAP7_75t_L g10474 ( 
.A(n_9970),
.Y(n_10474)
);

INVx2_ASAP7_75t_L g10475 ( 
.A(n_9972),
.Y(n_10475)
);

INVx1_ASAP7_75t_L g10476 ( 
.A(n_9973),
.Y(n_10476)
);

AND2x2_ASAP7_75t_L g10477 ( 
.A(n_10300),
.B(n_9918),
.Y(n_10477)
);

AND2x2_ASAP7_75t_L g10478 ( 
.A(n_10115),
.B(n_10124),
.Y(n_10478)
);

NAND2xp5_ASAP7_75t_L g10479 ( 
.A(n_10285),
.B(n_9918),
.Y(n_10479)
);

OR2x2_ASAP7_75t_L g10480 ( 
.A(n_10269),
.B(n_9787),
.Y(n_10480)
);

INVxp67_ASAP7_75t_SL g10481 ( 
.A(n_9989),
.Y(n_10481)
);

INVx1_ASAP7_75t_L g10482 ( 
.A(n_9973),
.Y(n_10482)
);

AND2x2_ASAP7_75t_L g10483 ( 
.A(n_10126),
.B(n_9843),
.Y(n_10483)
);

AND2x2_ASAP7_75t_L g10484 ( 
.A(n_10109),
.B(n_9843),
.Y(n_10484)
);

INVxp33_ASAP7_75t_L g10485 ( 
.A(n_10267),
.Y(n_10485)
);

OR2x2_ASAP7_75t_L g10486 ( 
.A(n_10279),
.B(n_9570),
.Y(n_10486)
);

HB1xp67_ASAP7_75t_L g10487 ( 
.A(n_9978),
.Y(n_10487)
);

BUFx2_ASAP7_75t_R g10488 ( 
.A(n_10212),
.Y(n_10488)
);

AND2x4_ASAP7_75t_SL g10489 ( 
.A(n_10018),
.B(n_9571),
.Y(n_10489)
);

AOI221x1_ASAP7_75t_L g10490 ( 
.A1(n_9987),
.A2(n_9586),
.B1(n_9593),
.B2(n_9575),
.C(n_9574),
.Y(n_10490)
);

HB1xp67_ASAP7_75t_L g10491 ( 
.A(n_9978),
.Y(n_10491)
);

BUFx2_ASAP7_75t_L g10492 ( 
.A(n_10052),
.Y(n_10492)
);

NOR2xp33_ASAP7_75t_L g10493 ( 
.A(n_10242),
.B(n_9608),
.Y(n_10493)
);

OR2x2_ASAP7_75t_L g10494 ( 
.A(n_10037),
.B(n_9796),
.Y(n_10494)
);

NAND2xp5_ASAP7_75t_L g10495 ( 
.A(n_10285),
.B(n_9524),
.Y(n_10495)
);

AND2x2_ASAP7_75t_L g10496 ( 
.A(n_10132),
.B(n_9929),
.Y(n_10496)
);

HB1xp67_ASAP7_75t_L g10497 ( 
.A(n_10238),
.Y(n_10497)
);

NAND2xp5_ASAP7_75t_L g10498 ( 
.A(n_10070),
.B(n_9532),
.Y(n_10498)
);

HB1xp67_ASAP7_75t_L g10499 ( 
.A(n_10268),
.Y(n_10499)
);

HB1xp67_ASAP7_75t_L g10500 ( 
.A(n_9981),
.Y(n_10500)
);

AND2x2_ASAP7_75t_L g10501 ( 
.A(n_10154),
.B(n_9933),
.Y(n_10501)
);

AND2x2_ASAP7_75t_L g10502 ( 
.A(n_10005),
.B(n_10165),
.Y(n_10502)
);

AND2x2_ASAP7_75t_L g10503 ( 
.A(n_10167),
.B(n_9934),
.Y(n_10503)
);

AND2x2_ASAP7_75t_L g10504 ( 
.A(n_10062),
.B(n_9935),
.Y(n_10504)
);

OR2x2_ASAP7_75t_L g10505 ( 
.A(n_10002),
.B(n_9796),
.Y(n_10505)
);

INVx1_ASAP7_75t_L g10506 ( 
.A(n_9981),
.Y(n_10506)
);

AND2x2_ASAP7_75t_L g10507 ( 
.A(n_10064),
.B(n_9939),
.Y(n_10507)
);

AND2x2_ASAP7_75t_L g10508 ( 
.A(n_10106),
.B(n_9801),
.Y(n_10508)
);

INVx1_ASAP7_75t_L g10509 ( 
.A(n_9985),
.Y(n_10509)
);

HB1xp67_ASAP7_75t_L g10510 ( 
.A(n_9985),
.Y(n_10510)
);

INVx1_ASAP7_75t_L g10511 ( 
.A(n_9975),
.Y(n_10511)
);

INVx2_ASAP7_75t_L g10512 ( 
.A(n_9963),
.Y(n_10512)
);

INVx1_ASAP7_75t_L g10513 ( 
.A(n_9975),
.Y(n_10513)
);

AND2x2_ASAP7_75t_L g10514 ( 
.A(n_10043),
.B(n_9801),
.Y(n_10514)
);

AND2x2_ASAP7_75t_L g10515 ( 
.A(n_10170),
.B(n_9803),
.Y(n_10515)
);

AND2x2_ASAP7_75t_L g10516 ( 
.A(n_10178),
.B(n_9803),
.Y(n_10516)
);

INVx2_ASAP7_75t_SL g10517 ( 
.A(n_10070),
.Y(n_10517)
);

INVx1_ASAP7_75t_L g10518 ( 
.A(n_9979),
.Y(n_10518)
);

OR2x2_ASAP7_75t_L g10519 ( 
.A(n_10169),
.B(n_9915),
.Y(n_10519)
);

AND2x2_ASAP7_75t_L g10520 ( 
.A(n_10245),
.B(n_9813),
.Y(n_10520)
);

OR2x2_ASAP7_75t_L g10521 ( 
.A(n_10146),
.B(n_9917),
.Y(n_10521)
);

AND2x4_ASAP7_75t_SL g10522 ( 
.A(n_10182),
.B(n_9539),
.Y(n_10522)
);

NOR2xp67_ASAP7_75t_L g10523 ( 
.A(n_10235),
.B(n_9860),
.Y(n_10523)
);

AND2x2_ASAP7_75t_L g10524 ( 
.A(n_10033),
.B(n_10047),
.Y(n_10524)
);

AND2x2_ASAP7_75t_L g10525 ( 
.A(n_10232),
.B(n_9813),
.Y(n_10525)
);

NOR2xp33_ASAP7_75t_L g10526 ( 
.A(n_10210),
.B(n_7874),
.Y(n_10526)
);

AND2x2_ASAP7_75t_L g10527 ( 
.A(n_10293),
.B(n_9545),
.Y(n_10527)
);

INVx1_ASAP7_75t_L g10528 ( 
.A(n_9979),
.Y(n_10528)
);

INVx2_ASAP7_75t_L g10529 ( 
.A(n_10078),
.Y(n_10529)
);

INVx1_ASAP7_75t_L g10530 ( 
.A(n_10057),
.Y(n_10530)
);

AND2x2_ASAP7_75t_L g10531 ( 
.A(n_10296),
.B(n_9552),
.Y(n_10531)
);

INVx1_ASAP7_75t_L g10532 ( 
.A(n_10061),
.Y(n_10532)
);

INVx2_ASAP7_75t_SL g10533 ( 
.A(n_10078),
.Y(n_10533)
);

AND2x2_ASAP7_75t_L g10534 ( 
.A(n_10297),
.B(n_10314),
.Y(n_10534)
);

HB1xp67_ASAP7_75t_L g10535 ( 
.A(n_10129),
.Y(n_10535)
);

AND2x2_ASAP7_75t_L g10536 ( 
.A(n_10315),
.B(n_9557),
.Y(n_10536)
);

AND2x2_ASAP7_75t_L g10537 ( 
.A(n_10316),
.B(n_9559),
.Y(n_10537)
);

NOR2x1p5_ASAP7_75t_L g10538 ( 
.A(n_10199),
.B(n_9704),
.Y(n_10538)
);

AND2x4_ASAP7_75t_SL g10539 ( 
.A(n_10090),
.B(n_9880),
.Y(n_10539)
);

NAND2xp5_ASAP7_75t_L g10540 ( 
.A(n_10085),
.B(n_9883),
.Y(n_10540)
);

AND2x2_ASAP7_75t_L g10541 ( 
.A(n_10237),
.B(n_10190),
.Y(n_10541)
);

AND2x2_ASAP7_75t_L g10542 ( 
.A(n_10292),
.B(n_9886),
.Y(n_10542)
);

INVx1_ASAP7_75t_L g10543 ( 
.A(n_10119),
.Y(n_10543)
);

NAND2xp5_ASAP7_75t_L g10544 ( 
.A(n_10085),
.B(n_9887),
.Y(n_10544)
);

INVx2_ASAP7_75t_SL g10545 ( 
.A(n_10159),
.Y(n_10545)
);

NAND2xp5_ASAP7_75t_L g10546 ( 
.A(n_10194),
.B(n_9890),
.Y(n_10546)
);

AND2x2_ASAP7_75t_L g10547 ( 
.A(n_10192),
.B(n_9905),
.Y(n_10547)
);

AND2x2_ASAP7_75t_L g10548 ( 
.A(n_10156),
.B(n_9928),
.Y(n_10548)
);

NAND2x1p5_ASAP7_75t_L g10549 ( 
.A(n_10235),
.B(n_9921),
.Y(n_10549)
);

INVx2_ASAP7_75t_L g10550 ( 
.A(n_9999),
.Y(n_10550)
);

NAND2xp5_ASAP7_75t_L g10551 ( 
.A(n_10201),
.B(n_9514),
.Y(n_10551)
);

AND2x4_ASAP7_75t_L g10552 ( 
.A(n_9999),
.B(n_9955),
.Y(n_10552)
);

INVx1_ASAP7_75t_L g10553 ( 
.A(n_10119),
.Y(n_10553)
);

AND2x2_ASAP7_75t_L g10554 ( 
.A(n_10158),
.B(n_9955),
.Y(n_10554)
);

INVx2_ASAP7_75t_L g10555 ( 
.A(n_10118),
.Y(n_10555)
);

AND2x2_ASAP7_75t_L g10556 ( 
.A(n_10259),
.B(n_9957),
.Y(n_10556)
);

AND2x2_ASAP7_75t_L g10557 ( 
.A(n_10251),
.B(n_9957),
.Y(n_10557)
);

AND2x2_ASAP7_75t_L g10558 ( 
.A(n_10291),
.B(n_9909),
.Y(n_10558)
);

OR2x2_ASAP7_75t_L g10559 ( 
.A(n_10161),
.B(n_9704),
.Y(n_10559)
);

AND2x4_ASAP7_75t_L g10560 ( 
.A(n_10159),
.B(n_9514),
.Y(n_10560)
);

INVx2_ASAP7_75t_L g10561 ( 
.A(n_10118),
.Y(n_10561)
);

NAND2xp5_ASAP7_75t_L g10562 ( 
.A(n_10234),
.B(n_9863),
.Y(n_10562)
);

AND2x2_ASAP7_75t_L g10563 ( 
.A(n_10208),
.B(n_9909),
.Y(n_10563)
);

INVx2_ASAP7_75t_L g10564 ( 
.A(n_10151),
.Y(n_10564)
);

INVx1_ASAP7_75t_L g10565 ( 
.A(n_10120),
.Y(n_10565)
);

NAND2xp5_ASAP7_75t_L g10566 ( 
.A(n_10234),
.B(n_10202),
.Y(n_10566)
);

INVx2_ASAP7_75t_L g10567 ( 
.A(n_10151),
.Y(n_10567)
);

NAND2xp5_ASAP7_75t_L g10568 ( 
.A(n_10108),
.B(n_9863),
.Y(n_10568)
);

INVx2_ASAP7_75t_L g10569 ( 
.A(n_10141),
.Y(n_10569)
);

INVx2_ASAP7_75t_L g10570 ( 
.A(n_10163),
.Y(n_10570)
);

AND2x2_ASAP7_75t_L g10571 ( 
.A(n_10130),
.B(n_9909),
.Y(n_10571)
);

NAND2xp5_ASAP7_75t_L g10572 ( 
.A(n_10125),
.B(n_9864),
.Y(n_10572)
);

INVx2_ASAP7_75t_L g10573 ( 
.A(n_10172),
.Y(n_10573)
);

NAND2x1p5_ASAP7_75t_L g10574 ( 
.A(n_10083),
.B(n_9265),
.Y(n_10574)
);

INVx1_ASAP7_75t_L g10575 ( 
.A(n_10120),
.Y(n_10575)
);

INVx1_ASAP7_75t_L g10576 ( 
.A(n_10121),
.Y(n_10576)
);

INVx1_ASAP7_75t_L g10577 ( 
.A(n_10121),
.Y(n_10577)
);

HB1xp67_ASAP7_75t_L g10578 ( 
.A(n_10129),
.Y(n_10578)
);

INVx2_ASAP7_75t_SL g10579 ( 
.A(n_9977),
.Y(n_10579)
);

AND2x2_ASAP7_75t_L g10580 ( 
.A(n_10260),
.B(n_9909),
.Y(n_10580)
);

AND2x2_ASAP7_75t_L g10581 ( 
.A(n_10306),
.B(n_9909),
.Y(n_10581)
);

OR2x2_ASAP7_75t_L g10582 ( 
.A(n_10015),
.B(n_9729),
.Y(n_10582)
);

INVx1_ASAP7_75t_L g10583 ( 
.A(n_10122),
.Y(n_10583)
);

INVx1_ASAP7_75t_L g10584 ( 
.A(n_10122),
.Y(n_10584)
);

NAND2xp5_ASAP7_75t_L g10585 ( 
.A(n_10191),
.B(n_9864),
.Y(n_10585)
);

AND2x2_ASAP7_75t_L g10586 ( 
.A(n_10133),
.B(n_9909),
.Y(n_10586)
);

AND2x4_ASAP7_75t_SL g10587 ( 
.A(n_10091),
.B(n_9888),
.Y(n_10587)
);

OR2x2_ASAP7_75t_L g10588 ( 
.A(n_10131),
.B(n_9729),
.Y(n_10588)
);

INVx2_ASAP7_75t_L g10589 ( 
.A(n_10206),
.Y(n_10589)
);

INVxp67_ASAP7_75t_L g10590 ( 
.A(n_10200),
.Y(n_10590)
);

AND2x2_ASAP7_75t_L g10591 ( 
.A(n_10219),
.B(n_9836),
.Y(n_10591)
);

AND2x2_ASAP7_75t_L g10592 ( 
.A(n_10265),
.B(n_9836),
.Y(n_10592)
);

AND2x2_ASAP7_75t_L g10593 ( 
.A(n_10287),
.B(n_9869),
.Y(n_10593)
);

AND2x2_ASAP7_75t_L g10594 ( 
.A(n_10149),
.B(n_9869),
.Y(n_10594)
);

INVx1_ASAP7_75t_L g10595 ( 
.A(n_10053),
.Y(n_10595)
);

AOI22xp33_ASAP7_75t_L g10596 ( 
.A1(n_9966),
.A2(n_9856),
.B1(n_9919),
.B2(n_9946),
.Y(n_10596)
);

NAND2xp5_ASAP7_75t_SL g10597 ( 
.A(n_10098),
.B(n_9946),
.Y(n_10597)
);

HB1xp67_ASAP7_75t_L g10598 ( 
.A(n_10136),
.Y(n_10598)
);

NAND2xp5_ASAP7_75t_L g10599 ( 
.A(n_10207),
.B(n_9893),
.Y(n_10599)
);

INVx2_ASAP7_75t_L g10600 ( 
.A(n_10103),
.Y(n_10600)
);

INVx1_ASAP7_75t_L g10601 ( 
.A(n_10054),
.Y(n_10601)
);

INVx1_ASAP7_75t_L g10602 ( 
.A(n_10065),
.Y(n_10602)
);

INVx2_ASAP7_75t_L g10603 ( 
.A(n_10103),
.Y(n_10603)
);

INVx2_ASAP7_75t_L g10604 ( 
.A(n_10140),
.Y(n_10604)
);

NAND2xp5_ASAP7_75t_L g10605 ( 
.A(n_10152),
.B(n_9893),
.Y(n_10605)
);

AND2x2_ASAP7_75t_L g10606 ( 
.A(n_10168),
.B(n_9631),
.Y(n_10606)
);

AND2x4_ASAP7_75t_L g10607 ( 
.A(n_10278),
.B(n_9601),
.Y(n_10607)
);

AND2x2_ASAP7_75t_L g10608 ( 
.A(n_10323),
.B(n_9631),
.Y(n_10608)
);

INVx1_ASAP7_75t_L g10609 ( 
.A(n_10066),
.Y(n_10609)
);

INVx2_ASAP7_75t_SL g10610 ( 
.A(n_10140),
.Y(n_10610)
);

AND2x2_ASAP7_75t_L g10611 ( 
.A(n_10336),
.B(n_9650),
.Y(n_10611)
);

AND2x2_ASAP7_75t_L g10612 ( 
.A(n_10216),
.B(n_9650),
.Y(n_10612)
);

AND2x2_ASAP7_75t_L g10613 ( 
.A(n_10256),
.B(n_9601),
.Y(n_10613)
);

INVx1_ASAP7_75t_SL g10614 ( 
.A(n_10174),
.Y(n_10614)
);

AND2x2_ASAP7_75t_L g10615 ( 
.A(n_10351),
.B(n_9603),
.Y(n_10615)
);

AND2x2_ASAP7_75t_L g10616 ( 
.A(n_10353),
.B(n_9603),
.Y(n_10616)
);

INVx2_ASAP7_75t_L g10617 ( 
.A(n_10215),
.Y(n_10617)
);

INVx1_ASAP7_75t_L g10618 ( 
.A(n_10073),
.Y(n_10618)
);

INVx2_ASAP7_75t_L g10619 ( 
.A(n_10227),
.Y(n_10619)
);

NAND2xp5_ASAP7_75t_L g10620 ( 
.A(n_10368),
.B(n_9920),
.Y(n_10620)
);

AND2x2_ASAP7_75t_L g10621 ( 
.A(n_10367),
.B(n_9800),
.Y(n_10621)
);

INVx1_ASAP7_75t_L g10622 ( 
.A(n_10077),
.Y(n_10622)
);

INVx2_ASAP7_75t_L g10623 ( 
.A(n_10229),
.Y(n_10623)
);

INVx2_ASAP7_75t_L g10624 ( 
.A(n_10262),
.Y(n_10624)
);

INVx1_ASAP7_75t_L g10625 ( 
.A(n_10082),
.Y(n_10625)
);

INVx6_ASAP7_75t_L g10626 ( 
.A(n_10240),
.Y(n_10626)
);

INVx1_ASAP7_75t_L g10627 ( 
.A(n_10084),
.Y(n_10627)
);

NAND2xp5_ASAP7_75t_L g10628 ( 
.A(n_9996),
.B(n_10273),
.Y(n_10628)
);

INVx2_ASAP7_75t_L g10629 ( 
.A(n_10299),
.Y(n_10629)
);

INVx2_ASAP7_75t_L g10630 ( 
.A(n_9996),
.Y(n_10630)
);

INVx2_ASAP7_75t_L g10631 ( 
.A(n_10344),
.Y(n_10631)
);

AND2x4_ASAP7_75t_L g10632 ( 
.A(n_9986),
.B(n_9920),
.Y(n_10632)
);

OR2x2_ASAP7_75t_L g10633 ( 
.A(n_10099),
.B(n_9841),
.Y(n_10633)
);

HB1xp67_ASAP7_75t_L g10634 ( 
.A(n_10136),
.Y(n_10634)
);

BUFx2_ASAP7_75t_L g10635 ( 
.A(n_10045),
.Y(n_10635)
);

INVx2_ASAP7_75t_L g10636 ( 
.A(n_10344),
.Y(n_10636)
);

INVx1_ASAP7_75t_L g10637 ( 
.A(n_10089),
.Y(n_10637)
);

AND2x2_ASAP7_75t_L g10638 ( 
.A(n_10342),
.B(n_9800),
.Y(n_10638)
);

INVx2_ASAP7_75t_L g10639 ( 
.A(n_10345),
.Y(n_10639)
);

OR2x2_ASAP7_75t_L g10640 ( 
.A(n_10004),
.B(n_9953),
.Y(n_10640)
);

OR2x2_ASAP7_75t_L g10641 ( 
.A(n_10007),
.B(n_9953),
.Y(n_10641)
);

INVx2_ASAP7_75t_L g10642 ( 
.A(n_10345),
.Y(n_10642)
);

INVx2_ASAP7_75t_L g10643 ( 
.A(n_10363),
.Y(n_10643)
);

NAND2xp5_ASAP7_75t_L g10644 ( 
.A(n_10195),
.B(n_9878),
.Y(n_10644)
);

AND2x2_ASAP7_75t_L g10645 ( 
.A(n_10359),
.B(n_9266),
.Y(n_10645)
);

INVx1_ASAP7_75t_L g10646 ( 
.A(n_10092),
.Y(n_10646)
);

AND2x2_ASAP7_75t_L g10647 ( 
.A(n_10346),
.B(n_9266),
.Y(n_10647)
);

INVx1_ASAP7_75t_L g10648 ( 
.A(n_10008),
.Y(n_10648)
);

NOR2xp33_ASAP7_75t_L g10649 ( 
.A(n_9959),
.B(n_7973),
.Y(n_10649)
);

NAND2xp5_ASAP7_75t_L g10650 ( 
.A(n_10240),
.B(n_9885),
.Y(n_10650)
);

OR2x2_ASAP7_75t_L g10651 ( 
.A(n_10284),
.B(n_9872),
.Y(n_10651)
);

INVx2_ASAP7_75t_L g10652 ( 
.A(n_10363),
.Y(n_10652)
);

OR2x2_ASAP7_75t_L g10653 ( 
.A(n_10302),
.B(n_10303),
.Y(n_10653)
);

AND2x2_ASAP7_75t_L g10654 ( 
.A(n_10038),
.B(n_9271),
.Y(n_10654)
);

INVxp67_ASAP7_75t_SL g10655 ( 
.A(n_10023),
.Y(n_10655)
);

NOR2xp33_ASAP7_75t_L g10656 ( 
.A(n_10153),
.B(n_9856),
.Y(n_10656)
);

INVx2_ASAP7_75t_L g10657 ( 
.A(n_10028),
.Y(n_10657)
);

AND2x2_ASAP7_75t_L g10658 ( 
.A(n_10253),
.B(n_9271),
.Y(n_10658)
);

NAND2xp5_ASAP7_75t_L g10659 ( 
.A(n_10013),
.B(n_9737),
.Y(n_10659)
);

INVx2_ASAP7_75t_SL g10660 ( 
.A(n_9994),
.Y(n_10660)
);

OR2x2_ASAP7_75t_L g10661 ( 
.A(n_10347),
.B(n_9529),
.Y(n_10661)
);

OR2x2_ASAP7_75t_L g10662 ( 
.A(n_9997),
.B(n_9529),
.Y(n_10662)
);

AND2x2_ASAP7_75t_L g10663 ( 
.A(n_10068),
.B(n_9272),
.Y(n_10663)
);

NAND2xp5_ASAP7_75t_L g10664 ( 
.A(n_10014),
.B(n_9744),
.Y(n_10664)
);

INVx2_ASAP7_75t_L g10665 ( 
.A(n_10035),
.Y(n_10665)
);

OR2x2_ASAP7_75t_L g10666 ( 
.A(n_10039),
.B(n_9549),
.Y(n_10666)
);

INVx1_ASAP7_75t_L g10667 ( 
.A(n_10042),
.Y(n_10667)
);

AND2x2_ASAP7_75t_L g10668 ( 
.A(n_10087),
.B(n_9272),
.Y(n_10668)
);

CKINVDCx16_ASAP7_75t_R g10669 ( 
.A(n_10157),
.Y(n_10669)
);

AND2x2_ASAP7_75t_L g10670 ( 
.A(n_10135),
.B(n_9277),
.Y(n_10670)
);

OR2x2_ASAP7_75t_L g10671 ( 
.A(n_10093),
.B(n_9549),
.Y(n_10671)
);

AND2x2_ASAP7_75t_L g10672 ( 
.A(n_10031),
.B(n_9277),
.Y(n_10672)
);

INVx1_ASAP7_75t_L g10673 ( 
.A(n_10044),
.Y(n_10673)
);

OR2x2_ASAP7_75t_L g10674 ( 
.A(n_10164),
.B(n_9751),
.Y(n_10674)
);

AND2x2_ASAP7_75t_L g10675 ( 
.A(n_10040),
.B(n_9283),
.Y(n_10675)
);

INVx2_ASAP7_75t_L g10676 ( 
.A(n_10254),
.Y(n_10676)
);

INVx1_ASAP7_75t_L g10677 ( 
.A(n_10340),
.Y(n_10677)
);

AND2x2_ASAP7_75t_L g10678 ( 
.A(n_10055),
.B(n_9283),
.Y(n_10678)
);

INVx1_ASAP7_75t_L g10679 ( 
.A(n_10348),
.Y(n_10679)
);

INVx1_ASAP7_75t_L g10680 ( 
.A(n_10361),
.Y(n_10680)
);

BUFx3_ASAP7_75t_L g10681 ( 
.A(n_10294),
.Y(n_10681)
);

INVx2_ASAP7_75t_L g10682 ( 
.A(n_10254),
.Y(n_10682)
);

NAND2xp5_ASAP7_75t_L g10683 ( 
.A(n_10123),
.B(n_9764),
.Y(n_10683)
);

INVx1_ASAP7_75t_L g10684 ( 
.A(n_10046),
.Y(n_10684)
);

AND2x2_ASAP7_75t_L g10685 ( 
.A(n_10056),
.B(n_9289),
.Y(n_10685)
);

INVx1_ASAP7_75t_L g10686 ( 
.A(n_10048),
.Y(n_10686)
);

INVx1_ASAP7_75t_L g10687 ( 
.A(n_10050),
.Y(n_10687)
);

AND2x2_ASAP7_75t_L g10688 ( 
.A(n_10059),
.B(n_9289),
.Y(n_10688)
);

NOR2xp33_ASAP7_75t_L g10689 ( 
.A(n_10009),
.B(n_9889),
.Y(n_10689)
);

INVx1_ASAP7_75t_L g10690 ( 
.A(n_10094),
.Y(n_10690)
);

INVx1_ASAP7_75t_L g10691 ( 
.A(n_10095),
.Y(n_10691)
);

NAND2xp5_ASAP7_75t_L g10692 ( 
.A(n_10270),
.B(n_9765),
.Y(n_10692)
);

AND2x2_ASAP7_75t_L g10693 ( 
.A(n_10063),
.B(n_9770),
.Y(n_10693)
);

AND2x2_ASAP7_75t_L g10694 ( 
.A(n_10071),
.B(n_9774),
.Y(n_10694)
);

AND2x2_ASAP7_75t_L g10695 ( 
.A(n_10270),
.B(n_9777),
.Y(n_10695)
);

AND2x2_ASAP7_75t_L g10696 ( 
.A(n_10277),
.B(n_9805),
.Y(n_10696)
);

INVx1_ASAP7_75t_L g10697 ( 
.A(n_10096),
.Y(n_10697)
);

BUFx3_ASAP7_75t_L g10698 ( 
.A(n_10016),
.Y(n_10698)
);

INVx1_ASAP7_75t_L g10699 ( 
.A(n_10104),
.Y(n_10699)
);

OR2x2_ASAP7_75t_L g10700 ( 
.A(n_10166),
.B(n_9807),
.Y(n_10700)
);

AND2x2_ASAP7_75t_L g10701 ( 
.A(n_10277),
.B(n_9808),
.Y(n_10701)
);

INVx2_ASAP7_75t_SL g10702 ( 
.A(n_10286),
.Y(n_10702)
);

AND2x4_ASAP7_75t_SL g10703 ( 
.A(n_9958),
.B(n_9892),
.Y(n_10703)
);

INVx1_ASAP7_75t_L g10704 ( 
.A(n_10110),
.Y(n_10704)
);

INVx1_ASAP7_75t_L g10705 ( 
.A(n_10116),
.Y(n_10705)
);

NAND2xp5_ASAP7_75t_L g10706 ( 
.A(n_10160),
.B(n_9809),
.Y(n_10706)
);

NAND2xp5_ASAP7_75t_L g10707 ( 
.A(n_10286),
.B(n_9810),
.Y(n_10707)
);

NAND2xp5_ASAP7_75t_L g10708 ( 
.A(n_10155),
.B(n_9819),
.Y(n_10708)
);

AND2x2_ASAP7_75t_L g10709 ( 
.A(n_10177),
.B(n_9821),
.Y(n_10709)
);

AND2x2_ASAP7_75t_L g10710 ( 
.A(n_10305),
.B(n_9822),
.Y(n_10710)
);

INVxp67_ASAP7_75t_L g10711 ( 
.A(n_10022),
.Y(n_10711)
);

AND2x2_ASAP7_75t_L g10712 ( 
.A(n_10313),
.B(n_9824),
.Y(n_10712)
);

INVx2_ASAP7_75t_L g10713 ( 
.A(n_9971),
.Y(n_10713)
);

AND2x2_ASAP7_75t_L g10714 ( 
.A(n_10321),
.B(n_9825),
.Y(n_10714)
);

NAND2x1p5_ASAP7_75t_L g10715 ( 
.A(n_10322),
.B(n_9387),
.Y(n_10715)
);

AND2x4_ASAP7_75t_L g10716 ( 
.A(n_10324),
.B(n_9827),
.Y(n_10716)
);

INVx1_ASAP7_75t_L g10717 ( 
.A(n_10176),
.Y(n_10717)
);

INVx4_ASAP7_75t_L g10718 ( 
.A(n_10325),
.Y(n_10718)
);

NAND2xp5_ASAP7_75t_L g10719 ( 
.A(n_10011),
.B(n_9829),
.Y(n_10719)
);

INVx1_ASAP7_75t_L g10720 ( 
.A(n_10176),
.Y(n_10720)
);

AND2x2_ASAP7_75t_L g10721 ( 
.A(n_10326),
.B(n_9830),
.Y(n_10721)
);

AND2x2_ASAP7_75t_L g10722 ( 
.A(n_10333),
.B(n_9832),
.Y(n_10722)
);

OR2x2_ASAP7_75t_L g10723 ( 
.A(n_10185),
.B(n_9849),
.Y(n_10723)
);

NAND2xp5_ASAP7_75t_L g10724 ( 
.A(n_10230),
.B(n_9851),
.Y(n_10724)
);

AND2x2_ASAP7_75t_L g10725 ( 
.A(n_10357),
.B(n_9852),
.Y(n_10725)
);

AND2x2_ASAP7_75t_L g10726 ( 
.A(n_10142),
.B(n_9857),
.Y(n_10726)
);

INVx2_ASAP7_75t_L g10727 ( 
.A(n_10026),
.Y(n_10727)
);

AND2x4_ASAP7_75t_L g10728 ( 
.A(n_10217),
.B(n_9859),
.Y(n_10728)
);

NAND2xp5_ASAP7_75t_L g10729 ( 
.A(n_10308),
.B(n_9865),
.Y(n_10729)
);

INVx1_ASAP7_75t_L g10730 ( 
.A(n_10180),
.Y(n_10730)
);

INVx2_ASAP7_75t_SL g10731 ( 
.A(n_10224),
.Y(n_10731)
);

NOR2xp67_ASAP7_75t_L g10732 ( 
.A(n_10029),
.B(n_9678),
.Y(n_10732)
);

AND2x2_ASAP7_75t_L g10733 ( 
.A(n_10247),
.B(n_9894),
.Y(n_10733)
);

INVx2_ASAP7_75t_L g10734 ( 
.A(n_10365),
.Y(n_10734)
);

INVx1_ASAP7_75t_SL g10735 ( 
.A(n_10188),
.Y(n_10735)
);

INVx1_ASAP7_75t_L g10736 ( 
.A(n_10180),
.Y(n_10736)
);

AND2x2_ASAP7_75t_L g10737 ( 
.A(n_10257),
.B(n_9904),
.Y(n_10737)
);

INVx2_ASAP7_75t_L g10738 ( 
.A(n_10369),
.Y(n_10738)
);

INVx2_ASAP7_75t_L g10739 ( 
.A(n_10370),
.Y(n_10739)
);

NOR2xp67_ASAP7_75t_L g10740 ( 
.A(n_10304),
.B(n_9678),
.Y(n_10740)
);

NAND2xp5_ASAP7_75t_L g10741 ( 
.A(n_10311),
.B(n_9906),
.Y(n_10741)
);

AND2x2_ASAP7_75t_L g10742 ( 
.A(n_10101),
.B(n_9907),
.Y(n_10742)
);

INVx1_ASAP7_75t_SL g10743 ( 
.A(n_10019),
.Y(n_10743)
);

AND2x2_ASAP7_75t_L g10744 ( 
.A(n_10318),
.B(n_9912),
.Y(n_10744)
);

INVx2_ASAP7_75t_L g10745 ( 
.A(n_10334),
.Y(n_10745)
);

INVx2_ASAP7_75t_L g10746 ( 
.A(n_10349),
.Y(n_10746)
);

AND2x4_ASAP7_75t_L g10747 ( 
.A(n_10218),
.B(n_9925),
.Y(n_10747)
);

INVx2_ASAP7_75t_L g10748 ( 
.A(n_10312),
.Y(n_10748)
);

INVx1_ASAP7_75t_L g10749 ( 
.A(n_10181),
.Y(n_10749)
);

INVx3_ASAP7_75t_L g10750 ( 
.A(n_10181),
.Y(n_10750)
);

NOR2xp33_ASAP7_75t_L g10751 ( 
.A(n_10012),
.B(n_9931),
.Y(n_10751)
);

OR2x2_ASAP7_75t_L g10752 ( 
.A(n_10239),
.B(n_9938),
.Y(n_10752)
);

HB1xp67_ASAP7_75t_L g10753 ( 
.A(n_10320),
.Y(n_10753)
);

NAND2xp5_ASAP7_75t_L g10754 ( 
.A(n_10328),
.B(n_9943),
.Y(n_10754)
);

NAND2xp5_ASAP7_75t_L g10755 ( 
.A(n_10329),
.B(n_9947),
.Y(n_10755)
);

INVx1_ASAP7_75t_L g10756 ( 
.A(n_10397),
.Y(n_10756)
);

NAND2x1_ASAP7_75t_L g10757 ( 
.A(n_10626),
.B(n_9919),
.Y(n_10757)
);

OR2x2_ASAP7_75t_L g10758 ( 
.A(n_10669),
.B(n_10034),
.Y(n_10758)
);

NAND2xp5_ASAP7_75t_L g10759 ( 
.A(n_10610),
.B(n_10274),
.Y(n_10759)
);

INVx1_ASAP7_75t_L g10760 ( 
.A(n_10397),
.Y(n_10760)
);

NAND2xp5_ASAP7_75t_L g10761 ( 
.A(n_10445),
.B(n_10069),
.Y(n_10761)
);

INVx1_ASAP7_75t_L g10762 ( 
.A(n_10398),
.Y(n_10762)
);

INVx1_ASAP7_75t_L g10763 ( 
.A(n_10398),
.Y(n_10763)
);

INVx1_ASAP7_75t_L g10764 ( 
.A(n_10492),
.Y(n_10764)
);

INVx2_ASAP7_75t_L g10765 ( 
.A(n_10626),
.Y(n_10765)
);

INVx2_ASAP7_75t_L g10766 ( 
.A(n_10456),
.Y(n_10766)
);

AND2x2_ASAP7_75t_L g10767 ( 
.A(n_10446),
.B(n_10244),
.Y(n_10767)
);

OR2x2_ASAP7_75t_L g10768 ( 
.A(n_10383),
.B(n_10036),
.Y(n_10768)
);

INVx1_ASAP7_75t_L g10769 ( 
.A(n_10487),
.Y(n_10769)
);

NAND2xp5_ASAP7_75t_L g10770 ( 
.A(n_10376),
.B(n_10221),
.Y(n_10770)
);

INVx4_ASAP7_75t_L g10771 ( 
.A(n_10453),
.Y(n_10771)
);

INVx2_ASAP7_75t_L g10772 ( 
.A(n_10456),
.Y(n_10772)
);

INVx2_ASAP7_75t_L g10773 ( 
.A(n_10459),
.Y(n_10773)
);

HB1xp67_ASAP7_75t_L g10774 ( 
.A(n_10491),
.Y(n_10774)
);

AND2x2_ASAP7_75t_L g10775 ( 
.A(n_10449),
.B(n_10222),
.Y(n_10775)
);

INVx1_ASAP7_75t_L g10776 ( 
.A(n_10408),
.Y(n_10776)
);

AND2x2_ASAP7_75t_L g10777 ( 
.A(n_10477),
.B(n_10225),
.Y(n_10777)
);

NAND2xp5_ASAP7_75t_L g10778 ( 
.A(n_10376),
.B(n_10226),
.Y(n_10778)
);

INVx2_ASAP7_75t_L g10779 ( 
.A(n_10459),
.Y(n_10779)
);

INVx1_ASAP7_75t_L g10780 ( 
.A(n_10500),
.Y(n_10780)
);

INVx2_ASAP7_75t_L g10781 ( 
.A(n_10549),
.Y(n_10781)
);

INVx3_ASAP7_75t_L g10782 ( 
.A(n_10552),
.Y(n_10782)
);

AND2x2_ASAP7_75t_L g10783 ( 
.A(n_10478),
.B(n_10231),
.Y(n_10783)
);

NAND2xp5_ASAP7_75t_L g10784 ( 
.A(n_10413),
.B(n_10233),
.Y(n_10784)
);

NAND2xp5_ASAP7_75t_L g10785 ( 
.A(n_10413),
.B(n_10236),
.Y(n_10785)
);

AND2x2_ASAP7_75t_L g10786 ( 
.A(n_10466),
.B(n_10331),
.Y(n_10786)
);

AND2x2_ASAP7_75t_L g10787 ( 
.A(n_10373),
.B(n_10298),
.Y(n_10787)
);

INVx1_ASAP7_75t_L g10788 ( 
.A(n_10510),
.Y(n_10788)
);

INVxp67_ASAP7_75t_SL g10789 ( 
.A(n_10523),
.Y(n_10789)
);

AND2x2_ASAP7_75t_L g10790 ( 
.A(n_10451),
.B(n_10350),
.Y(n_10790)
);

AND2x2_ASAP7_75t_L g10791 ( 
.A(n_10524),
.B(n_10350),
.Y(n_10791)
);

INVx1_ASAP7_75t_L g10792 ( 
.A(n_10535),
.Y(n_10792)
);

INVx1_ASAP7_75t_L g10793 ( 
.A(n_10578),
.Y(n_10793)
);

AND2x4_ASAP7_75t_L g10794 ( 
.A(n_10552),
.B(n_10184),
.Y(n_10794)
);

AND2x2_ASAP7_75t_L g10795 ( 
.A(n_10541),
.B(n_10356),
.Y(n_10795)
);

INVx1_ASAP7_75t_L g10796 ( 
.A(n_10598),
.Y(n_10796)
);

INVx1_ASAP7_75t_L g10797 ( 
.A(n_10634),
.Y(n_10797)
);

INVx2_ASAP7_75t_SL g10798 ( 
.A(n_10414),
.Y(n_10798)
);

INVx1_ASAP7_75t_L g10799 ( 
.A(n_10401),
.Y(n_10799)
);

AND2x4_ASAP7_75t_L g10800 ( 
.A(n_10414),
.B(n_10184),
.Y(n_10800)
);

AND2x4_ASAP7_75t_SL g10801 ( 
.A(n_10375),
.B(n_10241),
.Y(n_10801)
);

INVx1_ASAP7_75t_L g10802 ( 
.A(n_10436),
.Y(n_10802)
);

INVx2_ASAP7_75t_L g10803 ( 
.A(n_10574),
.Y(n_10803)
);

AND2x2_ASAP7_75t_L g10804 ( 
.A(n_10425),
.B(n_10356),
.Y(n_10804)
);

INVx1_ASAP7_75t_L g10805 ( 
.A(n_10454),
.Y(n_10805)
);

INVx1_ASAP7_75t_L g10806 ( 
.A(n_10481),
.Y(n_10806)
);

AND2x2_ASAP7_75t_L g10807 ( 
.A(n_10432),
.B(n_10470),
.Y(n_10807)
);

NAND2xp5_ASAP7_75t_L g10808 ( 
.A(n_10621),
.B(n_10341),
.Y(n_10808)
);

INVx2_ASAP7_75t_L g10809 ( 
.A(n_10715),
.Y(n_10809)
);

NAND2xp5_ASAP7_75t_L g10810 ( 
.A(n_10545),
.B(n_10266),
.Y(n_10810)
);

AND2x2_ASAP7_75t_L g10811 ( 
.A(n_10534),
.B(n_10111),
.Y(n_10811)
);

AND3x2_ASAP7_75t_L g10812 ( 
.A(n_10458),
.B(n_10197),
.C(n_10186),
.Y(n_10812)
);

NAND2xp5_ASAP7_75t_SL g10813 ( 
.A(n_10579),
.B(n_9599),
.Y(n_10813)
);

INVx1_ASAP7_75t_L g10814 ( 
.A(n_10411),
.Y(n_10814)
);

INVx2_ASAP7_75t_L g10815 ( 
.A(n_10448),
.Y(n_10815)
);

INVx3_ASAP7_75t_L g10816 ( 
.A(n_10448),
.Y(n_10816)
);

BUFx3_ASAP7_75t_L g10817 ( 
.A(n_10380),
.Y(n_10817)
);

INVx2_ASAP7_75t_L g10818 ( 
.A(n_10702),
.Y(n_10818)
);

INVx1_ASAP7_75t_L g10819 ( 
.A(n_10426),
.Y(n_10819)
);

INVx1_ASAP7_75t_L g10820 ( 
.A(n_10426),
.Y(n_10820)
);

AND2x2_ASAP7_75t_L g10821 ( 
.A(n_10384),
.B(n_10405),
.Y(n_10821)
);

AND2x2_ASAP7_75t_L g10822 ( 
.A(n_10422),
.B(n_10127),
.Y(n_10822)
);

AOI22xp5_ASAP7_75t_L g10823 ( 
.A1(n_10656),
.A2(n_10041),
.B1(n_9991),
.B2(n_10310),
.Y(n_10823)
);

NAND2xp5_ASAP7_75t_L g10824 ( 
.A(n_10517),
.B(n_10223),
.Y(n_10824)
);

INVx1_ASAP7_75t_L g10825 ( 
.A(n_10427),
.Y(n_10825)
);

HB1xp67_ASAP7_75t_L g10826 ( 
.A(n_10607),
.Y(n_10826)
);

AND2x2_ASAP7_75t_L g10827 ( 
.A(n_10461),
.B(n_10134),
.Y(n_10827)
);

INVx1_ASAP7_75t_L g10828 ( 
.A(n_10427),
.Y(n_10828)
);

INVx2_ASAP7_75t_L g10829 ( 
.A(n_10440),
.Y(n_10829)
);

OR2x2_ASAP7_75t_L g10830 ( 
.A(n_10420),
.B(n_10138),
.Y(n_10830)
);

AND2x2_ASAP7_75t_L g10831 ( 
.A(n_10431),
.B(n_10248),
.Y(n_10831)
);

INVx1_ASAP7_75t_L g10832 ( 
.A(n_10439),
.Y(n_10832)
);

OR2x2_ASAP7_75t_L g10833 ( 
.A(n_10457),
.B(n_10024),
.Y(n_10833)
);

INVx1_ASAP7_75t_L g10834 ( 
.A(n_10439),
.Y(n_10834)
);

INVx1_ASAP7_75t_L g10835 ( 
.A(n_10443),
.Y(n_10835)
);

INVx1_ASAP7_75t_L g10836 ( 
.A(n_10443),
.Y(n_10836)
);

INVx1_ASAP7_75t_L g10837 ( 
.A(n_10750),
.Y(n_10837)
);

AND2x2_ASAP7_75t_L g10838 ( 
.A(n_10404),
.B(n_10250),
.Y(n_10838)
);

INVx1_ASAP7_75t_L g10839 ( 
.A(n_10750),
.Y(n_10839)
);

OR2x2_ASAP7_75t_L g10840 ( 
.A(n_10533),
.B(n_10282),
.Y(n_10840)
);

INVx1_ASAP7_75t_L g10841 ( 
.A(n_10631),
.Y(n_10841)
);

INVx2_ASAP7_75t_L g10842 ( 
.A(n_10440),
.Y(n_10842)
);

AND2x2_ASAP7_75t_L g10843 ( 
.A(n_10514),
.B(n_10261),
.Y(n_10843)
);

NAND2xp5_ASAP7_75t_L g10844 ( 
.A(n_10638),
.B(n_10107),
.Y(n_10844)
);

AND2x2_ASAP7_75t_L g10845 ( 
.A(n_10382),
.B(n_10263),
.Y(n_10845)
);

INVx1_ASAP7_75t_L g10846 ( 
.A(n_10636),
.Y(n_10846)
);

OR2x2_ASAP7_75t_L g10847 ( 
.A(n_10562),
.B(n_10276),
.Y(n_10847)
);

NAND2xp5_ASAP7_75t_L g10848 ( 
.A(n_10560),
.B(n_10264),
.Y(n_10848)
);

AND2x2_ASAP7_75t_L g10849 ( 
.A(n_10502),
.B(n_10272),
.Y(n_10849)
);

NAND2xp5_ASAP7_75t_L g10850 ( 
.A(n_10560),
.B(n_10280),
.Y(n_10850)
);

NOR2xp33_ASAP7_75t_L g10851 ( 
.A(n_10488),
.B(n_10355),
.Y(n_10851)
);

AND2x2_ASAP7_75t_L g10852 ( 
.A(n_10423),
.B(n_10455),
.Y(n_10852)
);

NAND2xp5_ASAP7_75t_L g10853 ( 
.A(n_10591),
.B(n_10283),
.Y(n_10853)
);

INVx1_ASAP7_75t_L g10854 ( 
.A(n_10639),
.Y(n_10854)
);

AND2x2_ASAP7_75t_L g10855 ( 
.A(n_10483),
.B(n_10288),
.Y(n_10855)
);

OR2x2_ASAP7_75t_L g10856 ( 
.A(n_10438),
.B(n_10258),
.Y(n_10856)
);

NAND2xp5_ASAP7_75t_L g10857 ( 
.A(n_10508),
.B(n_10290),
.Y(n_10857)
);

OR2x2_ASAP7_75t_L g10858 ( 
.A(n_10403),
.B(n_10319),
.Y(n_10858)
);

AND2x2_ASAP7_75t_L g10859 ( 
.A(n_10394),
.B(n_10301),
.Y(n_10859)
);

INVxp67_ASAP7_75t_L g10860 ( 
.A(n_10497),
.Y(n_10860)
);

AND2x2_ASAP7_75t_L g10861 ( 
.A(n_10385),
.B(n_10309),
.Y(n_10861)
);

OR2x2_ASAP7_75t_L g10862 ( 
.A(n_10387),
.B(n_10330),
.Y(n_10862)
);

INVx1_ASAP7_75t_L g10863 ( 
.A(n_10642),
.Y(n_10863)
);

INVx1_ASAP7_75t_L g10864 ( 
.A(n_10643),
.Y(n_10864)
);

NAND2xp5_ASAP7_75t_L g10865 ( 
.A(n_10600),
.B(n_10360),
.Y(n_10865)
);

INVx1_ASAP7_75t_L g10866 ( 
.A(n_10652),
.Y(n_10866)
);

AND2x2_ASAP7_75t_L g10867 ( 
.A(n_10393),
.B(n_10360),
.Y(n_10867)
);

NAND2xp5_ASAP7_75t_L g10868 ( 
.A(n_10603),
.B(n_10362),
.Y(n_10868)
);

AND2x2_ASAP7_75t_L g10869 ( 
.A(n_10507),
.B(n_10362),
.Y(n_10869)
);

INVx1_ASAP7_75t_L g10870 ( 
.A(n_10412),
.Y(n_10870)
);

NOR2xp33_ASAP7_75t_L g10871 ( 
.A(n_10450),
.B(n_10252),
.Y(n_10871)
);

INVx2_ASAP7_75t_L g10872 ( 
.A(n_10607),
.Y(n_10872)
);

AND2x2_ASAP7_75t_L g10873 ( 
.A(n_10407),
.B(n_10366),
.Y(n_10873)
);

OR2x2_ASAP7_75t_L g10874 ( 
.A(n_10604),
.B(n_10335),
.Y(n_10874)
);

INVx2_ASAP7_75t_L g10875 ( 
.A(n_10453),
.Y(n_10875)
);

INVx1_ASAP7_75t_L g10876 ( 
.A(n_10495),
.Y(n_10876)
);

AND2x2_ASAP7_75t_L g10877 ( 
.A(n_10460),
.B(n_10366),
.Y(n_10877)
);

NAND2xp5_ASAP7_75t_L g10878 ( 
.A(n_10429),
.B(n_10371),
.Y(n_10878)
);

AND2x2_ASAP7_75t_L g10879 ( 
.A(n_10557),
.B(n_10371),
.Y(n_10879)
);

INVxp67_ASAP7_75t_L g10880 ( 
.A(n_10499),
.Y(n_10880)
);

INVx2_ASAP7_75t_L g10881 ( 
.A(n_10489),
.Y(n_10881)
);

AND2x2_ASAP7_75t_L g10882 ( 
.A(n_10378),
.B(n_10372),
.Y(n_10882)
);

INVxp67_ASAP7_75t_L g10883 ( 
.A(n_10526),
.Y(n_10883)
);

OR2x2_ASAP7_75t_L g10884 ( 
.A(n_10529),
.B(n_10337),
.Y(n_10884)
);

AND2x2_ASAP7_75t_L g10885 ( 
.A(n_10430),
.B(n_10372),
.Y(n_10885)
);

AND2x2_ASAP7_75t_L g10886 ( 
.A(n_10395),
.B(n_10186),
.Y(n_10886)
);

INVx1_ASAP7_75t_L g10887 ( 
.A(n_10550),
.Y(n_10887)
);

AND2x2_ASAP7_75t_L g10888 ( 
.A(n_10406),
.B(n_10197),
.Y(n_10888)
);

INVx1_ASAP7_75t_L g10889 ( 
.A(n_10536),
.Y(n_10889)
);

INVx1_ASAP7_75t_SL g10890 ( 
.A(n_10522),
.Y(n_10890)
);

AND2x2_ASAP7_75t_L g10891 ( 
.A(n_10592),
.B(n_10198),
.Y(n_10891)
);

HB1xp67_ASAP7_75t_L g10892 ( 
.A(n_10732),
.Y(n_10892)
);

INVx1_ASAP7_75t_L g10893 ( 
.A(n_10537),
.Y(n_10893)
);

HB1xp67_ASAP7_75t_L g10894 ( 
.A(n_10467),
.Y(n_10894)
);

INVx1_ASAP7_75t_L g10895 ( 
.A(n_10676),
.Y(n_10895)
);

INVx1_ASAP7_75t_L g10896 ( 
.A(n_10682),
.Y(n_10896)
);

OR2x2_ASAP7_75t_L g10897 ( 
.A(n_10391),
.B(n_10338),
.Y(n_10897)
);

NAND2xp5_ASAP7_75t_L g10898 ( 
.A(n_10520),
.B(n_10198),
.Y(n_10898)
);

OR2x2_ASAP7_75t_L g10899 ( 
.A(n_10498),
.B(n_10519),
.Y(n_10899)
);

INVx1_ASAP7_75t_L g10900 ( 
.A(n_10543),
.Y(n_10900)
);

INVx2_ASAP7_75t_L g10901 ( 
.A(n_10475),
.Y(n_10901)
);

NAND2xp5_ASAP7_75t_L g10902 ( 
.A(n_10525),
.B(n_10204),
.Y(n_10902)
);

AND2x2_ASAP7_75t_L g10903 ( 
.A(n_10421),
.B(n_10204),
.Y(n_10903)
);

INVx1_ASAP7_75t_SL g10904 ( 
.A(n_10614),
.Y(n_10904)
);

OR2x2_ASAP7_75t_L g10905 ( 
.A(n_10396),
.B(n_10352),
.Y(n_10905)
);

INVx3_ASAP7_75t_L g10906 ( 
.A(n_10718),
.Y(n_10906)
);

AND2x4_ASAP7_75t_L g10907 ( 
.A(n_10564),
.B(n_10213),
.Y(n_10907)
);

NAND2x1p5_ASAP7_75t_L g10908 ( 
.A(n_10558),
.B(n_10213),
.Y(n_10908)
);

INVx3_ASAP7_75t_L g10909 ( 
.A(n_10718),
.Y(n_10909)
);

AND2x4_ASAP7_75t_L g10910 ( 
.A(n_10567),
.B(n_10214),
.Y(n_10910)
);

NOR2xp33_ASAP7_75t_SL g10911 ( 
.A(n_10743),
.B(n_10442),
.Y(n_10911)
);

INVx1_ASAP7_75t_L g10912 ( 
.A(n_10543),
.Y(n_10912)
);

INVx1_ASAP7_75t_L g10913 ( 
.A(n_10553),
.Y(n_10913)
);

NAND2xp5_ASAP7_75t_L g10914 ( 
.A(n_10515),
.B(n_10214),
.Y(n_10914)
);

INVx2_ASAP7_75t_L g10915 ( 
.A(n_10402),
.Y(n_10915)
);

AOI22xp5_ASAP7_75t_L g10916 ( 
.A1(n_10596),
.A2(n_10740),
.B1(n_9599),
.B2(n_9634),
.Y(n_10916)
);

AND2x2_ASAP7_75t_L g10917 ( 
.A(n_10484),
.B(n_10354),
.Y(n_10917)
);

OAI21xp5_ASAP7_75t_L g10918 ( 
.A1(n_10490),
.A2(n_10597),
.B(n_10339),
.Y(n_10918)
);

BUFx2_ASAP7_75t_L g10919 ( 
.A(n_10433),
.Y(n_10919)
);

INVx1_ASAP7_75t_L g10920 ( 
.A(n_10553),
.Y(n_10920)
);

INVx1_ASAP7_75t_L g10921 ( 
.A(n_10565),
.Y(n_10921)
);

INVx2_ASAP7_75t_L g10922 ( 
.A(n_10419),
.Y(n_10922)
);

AND2x2_ASAP7_75t_L g10923 ( 
.A(n_10415),
.B(n_10358),
.Y(n_10923)
);

INVx3_ASAP7_75t_L g10924 ( 
.A(n_10381),
.Y(n_10924)
);

INVx2_ASAP7_75t_L g10925 ( 
.A(n_10516),
.Y(n_10925)
);

INVx1_ASAP7_75t_L g10926 ( 
.A(n_10565),
.Y(n_10926)
);

AOI22xp5_ASAP7_75t_L g10927 ( 
.A1(n_10726),
.A2(n_9634),
.B1(n_10249),
.B2(n_9675),
.Y(n_10927)
);

NOR3xp33_ASAP7_75t_L g10928 ( 
.A(n_10452),
.B(n_10364),
.C(n_9675),
.Y(n_10928)
);

INVx2_ASAP7_75t_L g10929 ( 
.A(n_10388),
.Y(n_10929)
);

OR2x2_ASAP7_75t_L g10930 ( 
.A(n_10386),
.B(n_9949),
.Y(n_10930)
);

INVx1_ASAP7_75t_SL g10931 ( 
.A(n_10424),
.Y(n_10931)
);

INVx3_ASAP7_75t_L g10932 ( 
.A(n_10390),
.Y(n_10932)
);

AND2x2_ASAP7_75t_L g10933 ( 
.A(n_10379),
.B(n_9954),
.Y(n_10933)
);

OR2x2_ASAP7_75t_L g10934 ( 
.A(n_10605),
.B(n_9155),
.Y(n_10934)
);

INVxp67_ASAP7_75t_SL g10935 ( 
.A(n_10418),
.Y(n_10935)
);

NOR2xp33_ASAP7_75t_L g10936 ( 
.A(n_10485),
.B(n_10698),
.Y(n_10936)
);

AND2x2_ASAP7_75t_L g10937 ( 
.A(n_10416),
.B(n_9156),
.Y(n_10937)
);

INVx1_ASAP7_75t_L g10938 ( 
.A(n_10575),
.Y(n_10938)
);

HB1xp67_ASAP7_75t_L g10939 ( 
.A(n_10479),
.Y(n_10939)
);

NAND2xp5_ASAP7_75t_L g10940 ( 
.A(n_10556),
.B(n_9182),
.Y(n_10940)
);

NOR2x1_ASAP7_75t_L g10941 ( 
.A(n_10680),
.B(n_9680),
.Y(n_10941)
);

NAND2xp5_ASAP7_75t_L g10942 ( 
.A(n_10554),
.B(n_9187),
.Y(n_10942)
);

INVx2_ASAP7_75t_L g10943 ( 
.A(n_10374),
.Y(n_10943)
);

NAND2xp5_ASAP7_75t_L g10944 ( 
.A(n_10527),
.B(n_9189),
.Y(n_10944)
);

INVxp67_ASAP7_75t_L g10945 ( 
.A(n_10463),
.Y(n_10945)
);

NAND2xp5_ASAP7_75t_L g10946 ( 
.A(n_10531),
.B(n_9195),
.Y(n_10946)
);

NOR2xp33_ASAP7_75t_L g10947 ( 
.A(n_10711),
.B(n_10392),
.Y(n_10947)
);

INVx1_ASAP7_75t_L g10948 ( 
.A(n_10575),
.Y(n_10948)
);

INVx1_ASAP7_75t_L g10949 ( 
.A(n_10576),
.Y(n_10949)
);

NAND2x1p5_ASAP7_75t_L g10950 ( 
.A(n_10580),
.B(n_9387),
.Y(n_10950)
);

AND2x4_ASAP7_75t_L g10951 ( 
.A(n_10695),
.B(n_9196),
.Y(n_10951)
);

OR2x2_ASAP7_75t_L g10952 ( 
.A(n_10464),
.B(n_10551),
.Y(n_10952)
);

NAND2x1p5_ASAP7_75t_L g10953 ( 
.A(n_10581),
.B(n_8741),
.Y(n_10953)
);

OR2x2_ASAP7_75t_L g10954 ( 
.A(n_10468),
.B(n_9203),
.Y(n_10954)
);

INVx1_ASAP7_75t_L g10955 ( 
.A(n_10576),
.Y(n_10955)
);

INVx1_ASAP7_75t_L g10956 ( 
.A(n_10577),
.Y(n_10956)
);

OR2x2_ASAP7_75t_L g10957 ( 
.A(n_10471),
.B(n_9218),
.Y(n_10957)
);

INVx1_ASAP7_75t_L g10958 ( 
.A(n_10577),
.Y(n_10958)
);

INVx1_ASAP7_75t_L g10959 ( 
.A(n_10583),
.Y(n_10959)
);

OR2x2_ASAP7_75t_L g10960 ( 
.A(n_10473),
.B(n_9221),
.Y(n_10960)
);

INVx1_ASAP7_75t_L g10961 ( 
.A(n_10583),
.Y(n_10961)
);

NOR2x1p5_ASAP7_75t_L g10962 ( 
.A(n_10566),
.B(n_9224),
.Y(n_10962)
);

AND2x2_ASAP7_75t_L g10963 ( 
.A(n_10504),
.B(n_9228),
.Y(n_10963)
);

INVx1_ASAP7_75t_L g10964 ( 
.A(n_10584),
.Y(n_10964)
);

INVx1_ASAP7_75t_L g10965 ( 
.A(n_10584),
.Y(n_10965)
);

AND2x2_ASAP7_75t_L g10966 ( 
.A(n_10608),
.B(n_9236),
.Y(n_10966)
);

AND2x4_ASAP7_75t_L g10967 ( 
.A(n_10696),
.B(n_9238),
.Y(n_10967)
);

AND2x2_ASAP7_75t_L g10968 ( 
.A(n_10611),
.B(n_9239),
.Y(n_10968)
);

NAND2xp5_ASAP7_75t_L g10969 ( 
.A(n_10615),
.B(n_9244),
.Y(n_10969)
);

OR2x2_ASAP7_75t_L g10970 ( 
.A(n_10480),
.B(n_9247),
.Y(n_10970)
);

AND2x2_ASAP7_75t_L g10971 ( 
.A(n_10593),
.B(n_10612),
.Y(n_10971)
);

AND2x2_ASAP7_75t_L g10972 ( 
.A(n_10606),
.B(n_9248),
.Y(n_10972)
);

NAND2xp5_ASAP7_75t_L g10973 ( 
.A(n_10616),
.B(n_9249),
.Y(n_10973)
);

INVx1_ASAP7_75t_L g10974 ( 
.A(n_10635),
.Y(n_10974)
);

INVx1_ASAP7_75t_L g10975 ( 
.A(n_10506),
.Y(n_10975)
);

INVx1_ASAP7_75t_L g10976 ( 
.A(n_10506),
.Y(n_10976)
);

AND2x2_ASAP7_75t_L g10977 ( 
.A(n_10496),
.B(n_9250),
.Y(n_10977)
);

NAND2xp5_ASAP7_75t_L g10978 ( 
.A(n_10647),
.B(n_9251),
.Y(n_10978)
);

INVxp67_ASAP7_75t_L g10979 ( 
.A(n_10447),
.Y(n_10979)
);

NAND2xp5_ASAP7_75t_L g10980 ( 
.A(n_10658),
.B(n_10645),
.Y(n_10980)
);

INVx1_ASAP7_75t_L g10981 ( 
.A(n_10509),
.Y(n_10981)
);

INVx2_ASAP7_75t_L g10982 ( 
.A(n_10681),
.Y(n_10982)
);

OAI22xp33_ASAP7_75t_L g10983 ( 
.A1(n_10683),
.A2(n_9680),
.B1(n_8631),
.B2(n_8638),
.Y(n_10983)
);

AND2x2_ASAP7_75t_L g10984 ( 
.A(n_10594),
.B(n_9261),
.Y(n_10984)
);

NAND2xp5_ASAP7_75t_SL g10985 ( 
.A(n_10512),
.B(n_9845),
.Y(n_10985)
);

INVx2_ASAP7_75t_L g10986 ( 
.A(n_10632),
.Y(n_10986)
);

AND2x2_ASAP7_75t_L g10987 ( 
.A(n_10501),
.B(n_9263),
.Y(n_10987)
);

INVx2_ASAP7_75t_L g10988 ( 
.A(n_10632),
.Y(n_10988)
);

AND2x2_ASAP7_75t_L g10989 ( 
.A(n_10503),
.B(n_9268),
.Y(n_10989)
);

INVx1_ASAP7_75t_SL g10990 ( 
.A(n_10539),
.Y(n_10990)
);

AND2x2_ASAP7_75t_SL g10991 ( 
.A(n_10582),
.B(n_9275),
.Y(n_10991)
);

INVx1_ASAP7_75t_L g10992 ( 
.A(n_10509),
.Y(n_10992)
);

OR2x2_ASAP7_75t_L g10993 ( 
.A(n_10444),
.B(n_9279),
.Y(n_10993)
);

AND2x2_ASAP7_75t_L g10994 ( 
.A(n_10547),
.B(n_9284),
.Y(n_10994)
);

INVx1_ASAP7_75t_L g10995 ( 
.A(n_10462),
.Y(n_10995)
);

AND2x4_ASAP7_75t_SL g10996 ( 
.A(n_10571),
.B(n_9286),
.Y(n_10996)
);

NAND2xp5_ASAP7_75t_L g10997 ( 
.A(n_10613),
.B(n_9290),
.Y(n_10997)
);

INVx1_ASAP7_75t_L g10998 ( 
.A(n_10462),
.Y(n_10998)
);

INVx1_ASAP7_75t_L g10999 ( 
.A(n_10465),
.Y(n_10999)
);

INVx1_ASAP7_75t_L g11000 ( 
.A(n_10465),
.Y(n_11000)
);

INVx1_ASAP7_75t_L g11001 ( 
.A(n_10472),
.Y(n_11001)
);

INVx1_ASAP7_75t_L g11002 ( 
.A(n_10472),
.Y(n_11002)
);

NAND2xp5_ASAP7_75t_L g11003 ( 
.A(n_10542),
.B(n_9292),
.Y(n_11003)
);

INVx3_ASAP7_75t_L g11004 ( 
.A(n_10716),
.Y(n_11004)
);

INVx1_ASAP7_75t_L g11005 ( 
.A(n_10474),
.Y(n_11005)
);

HB1xp67_ASAP7_75t_L g11006 ( 
.A(n_10400),
.Y(n_11006)
);

NOR2x1_ASAP7_75t_L g11007 ( 
.A(n_10680),
.B(n_9695),
.Y(n_11007)
);

AND2x2_ASAP7_75t_L g11008 ( 
.A(n_10548),
.B(n_10654),
.Y(n_11008)
);

INVx1_ASAP7_75t_L g11009 ( 
.A(n_10474),
.Y(n_11009)
);

INVx2_ASAP7_75t_L g11010 ( 
.A(n_10586),
.Y(n_11010)
);

NAND2xp5_ASAP7_75t_L g11011 ( 
.A(n_10660),
.B(n_9294),
.Y(n_11011)
);

INVx1_ASAP7_75t_L g11012 ( 
.A(n_10377),
.Y(n_11012)
);

INVx2_ASAP7_75t_L g11013 ( 
.A(n_10563),
.Y(n_11013)
);

AND2x2_ASAP7_75t_L g11014 ( 
.A(n_10663),
.B(n_9295),
.Y(n_11014)
);

HB1xp67_ASAP7_75t_L g11015 ( 
.A(n_10400),
.Y(n_11015)
);

INVx1_ASAP7_75t_L g11016 ( 
.A(n_10377),
.Y(n_11016)
);

INVx3_ASAP7_75t_L g11017 ( 
.A(n_10716),
.Y(n_11017)
);

HB1xp67_ASAP7_75t_L g11018 ( 
.A(n_10409),
.Y(n_11018)
);

INVx1_ASAP7_75t_L g11019 ( 
.A(n_10389),
.Y(n_11019)
);

INVx1_ASAP7_75t_L g11020 ( 
.A(n_10389),
.Y(n_11020)
);

CKINVDCx16_ASAP7_75t_R g11021 ( 
.A(n_10633),
.Y(n_11021)
);

AND2x2_ASAP7_75t_L g11022 ( 
.A(n_10668),
.B(n_9297),
.Y(n_11022)
);

NAND2xp5_ASAP7_75t_L g11023 ( 
.A(n_10555),
.B(n_9300),
.Y(n_11023)
);

AND2x2_ASAP7_75t_L g11024 ( 
.A(n_10649),
.B(n_9301),
.Y(n_11024)
);

INVx2_ASAP7_75t_SL g11025 ( 
.A(n_10703),
.Y(n_11025)
);

OR2x2_ASAP7_75t_L g11026 ( 
.A(n_10428),
.B(n_9310),
.Y(n_11026)
);

NAND2x1p5_ASAP7_75t_L g11027 ( 
.A(n_10435),
.B(n_10561),
.Y(n_11027)
);

AND2x2_ASAP7_75t_L g11028 ( 
.A(n_10735),
.B(n_9312),
.Y(n_11028)
);

INVx2_ASAP7_75t_L g11029 ( 
.A(n_10701),
.Y(n_11029)
);

INVx1_ASAP7_75t_L g11030 ( 
.A(n_10476),
.Y(n_11030)
);

INVx2_ASAP7_75t_SL g11031 ( 
.A(n_10587),
.Y(n_11031)
);

INVxp67_ASAP7_75t_L g11032 ( 
.A(n_10493),
.Y(n_11032)
);

AND2x2_ASAP7_75t_L g11033 ( 
.A(n_10670),
.B(n_9313),
.Y(n_11033)
);

AND2x2_ASAP7_75t_L g11034 ( 
.A(n_10727),
.B(n_9318),
.Y(n_11034)
);

OR2x2_ASAP7_75t_L g11035 ( 
.A(n_10540),
.B(n_9321),
.Y(n_11035)
);

NOR2xp33_ASAP7_75t_L g11036 ( 
.A(n_10590),
.B(n_9322),
.Y(n_11036)
);

NOR2xp33_ASAP7_75t_L g11037 ( 
.A(n_10417),
.B(n_9324),
.Y(n_11037)
);

NAND2xp5_ASAP7_75t_L g11038 ( 
.A(n_10630),
.B(n_9327),
.Y(n_11038)
);

INVx1_ASAP7_75t_L g11039 ( 
.A(n_10476),
.Y(n_11039)
);

INVx2_ASAP7_75t_L g11040 ( 
.A(n_10486),
.Y(n_11040)
);

INVxp67_ASAP7_75t_L g11041 ( 
.A(n_10399),
.Y(n_11041)
);

OR2x2_ASAP7_75t_L g11042 ( 
.A(n_10544),
.B(n_9335),
.Y(n_11042)
);

NAND2xp5_ASAP7_75t_L g11043 ( 
.A(n_10655),
.B(n_9695),
.Y(n_11043)
);

AND2x2_ASAP7_75t_L g11044 ( 
.A(n_10731),
.B(n_8985),
.Y(n_11044)
);

INVx2_ASAP7_75t_SL g11045 ( 
.A(n_10677),
.Y(n_11045)
);

AND2x2_ASAP7_75t_L g11046 ( 
.A(n_10538),
.B(n_8994),
.Y(n_11046)
);

AND2x2_ASAP7_75t_L g11047 ( 
.A(n_10672),
.B(n_8995),
.Y(n_11047)
);

AND2x2_ASAP7_75t_L g11048 ( 
.A(n_10675),
.B(n_9001),
.Y(n_11048)
);

OR2x2_ASAP7_75t_L g11049 ( 
.A(n_10588),
.B(n_9004),
.Y(n_11049)
);

INVx1_ASAP7_75t_L g11050 ( 
.A(n_10482),
.Y(n_11050)
);

AND2x2_ASAP7_75t_L g11051 ( 
.A(n_10678),
.B(n_9005),
.Y(n_11051)
);

AND2x2_ASAP7_75t_L g11052 ( 
.A(n_10746),
.B(n_9006),
.Y(n_11052)
);

AND2x2_ASAP7_75t_L g11053 ( 
.A(n_10569),
.B(n_9010),
.Y(n_11053)
);

INVx1_ASAP7_75t_SL g11054 ( 
.A(n_10653),
.Y(n_11054)
);

INVx1_ASAP7_75t_L g11055 ( 
.A(n_10482),
.Y(n_11055)
);

AND2x2_ASAP7_75t_L g11056 ( 
.A(n_10570),
.B(n_10573),
.Y(n_11056)
);

AND2x2_ASAP7_75t_L g11057 ( 
.A(n_10589),
.B(n_9014),
.Y(n_11057)
);

OR2x2_ASAP7_75t_L g11058 ( 
.A(n_10469),
.B(n_9015),
.Y(n_11058)
);

OR2x2_ASAP7_75t_L g11059 ( 
.A(n_10568),
.B(n_9017),
.Y(n_11059)
);

INVx2_ASAP7_75t_SL g11060 ( 
.A(n_10679),
.Y(n_11060)
);

NAND2xp5_ASAP7_75t_L g11061 ( 
.A(n_10685),
.B(n_9020),
.Y(n_11061)
);

AND2x2_ASAP7_75t_L g11062 ( 
.A(n_10617),
.B(n_9025),
.Y(n_11062)
);

AND2x2_ASAP7_75t_L g11063 ( 
.A(n_10619),
.B(n_9081),
.Y(n_11063)
);

INVx1_ASAP7_75t_L g11064 ( 
.A(n_10511),
.Y(n_11064)
);

NAND2xp5_ASAP7_75t_L g11065 ( 
.A(n_10688),
.B(n_9520),
.Y(n_11065)
);

INVx2_ASAP7_75t_L g11066 ( 
.A(n_10409),
.Y(n_11066)
);

INVx1_ASAP7_75t_L g11067 ( 
.A(n_10511),
.Y(n_11067)
);

OR2x2_ASAP7_75t_L g11068 ( 
.A(n_10572),
.B(n_9427),
.Y(n_11068)
);

NOR2xp33_ASAP7_75t_L g11069 ( 
.A(n_10628),
.B(n_8741),
.Y(n_11069)
);

AND2x2_ASAP7_75t_L g11070 ( 
.A(n_10623),
.B(n_10624),
.Y(n_11070)
);

INVx1_ASAP7_75t_L g11071 ( 
.A(n_10513),
.Y(n_11071)
);

NAND2xp5_ASAP7_75t_L g11072 ( 
.A(n_10713),
.B(n_9520),
.Y(n_11072)
);

INVx2_ASAP7_75t_L g11073 ( 
.A(n_10521),
.Y(n_11073)
);

INVxp67_ASAP7_75t_L g11074 ( 
.A(n_10620),
.Y(n_11074)
);

INVx1_ASAP7_75t_L g11075 ( 
.A(n_10513),
.Y(n_11075)
);

INVx2_ASAP7_75t_L g11076 ( 
.A(n_10518),
.Y(n_11076)
);

INVx2_ASAP7_75t_L g11077 ( 
.A(n_10518),
.Y(n_11077)
);

AND2x2_ASAP7_75t_L g11078 ( 
.A(n_10629),
.B(n_9081),
.Y(n_11078)
);

NOR2x1_ASAP7_75t_L g11079 ( 
.A(n_10528),
.B(n_9845),
.Y(n_11079)
);

AND2x2_ASAP7_75t_L g11080 ( 
.A(n_10739),
.B(n_9081),
.Y(n_11080)
);

INVx2_ASAP7_75t_L g11081 ( 
.A(n_10528),
.Y(n_11081)
);

OR2x2_ASAP7_75t_L g11082 ( 
.A(n_10661),
.B(n_9412),
.Y(n_11082)
);

OR2x2_ASAP7_75t_L g11083 ( 
.A(n_10585),
.B(n_9184),
.Y(n_11083)
);

INVx1_ASAP7_75t_L g11084 ( 
.A(n_10717),
.Y(n_11084)
);

NAND2xp5_ASAP7_75t_SL g11085 ( 
.A(n_10745),
.B(n_9855),
.Y(n_11085)
);

OR2x2_ASAP7_75t_L g11086 ( 
.A(n_10599),
.B(n_9341),
.Y(n_11086)
);

INVx1_ASAP7_75t_L g11087 ( 
.A(n_10826),
.Y(n_11087)
);

INVx2_ASAP7_75t_L g11088 ( 
.A(n_10782),
.Y(n_11088)
);

OR2x2_ASAP7_75t_L g11089 ( 
.A(n_11021),
.B(n_10640),
.Y(n_11089)
);

OR2x2_ASAP7_75t_L g11090 ( 
.A(n_10798),
.B(n_10641),
.Y(n_11090)
);

INVx2_ASAP7_75t_L g11091 ( 
.A(n_10782),
.Y(n_11091)
);

OR2x2_ASAP7_75t_L g11092 ( 
.A(n_10774),
.B(n_10559),
.Y(n_11092)
);

AND2x2_ASAP7_75t_L g11093 ( 
.A(n_10852),
.B(n_10748),
.Y(n_11093)
);

INVx1_ASAP7_75t_L g11094 ( 
.A(n_11007),
.Y(n_11094)
);

NAND2xp5_ASAP7_75t_L g11095 ( 
.A(n_10816),
.B(n_10657),
.Y(n_11095)
);

AND2x2_ASAP7_75t_L g11096 ( 
.A(n_10821),
.B(n_10737),
.Y(n_11096)
);

INVx2_ASAP7_75t_L g11097 ( 
.A(n_10816),
.Y(n_11097)
);

AND2x2_ASAP7_75t_L g11098 ( 
.A(n_10807),
.B(n_10734),
.Y(n_11098)
);

AND2x2_ASAP7_75t_L g11099 ( 
.A(n_10881),
.B(n_10738),
.Y(n_11099)
);

NOR2xp33_ASAP7_75t_L g11100 ( 
.A(n_10911),
.B(n_10494),
.Y(n_11100)
);

NAND2xp5_ASAP7_75t_L g11101 ( 
.A(n_10812),
.B(n_10665),
.Y(n_11101)
);

HB1xp67_ASAP7_75t_L g11102 ( 
.A(n_10892),
.Y(n_11102)
);

AND2x2_ASAP7_75t_L g11103 ( 
.A(n_11008),
.B(n_10733),
.Y(n_11103)
);

AND2x2_ASAP7_75t_L g11104 ( 
.A(n_10822),
.B(n_10817),
.Y(n_11104)
);

HB1xp67_ASAP7_75t_L g11105 ( 
.A(n_11004),
.Y(n_11105)
);

INVx2_ASAP7_75t_SL g11106 ( 
.A(n_10800),
.Y(n_11106)
);

AND2x2_ASAP7_75t_L g11107 ( 
.A(n_10767),
.B(n_10742),
.Y(n_11107)
);

AND2x2_ASAP7_75t_L g11108 ( 
.A(n_10845),
.B(n_10709),
.Y(n_11108)
);

AND2x2_ASAP7_75t_L g11109 ( 
.A(n_10890),
.B(n_10693),
.Y(n_11109)
);

AND2x2_ASAP7_75t_L g11110 ( 
.A(n_10827),
.B(n_10694),
.Y(n_11110)
);

AND2x2_ASAP7_75t_L g11111 ( 
.A(n_10990),
.B(n_10753),
.Y(n_11111)
);

INVx1_ASAP7_75t_L g11112 ( 
.A(n_10941),
.Y(n_11112)
);

INVx2_ASAP7_75t_SL g11113 ( 
.A(n_10800),
.Y(n_11113)
);

AND2x2_ASAP7_75t_L g11114 ( 
.A(n_10811),
.B(n_10410),
.Y(n_11114)
);

HB1xp67_ASAP7_75t_L g11115 ( 
.A(n_11004),
.Y(n_11115)
);

INVx4_ASAP7_75t_L g11116 ( 
.A(n_10771),
.Y(n_11116)
);

AND2x2_ASAP7_75t_L g11117 ( 
.A(n_11025),
.B(n_10546),
.Y(n_11117)
);

INVx1_ASAP7_75t_L g11118 ( 
.A(n_11017),
.Y(n_11118)
);

NAND2x1p5_ASAP7_75t_L g11119 ( 
.A(n_10771),
.B(n_10747),
.Y(n_11119)
);

INVx1_ASAP7_75t_L g11120 ( 
.A(n_11017),
.Y(n_11120)
);

AND2x4_ASAP7_75t_L g11121 ( 
.A(n_10794),
.B(n_10789),
.Y(n_11121)
);

HB1xp67_ASAP7_75t_L g11122 ( 
.A(n_11027),
.Y(n_11122)
);

AND2x2_ASAP7_75t_L g11123 ( 
.A(n_10971),
.B(n_10751),
.Y(n_11123)
);

INVx2_ASAP7_75t_L g11124 ( 
.A(n_10953),
.Y(n_11124)
);

INVx2_ASAP7_75t_L g11125 ( 
.A(n_10794),
.Y(n_11125)
);

OR2x2_ASAP7_75t_L g11126 ( 
.A(n_10810),
.B(n_10505),
.Y(n_11126)
);

AND2x4_ASAP7_75t_L g11127 ( 
.A(n_10766),
.B(n_10728),
.Y(n_11127)
);

INVx3_ASAP7_75t_L g11128 ( 
.A(n_10906),
.Y(n_11128)
);

INVx1_ASAP7_75t_L g11129 ( 
.A(n_11079),
.Y(n_11129)
);

INVx1_ASAP7_75t_L g11130 ( 
.A(n_10894),
.Y(n_11130)
);

NAND2xp5_ASAP7_75t_L g11131 ( 
.A(n_10829),
.B(n_10842),
.Y(n_11131)
);

NOR2xp33_ASAP7_75t_L g11132 ( 
.A(n_10904),
.B(n_10666),
.Y(n_11132)
);

AND2x4_ASAP7_75t_L g11133 ( 
.A(n_10772),
.B(n_10728),
.Y(n_11133)
);

AND2x2_ASAP7_75t_L g11134 ( 
.A(n_10765),
.B(n_10651),
.Y(n_11134)
);

HB1xp67_ASAP7_75t_L g11135 ( 
.A(n_10906),
.Y(n_11135)
);

AND2x2_ASAP7_75t_L g11136 ( 
.A(n_10787),
.B(n_10710),
.Y(n_11136)
);

NAND2xp5_ASAP7_75t_L g11137 ( 
.A(n_10891),
.B(n_10667),
.Y(n_11137)
);

INVx1_ASAP7_75t_L g11138 ( 
.A(n_10769),
.Y(n_11138)
);

NAND2xp5_ASAP7_75t_L g11139 ( 
.A(n_10764),
.B(n_10673),
.Y(n_11139)
);

INVx3_ASAP7_75t_L g11140 ( 
.A(n_10909),
.Y(n_11140)
);

OR2x2_ASAP7_75t_L g11141 ( 
.A(n_10856),
.B(n_10650),
.Y(n_11141)
);

INVx1_ASAP7_75t_L g11142 ( 
.A(n_10769),
.Y(n_11142)
);

AND2x2_ASAP7_75t_L g11143 ( 
.A(n_10831),
.B(n_10712),
.Y(n_11143)
);

AND2x2_ASAP7_75t_SL g11144 ( 
.A(n_10801),
.B(n_10441),
.Y(n_11144)
);

AND2x2_ASAP7_75t_L g11145 ( 
.A(n_11031),
.B(n_10714),
.Y(n_11145)
);

AND2x2_ASAP7_75t_L g11146 ( 
.A(n_10775),
.B(n_10721),
.Y(n_11146)
);

OR2x2_ASAP7_75t_L g11147 ( 
.A(n_10773),
.B(n_10671),
.Y(n_11147)
);

INVx2_ASAP7_75t_SL g11148 ( 
.A(n_10996),
.Y(n_11148)
);

INVx1_ASAP7_75t_L g11149 ( 
.A(n_10779),
.Y(n_11149)
);

INVx1_ASAP7_75t_L g11150 ( 
.A(n_10919),
.Y(n_11150)
);

INVx1_ASAP7_75t_L g11151 ( 
.A(n_10886),
.Y(n_11151)
);

INVx2_ASAP7_75t_L g11152 ( 
.A(n_10909),
.Y(n_11152)
);

AND2x2_ASAP7_75t_L g11153 ( 
.A(n_10849),
.B(n_10722),
.Y(n_11153)
);

NAND2xp5_ASAP7_75t_L g11154 ( 
.A(n_10764),
.B(n_10618),
.Y(n_11154)
);

NAND2xp5_ASAP7_75t_L g11155 ( 
.A(n_10815),
.B(n_10622),
.Y(n_11155)
);

NAND2xp5_ASAP7_75t_L g11156 ( 
.A(n_10924),
.B(n_10725),
.Y(n_11156)
);

NAND2xp5_ASAP7_75t_L g11157 ( 
.A(n_10924),
.B(n_10684),
.Y(n_11157)
);

INVx1_ASAP7_75t_L g11158 ( 
.A(n_10867),
.Y(n_11158)
);

NAND2xp5_ASAP7_75t_L g11159 ( 
.A(n_10932),
.B(n_10684),
.Y(n_11159)
);

INVx3_ASAP7_75t_R g11160 ( 
.A(n_10758),
.Y(n_11160)
);

NAND2xp5_ASAP7_75t_L g11161 ( 
.A(n_10932),
.B(n_10686),
.Y(n_11161)
);

AND2x2_ASAP7_75t_L g11162 ( 
.A(n_10777),
.B(n_10689),
.Y(n_11162)
);

AND2x2_ASAP7_75t_L g11163 ( 
.A(n_10791),
.B(n_10744),
.Y(n_11163)
);

AND2x2_ASAP7_75t_L g11164 ( 
.A(n_10790),
.B(n_10786),
.Y(n_11164)
);

INVx1_ASAP7_75t_L g11165 ( 
.A(n_10873),
.Y(n_11165)
);

INVx1_ASAP7_75t_L g11166 ( 
.A(n_10888),
.Y(n_11166)
);

INVxp67_ASAP7_75t_L g11167 ( 
.A(n_10851),
.Y(n_11167)
);

INVx1_ASAP7_75t_L g11168 ( 
.A(n_10903),
.Y(n_11168)
);

AND2x2_ASAP7_75t_L g11169 ( 
.A(n_10923),
.B(n_10686),
.Y(n_11169)
);

NAND2xp5_ASAP7_75t_L g11170 ( 
.A(n_10879),
.B(n_10687),
.Y(n_11170)
);

AND2x2_ASAP7_75t_L g11171 ( 
.A(n_10818),
.B(n_10687),
.Y(n_11171)
);

NAND2xp5_ASAP7_75t_SL g11172 ( 
.A(n_10918),
.B(n_10662),
.Y(n_11172)
);

AND2x2_ASAP7_75t_L g11173 ( 
.A(n_10859),
.B(n_10648),
.Y(n_11173)
);

OR2x2_ASAP7_75t_L g11174 ( 
.A(n_10840),
.B(n_10706),
.Y(n_11174)
);

OR2x2_ASAP7_75t_L g11175 ( 
.A(n_10759),
.B(n_10719),
.Y(n_11175)
);

NAND2xp5_ASAP7_75t_L g11176 ( 
.A(n_10872),
.B(n_10648),
.Y(n_11176)
);

AND2x2_ASAP7_75t_L g11177 ( 
.A(n_10861),
.B(n_10690),
.Y(n_11177)
);

AND2x2_ASAP7_75t_L g11178 ( 
.A(n_10783),
.B(n_10690),
.Y(n_11178)
);

INVx1_ASAP7_75t_L g11179 ( 
.A(n_11006),
.Y(n_11179)
);

NAND2xp5_ASAP7_75t_L g11180 ( 
.A(n_10885),
.B(n_10877),
.Y(n_11180)
);

AND2x4_ASAP7_75t_L g11181 ( 
.A(n_10803),
.B(n_10747),
.Y(n_11181)
);

INVx2_ASAP7_75t_L g11182 ( 
.A(n_10908),
.Y(n_11182)
);

INVx2_ASAP7_75t_SL g11183 ( 
.A(n_10907),
.Y(n_11183)
);

AND2x2_ASAP7_75t_L g11184 ( 
.A(n_10925),
.B(n_10691),
.Y(n_11184)
);

OR2x2_ASAP7_75t_L g11185 ( 
.A(n_10931),
.B(n_10692),
.Y(n_11185)
);

INVx1_ASAP7_75t_L g11186 ( 
.A(n_11015),
.Y(n_11186)
);

NOR2xp33_ASAP7_75t_L g11187 ( 
.A(n_11041),
.B(n_10860),
.Y(n_11187)
);

AND2x2_ASAP7_75t_L g11188 ( 
.A(n_10917),
.B(n_10691),
.Y(n_11188)
);

OR2x2_ASAP7_75t_L g11189 ( 
.A(n_11054),
.B(n_10729),
.Y(n_11189)
);

NAND2xp5_ASAP7_75t_L g11190 ( 
.A(n_10869),
.B(n_10697),
.Y(n_11190)
);

INVx1_ASAP7_75t_SL g11191 ( 
.A(n_10795),
.Y(n_11191)
);

AND2x2_ASAP7_75t_L g11192 ( 
.A(n_11029),
.B(n_10697),
.Y(n_11192)
);

INVx2_ASAP7_75t_L g11193 ( 
.A(n_10950),
.Y(n_11193)
);

INVx1_ASAP7_75t_L g11194 ( 
.A(n_11018),
.Y(n_11194)
);

AND2x2_ASAP7_75t_L g11195 ( 
.A(n_10889),
.B(n_10699),
.Y(n_11195)
);

AND2x2_ASAP7_75t_L g11196 ( 
.A(n_10893),
.B(n_10699),
.Y(n_11196)
);

INVx1_ASAP7_75t_L g11197 ( 
.A(n_10756),
.Y(n_11197)
);

OR2x2_ASAP7_75t_L g11198 ( 
.A(n_10768),
.B(n_10724),
.Y(n_11198)
);

INVx1_ASAP7_75t_L g11199 ( 
.A(n_10756),
.Y(n_11199)
);

NAND2xp5_ASAP7_75t_L g11200 ( 
.A(n_10986),
.B(n_10704),
.Y(n_11200)
);

AND2x2_ASAP7_75t_L g11201 ( 
.A(n_10781),
.B(n_10704),
.Y(n_11201)
);

AND2x4_ASAP7_75t_L g11202 ( 
.A(n_10988),
.B(n_10530),
.Y(n_11202)
);

INVx1_ASAP7_75t_L g11203 ( 
.A(n_10760),
.Y(n_11203)
);

INVx1_ASAP7_75t_L g11204 ( 
.A(n_10760),
.Y(n_11204)
);

INVx1_ASAP7_75t_L g11205 ( 
.A(n_10762),
.Y(n_11205)
);

INVx1_ASAP7_75t_L g11206 ( 
.A(n_10762),
.Y(n_11206)
);

OR2x6_ASAP7_75t_L g11207 ( 
.A(n_10982),
.B(n_10644),
.Y(n_11207)
);

INVx2_ASAP7_75t_L g11208 ( 
.A(n_10907),
.Y(n_11208)
);

INVx1_ASAP7_75t_L g11209 ( 
.A(n_10763),
.Y(n_11209)
);

OAI211xp5_ASAP7_75t_L g11210 ( 
.A1(n_10916),
.A2(n_10708),
.B(n_10664),
.C(n_10659),
.Y(n_11210)
);

INVx1_ASAP7_75t_L g11211 ( 
.A(n_10763),
.Y(n_11211)
);

AND2x2_ASAP7_75t_L g11212 ( 
.A(n_10843),
.B(n_10705),
.Y(n_11212)
);

INVx1_ASAP7_75t_L g11213 ( 
.A(n_10838),
.Y(n_11213)
);

AND2x2_ASAP7_75t_L g11214 ( 
.A(n_10935),
.B(n_10705),
.Y(n_11214)
);

AND2x2_ASAP7_75t_L g11215 ( 
.A(n_10855),
.B(n_10530),
.Y(n_11215)
);

OR2x2_ASAP7_75t_L g11216 ( 
.A(n_10899),
.B(n_10707),
.Y(n_11216)
);

AND2x2_ASAP7_75t_L g11217 ( 
.A(n_10804),
.B(n_10532),
.Y(n_11217)
);

NAND2x1_ASAP7_75t_L g11218 ( 
.A(n_10910),
.B(n_10837),
.Y(n_11218)
);

NAND2xp5_ASAP7_75t_L g11219 ( 
.A(n_10901),
.B(n_10882),
.Y(n_11219)
);

OR2x6_ASAP7_75t_L g11220 ( 
.A(n_11040),
.B(n_10532),
.Y(n_11220)
);

INVx2_ASAP7_75t_L g11221 ( 
.A(n_10910),
.Y(n_11221)
);

AND2x2_ASAP7_75t_L g11222 ( 
.A(n_10943),
.B(n_10595),
.Y(n_11222)
);

AND2x2_ASAP7_75t_L g11223 ( 
.A(n_10933),
.B(n_10595),
.Y(n_11223)
);

NAND2xp5_ASAP7_75t_L g11224 ( 
.A(n_10776),
.B(n_10601),
.Y(n_11224)
);

AND2x4_ASAP7_75t_L g11225 ( 
.A(n_10974),
.B(n_10601),
.Y(n_11225)
);

OR2x2_ASAP7_75t_L g11226 ( 
.A(n_10784),
.B(n_10752),
.Y(n_11226)
);

INVx2_ASAP7_75t_L g11227 ( 
.A(n_10809),
.Y(n_11227)
);

INVx1_ASAP7_75t_L g11228 ( 
.A(n_11030),
.Y(n_11228)
);

NAND2xp5_ASAP7_75t_L g11229 ( 
.A(n_10799),
.B(n_10602),
.Y(n_11229)
);

OR2x2_ASAP7_75t_L g11230 ( 
.A(n_10785),
.B(n_10674),
.Y(n_11230)
);

INVx2_ASAP7_75t_L g11231 ( 
.A(n_11010),
.Y(n_11231)
);

INVx1_ASAP7_75t_L g11232 ( 
.A(n_10770),
.Y(n_11232)
);

INVx2_ASAP7_75t_L g11233 ( 
.A(n_10874),
.Y(n_11233)
);

AND2x2_ASAP7_75t_L g11234 ( 
.A(n_10880),
.B(n_10602),
.Y(n_11234)
);

INVx1_ASAP7_75t_L g11235 ( 
.A(n_11030),
.Y(n_11235)
);

NAND2xp5_ASAP7_75t_L g11236 ( 
.A(n_10871),
.B(n_10609),
.Y(n_11236)
);

AOI22xp33_ASAP7_75t_L g11237 ( 
.A1(n_10928),
.A2(n_8478),
.B1(n_8448),
.B2(n_8801),
.Y(n_11237)
);

INVx1_ASAP7_75t_L g11238 ( 
.A(n_11039),
.Y(n_11238)
);

HB1xp67_ASAP7_75t_L g11239 ( 
.A(n_10839),
.Y(n_11239)
);

INVx2_ASAP7_75t_L g11240 ( 
.A(n_10830),
.Y(n_11240)
);

AND2x4_ASAP7_75t_L g11241 ( 
.A(n_10792),
.B(n_10609),
.Y(n_11241)
);

INVx2_ASAP7_75t_L g11242 ( 
.A(n_10858),
.Y(n_11242)
);

INVx2_ASAP7_75t_L g11243 ( 
.A(n_10875),
.Y(n_11243)
);

INVx1_ASAP7_75t_L g11244 ( 
.A(n_11039),
.Y(n_11244)
);

INVx1_ASAP7_75t_L g11245 ( 
.A(n_10778),
.Y(n_11245)
);

INVx1_ASAP7_75t_L g11246 ( 
.A(n_10898),
.Y(n_11246)
);

INVx1_ASAP7_75t_L g11247 ( 
.A(n_10902),
.Y(n_11247)
);

INVx1_ASAP7_75t_SL g11248 ( 
.A(n_11082),
.Y(n_11248)
);

INVx1_ASAP7_75t_L g11249 ( 
.A(n_10914),
.Y(n_11249)
);

INVx1_ASAP7_75t_L g11250 ( 
.A(n_10878),
.Y(n_11250)
);

NAND2xp5_ASAP7_75t_L g11251 ( 
.A(n_10802),
.B(n_10625),
.Y(n_11251)
);

NAND2xp5_ASAP7_75t_L g11252 ( 
.A(n_10805),
.B(n_10625),
.Y(n_11252)
);

NAND2xp5_ASAP7_75t_L g11253 ( 
.A(n_10806),
.B(n_10627),
.Y(n_11253)
);

INVx1_ASAP7_75t_L g11254 ( 
.A(n_11050),
.Y(n_11254)
);

INVx1_ASAP7_75t_L g11255 ( 
.A(n_11050),
.Y(n_11255)
);

INVx1_ASAP7_75t_L g11256 ( 
.A(n_11055),
.Y(n_11256)
);

AND2x2_ASAP7_75t_L g11257 ( 
.A(n_10979),
.B(n_10937),
.Y(n_11257)
);

AND2x2_ASAP7_75t_L g11258 ( 
.A(n_11073),
.B(n_10627),
.Y(n_11258)
);

INVx1_ASAP7_75t_L g11259 ( 
.A(n_11055),
.Y(n_11259)
);

INVx1_ASAP7_75t_L g11260 ( 
.A(n_11064),
.Y(n_11260)
);

NAND2xp5_ASAP7_75t_L g11261 ( 
.A(n_10793),
.B(n_10637),
.Y(n_11261)
);

NAND2xp5_ASAP7_75t_L g11262 ( 
.A(n_10796),
.B(n_10637),
.Y(n_11262)
);

INVx2_ASAP7_75t_L g11263 ( 
.A(n_10884),
.Y(n_11263)
);

NAND2xp5_ASAP7_75t_L g11264 ( 
.A(n_10797),
.B(n_10646),
.Y(n_11264)
);

INVx1_ASAP7_75t_L g11265 ( 
.A(n_11064),
.Y(n_11265)
);

AND2x4_ASAP7_75t_L g11266 ( 
.A(n_10780),
.B(n_10646),
.Y(n_11266)
);

OR2x2_ASAP7_75t_L g11267 ( 
.A(n_10844),
.B(n_10700),
.Y(n_11267)
);

NAND2xp5_ASAP7_75t_L g11268 ( 
.A(n_10870),
.B(n_10434),
.Y(n_11268)
);

NAND2xp5_ASAP7_75t_L g11269 ( 
.A(n_10788),
.B(n_10437),
.Y(n_11269)
);

INVx3_ASAP7_75t_L g11270 ( 
.A(n_10951),
.Y(n_11270)
);

AND2x2_ASAP7_75t_L g11271 ( 
.A(n_10939),
.B(n_11028),
.Y(n_11271)
);

AND2x2_ASAP7_75t_L g11272 ( 
.A(n_10977),
.B(n_10723),
.Y(n_11272)
);

NOR2xp33_ASAP7_75t_L g11273 ( 
.A(n_10761),
.B(n_10741),
.Y(n_11273)
);

AND2x2_ASAP7_75t_L g11274 ( 
.A(n_10915),
.B(n_10717),
.Y(n_11274)
);

INVx1_ASAP7_75t_L g11275 ( 
.A(n_11067),
.Y(n_11275)
);

AND2x2_ASAP7_75t_L g11276 ( 
.A(n_10922),
.B(n_10720),
.Y(n_11276)
);

INVx2_ASAP7_75t_L g11277 ( 
.A(n_11013),
.Y(n_11277)
);

AND2x2_ASAP7_75t_L g11278 ( 
.A(n_10929),
.B(n_10720),
.Y(n_11278)
);

INVx1_ASAP7_75t_L g11279 ( 
.A(n_11067),
.Y(n_11279)
);

INVx1_ASAP7_75t_L g11280 ( 
.A(n_11071),
.Y(n_11280)
);

INVx1_ASAP7_75t_L g11281 ( 
.A(n_11043),
.Y(n_11281)
);

OR2x2_ASAP7_75t_L g11282 ( 
.A(n_10847),
.B(n_10754),
.Y(n_11282)
);

BUFx3_ASAP7_75t_L g11283 ( 
.A(n_10887),
.Y(n_11283)
);

INVx1_ASAP7_75t_SL g11284 ( 
.A(n_10862),
.Y(n_11284)
);

INVx3_ASAP7_75t_L g11285 ( 
.A(n_10951),
.Y(n_11285)
);

INVx2_ASAP7_75t_L g11286 ( 
.A(n_10991),
.Y(n_11286)
);

NAND2xp5_ASAP7_75t_L g11287 ( 
.A(n_10895),
.B(n_10730),
.Y(n_11287)
);

INVx1_ASAP7_75t_L g11288 ( 
.A(n_11071),
.Y(n_11288)
);

INVx1_ASAP7_75t_L g11289 ( 
.A(n_11075),
.Y(n_11289)
);

INVx1_ASAP7_75t_L g11290 ( 
.A(n_11075),
.Y(n_11290)
);

NOR2xp33_ASAP7_75t_L g11291 ( 
.A(n_10980),
.B(n_10755),
.Y(n_11291)
);

INVx1_ASAP7_75t_L g11292 ( 
.A(n_10848),
.Y(n_11292)
);

AND2x2_ASAP7_75t_L g11293 ( 
.A(n_11014),
.B(n_10730),
.Y(n_11293)
);

INVx1_ASAP7_75t_SL g11294 ( 
.A(n_10833),
.Y(n_11294)
);

NAND2xp5_ASAP7_75t_L g11295 ( 
.A(n_10896),
.B(n_10736),
.Y(n_11295)
);

INVx2_ASAP7_75t_L g11296 ( 
.A(n_10905),
.Y(n_11296)
);

NAND2xp5_ASAP7_75t_L g11297 ( 
.A(n_10841),
.B(n_10736),
.Y(n_11297)
);

INVx2_ASAP7_75t_L g11298 ( 
.A(n_10967),
.Y(n_11298)
);

INVx2_ASAP7_75t_L g11299 ( 
.A(n_10967),
.Y(n_11299)
);

INVx2_ASAP7_75t_L g11300 ( 
.A(n_11066),
.Y(n_11300)
);

INVx1_ASAP7_75t_SL g11301 ( 
.A(n_11080),
.Y(n_11301)
);

INVx1_ASAP7_75t_L g11302 ( 
.A(n_10850),
.Y(n_11302)
);

INVx1_ASAP7_75t_L g11303 ( 
.A(n_10853),
.Y(n_11303)
);

AND2x2_ASAP7_75t_L g11304 ( 
.A(n_11022),
.B(n_10749),
.Y(n_11304)
);

OR2x2_ASAP7_75t_L g11305 ( 
.A(n_10824),
.B(n_10749),
.Y(n_11305)
);

INVx1_ASAP7_75t_SL g11306 ( 
.A(n_11063),
.Y(n_11306)
);

INVx1_ASAP7_75t_L g11307 ( 
.A(n_10865),
.Y(n_11307)
);

INVx2_ASAP7_75t_L g11308 ( 
.A(n_10962),
.Y(n_11308)
);

AND2x2_ASAP7_75t_L g11309 ( 
.A(n_11056),
.B(n_9081),
.Y(n_11309)
);

AND2x2_ASAP7_75t_L g11310 ( 
.A(n_11070),
.B(n_8768),
.Y(n_11310)
);

INVx2_ASAP7_75t_L g11311 ( 
.A(n_11047),
.Y(n_11311)
);

NOR2xp33_ASAP7_75t_L g11312 ( 
.A(n_11032),
.B(n_8768),
.Y(n_11312)
);

INVx1_ASAP7_75t_L g11313 ( 
.A(n_10868),
.Y(n_11313)
);

OR2x2_ASAP7_75t_L g11314 ( 
.A(n_10857),
.B(n_9359),
.Y(n_11314)
);

AND2x2_ASAP7_75t_L g11315 ( 
.A(n_11024),
.B(n_8782),
.Y(n_11315)
);

NOR2xp33_ASAP7_75t_SL g11316 ( 
.A(n_10936),
.B(n_8782),
.Y(n_11316)
);

NAND2xp5_ASAP7_75t_L g11317 ( 
.A(n_10846),
.B(n_8445),
.Y(n_11317)
);

INVx1_ASAP7_75t_L g11318 ( 
.A(n_11048),
.Y(n_11318)
);

INVx2_ASAP7_75t_L g11319 ( 
.A(n_11051),
.Y(n_11319)
);

INVx1_ASAP7_75t_L g11320 ( 
.A(n_11084),
.Y(n_11320)
);

INVx1_ASAP7_75t_L g11321 ( 
.A(n_11084),
.Y(n_11321)
);

OR2x2_ASAP7_75t_L g11322 ( 
.A(n_10854),
.B(n_9378),
.Y(n_11322)
);

AND2x2_ASAP7_75t_L g11323 ( 
.A(n_10863),
.B(n_8445),
.Y(n_11323)
);

NAND2xp5_ASAP7_75t_L g11324 ( 
.A(n_10864),
.B(n_8450),
.Y(n_11324)
);

INVx1_ASAP7_75t_L g11325 ( 
.A(n_11012),
.Y(n_11325)
);

AND2x2_ASAP7_75t_L g11326 ( 
.A(n_10866),
.B(n_8450),
.Y(n_11326)
);

NOR2xp33_ASAP7_75t_L g11327 ( 
.A(n_10945),
.B(n_10883),
.Y(n_11327)
);

INVx1_ASAP7_75t_L g11328 ( 
.A(n_11012),
.Y(n_11328)
);

OR2x2_ASAP7_75t_L g11329 ( 
.A(n_10757),
.B(n_10813),
.Y(n_11329)
);

NAND2xp5_ASAP7_75t_L g11330 ( 
.A(n_11045),
.B(n_9855),
.Y(n_11330)
);

INVx1_ASAP7_75t_L g11331 ( 
.A(n_11016),
.Y(n_11331)
);

OR2x2_ASAP7_75t_L g11332 ( 
.A(n_11060),
.B(n_9377),
.Y(n_11332)
);

INVx1_ASAP7_75t_L g11333 ( 
.A(n_11016),
.Y(n_11333)
);

INVx1_ASAP7_75t_L g11334 ( 
.A(n_11019),
.Y(n_11334)
);

INVx1_ASAP7_75t_L g11335 ( 
.A(n_11019),
.Y(n_11335)
);

AND2x2_ASAP7_75t_L g11336 ( 
.A(n_10963),
.B(n_8383),
.Y(n_11336)
);

NAND2xp5_ASAP7_75t_L g11337 ( 
.A(n_11069),
.B(n_8895),
.Y(n_11337)
);

AND2x2_ASAP7_75t_L g11338 ( 
.A(n_10987),
.B(n_8383),
.Y(n_11338)
);

OR2x2_ASAP7_75t_L g11339 ( 
.A(n_10952),
.B(n_9285),
.Y(n_11339)
);

NAND2xp5_ASAP7_75t_L g11340 ( 
.A(n_10823),
.B(n_10927),
.Y(n_11340)
);

INVx2_ASAP7_75t_L g11341 ( 
.A(n_11033),
.Y(n_11341)
);

INVx2_ASAP7_75t_L g11342 ( 
.A(n_10993),
.Y(n_11342)
);

INVx3_ASAP7_75t_SL g11343 ( 
.A(n_10930),
.Y(n_11343)
);

NAND2xp5_ASAP7_75t_L g11344 ( 
.A(n_11078),
.B(n_8362),
.Y(n_11344)
);

OR2x2_ASAP7_75t_L g11345 ( 
.A(n_11068),
.B(n_10897),
.Y(n_11345)
);

INVx2_ASAP7_75t_SL g11346 ( 
.A(n_11026),
.Y(n_11346)
);

NAND2xp5_ASAP7_75t_L g11347 ( 
.A(n_10989),
.B(n_8362),
.Y(n_11347)
);

INVx1_ASAP7_75t_SL g11348 ( 
.A(n_11046),
.Y(n_11348)
);

OR2x2_ASAP7_75t_L g11349 ( 
.A(n_10944),
.B(n_9430),
.Y(n_11349)
);

INVx1_ASAP7_75t_L g11350 ( 
.A(n_11020),
.Y(n_11350)
);

AND2x4_ASAP7_75t_L g11351 ( 
.A(n_10994),
.B(n_8831),
.Y(n_11351)
);

NAND2xp5_ASAP7_75t_L g11352 ( 
.A(n_10966),
.B(n_8364),
.Y(n_11352)
);

INVx1_ASAP7_75t_SL g11353 ( 
.A(n_10968),
.Y(n_11353)
);

INVx2_ASAP7_75t_L g11354 ( 
.A(n_11076),
.Y(n_11354)
);

AND2x2_ASAP7_75t_L g11355 ( 
.A(n_10972),
.B(n_8383),
.Y(n_11355)
);

AND2x2_ASAP7_75t_L g11356 ( 
.A(n_10984),
.B(n_8349),
.Y(n_11356)
);

INVx1_ASAP7_75t_SL g11357 ( 
.A(n_11044),
.Y(n_11357)
);

AOI21xp33_ASAP7_75t_L g11358 ( 
.A1(n_10808),
.A2(n_10947),
.B(n_10814),
.Y(n_11358)
);

AND2x2_ASAP7_75t_L g11359 ( 
.A(n_10876),
.B(n_8349),
.Y(n_11359)
);

INVx2_ASAP7_75t_L g11360 ( 
.A(n_11077),
.Y(n_11360)
);

INVx2_ASAP7_75t_L g11361 ( 
.A(n_11081),
.Y(n_11361)
);

INVx1_ASAP7_75t_L g11362 ( 
.A(n_11020),
.Y(n_11362)
);

INVx1_ASAP7_75t_L g11363 ( 
.A(n_10900),
.Y(n_11363)
);

NAND2xp5_ASAP7_75t_L g11364 ( 
.A(n_11052),
.B(n_8364),
.Y(n_11364)
);

INVx1_ASAP7_75t_L g11365 ( 
.A(n_10912),
.Y(n_11365)
);

INVx2_ASAP7_75t_L g11366 ( 
.A(n_11049),
.Y(n_11366)
);

NOR2xp33_ASAP7_75t_L g11367 ( 
.A(n_11074),
.B(n_8366),
.Y(n_11367)
);

NOR2xp33_ASAP7_75t_L g11368 ( 
.A(n_10946),
.B(n_8366),
.Y(n_11368)
);

INVx1_ASAP7_75t_SL g11369 ( 
.A(n_11058),
.Y(n_11369)
);

NAND2xp5_ASAP7_75t_L g11370 ( 
.A(n_11053),
.B(n_8367),
.Y(n_11370)
);

NAND2xp5_ASAP7_75t_L g11371 ( 
.A(n_11057),
.B(n_8367),
.Y(n_11371)
);

HB1xp67_ASAP7_75t_L g11372 ( 
.A(n_11065),
.Y(n_11372)
);

INVx3_ASAP7_75t_L g11373 ( 
.A(n_10957),
.Y(n_11373)
);

AND2x2_ASAP7_75t_L g11374 ( 
.A(n_11062),
.B(n_8349),
.Y(n_11374)
);

INVx1_ASAP7_75t_L g11375 ( 
.A(n_10913),
.Y(n_11375)
);

INVx1_ASAP7_75t_L g11376 ( 
.A(n_10920),
.Y(n_11376)
);

NAND2xp5_ASAP7_75t_L g11377 ( 
.A(n_11034),
.B(n_8921),
.Y(n_11377)
);

INVx1_ASAP7_75t_L g11378 ( 
.A(n_10921),
.Y(n_11378)
);

AOI32xp33_ASAP7_75t_L g11379 ( 
.A1(n_10983),
.A2(n_8903),
.A3(n_8916),
.B1(n_8896),
.B2(n_8885),
.Y(n_11379)
);

NAND2xp33_ASAP7_75t_SL g11380 ( 
.A(n_10960),
.B(n_8377),
.Y(n_11380)
);

INVx1_ASAP7_75t_L g11381 ( 
.A(n_10926),
.Y(n_11381)
);

INVx3_ASAP7_75t_L g11382 ( 
.A(n_10970),
.Y(n_11382)
);

NAND2xp5_ASAP7_75t_L g11383 ( 
.A(n_11036),
.B(n_8921),
.Y(n_11383)
);

NAND2xp5_ASAP7_75t_L g11384 ( 
.A(n_10985),
.B(n_8921),
.Y(n_11384)
);

INVx1_ASAP7_75t_L g11385 ( 
.A(n_10938),
.Y(n_11385)
);

OR2x2_ASAP7_75t_L g11386 ( 
.A(n_10940),
.B(n_8462),
.Y(n_11386)
);

NAND2xp5_ASAP7_75t_L g11387 ( 
.A(n_11037),
.B(n_11085),
.Y(n_11387)
);

NAND2xp5_ASAP7_75t_L g11388 ( 
.A(n_10942),
.B(n_10978),
.Y(n_11388)
);

INVx1_ASAP7_75t_SL g11389 ( 
.A(n_11086),
.Y(n_11389)
);

AND2x2_ASAP7_75t_L g11390 ( 
.A(n_11003),
.B(n_8668),
.Y(n_11390)
);

NAND2xp5_ASAP7_75t_L g11391 ( 
.A(n_11106),
.B(n_11061),
.Y(n_11391)
);

OAI21xp5_ASAP7_75t_L g11392 ( 
.A1(n_11172),
.A2(n_10973),
.B(n_10969),
.Y(n_11392)
);

OR2x2_ASAP7_75t_L g11393 ( 
.A(n_11113),
.B(n_11011),
.Y(n_11393)
);

NAND2xp5_ASAP7_75t_SL g11394 ( 
.A(n_11144),
.B(n_11083),
.Y(n_11394)
);

HB1xp67_ASAP7_75t_L g11395 ( 
.A(n_11218),
.Y(n_11395)
);

OAI22xp33_ASAP7_75t_L g11396 ( 
.A1(n_11089),
.A2(n_11329),
.B1(n_11112),
.B2(n_11122),
.Y(n_11396)
);

INVxp33_ASAP7_75t_L g11397 ( 
.A(n_11100),
.Y(n_11397)
);

NAND2xp5_ASAP7_75t_L g11398 ( 
.A(n_11121),
.B(n_10997),
.Y(n_11398)
);

NAND2xp5_ASAP7_75t_L g11399 ( 
.A(n_11121),
.B(n_11038),
.Y(n_11399)
);

NAND2xp5_ASAP7_75t_L g11400 ( 
.A(n_11183),
.B(n_10948),
.Y(n_11400)
);

INVx1_ASAP7_75t_L g11401 ( 
.A(n_11105),
.Y(n_11401)
);

INVx1_ASAP7_75t_L g11402 ( 
.A(n_11115),
.Y(n_11402)
);

AND2x2_ASAP7_75t_L g11403 ( 
.A(n_11164),
.B(n_10954),
.Y(n_11403)
);

AOI21xp33_ASAP7_75t_SL g11404 ( 
.A1(n_11119),
.A2(n_11059),
.B(n_11042),
.Y(n_11404)
);

NAND2xp5_ASAP7_75t_L g11405 ( 
.A(n_11125),
.B(n_10949),
.Y(n_11405)
);

INVx2_ASAP7_75t_SL g11406 ( 
.A(n_11218),
.Y(n_11406)
);

INVx2_ASAP7_75t_SL g11407 ( 
.A(n_11127),
.Y(n_11407)
);

HB1xp67_ASAP7_75t_L g11408 ( 
.A(n_11270),
.Y(n_11408)
);

INVx1_ASAP7_75t_L g11409 ( 
.A(n_11270),
.Y(n_11409)
);

NOR2xp33_ASAP7_75t_L g11410 ( 
.A(n_11343),
.B(n_11035),
.Y(n_11410)
);

NOR2x1_ASAP7_75t_SL g11411 ( 
.A(n_11220),
.B(n_10955),
.Y(n_11411)
);

AND2x2_ASAP7_75t_L g11412 ( 
.A(n_11096),
.B(n_11023),
.Y(n_11412)
);

NAND2x1p5_ASAP7_75t_L g11413 ( 
.A(n_11285),
.B(n_11116),
.Y(n_11413)
);

INVxp67_ASAP7_75t_SL g11414 ( 
.A(n_11285),
.Y(n_11414)
);

NAND2xp5_ASAP7_75t_L g11415 ( 
.A(n_11097),
.B(n_10956),
.Y(n_11415)
);

OR2x2_ASAP7_75t_L g11416 ( 
.A(n_11191),
.B(n_10934),
.Y(n_11416)
);

INVx1_ASAP7_75t_L g11417 ( 
.A(n_11135),
.Y(n_11417)
);

INVx1_ASAP7_75t_L g11418 ( 
.A(n_11129),
.Y(n_11418)
);

INVx2_ASAP7_75t_SL g11419 ( 
.A(n_11127),
.Y(n_11419)
);

INVx2_ASAP7_75t_L g11420 ( 
.A(n_11116),
.Y(n_11420)
);

AND2x2_ASAP7_75t_L g11421 ( 
.A(n_11103),
.B(n_10958),
.Y(n_11421)
);

AND2x2_ASAP7_75t_L g11422 ( 
.A(n_11136),
.B(n_10959),
.Y(n_11422)
);

INVx1_ASAP7_75t_L g11423 ( 
.A(n_11098),
.Y(n_11423)
);

AND2x4_ASAP7_75t_L g11424 ( 
.A(n_11133),
.B(n_10961),
.Y(n_11424)
);

INVx2_ASAP7_75t_L g11425 ( 
.A(n_11128),
.Y(n_11425)
);

OR2x2_ASAP7_75t_L g11426 ( 
.A(n_11092),
.B(n_11072),
.Y(n_11426)
);

OR2x2_ASAP7_75t_L g11427 ( 
.A(n_11248),
.B(n_10998),
.Y(n_11427)
);

INVx2_ASAP7_75t_L g11428 ( 
.A(n_11128),
.Y(n_11428)
);

INVxp67_ASAP7_75t_SL g11429 ( 
.A(n_11140),
.Y(n_11429)
);

OR2x2_ASAP7_75t_L g11430 ( 
.A(n_11180),
.B(n_10999),
.Y(n_11430)
);

INVx1_ASAP7_75t_L g11431 ( 
.A(n_11094),
.Y(n_11431)
);

INVx1_ASAP7_75t_SL g11432 ( 
.A(n_11163),
.Y(n_11432)
);

INVx2_ASAP7_75t_L g11433 ( 
.A(n_11140),
.Y(n_11433)
);

NOR2xp33_ASAP7_75t_L g11434 ( 
.A(n_11167),
.B(n_10964),
.Y(n_11434)
);

INVx1_ASAP7_75t_L g11435 ( 
.A(n_11102),
.Y(n_11435)
);

INVxp67_ASAP7_75t_L g11436 ( 
.A(n_11316),
.Y(n_11436)
);

INVx1_ASAP7_75t_L g11437 ( 
.A(n_11093),
.Y(n_11437)
);

OR2x2_ASAP7_75t_L g11438 ( 
.A(n_11088),
.B(n_11001),
.Y(n_11438)
);

NOR2xp33_ASAP7_75t_L g11439 ( 
.A(n_11353),
.B(n_11160),
.Y(n_11439)
);

OR2x2_ASAP7_75t_L g11440 ( 
.A(n_11091),
.B(n_11131),
.Y(n_11440)
);

AND2x4_ASAP7_75t_SL g11441 ( 
.A(n_11145),
.B(n_10819),
.Y(n_11441)
);

INVx1_ASAP7_75t_L g11442 ( 
.A(n_11217),
.Y(n_11442)
);

AND2x2_ASAP7_75t_L g11443 ( 
.A(n_11146),
.B(n_10965),
.Y(n_11443)
);

NAND2xp5_ASAP7_75t_L g11444 ( 
.A(n_11133),
.B(n_10995),
.Y(n_11444)
);

AND2x4_ASAP7_75t_L g11445 ( 
.A(n_11208),
.B(n_11000),
.Y(n_11445)
);

AND2x2_ASAP7_75t_L g11446 ( 
.A(n_11109),
.B(n_11002),
.Y(n_11446)
);

INVxp67_ASAP7_75t_SL g11447 ( 
.A(n_11373),
.Y(n_11447)
);

NAND2xp5_ASAP7_75t_L g11448 ( 
.A(n_11221),
.B(n_11005),
.Y(n_11448)
);

NAND2xp5_ASAP7_75t_L g11449 ( 
.A(n_11087),
.B(n_11009),
.Y(n_11449)
);

INVx1_ASAP7_75t_L g11450 ( 
.A(n_11178),
.Y(n_11450)
);

NAND2xp5_ASAP7_75t_L g11451 ( 
.A(n_11153),
.B(n_10820),
.Y(n_11451)
);

OR2x2_ASAP7_75t_L g11452 ( 
.A(n_11090),
.B(n_11095),
.Y(n_11452)
);

INVx1_ASAP7_75t_L g11453 ( 
.A(n_11212),
.Y(n_11453)
);

OAI21xp33_ASAP7_75t_L g11454 ( 
.A1(n_11132),
.A2(n_10828),
.B(n_10825),
.Y(n_11454)
);

INVx2_ASAP7_75t_L g11455 ( 
.A(n_11373),
.Y(n_11455)
);

INVx1_ASAP7_75t_L g11456 ( 
.A(n_11215),
.Y(n_11456)
);

AOI21xp33_ASAP7_75t_L g11457 ( 
.A1(n_11294),
.A2(n_10834),
.B(n_10832),
.Y(n_11457)
);

NAND2xp5_ASAP7_75t_L g11458 ( 
.A(n_11143),
.B(n_10835),
.Y(n_11458)
);

AND2x2_ASAP7_75t_L g11459 ( 
.A(n_11108),
.B(n_10836),
.Y(n_11459)
);

OR2x2_ASAP7_75t_L g11460 ( 
.A(n_11101),
.B(n_10975),
.Y(n_11460)
);

AND2x4_ASAP7_75t_L g11461 ( 
.A(n_11382),
.B(n_10976),
.Y(n_11461)
);

NAND2xp5_ASAP7_75t_L g11462 ( 
.A(n_11118),
.B(n_10981),
.Y(n_11462)
);

NAND2xp5_ASAP7_75t_L g11463 ( 
.A(n_11120),
.B(n_10992),
.Y(n_11463)
);

NOR2x1_ASAP7_75t_L g11464 ( 
.A(n_11094),
.B(n_8377),
.Y(n_11464)
);

INVx2_ASAP7_75t_L g11465 ( 
.A(n_11382),
.Y(n_11465)
);

INVx1_ASAP7_75t_L g11466 ( 
.A(n_11223),
.Y(n_11466)
);

INVx1_ASAP7_75t_L g11467 ( 
.A(n_11173),
.Y(n_11467)
);

INVx2_ASAP7_75t_L g11468 ( 
.A(n_11220),
.Y(n_11468)
);

INVx2_ASAP7_75t_L g11469 ( 
.A(n_11202),
.Y(n_11469)
);

AND2x2_ASAP7_75t_L g11470 ( 
.A(n_11110),
.B(n_8668),
.Y(n_11470)
);

INVx1_ASAP7_75t_L g11471 ( 
.A(n_11202),
.Y(n_11471)
);

OR2x2_ASAP7_75t_L g11472 ( 
.A(n_11185),
.B(n_8611),
.Y(n_11472)
);

OR2x2_ASAP7_75t_L g11473 ( 
.A(n_11147),
.B(n_9399),
.Y(n_11473)
);

NAND2xp5_ASAP7_75t_L g11474 ( 
.A(n_11181),
.B(n_9399),
.Y(n_11474)
);

AND2x2_ASAP7_75t_L g11475 ( 
.A(n_11117),
.B(n_8377),
.Y(n_11475)
);

AND2x2_ASAP7_75t_L g11476 ( 
.A(n_11099),
.B(n_9399),
.Y(n_11476)
);

AOI21xp33_ASAP7_75t_L g11477 ( 
.A1(n_11284),
.A2(n_8623),
.B(n_8615),
.Y(n_11477)
);

NAND2xp5_ASAP7_75t_L g11478 ( 
.A(n_11181),
.B(n_9399),
.Y(n_11478)
);

AND2x2_ASAP7_75t_L g11479 ( 
.A(n_11111),
.B(n_8615),
.Y(n_11479)
);

NAND2xp5_ASAP7_75t_L g11480 ( 
.A(n_11177),
.B(n_8842),
.Y(n_11480)
);

INVx1_ASAP7_75t_L g11481 ( 
.A(n_11293),
.Y(n_11481)
);

INVx1_ASAP7_75t_L g11482 ( 
.A(n_11304),
.Y(n_11482)
);

INVx1_ASAP7_75t_L g11483 ( 
.A(n_11239),
.Y(n_11483)
);

OR2x2_ASAP7_75t_L g11484 ( 
.A(n_11156),
.B(n_8676),
.Y(n_11484)
);

INVxp67_ASAP7_75t_L g11485 ( 
.A(n_11309),
.Y(n_11485)
);

NAND2xp5_ASAP7_75t_L g11486 ( 
.A(n_11310),
.B(n_8842),
.Y(n_11486)
);

NOR5xp2_ASAP7_75t_L g11487 ( 
.A(n_11210),
.B(n_8769),
.C(n_8804),
.D(n_8808),
.E(n_8802),
.Y(n_11487)
);

AND2x4_ASAP7_75t_L g11488 ( 
.A(n_11182),
.B(n_8817),
.Y(n_11488)
);

INVx1_ASAP7_75t_L g11489 ( 
.A(n_11188),
.Y(n_11489)
);

INVx1_ASAP7_75t_L g11490 ( 
.A(n_11169),
.Y(n_11490)
);

OR2x2_ASAP7_75t_L g11491 ( 
.A(n_11174),
.B(n_8689),
.Y(n_11491)
);

INVx3_ASAP7_75t_L g11492 ( 
.A(n_11225),
.Y(n_11492)
);

OAI32xp33_ASAP7_75t_L g11493 ( 
.A1(n_11340),
.A2(n_8885),
.A3(n_8882),
.B1(n_8846),
.B2(n_8503),
.Y(n_11493)
);

INVxp67_ASAP7_75t_L g11494 ( 
.A(n_11315),
.Y(n_11494)
);

INVx1_ASAP7_75t_L g11495 ( 
.A(n_11271),
.Y(n_11495)
);

INVx1_ASAP7_75t_L g11496 ( 
.A(n_11114),
.Y(n_11496)
);

NOR2xp33_ASAP7_75t_L g11497 ( 
.A(n_11348),
.B(n_11357),
.Y(n_11497)
);

NAND2xp5_ASAP7_75t_L g11498 ( 
.A(n_11225),
.B(n_8842),
.Y(n_11498)
);

INVx1_ASAP7_75t_L g11499 ( 
.A(n_11134),
.Y(n_11499)
);

HB1xp67_ASAP7_75t_L g11500 ( 
.A(n_11298),
.Y(n_11500)
);

NAND2xp5_ASAP7_75t_L g11501 ( 
.A(n_11104),
.B(n_8478),
.Y(n_11501)
);

NAND2xp5_ASAP7_75t_L g11502 ( 
.A(n_11148),
.B(n_8478),
.Y(n_11502)
);

NAND2xp5_ASAP7_75t_SL g11503 ( 
.A(n_11286),
.B(n_8623),
.Y(n_11503)
);

NOR2xp33_ASAP7_75t_L g11504 ( 
.A(n_11150),
.B(n_8626),
.Y(n_11504)
);

AND2x2_ASAP7_75t_L g11505 ( 
.A(n_11107),
.B(n_8626),
.Y(n_11505)
);

INVx2_ASAP7_75t_L g11506 ( 
.A(n_11152),
.Y(n_11506)
);

INVx1_ASAP7_75t_L g11507 ( 
.A(n_11170),
.Y(n_11507)
);

OAI21xp33_ASAP7_75t_L g11508 ( 
.A1(n_11187),
.A2(n_8831),
.B(n_8817),
.Y(n_11508)
);

NAND2xp33_ASAP7_75t_SL g11509 ( 
.A(n_11346),
.B(n_11345),
.Y(n_11509)
);

INVx2_ASAP7_75t_SL g11510 ( 
.A(n_11299),
.Y(n_11510)
);

BUFx2_ASAP7_75t_L g11511 ( 
.A(n_11124),
.Y(n_11511)
);

OR2x2_ASAP7_75t_SL g11512 ( 
.A(n_11189),
.B(n_8820),
.Y(n_11512)
);

NAND2xp5_ASAP7_75t_L g11513 ( 
.A(n_11123),
.B(n_8856),
.Y(n_11513)
);

BUFx2_ASAP7_75t_L g11514 ( 
.A(n_11241),
.Y(n_11514)
);

NAND2xp5_ASAP7_75t_L g11515 ( 
.A(n_11151),
.B(n_8856),
.Y(n_11515)
);

OAI21xp33_ASAP7_75t_SL g11516 ( 
.A1(n_11237),
.A2(n_8372),
.B(n_8882),
.Y(n_11516)
);

INVx1_ASAP7_75t_L g11517 ( 
.A(n_11157),
.Y(n_11517)
);

OAI21xp5_ASAP7_75t_L g11518 ( 
.A1(n_11130),
.A2(n_8826),
.B(n_8777),
.Y(n_11518)
);

OR2x2_ASAP7_75t_L g11519 ( 
.A(n_11141),
.B(n_8703),
.Y(n_11519)
);

NAND2xp5_ASAP7_75t_L g11520 ( 
.A(n_11158),
.B(n_8856),
.Y(n_11520)
);

INVx1_ASAP7_75t_L g11521 ( 
.A(n_11159),
.Y(n_11521)
);

AND2x2_ASAP7_75t_L g11522 ( 
.A(n_11162),
.B(n_8640),
.Y(n_11522)
);

BUFx2_ASAP7_75t_L g11523 ( 
.A(n_11241),
.Y(n_11523)
);

HB1xp67_ASAP7_75t_L g11524 ( 
.A(n_11356),
.Y(n_11524)
);

INVxp67_ASAP7_75t_L g11525 ( 
.A(n_11312),
.Y(n_11525)
);

INVx1_ASAP7_75t_L g11526 ( 
.A(n_11161),
.Y(n_11526)
);

AND2x2_ASAP7_75t_L g11527 ( 
.A(n_11257),
.B(n_8640),
.Y(n_11527)
);

AND2x2_ASAP7_75t_L g11528 ( 
.A(n_11272),
.B(n_8645),
.Y(n_11528)
);

INVx2_ASAP7_75t_L g11529 ( 
.A(n_11266),
.Y(n_11529)
);

INVx1_ASAP7_75t_L g11530 ( 
.A(n_11190),
.Y(n_11530)
);

NOR2xp33_ASAP7_75t_L g11531 ( 
.A(n_11369),
.B(n_8645),
.Y(n_11531)
);

AND2x2_ASAP7_75t_L g11532 ( 
.A(n_11213),
.B(n_8646),
.Y(n_11532)
);

INVx1_ASAP7_75t_L g11533 ( 
.A(n_11171),
.Y(n_11533)
);

NAND2xp5_ASAP7_75t_L g11534 ( 
.A(n_11165),
.B(n_8646),
.Y(n_11534)
);

INVx1_ASAP7_75t_L g11535 ( 
.A(n_11192),
.Y(n_11535)
);

AND2x2_ASAP7_75t_L g11536 ( 
.A(n_11227),
.B(n_8655),
.Y(n_11536)
);

INVx1_ASAP7_75t_L g11537 ( 
.A(n_11214),
.Y(n_11537)
);

NOR3xp33_ASAP7_75t_L g11538 ( 
.A(n_11358),
.B(n_8655),
.C(n_8777),
.Y(n_11538)
);

INVx2_ASAP7_75t_SL g11539 ( 
.A(n_11266),
.Y(n_11539)
);

OR2x2_ASAP7_75t_L g11540 ( 
.A(n_11166),
.B(n_8737),
.Y(n_11540)
);

INVx1_ASAP7_75t_L g11541 ( 
.A(n_11234),
.Y(n_11541)
);

INVx1_ASAP7_75t_L g11542 ( 
.A(n_11323),
.Y(n_11542)
);

HB1xp67_ASAP7_75t_L g11543 ( 
.A(n_11179),
.Y(n_11543)
);

INVxp67_ASAP7_75t_L g11544 ( 
.A(n_11367),
.Y(n_11544)
);

INVx1_ASAP7_75t_L g11545 ( 
.A(n_11326),
.Y(n_11545)
);

AND2x2_ASAP7_75t_L g11546 ( 
.A(n_11193),
.B(n_8820),
.Y(n_11546)
);

INVx1_ASAP7_75t_L g11547 ( 
.A(n_11137),
.Y(n_11547)
);

INVx1_ASAP7_75t_L g11548 ( 
.A(n_11219),
.Y(n_11548)
);

INVx1_ASAP7_75t_L g11549 ( 
.A(n_11222),
.Y(n_11549)
);

NOR2xp33_ASAP7_75t_SL g11550 ( 
.A(n_11389),
.B(n_8039),
.Y(n_11550)
);

OR2x2_ASAP7_75t_L g11551 ( 
.A(n_11168),
.B(n_11216),
.Y(n_11551)
);

INVx1_ASAP7_75t_L g11552 ( 
.A(n_11258),
.Y(n_11552)
);

INVx1_ASAP7_75t_SL g11553 ( 
.A(n_11332),
.Y(n_11553)
);

NOR2xp33_ASAP7_75t_L g11554 ( 
.A(n_11318),
.B(n_7178),
.Y(n_11554)
);

OR2x2_ASAP7_75t_L g11555 ( 
.A(n_11352),
.B(n_8472),
.Y(n_11555)
);

INVx2_ASAP7_75t_SL g11556 ( 
.A(n_11351),
.Y(n_11556)
);

INVx1_ASAP7_75t_L g11557 ( 
.A(n_11195),
.Y(n_11557)
);

INVx3_ASAP7_75t_L g11558 ( 
.A(n_11351),
.Y(n_11558)
);

INVx2_ASAP7_75t_SL g11559 ( 
.A(n_11184),
.Y(n_11559)
);

HB1xp67_ASAP7_75t_L g11560 ( 
.A(n_11186),
.Y(n_11560)
);

NAND2xp5_ASAP7_75t_L g11561 ( 
.A(n_11194),
.B(n_8571),
.Y(n_11561)
);

AND2x2_ASAP7_75t_L g11562 ( 
.A(n_11207),
.B(n_8820),
.Y(n_11562)
);

INVxp67_ASAP7_75t_L g11563 ( 
.A(n_11368),
.Y(n_11563)
);

AND2x2_ASAP7_75t_L g11564 ( 
.A(n_11207),
.B(n_8827),
.Y(n_11564)
);

OR2x2_ASAP7_75t_L g11565 ( 
.A(n_11126),
.B(n_8827),
.Y(n_11565)
);

OR2x2_ASAP7_75t_L g11566 ( 
.A(n_11347),
.B(n_8827),
.Y(n_11566)
);

INVx1_ASAP7_75t_L g11567 ( 
.A(n_11196),
.Y(n_11567)
);

INVx2_ASAP7_75t_SL g11568 ( 
.A(n_11283),
.Y(n_11568)
);

INVx1_ASAP7_75t_L g11569 ( 
.A(n_11197),
.Y(n_11569)
);

NAND2xp5_ASAP7_75t_L g11570 ( 
.A(n_11149),
.B(n_8571),
.Y(n_11570)
);

INVx1_ASAP7_75t_L g11571 ( 
.A(n_11199),
.Y(n_11571)
);

NAND2xp5_ASAP7_75t_L g11572 ( 
.A(n_11138),
.B(n_8571),
.Y(n_11572)
);

NAND2xp5_ASAP7_75t_L g11573 ( 
.A(n_11142),
.B(n_8850),
.Y(n_11573)
);

INVx2_ASAP7_75t_L g11574 ( 
.A(n_11311),
.Y(n_11574)
);

INVx1_ASAP7_75t_L g11575 ( 
.A(n_11203),
.Y(n_11575)
);

AND2x2_ASAP7_75t_L g11576 ( 
.A(n_11242),
.B(n_8841),
.Y(n_11576)
);

INVxp67_ASAP7_75t_L g11577 ( 
.A(n_11273),
.Y(n_11577)
);

AND2x4_ASAP7_75t_L g11578 ( 
.A(n_11233),
.B(n_8783),
.Y(n_11578)
);

NAND3xp33_ASAP7_75t_L g11579 ( 
.A(n_11327),
.B(n_8841),
.C(n_8263),
.Y(n_11579)
);

INVx2_ASAP7_75t_L g11580 ( 
.A(n_11319),
.Y(n_11580)
);

AND2x2_ASAP7_75t_L g11581 ( 
.A(n_11231),
.B(n_8841),
.Y(n_11581)
);

INVxp67_ASAP7_75t_L g11582 ( 
.A(n_11201),
.Y(n_11582)
);

OR2x2_ASAP7_75t_L g11583 ( 
.A(n_11198),
.B(n_8562),
.Y(n_11583)
);

NAND2xp5_ASAP7_75t_L g11584 ( 
.A(n_11341),
.B(n_8850),
.Y(n_11584)
);

NAND3xp33_ASAP7_75t_SL g11585 ( 
.A(n_11387),
.B(n_11282),
.C(n_11301),
.Y(n_11585)
);

NOR2xp33_ASAP7_75t_L g11586 ( 
.A(n_11243),
.B(n_11366),
.Y(n_11586)
);

INVx1_ASAP7_75t_L g11587 ( 
.A(n_11204),
.Y(n_11587)
);

INVx2_ASAP7_75t_L g11588 ( 
.A(n_11322),
.Y(n_11588)
);

NAND2xp5_ASAP7_75t_L g11589 ( 
.A(n_11306),
.B(n_8850),
.Y(n_11589)
);

OAI211xp5_ASAP7_75t_L g11590 ( 
.A1(n_11236),
.A2(n_11155),
.B(n_11154),
.C(n_11139),
.Y(n_11590)
);

INVx1_ASAP7_75t_L g11591 ( 
.A(n_11205),
.Y(n_11591)
);

INVx1_ASAP7_75t_L g11592 ( 
.A(n_11206),
.Y(n_11592)
);

AND2x2_ASAP7_75t_L g11593 ( 
.A(n_11263),
.B(n_8783),
.Y(n_11593)
);

AOI22xp5_ASAP7_75t_L g11594 ( 
.A1(n_11291),
.A2(n_8448),
.B1(n_8495),
.B2(n_8239),
.Y(n_11594)
);

NAND2xp5_ASAP7_75t_L g11595 ( 
.A(n_11277),
.B(n_8304),
.Y(n_11595)
);

INVx1_ASAP7_75t_L g11596 ( 
.A(n_11209),
.Y(n_11596)
);

HB1xp67_ASAP7_75t_L g11597 ( 
.A(n_11374),
.Y(n_11597)
);

INVx2_ASAP7_75t_L g11598 ( 
.A(n_11274),
.Y(n_11598)
);

INVx1_ASAP7_75t_L g11599 ( 
.A(n_11211),
.Y(n_11599)
);

INVx1_ASAP7_75t_L g11600 ( 
.A(n_11330),
.Y(n_11600)
);

NAND4xp25_ASAP7_75t_L g11601 ( 
.A(n_11175),
.B(n_7885),
.C(n_7893),
.D(n_7884),
.Y(n_11601)
);

INVx1_ASAP7_75t_L g11602 ( 
.A(n_11176),
.Y(n_11602)
);

INVx2_ASAP7_75t_L g11603 ( 
.A(n_11276),
.Y(n_11603)
);

INVx1_ASAP7_75t_L g11604 ( 
.A(n_11200),
.Y(n_11604)
);

AND2x2_ASAP7_75t_L g11605 ( 
.A(n_11296),
.B(n_8388),
.Y(n_11605)
);

INVx1_ASAP7_75t_L g11606 ( 
.A(n_11228),
.Y(n_11606)
);

INVx2_ASAP7_75t_L g11607 ( 
.A(n_11278),
.Y(n_11607)
);

AND2x2_ASAP7_75t_L g11608 ( 
.A(n_11240),
.B(n_8388),
.Y(n_11608)
);

INVx1_ASAP7_75t_L g11609 ( 
.A(n_11228),
.Y(n_11609)
);

HB1xp67_ASAP7_75t_L g11610 ( 
.A(n_11355),
.Y(n_11610)
);

AND2x2_ASAP7_75t_L g11611 ( 
.A(n_11342),
.B(n_8388),
.Y(n_11611)
);

INVx1_ASAP7_75t_L g11612 ( 
.A(n_11235),
.Y(n_11612)
);

HB1xp67_ASAP7_75t_L g11613 ( 
.A(n_11336),
.Y(n_11613)
);

NAND2xp5_ASAP7_75t_L g11614 ( 
.A(n_11300),
.B(n_8304),
.Y(n_11614)
);

OR2x2_ASAP7_75t_L g11615 ( 
.A(n_11364),
.B(n_8562),
.Y(n_11615)
);

INVxp67_ASAP7_75t_L g11616 ( 
.A(n_11344),
.Y(n_11616)
);

INVx1_ASAP7_75t_L g11617 ( 
.A(n_11235),
.Y(n_11617)
);

INVx1_ASAP7_75t_L g11618 ( 
.A(n_11238),
.Y(n_11618)
);

INVx2_ASAP7_75t_L g11619 ( 
.A(n_11226),
.Y(n_11619)
);

AND2x2_ASAP7_75t_L g11620 ( 
.A(n_11308),
.B(n_11232),
.Y(n_11620)
);

INVx1_ASAP7_75t_L g11621 ( 
.A(n_11238),
.Y(n_11621)
);

HB1xp67_ASAP7_75t_L g11622 ( 
.A(n_11338),
.Y(n_11622)
);

INVx2_ASAP7_75t_L g11623 ( 
.A(n_11230),
.Y(n_11623)
);

INVx2_ASAP7_75t_L g11624 ( 
.A(n_11325),
.Y(n_11624)
);

INVx1_ASAP7_75t_L g11625 ( 
.A(n_11244),
.Y(n_11625)
);

AND2x2_ASAP7_75t_L g11626 ( 
.A(n_11245),
.B(n_8259),
.Y(n_11626)
);

AND2x4_ASAP7_75t_L g11627 ( 
.A(n_11354),
.B(n_8833),
.Y(n_11627)
);

OR2x2_ASAP7_75t_L g11628 ( 
.A(n_11370),
.B(n_8562),
.Y(n_11628)
);

NAND2xp5_ASAP7_75t_L g11629 ( 
.A(n_11390),
.B(n_8868),
.Y(n_11629)
);

INVxp67_ASAP7_75t_SL g11630 ( 
.A(n_11384),
.Y(n_11630)
);

OAI21xp33_ASAP7_75t_L g11631 ( 
.A1(n_11337),
.A2(n_8839),
.B(n_8838),
.Y(n_11631)
);

OR2x2_ASAP7_75t_L g11632 ( 
.A(n_11371),
.B(n_8570),
.Y(n_11632)
);

INVx1_ASAP7_75t_L g11633 ( 
.A(n_11244),
.Y(n_11633)
);

CKINVDCx16_ASAP7_75t_R g11634 ( 
.A(n_11267),
.Y(n_11634)
);

INVx1_ASAP7_75t_L g11635 ( 
.A(n_11224),
.Y(n_11635)
);

NAND3xp33_ASAP7_75t_L g11636 ( 
.A(n_11380),
.B(n_8257),
.C(n_8354),
.Y(n_11636)
);

INVx2_ASAP7_75t_L g11637 ( 
.A(n_11328),
.Y(n_11637)
);

BUFx2_ASAP7_75t_L g11638 ( 
.A(n_11360),
.Y(n_11638)
);

OR2x2_ASAP7_75t_L g11639 ( 
.A(n_11305),
.B(n_8570),
.Y(n_11639)
);

NAND2xp5_ASAP7_75t_L g11640 ( 
.A(n_11361),
.B(n_8868),
.Y(n_11640)
);

AND2x2_ASAP7_75t_L g11641 ( 
.A(n_11292),
.B(n_8868),
.Y(n_11641)
);

OR2x2_ASAP7_75t_L g11642 ( 
.A(n_11339),
.B(n_8570),
.Y(n_11642)
);

NOR2xp67_ASAP7_75t_L g11643 ( 
.A(n_11229),
.B(n_8334),
.Y(n_11643)
);

OAI22xp5_ASAP7_75t_L g11644 ( 
.A1(n_11314),
.A2(n_8278),
.B1(n_7962),
.B2(n_7944),
.Y(n_11644)
);

INVx2_ASAP7_75t_L g11645 ( 
.A(n_11331),
.Y(n_11645)
);

AND2x2_ASAP7_75t_L g11646 ( 
.A(n_11407),
.B(n_11302),
.Y(n_11646)
);

INVx1_ASAP7_75t_SL g11647 ( 
.A(n_11514),
.Y(n_11647)
);

NAND2xp5_ASAP7_75t_L g11648 ( 
.A(n_11419),
.B(n_11359),
.Y(n_11648)
);

INVx1_ASAP7_75t_L g11649 ( 
.A(n_11395),
.Y(n_11649)
);

INVx2_ASAP7_75t_L g11650 ( 
.A(n_11492),
.Y(n_11650)
);

INVx2_ASAP7_75t_L g11651 ( 
.A(n_11492),
.Y(n_11651)
);

OR2x2_ASAP7_75t_L g11652 ( 
.A(n_11634),
.B(n_11317),
.Y(n_11652)
);

AND2x2_ASAP7_75t_L g11653 ( 
.A(n_11403),
.B(n_11303),
.Y(n_11653)
);

OA21x2_ASAP7_75t_L g11654 ( 
.A1(n_11523),
.A2(n_11334),
.B(n_11333),
.Y(n_11654)
);

INVx1_ASAP7_75t_SL g11655 ( 
.A(n_11509),
.Y(n_11655)
);

INVx1_ASAP7_75t_L g11656 ( 
.A(n_11411),
.Y(n_11656)
);

OR2x2_ASAP7_75t_L g11657 ( 
.A(n_11539),
.B(n_11447),
.Y(n_11657)
);

INVx1_ASAP7_75t_L g11658 ( 
.A(n_11411),
.Y(n_11658)
);

OAI221xp5_ASAP7_75t_L g11659 ( 
.A1(n_11550),
.A2(n_11379),
.B1(n_11268),
.B2(n_11252),
.C(n_11251),
.Y(n_11659)
);

CKINVDCx16_ASAP7_75t_R g11660 ( 
.A(n_11585),
.Y(n_11660)
);

AND2x2_ASAP7_75t_L g11661 ( 
.A(n_11432),
.B(n_11246),
.Y(n_11661)
);

OAI32xp33_ASAP7_75t_L g11662 ( 
.A1(n_11516),
.A2(n_11269),
.A3(n_11383),
.B1(n_11262),
.B2(n_11264),
.Y(n_11662)
);

INVx1_ASAP7_75t_L g11663 ( 
.A(n_11408),
.Y(n_11663)
);

INVx1_ASAP7_75t_L g11664 ( 
.A(n_11414),
.Y(n_11664)
);

NAND2x1p5_ASAP7_75t_L g11665 ( 
.A(n_11553),
.B(n_11558),
.Y(n_11665)
);

AND2x2_ASAP7_75t_L g11666 ( 
.A(n_11446),
.B(n_11247),
.Y(n_11666)
);

INVx2_ASAP7_75t_L g11667 ( 
.A(n_11406),
.Y(n_11667)
);

INVx1_ASAP7_75t_L g11668 ( 
.A(n_11413),
.Y(n_11668)
);

INVx1_ASAP7_75t_L g11669 ( 
.A(n_11429),
.Y(n_11669)
);

NAND2xp5_ASAP7_75t_L g11670 ( 
.A(n_11424),
.B(n_11249),
.Y(n_11670)
);

OR2x2_ASAP7_75t_L g11671 ( 
.A(n_11529),
.B(n_11324),
.Y(n_11671)
);

INVx2_ASAP7_75t_L g11672 ( 
.A(n_11424),
.Y(n_11672)
);

AOI21xp33_ASAP7_75t_L g11673 ( 
.A1(n_11397),
.A2(n_11253),
.B(n_11372),
.Y(n_11673)
);

INVx1_ASAP7_75t_L g11674 ( 
.A(n_11471),
.Y(n_11674)
);

INVxp67_ASAP7_75t_SL g11675 ( 
.A(n_11487),
.Y(n_11675)
);

NAND2xp5_ASAP7_75t_L g11676 ( 
.A(n_11469),
.B(n_11250),
.Y(n_11676)
);

OR2x2_ASAP7_75t_L g11677 ( 
.A(n_11455),
.B(n_11261),
.Y(n_11677)
);

NAND2x1_ASAP7_75t_L g11678 ( 
.A(n_11461),
.B(n_11335),
.Y(n_11678)
);

INVx1_ASAP7_75t_L g11679 ( 
.A(n_11471),
.Y(n_11679)
);

AND2x2_ASAP7_75t_L g11680 ( 
.A(n_11412),
.B(n_11307),
.Y(n_11680)
);

INVx2_ASAP7_75t_L g11681 ( 
.A(n_11461),
.Y(n_11681)
);

O2A1O1Ixp33_ASAP7_75t_SL g11682 ( 
.A1(n_11474),
.A2(n_11295),
.B(n_11297),
.C(n_11287),
.Y(n_11682)
);

AND2x4_ASAP7_75t_L g11683 ( 
.A(n_11465),
.B(n_11350),
.Y(n_11683)
);

AND2x2_ASAP7_75t_L g11684 ( 
.A(n_11459),
.B(n_11313),
.Y(n_11684)
);

OAI22xp33_ASAP7_75t_L g11685 ( 
.A1(n_11594),
.A2(n_11349),
.B1(n_11388),
.B2(n_11386),
.Y(n_11685)
);

NAND2x1_ASAP7_75t_L g11686 ( 
.A(n_11464),
.B(n_11362),
.Y(n_11686)
);

INVx2_ASAP7_75t_L g11687 ( 
.A(n_11512),
.Y(n_11687)
);

NOR4xp25_ASAP7_75t_L g11688 ( 
.A(n_11396),
.B(n_11281),
.C(n_11365),
.D(n_11363),
.Y(n_11688)
);

INVx1_ASAP7_75t_L g11689 ( 
.A(n_11500),
.Y(n_11689)
);

AOI32xp33_ASAP7_75t_L g11690 ( 
.A1(n_11439),
.A2(n_11281),
.A3(n_11385),
.B1(n_11376),
.B2(n_11378),
.Y(n_11690)
);

NAND2xp5_ASAP7_75t_L g11691 ( 
.A(n_11409),
.B(n_11375),
.Y(n_11691)
);

AOI21xp5_ASAP7_75t_L g11692 ( 
.A1(n_11394),
.A2(n_11377),
.B(n_11376),
.Y(n_11692)
);

INVx1_ASAP7_75t_L g11693 ( 
.A(n_11421),
.Y(n_11693)
);

AND2x2_ASAP7_75t_L g11694 ( 
.A(n_11496),
.B(n_11375),
.Y(n_11694)
);

OAI31xp33_ASAP7_75t_L g11695 ( 
.A1(n_11579),
.A2(n_11381),
.A3(n_11378),
.B(n_11288),
.Y(n_11695)
);

AND2x2_ASAP7_75t_L g11696 ( 
.A(n_11423),
.B(n_11381),
.Y(n_11696)
);

AOI21xp5_ASAP7_75t_L g11697 ( 
.A1(n_11398),
.A2(n_11255),
.B(n_11254),
.Y(n_11697)
);

NOR2xp67_ASAP7_75t_L g11698 ( 
.A(n_11404),
.B(n_11256),
.Y(n_11698)
);

INVx1_ASAP7_75t_L g11699 ( 
.A(n_11422),
.Y(n_11699)
);

INVx1_ASAP7_75t_L g11700 ( 
.A(n_11444),
.Y(n_11700)
);

INVx1_ASAP7_75t_L g11701 ( 
.A(n_11443),
.Y(n_11701)
);

INVx1_ASAP7_75t_L g11702 ( 
.A(n_11478),
.Y(n_11702)
);

AND2x2_ASAP7_75t_L g11703 ( 
.A(n_11437),
.B(n_11259),
.Y(n_11703)
);

OR2x2_ASAP7_75t_L g11704 ( 
.A(n_11510),
.B(n_11260),
.Y(n_11704)
);

INVxp67_ASAP7_75t_L g11705 ( 
.A(n_11475),
.Y(n_11705)
);

NAND2xp5_ASAP7_75t_L g11706 ( 
.A(n_11558),
.B(n_11265),
.Y(n_11706)
);

INVx1_ASAP7_75t_L g11707 ( 
.A(n_11441),
.Y(n_11707)
);

INVx1_ASAP7_75t_SL g11708 ( 
.A(n_11427),
.Y(n_11708)
);

INVx1_ASAP7_75t_SL g11709 ( 
.A(n_11393),
.Y(n_11709)
);

INVx3_ASAP7_75t_L g11710 ( 
.A(n_11445),
.Y(n_11710)
);

INVx1_ASAP7_75t_L g11711 ( 
.A(n_11543),
.Y(n_11711)
);

INVx1_ASAP7_75t_L g11712 ( 
.A(n_11560),
.Y(n_11712)
);

INVx2_ASAP7_75t_L g11713 ( 
.A(n_11425),
.Y(n_11713)
);

OR2x2_ASAP7_75t_L g11714 ( 
.A(n_11401),
.B(n_11402),
.Y(n_11714)
);

AND2x2_ASAP7_75t_L g11715 ( 
.A(n_11499),
.B(n_11275),
.Y(n_11715)
);

NOR2x2_ASAP7_75t_L g11716 ( 
.A(n_11588),
.B(n_11279),
.Y(n_11716)
);

OR2x2_ASAP7_75t_L g11717 ( 
.A(n_11428),
.B(n_11280),
.Y(n_11717)
);

INVx1_ASAP7_75t_L g11718 ( 
.A(n_11473),
.Y(n_11718)
);

INVx2_ASAP7_75t_SL g11719 ( 
.A(n_11445),
.Y(n_11719)
);

AND2x2_ASAP7_75t_SL g11720 ( 
.A(n_11452),
.B(n_11289),
.Y(n_11720)
);

AND2x4_ASAP7_75t_L g11721 ( 
.A(n_11556),
.B(n_11290),
.Y(n_11721)
);

AND2x2_ASAP7_75t_L g11722 ( 
.A(n_11495),
.B(n_11320),
.Y(n_11722)
);

NOR2xp33_ASAP7_75t_L g11723 ( 
.A(n_11494),
.B(n_11321),
.Y(n_11723)
);

INVx2_ASAP7_75t_SL g11724 ( 
.A(n_11433),
.Y(n_11724)
);

BUFx2_ASAP7_75t_L g11725 ( 
.A(n_11476),
.Y(n_11725)
);

INVx1_ASAP7_75t_L g11726 ( 
.A(n_11610),
.Y(n_11726)
);

INVx1_ASAP7_75t_L g11727 ( 
.A(n_11613),
.Y(n_11727)
);

AND2x2_ASAP7_75t_L g11728 ( 
.A(n_11466),
.B(n_8874),
.Y(n_11728)
);

OR2x2_ASAP7_75t_L g11729 ( 
.A(n_11468),
.B(n_8874),
.Y(n_11729)
);

INVx2_ASAP7_75t_L g11730 ( 
.A(n_11420),
.Y(n_11730)
);

OR2x2_ASAP7_75t_L g11731 ( 
.A(n_11399),
.B(n_8874),
.Y(n_11731)
);

NAND2xp5_ASAP7_75t_L g11732 ( 
.A(n_11559),
.B(n_11417),
.Y(n_11732)
);

INVx1_ASAP7_75t_SL g11733 ( 
.A(n_11551),
.Y(n_11733)
);

AND2x2_ASAP7_75t_L g11734 ( 
.A(n_11489),
.B(n_8495),
.Y(n_11734)
);

INVx1_ASAP7_75t_L g11735 ( 
.A(n_11622),
.Y(n_11735)
);

NAND2x1_ASAP7_75t_L g11736 ( 
.A(n_11562),
.B(n_8334),
.Y(n_11736)
);

AND2x2_ASAP7_75t_L g11737 ( 
.A(n_11490),
.B(n_8495),
.Y(n_11737)
);

INVx2_ASAP7_75t_SL g11738 ( 
.A(n_11438),
.Y(n_11738)
);

AOI211x1_ASAP7_75t_SL g11739 ( 
.A1(n_11457),
.A2(n_8338),
.B(n_8343),
.C(n_8340),
.Y(n_11739)
);

INVx1_ASAP7_75t_L g11740 ( 
.A(n_11524),
.Y(n_11740)
);

INVx1_ASAP7_75t_L g11741 ( 
.A(n_11440),
.Y(n_11741)
);

NAND2xp5_ASAP7_75t_SL g11742 ( 
.A(n_11435),
.B(n_8338),
.Y(n_11742)
);

INVx1_ASAP7_75t_L g11743 ( 
.A(n_11597),
.Y(n_11743)
);

NAND2xp5_ASAP7_75t_L g11744 ( 
.A(n_11481),
.B(n_7181),
.Y(n_11744)
);

AND2x2_ASAP7_75t_L g11745 ( 
.A(n_11511),
.B(n_11450),
.Y(n_11745)
);

INVx1_ASAP7_75t_L g11746 ( 
.A(n_11482),
.Y(n_11746)
);

NOR2xp33_ASAP7_75t_SL g11747 ( 
.A(n_11436),
.B(n_7941),
.Y(n_11747)
);

AND2x2_ASAP7_75t_L g11748 ( 
.A(n_11453),
.B(n_8372),
.Y(n_11748)
);

A2O1A1Ixp33_ASAP7_75t_R g11749 ( 
.A1(n_11626),
.A2(n_8845),
.B(n_8854),
.C(n_8848),
.Y(n_11749)
);

INVx1_ASAP7_75t_L g11750 ( 
.A(n_11391),
.Y(n_11750)
);

NAND2xp5_ASAP7_75t_L g11751 ( 
.A(n_11442),
.B(n_11456),
.Y(n_11751)
);

AND2x2_ASAP7_75t_L g11752 ( 
.A(n_11467),
.B(n_8354),
.Y(n_11752)
);

INVx1_ASAP7_75t_L g11753 ( 
.A(n_11400),
.Y(n_11753)
);

INVx2_ASAP7_75t_L g11754 ( 
.A(n_11564),
.Y(n_11754)
);

OR2x2_ASAP7_75t_L g11755 ( 
.A(n_11542),
.B(n_7779),
.Y(n_11755)
);

NAND2xp5_ASAP7_75t_L g11756 ( 
.A(n_11545),
.B(n_7181),
.Y(n_11756)
);

INVx1_ASAP7_75t_SL g11757 ( 
.A(n_11416),
.Y(n_11757)
);

INVx2_ASAP7_75t_L g11758 ( 
.A(n_11470),
.Y(n_11758)
);

OAI322xp33_ASAP7_75t_SL g11759 ( 
.A1(n_11451),
.A2(n_8340),
.A3(n_8343),
.B1(n_8352),
.B2(n_8353),
.C1(n_8351),
.C2(n_8346),
.Y(n_11759)
);

NOR2xp67_ASAP7_75t_L g11760 ( 
.A(n_11568),
.B(n_8346),
.Y(n_11760)
);

OR2x2_ASAP7_75t_L g11761 ( 
.A(n_11458),
.B(n_7779),
.Y(n_11761)
);

HB1xp67_ASAP7_75t_L g11762 ( 
.A(n_11643),
.Y(n_11762)
);

INVx1_ASAP7_75t_SL g11763 ( 
.A(n_11472),
.Y(n_11763)
);

INVx1_ASAP7_75t_L g11764 ( 
.A(n_11405),
.Y(n_11764)
);

AND2x2_ASAP7_75t_L g11765 ( 
.A(n_11574),
.B(n_11580),
.Y(n_11765)
);

AND2x2_ASAP7_75t_L g11766 ( 
.A(n_11506),
.B(n_8354),
.Y(n_11766)
);

INVx1_ASAP7_75t_L g11767 ( 
.A(n_11483),
.Y(n_11767)
);

NOR2xp33_ASAP7_75t_SL g11768 ( 
.A(n_11410),
.B(n_11619),
.Y(n_11768)
);

NOR2x1_ASAP7_75t_L g11769 ( 
.A(n_11392),
.B(n_8801),
.Y(n_11769)
);

AND2x2_ASAP7_75t_L g11770 ( 
.A(n_11623),
.B(n_7280),
.Y(n_11770)
);

INVx1_ASAP7_75t_SL g11771 ( 
.A(n_11638),
.Y(n_11771)
);

NAND2xp5_ASAP7_75t_L g11772 ( 
.A(n_11537),
.B(n_7181),
.Y(n_11772)
);

INVx1_ASAP7_75t_L g11773 ( 
.A(n_11557),
.Y(n_11773)
);

OAI221xp5_ASAP7_75t_L g11774 ( 
.A1(n_11454),
.A2(n_8265),
.B1(n_8262),
.B2(n_8311),
.C(n_8284),
.Y(n_11774)
);

INVx2_ASAP7_75t_SL g11775 ( 
.A(n_11488),
.Y(n_11775)
);

INVx1_ASAP7_75t_L g11776 ( 
.A(n_11567),
.Y(n_11776)
);

NOR2xp33_ASAP7_75t_L g11777 ( 
.A(n_11582),
.B(n_7181),
.Y(n_11777)
);

AND2x2_ASAP7_75t_L g11778 ( 
.A(n_11541),
.B(n_11598),
.Y(n_11778)
);

NAND2x1_ASAP7_75t_L g11779 ( 
.A(n_11488),
.B(n_8351),
.Y(n_11779)
);

OR2x2_ASAP7_75t_L g11780 ( 
.A(n_11460),
.B(n_7813),
.Y(n_11780)
);

NAND2xp5_ASAP7_75t_L g11781 ( 
.A(n_11479),
.B(n_7226),
.Y(n_11781)
);

AOI21xp33_ASAP7_75t_L g11782 ( 
.A1(n_11497),
.A2(n_8862),
.B(n_8859),
.Y(n_11782)
);

OR2x2_ASAP7_75t_L g11783 ( 
.A(n_11552),
.B(n_7813),
.Y(n_11783)
);

INVx1_ASAP7_75t_L g11784 ( 
.A(n_11448),
.Y(n_11784)
);

AND2x2_ASAP7_75t_L g11785 ( 
.A(n_11603),
.B(n_7280),
.Y(n_11785)
);

OR2x2_ASAP7_75t_L g11786 ( 
.A(n_11513),
.B(n_8864),
.Y(n_11786)
);

NAND2xp5_ASAP7_75t_L g11787 ( 
.A(n_11535),
.B(n_7226),
.Y(n_11787)
);

NAND2xp5_ASAP7_75t_L g11788 ( 
.A(n_11528),
.B(n_7226),
.Y(n_11788)
);

INVx1_ASAP7_75t_L g11789 ( 
.A(n_11533),
.Y(n_11789)
);

INVx1_ASAP7_75t_L g11790 ( 
.A(n_11415),
.Y(n_11790)
);

INVx1_ASAP7_75t_L g11791 ( 
.A(n_11426),
.Y(n_11791)
);

AND2x4_ASAP7_75t_L g11792 ( 
.A(n_11607),
.B(n_11549),
.Y(n_11792)
);

INVxp67_ASAP7_75t_L g11793 ( 
.A(n_11586),
.Y(n_11793)
);

AND2x2_ASAP7_75t_L g11794 ( 
.A(n_11620),
.B(n_8499),
.Y(n_11794)
);

INVx2_ASAP7_75t_L g11795 ( 
.A(n_11546),
.Y(n_11795)
);

INVx1_ASAP7_75t_L g11796 ( 
.A(n_11527),
.Y(n_11796)
);

INVx1_ASAP7_75t_L g11797 ( 
.A(n_11536),
.Y(n_11797)
);

OAI22xp5_ASAP7_75t_L g11798 ( 
.A1(n_11577),
.A2(n_8905),
.B1(n_8884),
.B2(n_8887),
.Y(n_11798)
);

NAND2xp5_ASAP7_75t_L g11799 ( 
.A(n_11505),
.B(n_7226),
.Y(n_11799)
);

NAND4xp25_ASAP7_75t_L g11800 ( 
.A(n_11434),
.B(n_7875),
.C(n_7800),
.D(n_7945),
.Y(n_11800)
);

NAND2x1_ASAP7_75t_L g11801 ( 
.A(n_11581),
.B(n_8352),
.Y(n_11801)
);

INVx2_ASAP7_75t_L g11802 ( 
.A(n_11522),
.Y(n_11802)
);

NAND2xp33_ASAP7_75t_SL g11803 ( 
.A(n_11565),
.B(n_8353),
.Y(n_11803)
);

NAND3xp33_ASAP7_75t_SL g11804 ( 
.A(n_11590),
.B(n_8035),
.C(n_8033),
.Y(n_11804)
);

HB1xp67_ASAP7_75t_L g11805 ( 
.A(n_11498),
.Y(n_11805)
);

NAND2x1_ASAP7_75t_L g11806 ( 
.A(n_11627),
.B(n_8358),
.Y(n_11806)
);

OR2x2_ASAP7_75t_L g11807 ( 
.A(n_11430),
.B(n_8918),
.Y(n_11807)
);

AND2x2_ASAP7_75t_L g11808 ( 
.A(n_11563),
.B(n_8499),
.Y(n_11808)
);

INVx1_ASAP7_75t_L g11809 ( 
.A(n_11449),
.Y(n_11809)
);

OR2x2_ASAP7_75t_L g11810 ( 
.A(n_11595),
.B(n_11462),
.Y(n_11810)
);

INVx1_ASAP7_75t_L g11811 ( 
.A(n_11463),
.Y(n_11811)
);

AND2x2_ASAP7_75t_L g11812 ( 
.A(n_11525),
.B(n_8499),
.Y(n_11812)
);

AND2x2_ASAP7_75t_L g11813 ( 
.A(n_11544),
.B(n_11548),
.Y(n_11813)
);

INVx1_ASAP7_75t_L g11814 ( 
.A(n_11532),
.Y(n_11814)
);

INVx1_ASAP7_75t_L g11815 ( 
.A(n_11502),
.Y(n_11815)
);

AOI22xp5_ASAP7_75t_L g11816 ( 
.A1(n_11601),
.A2(n_8801),
.B1(n_8892),
.B2(n_8873),
.Y(n_11816)
);

INVx1_ASAP7_75t_L g11817 ( 
.A(n_11606),
.Y(n_11817)
);

INVx2_ASAP7_75t_L g11818 ( 
.A(n_11576),
.Y(n_11818)
);

INVx2_ASAP7_75t_L g11819 ( 
.A(n_11566),
.Y(n_11819)
);

INVx1_ASAP7_75t_L g11820 ( 
.A(n_11609),
.Y(n_11820)
);

INVx1_ASAP7_75t_L g11821 ( 
.A(n_11612),
.Y(n_11821)
);

AND2x2_ASAP7_75t_L g11822 ( 
.A(n_11616),
.B(n_8152),
.Y(n_11822)
);

INVx1_ASAP7_75t_SL g11823 ( 
.A(n_11614),
.Y(n_11823)
);

OAI21xp33_ASAP7_75t_SL g11824 ( 
.A1(n_11518),
.A2(n_11480),
.B(n_11486),
.Y(n_11824)
);

INVx1_ASAP7_75t_SL g11825 ( 
.A(n_11491),
.Y(n_11825)
);

INVx1_ASAP7_75t_L g11826 ( 
.A(n_11617),
.Y(n_11826)
);

INVx2_ASAP7_75t_L g11827 ( 
.A(n_11627),
.Y(n_11827)
);

OR2x2_ASAP7_75t_L g11828 ( 
.A(n_11515),
.B(n_8904),
.Y(n_11828)
);

NAND2xp5_ASAP7_75t_L g11829 ( 
.A(n_11485),
.B(n_7228),
.Y(n_11829)
);

NAND2xp5_ASAP7_75t_L g11830 ( 
.A(n_11418),
.B(n_11531),
.Y(n_11830)
);

NAND2xp5_ASAP7_75t_L g11831 ( 
.A(n_11554),
.B(n_7228),
.Y(n_11831)
);

INVx1_ASAP7_75t_L g11832 ( 
.A(n_11618),
.Y(n_11832)
);

INVx1_ASAP7_75t_L g11833 ( 
.A(n_11621),
.Y(n_11833)
);

INVx1_ASAP7_75t_L g11834 ( 
.A(n_11625),
.Y(n_11834)
);

INVx1_ASAP7_75t_L g11835 ( 
.A(n_11633),
.Y(n_11835)
);

AND2x2_ASAP7_75t_L g11836 ( 
.A(n_11547),
.B(n_8908),
.Y(n_11836)
);

AND2x2_ASAP7_75t_L g11837 ( 
.A(n_11507),
.B(n_8909),
.Y(n_11837)
);

INVxp67_ASAP7_75t_SL g11838 ( 
.A(n_11589),
.Y(n_11838)
);

OR2x6_ASAP7_75t_L g11839 ( 
.A(n_11530),
.B(n_7228),
.Y(n_11839)
);

OR2x2_ASAP7_75t_L g11840 ( 
.A(n_11520),
.B(n_8919),
.Y(n_11840)
);

INVx2_ASAP7_75t_L g11841 ( 
.A(n_11642),
.Y(n_11841)
);

INVx1_ASAP7_75t_L g11842 ( 
.A(n_11431),
.Y(n_11842)
);

NOR2xp33_ASAP7_75t_L g11843 ( 
.A(n_11600),
.B(n_7228),
.Y(n_11843)
);

INVx1_ASAP7_75t_L g11844 ( 
.A(n_11431),
.Y(n_11844)
);

INVx2_ASAP7_75t_SL g11845 ( 
.A(n_11624),
.Y(n_11845)
);

OAI22xp5_ASAP7_75t_L g11846 ( 
.A1(n_11636),
.A2(n_8920),
.B1(n_7307),
.B2(n_7345),
.Y(n_11846)
);

INVx1_ASAP7_75t_L g11847 ( 
.A(n_11501),
.Y(n_11847)
);

INVxp67_ASAP7_75t_L g11848 ( 
.A(n_11504),
.Y(n_11848)
);

OAI21xp33_ASAP7_75t_L g11849 ( 
.A1(n_11644),
.A2(n_8358),
.B(n_8889),
.Y(n_11849)
);

AND2x2_ASAP7_75t_L g11850 ( 
.A(n_11602),
.B(n_7307),
.Y(n_11850)
);

INVx2_ASAP7_75t_L g11851 ( 
.A(n_11583),
.Y(n_11851)
);

INVx2_ASAP7_75t_SL g11852 ( 
.A(n_11637),
.Y(n_11852)
);

AND2x2_ASAP7_75t_L g11853 ( 
.A(n_11604),
.B(n_7307),
.Y(n_11853)
);

AND2x2_ASAP7_75t_L g11854 ( 
.A(n_11517),
.B(n_11521),
.Y(n_11854)
);

AND2x2_ASAP7_75t_L g11855 ( 
.A(n_11526),
.B(n_7312),
.Y(n_11855)
);

NAND2xp5_ASAP7_75t_L g11856 ( 
.A(n_11645),
.B(n_7312),
.Y(n_11856)
);

INVx1_ASAP7_75t_L g11857 ( 
.A(n_11540),
.Y(n_11857)
);

INVx2_ASAP7_75t_L g11858 ( 
.A(n_11593),
.Y(n_11858)
);

INVx3_ASAP7_75t_L g11859 ( 
.A(n_11569),
.Y(n_11859)
);

AND2x2_ASAP7_75t_L g11860 ( 
.A(n_11635),
.B(n_7312),
.Y(n_11860)
);

NAND2xp33_ASAP7_75t_SL g11861 ( 
.A(n_11519),
.B(n_8891),
.Y(n_11861)
);

AOI322xp5_ASAP7_75t_L g11862 ( 
.A1(n_11608),
.A2(n_8102),
.A3(n_8071),
.B1(n_8288),
.B2(n_8291),
.C1(n_8283),
.C2(n_7965),
.Y(n_11862)
);

NAND2xp5_ASAP7_75t_L g11863 ( 
.A(n_11605),
.B(n_7312),
.Y(n_11863)
);

INVx1_ASAP7_75t_L g11864 ( 
.A(n_11534),
.Y(n_11864)
);

NAND3xp33_ASAP7_75t_L g11865 ( 
.A(n_11573),
.B(n_8889),
.C(n_8891),
.Y(n_11865)
);

INVx1_ASAP7_75t_L g11866 ( 
.A(n_11570),
.Y(n_11866)
);

OAI32xp33_ASAP7_75t_L g11867 ( 
.A1(n_11629),
.A2(n_8846),
.A3(n_8899),
.B1(n_8893),
.B2(n_7989),
.Y(n_11867)
);

INVx2_ASAP7_75t_L g11868 ( 
.A(n_11639),
.Y(n_11868)
);

NOR2xp33_ASAP7_75t_L g11869 ( 
.A(n_11508),
.B(n_7345),
.Y(n_11869)
);

OR2x2_ASAP7_75t_L g11870 ( 
.A(n_11584),
.B(n_8279),
.Y(n_11870)
);

INVx1_ASAP7_75t_L g11871 ( 
.A(n_11561),
.Y(n_11871)
);

OR2x2_ASAP7_75t_L g11872 ( 
.A(n_11555),
.B(n_8518),
.Y(n_11872)
);

AOI311xp33_ASAP7_75t_L g11873 ( 
.A1(n_11477),
.A2(n_7969),
.A3(n_7968),
.B(n_7940),
.C(n_8080),
.Y(n_11873)
);

AND2x4_ASAP7_75t_L g11874 ( 
.A(n_11571),
.B(n_8750),
.Y(n_11874)
);

INVx2_ASAP7_75t_L g11875 ( 
.A(n_11615),
.Y(n_11875)
);

NAND2xp5_ASAP7_75t_L g11876 ( 
.A(n_11641),
.B(n_7345),
.Y(n_11876)
);

AND2x4_ASAP7_75t_L g11877 ( 
.A(n_11575),
.B(n_8750),
.Y(n_11877)
);

OR2x2_ASAP7_75t_L g11878 ( 
.A(n_11484),
.B(n_8518),
.Y(n_11878)
);

INVxp67_ASAP7_75t_SL g11879 ( 
.A(n_11640),
.Y(n_11879)
);

INVx1_ASAP7_75t_SL g11880 ( 
.A(n_11611),
.Y(n_11880)
);

INVx2_ASAP7_75t_L g11881 ( 
.A(n_11628),
.Y(n_11881)
);

OR2x2_ASAP7_75t_L g11882 ( 
.A(n_11503),
.B(n_11587),
.Y(n_11882)
);

AND3x2_ASAP7_75t_L g11883 ( 
.A(n_11591),
.B(n_8899),
.C(n_8893),
.Y(n_11883)
);

INVx1_ASAP7_75t_L g11884 ( 
.A(n_11572),
.Y(n_11884)
);

INVx1_ASAP7_75t_L g11885 ( 
.A(n_11592),
.Y(n_11885)
);

AOI22xp5_ASAP7_75t_L g11886 ( 
.A1(n_11538),
.A2(n_7393),
.B1(n_7396),
.B2(n_7345),
.Y(n_11886)
);

AOI22xp5_ASAP7_75t_L g11887 ( 
.A1(n_11660),
.A2(n_11631),
.B1(n_11596),
.B2(n_11599),
.Y(n_11887)
);

INVx1_ASAP7_75t_L g11888 ( 
.A(n_11678),
.Y(n_11888)
);

OAI221xp5_ASAP7_75t_L g11889 ( 
.A1(n_11655),
.A2(n_11630),
.B1(n_11632),
.B2(n_8267),
.C(n_7822),
.Y(n_11889)
);

INVx2_ASAP7_75t_L g11890 ( 
.A(n_11665),
.Y(n_11890)
);

NAND2xp5_ASAP7_75t_L g11891 ( 
.A(n_11710),
.B(n_11493),
.Y(n_11891)
);

NAND2xp5_ASAP7_75t_L g11892 ( 
.A(n_11719),
.B(n_11493),
.Y(n_11892)
);

NAND2xp5_ASAP7_75t_L g11893 ( 
.A(n_11647),
.B(n_11578),
.Y(n_11893)
);

INVx1_ASAP7_75t_L g11894 ( 
.A(n_11678),
.Y(n_11894)
);

INVx1_ASAP7_75t_L g11895 ( 
.A(n_11654),
.Y(n_11895)
);

INVx1_ASAP7_75t_L g11896 ( 
.A(n_11654),
.Y(n_11896)
);

OAI21xp5_ASAP7_75t_L g11897 ( 
.A1(n_11698),
.A2(n_11578),
.B(n_8701),
.Y(n_11897)
);

AO21x1_ASAP7_75t_SL g11898 ( 
.A1(n_11656),
.A2(n_7817),
.B(n_7812),
.Y(n_11898)
);

INVxp67_ASAP7_75t_L g11899 ( 
.A(n_11658),
.Y(n_11899)
);

INVx3_ASAP7_75t_L g11900 ( 
.A(n_11721),
.Y(n_11900)
);

INVx1_ASAP7_75t_L g11901 ( 
.A(n_11657),
.Y(n_11901)
);

NAND2xp5_ASAP7_75t_SL g11902 ( 
.A(n_11721),
.B(n_11720),
.Y(n_11902)
);

NAND3x2_ASAP7_75t_L g11903 ( 
.A(n_11725),
.B(n_7943),
.C(n_8518),
.Y(n_11903)
);

NAND3xp33_ASAP7_75t_L g11904 ( 
.A(n_11695),
.B(n_8437),
.C(n_8359),
.Y(n_11904)
);

INVx2_ASAP7_75t_L g11905 ( 
.A(n_11716),
.Y(n_11905)
);

INVx1_ASAP7_75t_L g11906 ( 
.A(n_11672),
.Y(n_11906)
);

INVx1_ASAP7_75t_L g11907 ( 
.A(n_11650),
.Y(n_11907)
);

INVx1_ASAP7_75t_L g11908 ( 
.A(n_11651),
.Y(n_11908)
);

AOI21xp33_ASAP7_75t_SL g11909 ( 
.A1(n_11652),
.A2(n_8437),
.B(n_8536),
.Y(n_11909)
);

INVx1_ASAP7_75t_L g11910 ( 
.A(n_11745),
.Y(n_11910)
);

INVx2_ASAP7_75t_L g11911 ( 
.A(n_11681),
.Y(n_11911)
);

NOR2xp33_ASAP7_75t_L g11912 ( 
.A(n_11667),
.B(n_11771),
.Y(n_11912)
);

OR2x2_ASAP7_75t_L g11913 ( 
.A(n_11733),
.B(n_8437),
.Y(n_11913)
);

INVx1_ASAP7_75t_L g11914 ( 
.A(n_11649),
.Y(n_11914)
);

INVx1_ASAP7_75t_L g11915 ( 
.A(n_11762),
.Y(n_11915)
);

NAND2xp5_ASAP7_75t_SL g11916 ( 
.A(n_11688),
.B(n_7393),
.Y(n_11916)
);

NOR2xp67_ASAP7_75t_SL g11917 ( 
.A(n_11707),
.B(n_7393),
.Y(n_11917)
);

INVx1_ASAP7_75t_L g11918 ( 
.A(n_11706),
.Y(n_11918)
);

AOI22x1_ASAP7_75t_SL g11919 ( 
.A1(n_11693),
.A2(n_7396),
.B1(n_7463),
.B2(n_7393),
.Y(n_11919)
);

NOR2xp33_ASAP7_75t_L g11920 ( 
.A(n_11663),
.B(n_7396),
.Y(n_11920)
);

AOI22xp33_ASAP7_75t_L g11921 ( 
.A1(n_11804),
.A2(n_8359),
.B1(n_8761),
.B2(n_8759),
.Y(n_11921)
);

OR2x2_ASAP7_75t_L g11922 ( 
.A(n_11704),
.B(n_8359),
.Y(n_11922)
);

OAI22xp5_ASAP7_75t_L g11923 ( 
.A1(n_11757),
.A2(n_7463),
.B1(n_7396),
.B2(n_8275),
.Y(n_11923)
);

INVx1_ASAP7_75t_L g11924 ( 
.A(n_11686),
.Y(n_11924)
);

INVx1_ASAP7_75t_L g11925 ( 
.A(n_11686),
.Y(n_11925)
);

OAI32xp33_ASAP7_75t_L g11926 ( 
.A1(n_11739),
.A2(n_7463),
.A3(n_8316),
.B1(n_8078),
.B2(n_7741),
.Y(n_11926)
);

INVx1_ASAP7_75t_L g11927 ( 
.A(n_11664),
.Y(n_11927)
);

NAND2xp5_ASAP7_75t_L g11928 ( 
.A(n_11775),
.B(n_7463),
.Y(n_11928)
);

OAI22xp33_ASAP7_75t_L g11929 ( 
.A1(n_11747),
.A2(n_8282),
.B1(n_8776),
.B2(n_8705),
.Y(n_11929)
);

NAND2xp5_ASAP7_75t_SL g11930 ( 
.A(n_11708),
.B(n_8701),
.Y(n_11930)
);

AOI22xp5_ASAP7_75t_L g11931 ( 
.A1(n_11768),
.A2(n_8241),
.B1(n_8219),
.B2(n_8535),
.Y(n_11931)
);

INVx1_ASAP7_75t_SL g11932 ( 
.A(n_11709),
.Y(n_11932)
);

AOI21xp5_ASAP7_75t_L g11933 ( 
.A1(n_11692),
.A2(n_8761),
.B(n_8759),
.Y(n_11933)
);

INVx1_ASAP7_75t_L g11934 ( 
.A(n_11694),
.Y(n_11934)
);

OAI32xp33_ASAP7_75t_L g11935 ( 
.A1(n_11711),
.A2(n_7764),
.A3(n_7799),
.B1(n_7741),
.B2(n_7740),
.Y(n_11935)
);

INVx1_ASAP7_75t_L g11936 ( 
.A(n_11646),
.Y(n_11936)
);

OAI22xp5_ASAP7_75t_L g11937 ( 
.A1(n_11774),
.A2(n_8312),
.B1(n_8307),
.B2(n_7980),
.Y(n_11937)
);

INVx2_ASAP7_75t_L g11938 ( 
.A(n_11883),
.Y(n_11938)
);

NAND2xp5_ASAP7_75t_L g11939 ( 
.A(n_11760),
.B(n_8535),
.Y(n_11939)
);

NAND2xp5_ASAP7_75t_SL g11940 ( 
.A(n_11738),
.B(n_8256),
.Y(n_11940)
);

OAI211xp5_ASAP7_75t_L g11941 ( 
.A1(n_11673),
.A2(n_8206),
.B(n_7979),
.C(n_8776),
.Y(n_11941)
);

INVx1_ASAP7_75t_L g11942 ( 
.A(n_11736),
.Y(n_11942)
);

HB1xp67_ASAP7_75t_L g11943 ( 
.A(n_11779),
.Y(n_11943)
);

NAND2xp5_ASAP7_75t_L g11944 ( 
.A(n_11683),
.B(n_8535),
.Y(n_11944)
);

INVx1_ASAP7_75t_L g11945 ( 
.A(n_11736),
.Y(n_11945)
);

INVx1_ASAP7_75t_L g11946 ( 
.A(n_11714),
.Y(n_11946)
);

INVx1_ASAP7_75t_L g11947 ( 
.A(n_11671),
.Y(n_11947)
);

AOI21xp5_ASAP7_75t_L g11948 ( 
.A1(n_11769),
.A2(n_8761),
.B(n_8759),
.Y(n_11948)
);

INVx2_ASAP7_75t_SL g11949 ( 
.A(n_11683),
.Y(n_11949)
);

AOI32xp33_ASAP7_75t_L g11950 ( 
.A1(n_11873),
.A2(n_8301),
.A3(n_8298),
.B1(n_8303),
.B2(n_8200),
.Y(n_11950)
);

A2O1A1Ixp33_ASAP7_75t_L g11951 ( 
.A1(n_11675),
.A2(n_8172),
.B(n_7082),
.C(n_7090),
.Y(n_11951)
);

INVx2_ASAP7_75t_L g11952 ( 
.A(n_11874),
.Y(n_11952)
);

INVx1_ASAP7_75t_L g11953 ( 
.A(n_11687),
.Y(n_11953)
);

OAI211xp5_ASAP7_75t_L g11954 ( 
.A1(n_11690),
.A2(n_8776),
.B(n_8705),
.C(n_7802),
.Y(n_11954)
);

NOR2xp33_ASAP7_75t_SL g11955 ( 
.A(n_11659),
.B(n_8201),
.Y(n_11955)
);

AND2x2_ASAP7_75t_L g11956 ( 
.A(n_11653),
.B(n_7565),
.Y(n_11956)
);

HB1xp67_ASAP7_75t_L g11957 ( 
.A(n_11801),
.Y(n_11957)
);

NAND2xp5_ASAP7_75t_L g11958 ( 
.A(n_11674),
.B(n_8439),
.Y(n_11958)
);

OAI22xp5_ASAP7_75t_L g11959 ( 
.A1(n_11668),
.A2(n_7807),
.B1(n_8705),
.B2(n_8591),
.Y(n_11959)
);

OAI22xp5_ASAP7_75t_L g11960 ( 
.A1(n_11689),
.A2(n_8591),
.B1(n_7907),
.B2(n_7914),
.Y(n_11960)
);

INVx1_ASAP7_75t_L g11961 ( 
.A(n_11679),
.Y(n_11961)
);

OR2x2_ASAP7_75t_L g11962 ( 
.A(n_11699),
.B(n_8439),
.Y(n_11962)
);

INVx1_ASAP7_75t_L g11963 ( 
.A(n_11669),
.Y(n_11963)
);

AND2x4_ASAP7_75t_L g11964 ( 
.A(n_11792),
.B(n_8897),
.Y(n_11964)
);

AOI22xp5_ASAP7_75t_L g11965 ( 
.A1(n_11661),
.A2(n_8721),
.B1(n_8439),
.B2(n_8766),
.Y(n_11965)
);

INVx1_ASAP7_75t_L g11966 ( 
.A(n_11670),
.Y(n_11966)
);

INVx2_ASAP7_75t_L g11967 ( 
.A(n_11874),
.Y(n_11967)
);

AOI22xp33_ASAP7_75t_L g11968 ( 
.A1(n_11701),
.A2(n_8766),
.B1(n_8721),
.B2(n_8731),
.Y(n_11968)
);

NAND2xp5_ASAP7_75t_L g11969 ( 
.A(n_11792),
.B(n_11724),
.Y(n_11969)
);

INVx1_ASAP7_75t_L g11970 ( 
.A(n_11648),
.Y(n_11970)
);

OAI21xp33_ASAP7_75t_L g11971 ( 
.A1(n_11800),
.A2(n_8329),
.B(n_8323),
.Y(n_11971)
);

OAI22xp5_ASAP7_75t_L g11972 ( 
.A1(n_11793),
.A2(n_8591),
.B1(n_7916),
.B2(n_7905),
.Y(n_11972)
);

NAND2xp5_ASAP7_75t_L g11973 ( 
.A(n_11712),
.B(n_8721),
.Y(n_11973)
);

INVx1_ASAP7_75t_L g11974 ( 
.A(n_11696),
.Y(n_11974)
);

INVx1_ASAP7_75t_L g11975 ( 
.A(n_11770),
.Y(n_11975)
);

OAI31xp33_ASAP7_75t_L g11976 ( 
.A1(n_11763),
.A2(n_8060),
.A3(n_8061),
.B(n_6859),
.Y(n_11976)
);

INVx2_ASAP7_75t_L g11977 ( 
.A(n_11877),
.Y(n_11977)
);

AOI221xp5_ASAP7_75t_L g11978 ( 
.A1(n_11662),
.A2(n_8766),
.B1(n_8722),
.B2(n_8902),
.C(n_8897),
.Y(n_11978)
);

OAI21xp5_ASAP7_75t_L g11979 ( 
.A1(n_11732),
.A2(n_8731),
.B(n_8857),
.Y(n_11979)
);

INVx1_ASAP7_75t_L g11980 ( 
.A(n_11765),
.Y(n_11980)
);

O2A1O1Ixp5_ASAP7_75t_L g11981 ( 
.A1(n_11801),
.A2(n_7764),
.B(n_7799),
.C(n_7740),
.Y(n_11981)
);

NAND2xp5_ASAP7_75t_L g11982 ( 
.A(n_11726),
.B(n_8722),
.Y(n_11982)
);

NAND3xp33_ASAP7_75t_L g11983 ( 
.A(n_11727),
.B(n_8731),
.C(n_8857),
.Y(n_11983)
);

INVx1_ASAP7_75t_L g11984 ( 
.A(n_11722),
.Y(n_11984)
);

HB1xp67_ASAP7_75t_L g11985 ( 
.A(n_11806),
.Y(n_11985)
);

OAI22xp5_ASAP7_75t_L g11986 ( 
.A1(n_11825),
.A2(n_7359),
.B1(n_7022),
.B2(n_6859),
.Y(n_11986)
);

INVx1_ASAP7_75t_L g11987 ( 
.A(n_11715),
.Y(n_11987)
);

AND2x4_ASAP7_75t_L g11988 ( 
.A(n_11827),
.B(n_8897),
.Y(n_11988)
);

INVx2_ASAP7_75t_L g11989 ( 
.A(n_11877),
.Y(n_11989)
);

NOR2xp33_ASAP7_75t_L g11990 ( 
.A(n_11796),
.B(n_8722),
.Y(n_11990)
);

HB1xp67_ASAP7_75t_L g11991 ( 
.A(n_11794),
.Y(n_11991)
);

OAI22xp33_ASAP7_75t_L g11992 ( 
.A1(n_11886),
.A2(n_11740),
.B1(n_11743),
.B2(n_11735),
.Y(n_11992)
);

INVx2_ASAP7_75t_L g11993 ( 
.A(n_11729),
.Y(n_11993)
);

OAI21xp5_ASAP7_75t_SL g11994 ( 
.A1(n_11791),
.A2(n_8055),
.B(n_8092),
.Y(n_11994)
);

AND2x2_ASAP7_75t_L g11995 ( 
.A(n_11666),
.B(n_11684),
.Y(n_11995)
);

AND2x2_ASAP7_75t_L g11996 ( 
.A(n_11778),
.B(n_7565),
.Y(n_11996)
);

INVx2_ASAP7_75t_L g11997 ( 
.A(n_11717),
.Y(n_11997)
);

OAI22xp5_ASAP7_75t_SL g11998 ( 
.A1(n_11741),
.A2(n_11852),
.B1(n_11845),
.B2(n_11713),
.Y(n_11998)
);

OAI21xp33_ASAP7_75t_SL g11999 ( 
.A1(n_11862),
.A2(n_7809),
.B(n_7803),
.Y(n_11999)
);

INVx1_ASAP7_75t_L g12000 ( 
.A(n_11703),
.Y(n_12000)
);

NOR3xp33_ASAP7_75t_L g12001 ( 
.A(n_11685),
.B(n_6946),
.C(n_7077),
.Y(n_12001)
);

NAND2xp5_ASAP7_75t_L g12002 ( 
.A(n_11748),
.B(n_6820),
.Y(n_12002)
);

NAND2xp5_ASAP7_75t_L g12003 ( 
.A(n_11802),
.B(n_6820),
.Y(n_12003)
);

OAI22xp5_ASAP7_75t_L g12004 ( 
.A1(n_11758),
.A2(n_7359),
.B1(n_7022),
.B2(n_8911),
.Y(n_12004)
);

NOR2xp33_ASAP7_75t_L g12005 ( 
.A(n_11730),
.B(n_8902),
.Y(n_12005)
);

INVx1_ASAP7_75t_L g12006 ( 
.A(n_11752),
.Y(n_12006)
);

INVx2_ASAP7_75t_SL g12007 ( 
.A(n_11882),
.Y(n_12007)
);

OAI22xp5_ASAP7_75t_L g12008 ( 
.A1(n_11751),
.A2(n_8857),
.B1(n_8911),
.B2(n_7532),
.Y(n_12008)
);

NAND3xp33_ASAP7_75t_L g12009 ( 
.A(n_11723),
.B(n_8911),
.C(n_6829),
.Y(n_12009)
);

OAI21xp5_ASAP7_75t_SL g12010 ( 
.A1(n_11823),
.A2(n_8095),
.B(n_8104),
.Y(n_12010)
);

INVx1_ASAP7_75t_L g12011 ( 
.A(n_11677),
.Y(n_12011)
);

INVx1_ASAP7_75t_L g12012 ( 
.A(n_11691),
.Y(n_12012)
);

NOR2xp33_ASAP7_75t_L g12013 ( 
.A(n_11814),
.B(n_8902),
.Y(n_12013)
);

INVx2_ASAP7_75t_L g12014 ( 
.A(n_11728),
.Y(n_12014)
);

NAND2xp5_ASAP7_75t_L g12015 ( 
.A(n_11795),
.B(n_7034),
.Y(n_12015)
);

NAND3xp33_ASAP7_75t_SL g12016 ( 
.A(n_11697),
.B(n_8112),
.C(n_8109),
.Y(n_12016)
);

NOR2xp33_ASAP7_75t_L g12017 ( 
.A(n_11746),
.B(n_8603),
.Y(n_12017)
);

INVx2_ASAP7_75t_L g12018 ( 
.A(n_11766),
.Y(n_12018)
);

INVx1_ASAP7_75t_L g12019 ( 
.A(n_11822),
.Y(n_12019)
);

INVx1_ASAP7_75t_L g12020 ( 
.A(n_11818),
.Y(n_12020)
);

INVx2_ASAP7_75t_SL g12021 ( 
.A(n_11807),
.Y(n_12021)
);

OR2x2_ASAP7_75t_L g12022 ( 
.A(n_11772),
.B(n_7034),
.Y(n_12022)
);

NAND2xp5_ASAP7_75t_L g12023 ( 
.A(n_11785),
.B(n_7034),
.Y(n_12023)
);

AND2x2_ASAP7_75t_L g12024 ( 
.A(n_11680),
.B(n_7583),
.Y(n_12024)
);

INVxp67_ASAP7_75t_L g12025 ( 
.A(n_11777),
.Y(n_12025)
);

AO21x1_ASAP7_75t_L g12026 ( 
.A1(n_11803),
.A2(n_7809),
.B(n_7803),
.Y(n_12026)
);

AOI211xp5_ASAP7_75t_SL g12027 ( 
.A1(n_11682),
.A2(n_8270),
.B(n_7549),
.C(n_7529),
.Y(n_12027)
);

A2O1A1Ixp33_ASAP7_75t_R g12028 ( 
.A1(n_11813),
.A2(n_7568),
.B(n_7579),
.C(n_7583),
.Y(n_12028)
);

AOI221xp5_ASAP7_75t_L g12029 ( 
.A1(n_11782),
.A2(n_11759),
.B1(n_11849),
.B2(n_11867),
.C(n_11798),
.Y(n_12029)
);

INVx2_ASAP7_75t_SL g12030 ( 
.A(n_11839),
.Y(n_12030)
);

NOR3xp33_ASAP7_75t_L g12031 ( 
.A(n_11676),
.B(n_7082),
.C(n_7077),
.Y(n_12031)
);

OAI221xp5_ASAP7_75t_SL g12032 ( 
.A1(n_11816),
.A2(n_11824),
.B1(n_11767),
.B2(n_11848),
.C(n_11810),
.Y(n_12032)
);

AND2x2_ASAP7_75t_L g12033 ( 
.A(n_11700),
.B(n_7617),
.Y(n_12033)
);

INVx1_ASAP7_75t_L g12034 ( 
.A(n_11754),
.Y(n_12034)
);

OAI22xp5_ASAP7_75t_L g12035 ( 
.A1(n_11789),
.A2(n_8120),
.B1(n_7568),
.B2(n_7579),
.Y(n_12035)
);

NAND2xp5_ASAP7_75t_L g12036 ( 
.A(n_11859),
.B(n_7034),
.Y(n_12036)
);

OAI21xp33_ASAP7_75t_L g12037 ( 
.A1(n_11869),
.A2(n_8096),
.B(n_7865),
.Y(n_12037)
);

OAI21xp5_ASAP7_75t_L g12038 ( 
.A1(n_11773),
.A2(n_7098),
.B(n_7090),
.Y(n_12038)
);

NAND2xp5_ASAP7_75t_L g12039 ( 
.A(n_11776),
.B(n_7034),
.Y(n_12039)
);

AND2x2_ASAP7_75t_L g12040 ( 
.A(n_11753),
.B(n_7617),
.Y(n_12040)
);

INVxp67_ASAP7_75t_L g12041 ( 
.A(n_11843),
.Y(n_12041)
);

NAND2xp5_ASAP7_75t_L g12042 ( 
.A(n_11797),
.B(n_7034),
.Y(n_12042)
);

OAI22xp33_ASAP7_75t_L g12043 ( 
.A1(n_11731),
.A2(n_7865),
.B1(n_7868),
.B2(n_7863),
.Y(n_12043)
);

AOI211xp5_ASAP7_75t_L g12044 ( 
.A1(n_11857),
.A2(n_7615),
.B(n_7098),
.C(n_7105),
.Y(n_12044)
);

INVx1_ASAP7_75t_SL g12045 ( 
.A(n_11734),
.Y(n_12045)
);

OR2x2_ASAP7_75t_L g12046 ( 
.A(n_11744),
.B(n_7136),
.Y(n_12046)
);

INVx2_ASAP7_75t_L g12047 ( 
.A(n_11839),
.Y(n_12047)
);

INVx1_ASAP7_75t_L g12048 ( 
.A(n_11842),
.Y(n_12048)
);

INVx1_ASAP7_75t_L g12049 ( 
.A(n_11844),
.Y(n_12049)
);

INVxp67_ASAP7_75t_L g12050 ( 
.A(n_11742),
.Y(n_12050)
);

INVx1_ASAP7_75t_L g12051 ( 
.A(n_11787),
.Y(n_12051)
);

AND2x4_ASAP7_75t_L g12052 ( 
.A(n_11837),
.B(n_8603),
.Y(n_12052)
);

OAI22xp5_ASAP7_75t_L g12053 ( 
.A1(n_11750),
.A2(n_7868),
.B1(n_7877),
.B2(n_7863),
.Y(n_12053)
);

OAI21xp33_ASAP7_75t_L g12054 ( 
.A1(n_11830),
.A2(n_7896),
.B(n_7877),
.Y(n_12054)
);

OAI22xp5_ASAP7_75t_L g12055 ( 
.A1(n_11764),
.A2(n_7897),
.B1(n_7896),
.B2(n_8065),
.Y(n_12055)
);

INVx1_ASAP7_75t_L g12056 ( 
.A(n_11756),
.Y(n_12056)
);

INVx3_ASAP7_75t_L g12057 ( 
.A(n_11855),
.Y(n_12057)
);

OAI22xp33_ASAP7_75t_L g12058 ( 
.A1(n_11829),
.A2(n_7897),
.B1(n_7543),
.B2(n_7591),
.Y(n_12058)
);

INVxp67_ASAP7_75t_SL g12059 ( 
.A(n_11737),
.Y(n_12059)
);

OAI22xp5_ASAP7_75t_L g12060 ( 
.A1(n_11784),
.A2(n_11790),
.B1(n_11809),
.B2(n_11811),
.Y(n_12060)
);

HB1xp67_ASAP7_75t_L g12061 ( 
.A(n_11808),
.Y(n_12061)
);

OAI21xp33_ASAP7_75t_L g12062 ( 
.A1(n_11854),
.A2(n_7543),
.B(n_8047),
.Y(n_12062)
);

AND2x2_ASAP7_75t_L g12063 ( 
.A(n_11850),
.B(n_11853),
.Y(n_12063)
);

INVx2_ASAP7_75t_L g12064 ( 
.A(n_11783),
.Y(n_12064)
);

A2O1A1Ixp33_ASAP7_75t_L g12065 ( 
.A1(n_11705),
.A2(n_7105),
.B(n_7107),
.C(n_7100),
.Y(n_12065)
);

NAND2xp5_ASAP7_75t_L g12066 ( 
.A(n_11858),
.B(n_7358),
.Y(n_12066)
);

AOI21xp33_ASAP7_75t_L g12067 ( 
.A1(n_11749),
.A2(n_8632),
.B(n_8603),
.Y(n_12067)
);

INVx1_ASAP7_75t_L g12068 ( 
.A(n_11856),
.Y(n_12068)
);

INVx1_ASAP7_75t_L g12069 ( 
.A(n_11780),
.Y(n_12069)
);

NAND2x1p5_ASAP7_75t_L g12070 ( 
.A(n_11885),
.B(n_7100),
.Y(n_12070)
);

NOR2xp33_ASAP7_75t_L g12071 ( 
.A(n_11761),
.B(n_8632),
.Y(n_12071)
);

NAND2xp5_ASAP7_75t_L g12072 ( 
.A(n_11860),
.B(n_7358),
.Y(n_12072)
);

INVx1_ASAP7_75t_L g12073 ( 
.A(n_11836),
.Y(n_12073)
);

A2O1A1Ixp33_ASAP7_75t_L g12074 ( 
.A1(n_11819),
.A2(n_7117),
.B(n_7132),
.C(n_7107),
.Y(n_12074)
);

NAND2xp5_ASAP7_75t_L g12075 ( 
.A(n_11880),
.B(n_7358),
.Y(n_12075)
);

OAI221xp5_ASAP7_75t_L g12076 ( 
.A1(n_11955),
.A2(n_11838),
.B1(n_11831),
.B2(n_11876),
.C(n_11781),
.Y(n_12076)
);

INVx2_ASAP7_75t_SL g12077 ( 
.A(n_11900),
.Y(n_12077)
);

AOI222xp33_ASAP7_75t_L g12078 ( 
.A1(n_11904),
.A2(n_11812),
.B1(n_11861),
.B2(n_11820),
.C1(n_11826),
.C2(n_11821),
.Y(n_12078)
);

AOI22xp33_ASAP7_75t_L g12079 ( 
.A1(n_11890),
.A2(n_11846),
.B1(n_11832),
.B2(n_11833),
.Y(n_12079)
);

OAI22xp33_ASAP7_75t_L g12080 ( 
.A1(n_12027),
.A2(n_11900),
.B1(n_11896),
.B2(n_11895),
.Y(n_12080)
);

AOI32xp33_ASAP7_75t_L g12081 ( 
.A1(n_11932),
.A2(n_11817),
.A3(n_11835),
.B1(n_11834),
.B2(n_11864),
.Y(n_12081)
);

INVx1_ASAP7_75t_L g12082 ( 
.A(n_11957),
.Y(n_12082)
);

AOI33xp33_ASAP7_75t_L g12083 ( 
.A1(n_11992),
.A2(n_11718),
.A3(n_11847),
.B1(n_11702),
.B2(n_11815),
.B3(n_11871),
.Y(n_12083)
);

AOI22xp5_ASAP7_75t_L g12084 ( 
.A1(n_11912),
.A2(n_11788),
.B1(n_11799),
.B2(n_11879),
.Y(n_12084)
);

INVx2_ASAP7_75t_L g12085 ( 
.A(n_11888),
.Y(n_12085)
);

NAND2xp5_ASAP7_75t_L g12086 ( 
.A(n_11949),
.B(n_11841),
.Y(n_12086)
);

OA211x2_ASAP7_75t_L g12087 ( 
.A1(n_11916),
.A2(n_11863),
.B(n_11865),
.C(n_11805),
.Y(n_12087)
);

NOR2xp33_ASAP7_75t_L g12088 ( 
.A(n_11902),
.B(n_11899),
.Y(n_12088)
);

AOI322xp5_ASAP7_75t_L g12089 ( 
.A1(n_11940),
.A2(n_11910),
.A3(n_12007),
.B1(n_11936),
.B2(n_11901),
.C1(n_11905),
.C2(n_11906),
.Y(n_12089)
);

AOI21xp5_ASAP7_75t_L g12090 ( 
.A1(n_11930),
.A2(n_11969),
.B(n_11897),
.Y(n_12090)
);

INVx1_ASAP7_75t_L g12091 ( 
.A(n_11943),
.Y(n_12091)
);

AND2x4_ASAP7_75t_L g12092 ( 
.A(n_11894),
.B(n_11868),
.Y(n_12092)
);

INVx1_ASAP7_75t_L g12093 ( 
.A(n_11985),
.Y(n_12093)
);

AOI221xp5_ASAP7_75t_L g12094 ( 
.A1(n_11889),
.A2(n_11884),
.B1(n_11866),
.B2(n_11851),
.C(n_11881),
.Y(n_12094)
);

INVx1_ASAP7_75t_L g12095 ( 
.A(n_11995),
.Y(n_12095)
);

NOR2xp33_ASAP7_75t_L g12096 ( 
.A(n_11911),
.B(n_11755),
.Y(n_12096)
);

OAI31xp33_ASAP7_75t_L g12097 ( 
.A1(n_11954),
.A2(n_11878),
.A3(n_11872),
.B(n_11786),
.Y(n_12097)
);

OR2x2_ASAP7_75t_L g12098 ( 
.A(n_11913),
.B(n_11870),
.Y(n_12098)
);

INVx1_ASAP7_75t_L g12099 ( 
.A(n_11942),
.Y(n_12099)
);

NAND2xp5_ASAP7_75t_L g12100 ( 
.A(n_11956),
.B(n_11875),
.Y(n_12100)
);

NAND2xp5_ASAP7_75t_L g12101 ( 
.A(n_11996),
.B(n_11828),
.Y(n_12101)
);

INVx1_ASAP7_75t_L g12102 ( 
.A(n_11945),
.Y(n_12102)
);

INVx1_ASAP7_75t_L g12103 ( 
.A(n_11893),
.Y(n_12103)
);

NAND2xp5_ASAP7_75t_L g12104 ( 
.A(n_12024),
.B(n_11840),
.Y(n_12104)
);

AOI321xp33_ASAP7_75t_L g12105 ( 
.A1(n_11946),
.A2(n_8085),
.A3(n_8066),
.B1(n_8048),
.B2(n_8049),
.C(n_7131),
.Y(n_12105)
);

INVx1_ASAP7_75t_SL g12106 ( 
.A(n_11892),
.Y(n_12106)
);

NOR2xp33_ASAP7_75t_L g12107 ( 
.A(n_11934),
.B(n_8632),
.Y(n_12107)
);

NAND2xp5_ASAP7_75t_L g12108 ( 
.A(n_12006),
.B(n_8672),
.Y(n_12108)
);

NAND2x1_ASAP7_75t_L g12109 ( 
.A(n_11917),
.B(n_7543),
.Y(n_12109)
);

AOI221xp5_ASAP7_75t_L g12110 ( 
.A1(n_12032),
.A2(n_8672),
.B1(n_7615),
.B2(n_7165),
.C(n_7254),
.Y(n_12110)
);

OR4x1_ASAP7_75t_L g12111 ( 
.A(n_12030),
.B(n_6689),
.C(n_6729),
.D(n_6616),
.Y(n_12111)
);

NAND2xp5_ASAP7_75t_L g12112 ( 
.A(n_11974),
.B(n_8672),
.Y(n_12112)
);

OR2x2_ASAP7_75t_L g12113 ( 
.A(n_11891),
.B(n_7118),
.Y(n_12113)
);

OAI32xp33_ASAP7_75t_L g12114 ( 
.A1(n_11953),
.A2(n_7591),
.A3(n_7262),
.B1(n_7266),
.B2(n_7254),
.Y(n_12114)
);

INVx1_ASAP7_75t_L g12115 ( 
.A(n_11991),
.Y(n_12115)
);

INVx1_ASAP7_75t_L g12116 ( 
.A(n_11998),
.Y(n_12116)
);

OR2x2_ASAP7_75t_L g12117 ( 
.A(n_11928),
.B(n_7101),
.Y(n_12117)
);

NAND2xp5_ASAP7_75t_L g12118 ( 
.A(n_11984),
.B(n_7134),
.Y(n_12118)
);

AOI22xp5_ASAP7_75t_L g12119 ( 
.A1(n_12016),
.A2(n_7543),
.B1(n_6829),
.B2(n_7254),
.Y(n_12119)
);

INVx1_ASAP7_75t_L g12120 ( 
.A(n_12033),
.Y(n_12120)
);

OAI21xp33_ASAP7_75t_L g12121 ( 
.A1(n_11971),
.A2(n_12062),
.B(n_11994),
.Y(n_12121)
);

NAND3xp33_ASAP7_75t_L g12122 ( 
.A(n_12029),
.B(n_6829),
.C(n_7043),
.Y(n_12122)
);

OAI22xp5_ASAP7_75t_L g12123 ( 
.A1(n_11887),
.A2(n_7591),
.B1(n_7525),
.B2(n_7538),
.Y(n_12123)
);

O2A1O1Ixp33_ASAP7_75t_L g12124 ( 
.A1(n_11924),
.A2(n_7047),
.B(n_7255),
.C(n_7043),
.Y(n_12124)
);

AND2x4_ASAP7_75t_L g12125 ( 
.A(n_12021),
.B(n_7512),
.Y(n_12125)
);

INVx1_ASAP7_75t_L g12126 ( 
.A(n_11952),
.Y(n_12126)
);

INVx1_ASAP7_75t_L g12127 ( 
.A(n_11967),
.Y(n_12127)
);

NOR3xp33_ASAP7_75t_L g12128 ( 
.A(n_11947),
.B(n_7132),
.C(n_7117),
.Y(n_12128)
);

A2O1A1Ixp33_ASAP7_75t_L g12129 ( 
.A1(n_11920),
.A2(n_11909),
.B(n_12050),
.C(n_11990),
.Y(n_12129)
);

INVx1_ASAP7_75t_L g12130 ( 
.A(n_11977),
.Y(n_12130)
);

AND2x2_ASAP7_75t_L g12131 ( 
.A(n_12040),
.B(n_7139),
.Y(n_12131)
);

AOI21xp5_ASAP7_75t_L g12132 ( 
.A1(n_11944),
.A2(n_7525),
.B(n_7512),
.Y(n_12132)
);

INVx1_ASAP7_75t_L g12133 ( 
.A(n_11989),
.Y(n_12133)
);

INVx1_ASAP7_75t_L g12134 ( 
.A(n_11925),
.Y(n_12134)
);

INVx1_ASAP7_75t_L g12135 ( 
.A(n_11987),
.Y(n_12135)
);

NAND4xp25_ASAP7_75t_SL g12136 ( 
.A(n_11907),
.B(n_11908),
.C(n_12020),
.D(n_12000),
.Y(n_12136)
);

OAI22xp5_ASAP7_75t_L g12137 ( 
.A1(n_11931),
.A2(n_7525),
.B1(n_7538),
.B2(n_7512),
.Y(n_12137)
);

INVx1_ASAP7_75t_L g12138 ( 
.A(n_12059),
.Y(n_12138)
);

INVx1_ASAP7_75t_L g12139 ( 
.A(n_11980),
.Y(n_12139)
);

HB1xp67_ASAP7_75t_L g12140 ( 
.A(n_11939),
.Y(n_12140)
);

OAI22xp33_ASAP7_75t_L g12141 ( 
.A1(n_11914),
.A2(n_7262),
.B1(n_7266),
.B2(n_7243),
.Y(n_12141)
);

OAI21xp5_ASAP7_75t_SL g12142 ( 
.A1(n_12034),
.A2(n_7255),
.B(n_7047),
.Y(n_12142)
);

NAND3xp33_ASAP7_75t_L g12143 ( 
.A(n_11915),
.B(n_7043),
.C(n_7063),
.Y(n_12143)
);

AOI22xp5_ASAP7_75t_L g12144 ( 
.A1(n_11972),
.A2(n_7262),
.B1(n_7266),
.B2(n_7243),
.Y(n_12144)
);

NAND2xp5_ASAP7_75t_SL g12145 ( 
.A(n_11997),
.B(n_6889),
.Y(n_12145)
);

AND2x4_ASAP7_75t_L g12146 ( 
.A(n_12064),
.B(n_7538),
.Y(n_12146)
);

O2A1O1Ixp33_ASAP7_75t_L g12147 ( 
.A1(n_11938),
.A2(n_7255),
.B(n_7047),
.C(n_7063),
.Y(n_12147)
);

INVx2_ASAP7_75t_L g12148 ( 
.A(n_12057),
.Y(n_12148)
);

AND2x2_ASAP7_75t_L g12149 ( 
.A(n_12019),
.B(n_12011),
.Y(n_12149)
);

OAI22xp5_ASAP7_75t_L g12150 ( 
.A1(n_11966),
.A2(n_7586),
.B1(n_7588),
.B2(n_7548),
.Y(n_12150)
);

BUFx3_ASAP7_75t_L g12151 ( 
.A(n_11975),
.Y(n_12151)
);

AOI22xp5_ASAP7_75t_L g12152 ( 
.A1(n_11960),
.A2(n_7313),
.B1(n_7315),
.B2(n_7278),
.Y(n_12152)
);

NAND2xp5_ASAP7_75t_L g12153 ( 
.A(n_12057),
.B(n_7134),
.Y(n_12153)
);

NAND2xp5_ASAP7_75t_L g12154 ( 
.A(n_12018),
.B(n_7134),
.Y(n_12154)
);

INVx1_ASAP7_75t_L g12155 ( 
.A(n_12061),
.Y(n_12155)
);

INVx2_ASAP7_75t_SL g12156 ( 
.A(n_12063),
.Y(n_12156)
);

AOI221xp5_ASAP7_75t_L g12157 ( 
.A1(n_12060),
.A2(n_7165),
.B1(n_7313),
.B2(n_7315),
.C(n_7278),
.Y(n_12157)
);

AND2x2_ASAP7_75t_L g12158 ( 
.A(n_11898),
.B(n_11970),
.Y(n_12158)
);

AND2x2_ASAP7_75t_L g12159 ( 
.A(n_11918),
.B(n_7149),
.Y(n_12159)
);

AND2x2_ASAP7_75t_L g12160 ( 
.A(n_11927),
.B(n_7134),
.Y(n_12160)
);

INVx1_ASAP7_75t_L g12161 ( 
.A(n_11961),
.Y(n_12161)
);

NAND2xp5_ASAP7_75t_L g12162 ( 
.A(n_12045),
.B(n_12014),
.Y(n_12162)
);

AOI22xp33_ASAP7_75t_L g12163 ( 
.A1(n_12001),
.A2(n_7276),
.B1(n_7328),
.B2(n_7165),
.Y(n_12163)
);

AOI21xp5_ASAP7_75t_L g12164 ( 
.A1(n_11933),
.A2(n_7586),
.B(n_7548),
.Y(n_12164)
);

NOR2xp33_ASAP7_75t_L g12165 ( 
.A(n_12069),
.B(n_7103),
.Y(n_12165)
);

O2A1O1Ixp33_ASAP7_75t_L g12166 ( 
.A1(n_11958),
.A2(n_7063),
.B(n_7064),
.C(n_7278),
.Y(n_12166)
);

AND2x2_ASAP7_75t_L g12167 ( 
.A(n_11963),
.B(n_7134),
.Y(n_12167)
);

INVx2_ASAP7_75t_L g12168 ( 
.A(n_11922),
.Y(n_12168)
);

INVx1_ASAP7_75t_L g12169 ( 
.A(n_12048),
.Y(n_12169)
);

INVx1_ASAP7_75t_L g12170 ( 
.A(n_12049),
.Y(n_12170)
);

AOI22xp5_ASAP7_75t_L g12171 ( 
.A1(n_12010),
.A2(n_11937),
.B1(n_11941),
.B2(n_11923),
.Y(n_12171)
);

INVx1_ASAP7_75t_L g12172 ( 
.A(n_11973),
.Y(n_12172)
);

AOI21xp5_ASAP7_75t_L g12173 ( 
.A1(n_11982),
.A2(n_7588),
.B(n_7586),
.Y(n_12173)
);

NAND2xp5_ASAP7_75t_L g12174 ( 
.A(n_12073),
.B(n_7134),
.Y(n_12174)
);

AND2x2_ASAP7_75t_L g12175 ( 
.A(n_12025),
.B(n_7176),
.Y(n_12175)
);

OAI21xp33_ASAP7_75t_L g12176 ( 
.A1(n_11950),
.A2(n_7315),
.B(n_7313),
.Y(n_12176)
);

NOR2xp33_ASAP7_75t_L g12177 ( 
.A(n_12041),
.B(n_7155),
.Y(n_12177)
);

XNOR2x2_ASAP7_75t_L g12178 ( 
.A(n_12012),
.B(n_7133),
.Y(n_12178)
);

OAI21xp5_ASAP7_75t_L g12179 ( 
.A1(n_11903),
.A2(n_7135),
.B(n_7133),
.Y(n_12179)
);

XOR2x2_ASAP7_75t_L g12180 ( 
.A(n_12039),
.B(n_7000),
.Y(n_12180)
);

OAI21xp5_ASAP7_75t_L g12181 ( 
.A1(n_11951),
.A2(n_7137),
.B(n_7135),
.Y(n_12181)
);

NAND2xp5_ASAP7_75t_L g12182 ( 
.A(n_12047),
.B(n_7358),
.Y(n_12182)
);

XNOR2xp5_ASAP7_75t_L g12183 ( 
.A(n_12051),
.B(n_7000),
.Y(n_12183)
);

AND2x2_ASAP7_75t_L g12184 ( 
.A(n_12056),
.B(n_7176),
.Y(n_12184)
);

AND2x2_ASAP7_75t_L g12185 ( 
.A(n_12068),
.B(n_7176),
.Y(n_12185)
);

AOI221xp5_ASAP7_75t_L g12186 ( 
.A1(n_12067),
.A2(n_7431),
.B1(n_7449),
.B2(n_7357),
.C(n_7316),
.Y(n_12186)
);

NAND2xp5_ASAP7_75t_L g12187 ( 
.A(n_11993),
.B(n_7146),
.Y(n_12187)
);

NAND2xp5_ASAP7_75t_L g12188 ( 
.A(n_12015),
.B(n_7147),
.Y(n_12188)
);

OAI21xp33_ASAP7_75t_L g12189 ( 
.A1(n_12037),
.A2(n_7357),
.B(n_7316),
.Y(n_12189)
);

INVx1_ASAP7_75t_SL g12190 ( 
.A(n_12036),
.Y(n_12190)
);

A2O1A1Ixp33_ASAP7_75t_L g12191 ( 
.A1(n_11999),
.A2(n_7137),
.B(n_7183),
.C(n_7179),
.Y(n_12191)
);

OAI22xp5_ASAP7_75t_L g12192 ( 
.A1(n_11921),
.A2(n_7588),
.B1(n_7590),
.B2(n_7548),
.Y(n_12192)
);

INVx1_ASAP7_75t_L g12193 ( 
.A(n_11962),
.Y(n_12193)
);

AND2x2_ASAP7_75t_L g12194 ( 
.A(n_12046),
.B(n_7176),
.Y(n_12194)
);

O2A1O1Ixp33_ASAP7_75t_L g12195 ( 
.A1(n_12005),
.A2(n_7064),
.B(n_7357),
.C(n_7316),
.Y(n_12195)
);

AOI22xp5_ASAP7_75t_L g12196 ( 
.A1(n_11959),
.A2(n_7449),
.B1(n_7487),
.B2(n_7431),
.Y(n_12196)
);

AOI21xp5_ASAP7_75t_L g12197 ( 
.A1(n_12013),
.A2(n_7621),
.B(n_7590),
.Y(n_12197)
);

OAI33xp33_ASAP7_75t_L g12198 ( 
.A1(n_12042),
.A2(n_6970),
.A3(n_6964),
.B1(n_6987),
.B2(n_6971),
.B3(n_6913),
.Y(n_12198)
);

INVx1_ASAP7_75t_L g12199 ( 
.A(n_12017),
.Y(n_12199)
);

INVxp67_ASAP7_75t_L g12200 ( 
.A(n_12071),
.Y(n_12200)
);

AOI22xp33_ASAP7_75t_L g12201 ( 
.A1(n_11976),
.A2(n_7276),
.B1(n_7328),
.B2(n_7064),
.Y(n_12201)
);

NAND3xp33_ASAP7_75t_L g12202 ( 
.A(n_11983),
.B(n_7064),
.C(n_7276),
.Y(n_12202)
);

NOR2xp33_ASAP7_75t_L g12203 ( 
.A(n_12003),
.B(n_12002),
.Y(n_12203)
);

INVx2_ASAP7_75t_L g12204 ( 
.A(n_11964),
.Y(n_12204)
);

NAND2xp5_ASAP7_75t_L g12205 ( 
.A(n_12023),
.B(n_7147),
.Y(n_12205)
);

NOR2xp33_ASAP7_75t_L g12206 ( 
.A(n_12022),
.B(n_7164),
.Y(n_12206)
);

OAI21xp33_ASAP7_75t_SL g12207 ( 
.A1(n_11978),
.A2(n_7183),
.B(n_7179),
.Y(n_12207)
);

INVx2_ASAP7_75t_L g12208 ( 
.A(n_11964),
.Y(n_12208)
);

NAND2xp5_ASAP7_75t_L g12209 ( 
.A(n_12075),
.B(n_7156),
.Y(n_12209)
);

INVx1_ASAP7_75t_L g12210 ( 
.A(n_11919),
.Y(n_12210)
);

NAND2xp5_ASAP7_75t_L g12211 ( 
.A(n_12066),
.B(n_7156),
.Y(n_12211)
);

INVx1_ASAP7_75t_L g12212 ( 
.A(n_11926),
.Y(n_12212)
);

AOI221xp5_ASAP7_75t_L g12213 ( 
.A1(n_11979),
.A2(n_7487),
.B1(n_7449),
.B2(n_7431),
.C(n_6964),
.Y(n_12213)
);

NAND2xp33_ASAP7_75t_L g12214 ( 
.A(n_12054),
.B(n_7590),
.Y(n_12214)
);

AOI311xp33_ASAP7_75t_L g12215 ( 
.A1(n_12053),
.A2(n_7629),
.A3(n_7166),
.B(n_7182),
.C(n_7161),
.Y(n_12215)
);

INVx1_ASAP7_75t_L g12216 ( 
.A(n_12026),
.Y(n_12216)
);

AOI221xp5_ASAP7_75t_L g12217 ( 
.A1(n_11929),
.A2(n_7487),
.B1(n_6970),
.B2(n_6987),
.C(n_6971),
.Y(n_12217)
);

INVx1_ASAP7_75t_L g12218 ( 
.A(n_12052),
.Y(n_12218)
);

HB1xp67_ASAP7_75t_L g12219 ( 
.A(n_12052),
.Y(n_12219)
);

NAND2xp5_ASAP7_75t_L g12220 ( 
.A(n_11986),
.B(n_7158),
.Y(n_12220)
);

OAI21xp33_ASAP7_75t_L g12221 ( 
.A1(n_12072),
.A2(n_6990),
.B(n_6970),
.Y(n_12221)
);

NOR2x1_ASAP7_75t_L g12222 ( 
.A(n_11988),
.B(n_6913),
.Y(n_12222)
);

INVx1_ASAP7_75t_L g12223 ( 
.A(n_11988),
.Y(n_12223)
);

OAI22xp5_ASAP7_75t_L g12224 ( 
.A1(n_12009),
.A2(n_7623),
.B1(n_7621),
.B2(n_6971),
.Y(n_12224)
);

NAND2xp33_ASAP7_75t_L g12225 ( 
.A(n_11965),
.B(n_7621),
.Y(n_12225)
);

INVx2_ASAP7_75t_L g12226 ( 
.A(n_12070),
.Y(n_12226)
);

NAND3xp33_ASAP7_75t_L g12227 ( 
.A(n_11948),
.B(n_7276),
.C(n_7153),
.Y(n_12227)
);

AOI22xp5_ASAP7_75t_L g12228 ( 
.A1(n_12058),
.A2(n_12055),
.B1(n_12004),
.B2(n_12008),
.Y(n_12228)
);

INVx1_ASAP7_75t_L g12229 ( 
.A(n_11981),
.Y(n_12229)
);

AOI31xp33_ASAP7_75t_L g12230 ( 
.A1(n_11968),
.A2(n_6958),
.A3(n_6689),
.B(n_6729),
.Y(n_12230)
);

INVxp67_ASAP7_75t_L g12231 ( 
.A(n_12038),
.Y(n_12231)
);

NAND2xp5_ASAP7_75t_L g12232 ( 
.A(n_12044),
.B(n_7158),
.Y(n_12232)
);

AND2x2_ASAP7_75t_L g12233 ( 
.A(n_12031),
.B(n_7176),
.Y(n_12233)
);

NAND2xp5_ASAP7_75t_L g12234 ( 
.A(n_12035),
.B(n_7161),
.Y(n_12234)
);

INVx1_ASAP7_75t_L g12235 ( 
.A(n_12077),
.Y(n_12235)
);

INVx1_ASAP7_75t_L g12236 ( 
.A(n_12095),
.Y(n_12236)
);

INVx2_ASAP7_75t_SL g12237 ( 
.A(n_12092),
.Y(n_12237)
);

AND2x2_ASAP7_75t_L g12238 ( 
.A(n_12156),
.B(n_12028),
.Y(n_12238)
);

INVx1_ASAP7_75t_L g12239 ( 
.A(n_12219),
.Y(n_12239)
);

AOI222xp33_ASAP7_75t_L g12240 ( 
.A1(n_12110),
.A2(n_12043),
.B1(n_11935),
.B2(n_12065),
.C1(n_12074),
.C2(n_6987),
.Y(n_12240)
);

NOR2xp33_ASAP7_75t_L g12241 ( 
.A(n_12106),
.B(n_7623),
.Y(n_12241)
);

INVx2_ASAP7_75t_L g12242 ( 
.A(n_12092),
.Y(n_12242)
);

INVx2_ASAP7_75t_L g12243 ( 
.A(n_12151),
.Y(n_12243)
);

INVx1_ASAP7_75t_SL g12244 ( 
.A(n_12158),
.Y(n_12244)
);

INVx1_ASAP7_75t_L g12245 ( 
.A(n_12082),
.Y(n_12245)
);

INVx1_ASAP7_75t_L g12246 ( 
.A(n_12086),
.Y(n_12246)
);

INVx2_ASAP7_75t_L g12247 ( 
.A(n_12148),
.Y(n_12247)
);

OR2x2_ASAP7_75t_L g12248 ( 
.A(n_12091),
.B(n_6913),
.Y(n_12248)
);

INVxp67_ASAP7_75t_L g12249 ( 
.A(n_12096),
.Y(n_12249)
);

OAI21xp33_ASAP7_75t_SL g12250 ( 
.A1(n_12097),
.A2(n_7188),
.B(n_7185),
.Y(n_12250)
);

INVx1_ASAP7_75t_L g12251 ( 
.A(n_12093),
.Y(n_12251)
);

NAND2xp5_ASAP7_75t_L g12252 ( 
.A(n_12085),
.B(n_7176),
.Y(n_12252)
);

AOI21xp33_ASAP7_75t_L g12253 ( 
.A1(n_12088),
.A2(n_12080),
.B(n_12078),
.Y(n_12253)
);

INVx1_ASAP7_75t_L g12254 ( 
.A(n_12149),
.Y(n_12254)
);

INVx1_ASAP7_75t_L g12255 ( 
.A(n_12115),
.Y(n_12255)
);

NOR2xp33_ASAP7_75t_L g12256 ( 
.A(n_12126),
.B(n_7623),
.Y(n_12256)
);

INVx1_ASAP7_75t_L g12257 ( 
.A(n_12127),
.Y(n_12257)
);

INVx1_ASAP7_75t_SL g12258 ( 
.A(n_12098),
.Y(n_12258)
);

AOI211x1_ASAP7_75t_L g12259 ( 
.A1(n_12090),
.A2(n_7182),
.B(n_7184),
.C(n_7166),
.Y(n_12259)
);

NOR4xp25_ASAP7_75t_L g12260 ( 
.A(n_12136),
.B(n_6990),
.C(n_6997),
.D(n_6992),
.Y(n_12260)
);

INVx1_ASAP7_75t_L g12261 ( 
.A(n_12130),
.Y(n_12261)
);

OAI21xp33_ASAP7_75t_L g12262 ( 
.A1(n_12089),
.A2(n_6992),
.B(n_6990),
.Y(n_12262)
);

INVx1_ASAP7_75t_L g12263 ( 
.A(n_12133),
.Y(n_12263)
);

INVxp67_ASAP7_75t_L g12264 ( 
.A(n_12134),
.Y(n_12264)
);

INVx1_ASAP7_75t_L g12265 ( 
.A(n_12099),
.Y(n_12265)
);

INVx1_ASAP7_75t_L g12266 ( 
.A(n_12102),
.Y(n_12266)
);

INVx1_ASAP7_75t_L g12267 ( 
.A(n_12113),
.Y(n_12267)
);

NAND2xp5_ASAP7_75t_L g12268 ( 
.A(n_12116),
.B(n_7116),
.Y(n_12268)
);

OAI22xp5_ASAP7_75t_L g12269 ( 
.A1(n_12079),
.A2(n_6992),
.B1(n_7023),
.B2(n_6997),
.Y(n_12269)
);

INVx2_ASAP7_75t_L g12270 ( 
.A(n_12111),
.Y(n_12270)
);

INVxp67_ASAP7_75t_L g12271 ( 
.A(n_12100),
.Y(n_12271)
);

AND2x2_ASAP7_75t_L g12272 ( 
.A(n_12159),
.B(n_12120),
.Y(n_12272)
);

NAND2xp5_ASAP7_75t_L g12273 ( 
.A(n_12155),
.B(n_7116),
.Y(n_12273)
);

NAND2x1_ASAP7_75t_L g12274 ( 
.A(n_12125),
.B(n_6997),
.Y(n_12274)
);

INVxp33_ASAP7_75t_L g12275 ( 
.A(n_12162),
.Y(n_12275)
);

A2O1A1Ixp33_ASAP7_75t_L g12276 ( 
.A1(n_12081),
.A2(n_7185),
.B(n_7202),
.C(n_7188),
.Y(n_12276)
);

AOI21xp33_ASAP7_75t_L g12277 ( 
.A1(n_12138),
.A2(n_7153),
.B(n_7067),
.Y(n_12277)
);

INVx1_ASAP7_75t_L g12278 ( 
.A(n_12216),
.Y(n_12278)
);

INVx2_ASAP7_75t_L g12279 ( 
.A(n_12178),
.Y(n_12279)
);

INVx1_ASAP7_75t_L g12280 ( 
.A(n_12139),
.Y(n_12280)
);

INVx1_ASAP7_75t_L g12281 ( 
.A(n_12135),
.Y(n_12281)
);

AND2x2_ASAP7_75t_L g12282 ( 
.A(n_12165),
.B(n_7202),
.Y(n_12282)
);

NOR2xp33_ASAP7_75t_L g12283 ( 
.A(n_12076),
.B(n_7023),
.Y(n_12283)
);

AOI31xp33_ASAP7_75t_SL g12284 ( 
.A1(n_12094),
.A2(n_7023),
.A3(n_7089),
.B(n_6921),
.Y(n_12284)
);

INVx1_ASAP7_75t_L g12285 ( 
.A(n_12204),
.Y(n_12285)
);

AOI221xp5_ASAP7_75t_L g12286 ( 
.A1(n_12212),
.A2(n_7203),
.B1(n_7206),
.B2(n_7175),
.C(n_7196),
.Y(n_12286)
);

INVx1_ASAP7_75t_L g12287 ( 
.A(n_12208),
.Y(n_12287)
);

INVx1_ASAP7_75t_SL g12288 ( 
.A(n_12101),
.Y(n_12288)
);

OAI21xp5_ASAP7_75t_SL g12289 ( 
.A1(n_12171),
.A2(n_6958),
.B(n_6742),
.Y(n_12289)
);

HB1xp67_ASAP7_75t_L g12290 ( 
.A(n_12125),
.Y(n_12290)
);

OAI22xp5_ASAP7_75t_L g12291 ( 
.A1(n_12119),
.A2(n_7089),
.B1(n_7109),
.B2(n_6921),
.Y(n_12291)
);

AOI322xp5_ASAP7_75t_L g12292 ( 
.A1(n_12103),
.A2(n_6770),
.A3(n_6689),
.B1(n_6729),
.B2(n_6616),
.C1(n_7187),
.C2(n_7109),
.Y(n_12292)
);

NAND2xp5_ASAP7_75t_L g12293 ( 
.A(n_12168),
.B(n_7116),
.Y(n_12293)
);

AOI222xp33_ASAP7_75t_L g12294 ( 
.A1(n_12207),
.A2(n_7042),
.B1(n_7184),
.B2(n_7194),
.C1(n_7189),
.C2(n_7186),
.Y(n_12294)
);

NOR2xp33_ASAP7_75t_L g12295 ( 
.A(n_12161),
.B(n_7212),
.Y(n_12295)
);

AND2x2_ASAP7_75t_L g12296 ( 
.A(n_12131),
.B(n_7212),
.Y(n_12296)
);

AOI221xp5_ASAP7_75t_L g12297 ( 
.A1(n_12121),
.A2(n_7175),
.B1(n_7206),
.B2(n_7203),
.C(n_7602),
.Y(n_12297)
);

NOR2xp33_ASAP7_75t_L g12298 ( 
.A(n_12169),
.B(n_7217),
.Y(n_12298)
);

NOR2xp33_ASAP7_75t_SL g12299 ( 
.A(n_12210),
.B(n_12170),
.Y(n_12299)
);

INVxp67_ASAP7_75t_L g12300 ( 
.A(n_12104),
.Y(n_12300)
);

AND2x2_ASAP7_75t_L g12301 ( 
.A(n_12177),
.B(n_7217),
.Y(n_12301)
);

INVx1_ASAP7_75t_L g12302 ( 
.A(n_12218),
.Y(n_12302)
);

OAI22xp5_ASAP7_75t_L g12303 ( 
.A1(n_12228),
.A2(n_7191),
.B1(n_7196),
.B2(n_7187),
.Y(n_12303)
);

AOI22xp33_ASAP7_75t_L g12304 ( 
.A1(n_12087),
.A2(n_7203),
.B1(n_7206),
.B2(n_7175),
.Y(n_12304)
);

INVx1_ASAP7_75t_L g12305 ( 
.A(n_12083),
.Y(n_12305)
);

NAND2xp5_ASAP7_75t_L g12306 ( 
.A(n_12146),
.B(n_7116),
.Y(n_12306)
);

OR2x2_ASAP7_75t_L g12307 ( 
.A(n_12117),
.B(n_7567),
.Y(n_12307)
);

INVx1_ASAP7_75t_SL g12308 ( 
.A(n_12146),
.Y(n_12308)
);

AOI221x1_ASAP7_75t_L g12309 ( 
.A1(n_12129),
.A2(n_7292),
.B1(n_7596),
.B2(n_7592),
.C(n_7191),
.Y(n_12309)
);

INVx1_ASAP7_75t_L g12310 ( 
.A(n_12223),
.Y(n_12310)
);

INVx1_ASAP7_75t_L g12311 ( 
.A(n_12108),
.Y(n_12311)
);

INVx2_ASAP7_75t_L g12312 ( 
.A(n_12109),
.Y(n_12312)
);

INVx1_ASAP7_75t_L g12313 ( 
.A(n_12112),
.Y(n_12313)
);

AOI22xp33_ASAP7_75t_SL g12314 ( 
.A1(n_12175),
.A2(n_7218),
.B1(n_7220),
.B2(n_7219),
.Y(n_12314)
);

INVx1_ASAP7_75t_L g12315 ( 
.A(n_12229),
.Y(n_12315)
);

INVx1_ASAP7_75t_L g12316 ( 
.A(n_12140),
.Y(n_12316)
);

INVxp67_ASAP7_75t_L g12317 ( 
.A(n_12203),
.Y(n_12317)
);

NOR2xp33_ASAP7_75t_L g12318 ( 
.A(n_12084),
.B(n_7218),
.Y(n_12318)
);

INVx1_ASAP7_75t_L g12319 ( 
.A(n_12226),
.Y(n_12319)
);

INVx1_ASAP7_75t_L g12320 ( 
.A(n_12107),
.Y(n_12320)
);

INVx3_ASAP7_75t_L g12321 ( 
.A(n_12160),
.Y(n_12321)
);

AOI221xp5_ASAP7_75t_L g12322 ( 
.A1(n_12231),
.A2(n_7592),
.B1(n_7602),
.B2(n_7596),
.C(n_7292),
.Y(n_12322)
);

AND2x4_ASAP7_75t_L g12323 ( 
.A(n_12199),
.B(n_7219),
.Y(n_12323)
);

OAI221xp5_ASAP7_75t_L g12324 ( 
.A1(n_12176),
.A2(n_6958),
.B1(n_7000),
.B2(n_6770),
.C(n_6616),
.Y(n_12324)
);

INVx1_ASAP7_75t_L g12325 ( 
.A(n_12187),
.Y(n_12325)
);

INVx3_ASAP7_75t_L g12326 ( 
.A(n_12167),
.Y(n_12326)
);

AO22x2_ASAP7_75t_L g12327 ( 
.A1(n_12193),
.A2(n_7224),
.B1(n_6568),
.B2(n_6530),
.Y(n_12327)
);

INVx1_ASAP7_75t_L g12328 ( 
.A(n_12145),
.Y(n_12328)
);

NAND2xp5_ASAP7_75t_SL g12329 ( 
.A(n_12122),
.B(n_12153),
.Y(n_12329)
);

NAND2xp5_ASAP7_75t_SL g12330 ( 
.A(n_12183),
.B(n_7220),
.Y(n_12330)
);

INVx1_ASAP7_75t_L g12331 ( 
.A(n_12118),
.Y(n_12331)
);

OR2x2_ASAP7_75t_L g12332 ( 
.A(n_12154),
.B(n_7567),
.Y(n_12332)
);

OAI21xp5_ASAP7_75t_L g12333 ( 
.A1(n_12174),
.A2(n_7237),
.B(n_7222),
.Y(n_12333)
);

AOI221xp5_ASAP7_75t_L g12334 ( 
.A1(n_12206),
.A2(n_7224),
.B1(n_7194),
.B2(n_7195),
.C(n_7189),
.Y(n_12334)
);

OAI221xp5_ASAP7_75t_SL g12335 ( 
.A1(n_12190),
.A2(n_12182),
.B1(n_12142),
.B2(n_12232),
.C(n_12191),
.Y(n_12335)
);

NAND2xp33_ASAP7_75t_L g12336 ( 
.A(n_12222),
.B(n_7186),
.Y(n_12336)
);

AND2x2_ASAP7_75t_L g12337 ( 
.A(n_12185),
.B(n_7222),
.Y(n_12337)
);

OAI211xp5_ASAP7_75t_L g12338 ( 
.A1(n_12200),
.A2(n_7247),
.B(n_7253),
.C(n_7237),
.Y(n_12338)
);

OAI22xp5_ASAP7_75t_L g12339 ( 
.A1(n_12144),
.A2(n_6770),
.B1(n_7199),
.B2(n_7195),
.Y(n_12339)
);

NAND2xp5_ASAP7_75t_L g12340 ( 
.A(n_12184),
.B(n_7116),
.Y(n_12340)
);

NAND2x1p5_ASAP7_75t_L g12341 ( 
.A(n_12172),
.B(n_7247),
.Y(n_12341)
);

INVx1_ASAP7_75t_L g12342 ( 
.A(n_12188),
.Y(n_12342)
);

OAI22xp5_ASAP7_75t_L g12343 ( 
.A1(n_12152),
.A2(n_7208),
.B1(n_7213),
.B2(n_7199),
.Y(n_12343)
);

NAND3xp33_ASAP7_75t_L g12344 ( 
.A(n_12225),
.B(n_7153),
.C(n_7067),
.Y(n_12344)
);

AOI211xp5_ASAP7_75t_L g12345 ( 
.A1(n_12137),
.A2(n_7259),
.B(n_7283),
.C(n_7253),
.Y(n_12345)
);

A2O1A1Ixp33_ASAP7_75t_L g12346 ( 
.A1(n_12234),
.A2(n_12230),
.B(n_12220),
.C(n_12233),
.Y(n_12346)
);

AOI221xp5_ASAP7_75t_L g12347 ( 
.A1(n_12123),
.A2(n_7208),
.B1(n_7232),
.B2(n_7225),
.C(n_7213),
.Y(n_12347)
);

INVx1_ASAP7_75t_L g12348 ( 
.A(n_12205),
.Y(n_12348)
);

A2O1A1Ixp33_ASAP7_75t_L g12349 ( 
.A1(n_12209),
.A2(n_12194),
.B(n_12211),
.C(n_12214),
.Y(n_12349)
);

NAND2xp5_ASAP7_75t_SL g12350 ( 
.A(n_12141),
.B(n_7259),
.Y(n_12350)
);

NAND2xp5_ASAP7_75t_L g12351 ( 
.A(n_12180),
.B(n_7116),
.Y(n_12351)
);

INVx1_ASAP7_75t_L g12352 ( 
.A(n_12196),
.Y(n_12352)
);

INVxp67_ASAP7_75t_L g12353 ( 
.A(n_12198),
.Y(n_12353)
);

INVx2_ASAP7_75t_SL g12354 ( 
.A(n_12150),
.Y(n_12354)
);

NAND2xp5_ASAP7_75t_L g12355 ( 
.A(n_12189),
.B(n_7225),
.Y(n_12355)
);

INVxp67_ASAP7_75t_SL g12356 ( 
.A(n_12132),
.Y(n_12356)
);

INVx1_ASAP7_75t_L g12357 ( 
.A(n_12114),
.Y(n_12357)
);

NAND2xp5_ASAP7_75t_L g12358 ( 
.A(n_12179),
.B(n_12181),
.Y(n_12358)
);

INVx1_ASAP7_75t_L g12359 ( 
.A(n_12221),
.Y(n_12359)
);

AND2x2_ASAP7_75t_L g12360 ( 
.A(n_12215),
.B(n_12128),
.Y(n_12360)
);

OAI22xp5_ASAP7_75t_L g12361 ( 
.A1(n_12186),
.A2(n_7236),
.B1(n_7240),
.B2(n_7232),
.Y(n_12361)
);

OAI22xp5_ASAP7_75t_L g12362 ( 
.A1(n_12157),
.A2(n_7240),
.B1(n_7245),
.B2(n_7236),
.Y(n_12362)
);

AOI22xp5_ASAP7_75t_L g12363 ( 
.A1(n_12192),
.A2(n_7283),
.B1(n_6742),
.B2(n_6659),
.Y(n_12363)
);

OAI21xp33_ASAP7_75t_L g12364 ( 
.A1(n_12173),
.A2(n_6742),
.B(n_6659),
.Y(n_12364)
);

AOI221xp5_ASAP7_75t_L g12365 ( 
.A1(n_12197),
.A2(n_7245),
.B1(n_7260),
.B2(n_7248),
.C(n_7246),
.Y(n_12365)
);

AOI22xp5_ASAP7_75t_L g12366 ( 
.A1(n_12224),
.A2(n_6742),
.B1(n_6659),
.B2(n_7067),
.Y(n_12366)
);

INVx2_ASAP7_75t_L g12367 ( 
.A(n_12143),
.Y(n_12367)
);

AOI222xp33_ASAP7_75t_L g12368 ( 
.A1(n_12202),
.A2(n_7246),
.B1(n_7248),
.B2(n_7264),
.C1(n_7263),
.C2(n_7260),
.Y(n_12368)
);

HB1xp67_ASAP7_75t_L g12369 ( 
.A(n_12164),
.Y(n_12369)
);

INVx1_ASAP7_75t_L g12370 ( 
.A(n_12105),
.Y(n_12370)
);

OAI22xp33_ASAP7_75t_SL g12371 ( 
.A1(n_12147),
.A2(n_12217),
.B1(n_12195),
.B2(n_12227),
.Y(n_12371)
);

AOI32xp33_ASAP7_75t_L g12372 ( 
.A1(n_12213),
.A2(n_7407),
.A3(n_7482),
.B1(n_7480),
.B2(n_7389),
.Y(n_12372)
);

OR2x2_ASAP7_75t_L g12373 ( 
.A(n_12163),
.B(n_7567),
.Y(n_12373)
);

AND2x2_ASAP7_75t_L g12374 ( 
.A(n_12201),
.B(n_7198),
.Y(n_12374)
);

OAI22xp5_ASAP7_75t_L g12375 ( 
.A1(n_12124),
.A2(n_7264),
.B1(n_7265),
.B2(n_7263),
.Y(n_12375)
);

AOI22x1_ASAP7_75t_L g12376 ( 
.A1(n_12166),
.A2(n_7267),
.B1(n_7270),
.B2(n_7265),
.Y(n_12376)
);

INVx2_ASAP7_75t_L g12377 ( 
.A(n_12077),
.Y(n_12377)
);

INVxp67_ASAP7_75t_SL g12378 ( 
.A(n_12080),
.Y(n_12378)
);

AOI221xp5_ASAP7_75t_L g12379 ( 
.A1(n_12253),
.A2(n_7267),
.B1(n_7274),
.B2(n_7272),
.C(n_7270),
.Y(n_12379)
);

OAI322xp33_ASAP7_75t_L g12380 ( 
.A1(n_12299),
.A2(n_12353),
.A3(n_12264),
.B1(n_12244),
.B2(n_12239),
.C1(n_12305),
.C2(n_12278),
.Y(n_12380)
);

AOI322xp5_ASAP7_75t_L g12381 ( 
.A1(n_12378),
.A2(n_6530),
.A3(n_6545),
.B1(n_6537),
.B2(n_6568),
.C1(n_6567),
.C2(n_6529),
.Y(n_12381)
);

INVx1_ASAP7_75t_L g12382 ( 
.A(n_12290),
.Y(n_12382)
);

NAND2xp5_ASAP7_75t_SL g12383 ( 
.A(n_12237),
.B(n_7272),
.Y(n_12383)
);

INVx1_ASAP7_75t_L g12384 ( 
.A(n_12242),
.Y(n_12384)
);

O2A1O1Ixp33_ASAP7_75t_L g12385 ( 
.A1(n_12279),
.A2(n_7277),
.B(n_7285),
.C(n_7274),
.Y(n_12385)
);

INVx2_ASAP7_75t_L g12386 ( 
.A(n_12377),
.Y(n_12386)
);

AOI211xp5_ASAP7_75t_SL g12387 ( 
.A1(n_12271),
.A2(n_6742),
.B(n_6659),
.C(n_7277),
.Y(n_12387)
);

NAND2xp5_ASAP7_75t_L g12388 ( 
.A(n_12254),
.B(n_7198),
.Y(n_12388)
);

AOI22xp5_ASAP7_75t_L g12389 ( 
.A1(n_12258),
.A2(n_12235),
.B1(n_12288),
.B2(n_12236),
.Y(n_12389)
);

INVx4_ASAP7_75t_L g12390 ( 
.A(n_12243),
.Y(n_12390)
);

AOI221xp5_ASAP7_75t_L g12391 ( 
.A1(n_12262),
.A2(n_7286),
.B1(n_7301),
.B2(n_7298),
.C(n_7285),
.Y(n_12391)
);

O2A1O1Ixp5_ASAP7_75t_L g12392 ( 
.A1(n_12329),
.A2(n_7298),
.B(n_7301),
.C(n_7286),
.Y(n_12392)
);

O2A1O1Ixp33_ASAP7_75t_SL g12393 ( 
.A1(n_12346),
.A2(n_7351),
.B(n_7361),
.C(n_7306),
.Y(n_12393)
);

INVx1_ASAP7_75t_L g12394 ( 
.A(n_12272),
.Y(n_12394)
);

O2A1O1Ixp33_ASAP7_75t_SL g12395 ( 
.A1(n_12308),
.A2(n_7351),
.B(n_7361),
.C(n_7306),
.Y(n_12395)
);

AOI22xp5_ASAP7_75t_L g12396 ( 
.A1(n_12238),
.A2(n_12255),
.B1(n_12247),
.B2(n_12246),
.Y(n_12396)
);

AOI211xp5_ASAP7_75t_SL g12397 ( 
.A1(n_12249),
.A2(n_6659),
.B(n_7364),
.C(n_7362),
.Y(n_12397)
);

OAI22xp33_ASAP7_75t_L g12398 ( 
.A1(n_12275),
.A2(n_7364),
.B1(n_7365),
.B2(n_7362),
.Y(n_12398)
);

AND2x2_ASAP7_75t_L g12399 ( 
.A(n_12251),
.B(n_7198),
.Y(n_12399)
);

OAI221xp5_ASAP7_75t_L g12400 ( 
.A1(n_12250),
.A2(n_7365),
.B1(n_7377),
.B2(n_7375),
.C(n_7367),
.Y(n_12400)
);

O2A1O1Ixp33_ASAP7_75t_L g12401 ( 
.A1(n_12312),
.A2(n_7375),
.B(n_7377),
.C(n_7367),
.Y(n_12401)
);

OAI32xp33_ASAP7_75t_L g12402 ( 
.A1(n_12315),
.A2(n_7595),
.A3(n_7398),
.B1(n_7405),
.B2(n_7391),
.Y(n_12402)
);

AOI322xp5_ASAP7_75t_L g12403 ( 
.A1(n_12370),
.A2(n_6530),
.A3(n_6545),
.B1(n_6537),
.B2(n_6568),
.C1(n_6567),
.C2(n_6529),
.Y(n_12403)
);

AOI22xp5_ASAP7_75t_L g12404 ( 
.A1(n_12245),
.A2(n_7153),
.B1(n_7067),
.B2(n_7387),
.Y(n_12404)
);

OAI211xp5_ASAP7_75t_L g12405 ( 
.A1(n_12285),
.A2(n_7387),
.B(n_7398),
.C(n_7391),
.Y(n_12405)
);

NAND2xp5_ASAP7_75t_L g12406 ( 
.A(n_12287),
.B(n_7198),
.Y(n_12406)
);

INVx1_ASAP7_75t_L g12407 ( 
.A(n_12302),
.Y(n_12407)
);

OAI22xp5_ASAP7_75t_SL g12408 ( 
.A1(n_12257),
.A2(n_7408),
.B1(n_7412),
.B2(n_7405),
.Y(n_12408)
);

NAND3x2_ASAP7_75t_L g12409 ( 
.A(n_12248),
.B(n_7412),
.C(n_7408),
.Y(n_12409)
);

O2A1O1Ixp33_ASAP7_75t_L g12410 ( 
.A1(n_12261),
.A2(n_7419),
.B(n_7435),
.C(n_7418),
.Y(n_12410)
);

INVx1_ASAP7_75t_L g12411 ( 
.A(n_12263),
.Y(n_12411)
);

OAI22xp33_ASAP7_75t_L g12412 ( 
.A1(n_12268),
.A2(n_7419),
.B1(n_7435),
.B2(n_7418),
.Y(n_12412)
);

AOI21xp5_ASAP7_75t_L g12413 ( 
.A1(n_12358),
.A2(n_7436),
.B(n_7440),
.Y(n_12413)
);

AOI222xp33_ASAP7_75t_L g12414 ( 
.A1(n_12350),
.A2(n_7448),
.B1(n_7440),
.B2(n_7468),
.C1(n_7460),
.C2(n_7450),
.Y(n_12414)
);

OAI322xp33_ASAP7_75t_SL g12415 ( 
.A1(n_12319),
.A2(n_7468),
.A3(n_7450),
.B1(n_7472),
.B2(n_7483),
.C1(n_7460),
.C2(n_7448),
.Y(n_12415)
);

OAI221xp5_ASAP7_75t_SL g12416 ( 
.A1(n_12289),
.A2(n_7484),
.B1(n_7488),
.B2(n_7483),
.C(n_7472),
.Y(n_12416)
);

AOI222xp33_ASAP7_75t_L g12417 ( 
.A1(n_12374),
.A2(n_7488),
.B1(n_7484),
.B2(n_7503),
.C1(n_7500),
.C2(n_7498),
.Y(n_12417)
);

NOR2xp33_ASAP7_75t_L g12418 ( 
.A(n_12265),
.B(n_7227),
.Y(n_12418)
);

INVx1_ASAP7_75t_SL g12419 ( 
.A(n_12266),
.Y(n_12419)
);

AOI221xp5_ASAP7_75t_L g12420 ( 
.A1(n_12335),
.A2(n_12371),
.B1(n_12318),
.B2(n_12357),
.C(n_12260),
.Y(n_12420)
);

OAI21xp5_ASAP7_75t_L g12421 ( 
.A1(n_12300),
.A2(n_7407),
.B(n_7044),
.Y(n_12421)
);

O2A1O1Ixp33_ASAP7_75t_SL g12422 ( 
.A1(n_12349),
.A2(n_7500),
.B(n_7503),
.C(n_7498),
.Y(n_12422)
);

NAND2xp33_ASAP7_75t_L g12423 ( 
.A(n_12310),
.B(n_7515),
.Y(n_12423)
);

AOI21xp33_ASAP7_75t_L g12424 ( 
.A1(n_12280),
.A2(n_7436),
.B(n_7227),
.Y(n_12424)
);

NOR2x1_ASAP7_75t_L g12425 ( 
.A(n_12321),
.B(n_7515),
.Y(n_12425)
);

OAI321xp33_ASAP7_75t_L g12426 ( 
.A1(n_12281),
.A2(n_7566),
.A3(n_7275),
.B1(n_7338),
.B2(n_7564),
.C(n_7534),
.Y(n_12426)
);

OAI22xp5_ASAP7_75t_L g12427 ( 
.A1(n_12317),
.A2(n_7524),
.B1(n_7527),
.B2(n_7522),
.Y(n_12427)
);

OR2x2_ASAP7_75t_L g12428 ( 
.A(n_12267),
.B(n_7567),
.Y(n_12428)
);

INVxp67_ASAP7_75t_L g12429 ( 
.A(n_12241),
.Y(n_12429)
);

AOI221xp5_ASAP7_75t_L g12430 ( 
.A1(n_12283),
.A2(n_7527),
.B1(n_7547),
.B2(n_7524),
.C(n_7522),
.Y(n_12430)
);

AOI21xp33_ASAP7_75t_L g12431 ( 
.A1(n_12316),
.A2(n_7436),
.B(n_7227),
.Y(n_12431)
);

AND2x2_ASAP7_75t_L g12432 ( 
.A(n_12360),
.B(n_7198),
.Y(n_12432)
);

OAI31xp33_ASAP7_75t_L g12433 ( 
.A1(n_12328),
.A2(n_7555),
.A3(n_7578),
.B(n_7547),
.Y(n_12433)
);

NAND2xp5_ASAP7_75t_L g12434 ( 
.A(n_12256),
.B(n_7198),
.Y(n_12434)
);

INVx2_ASAP7_75t_L g12435 ( 
.A(n_12321),
.Y(n_12435)
);

NOR3xp33_ASAP7_75t_L g12436 ( 
.A(n_12325),
.B(n_7044),
.C(n_7379),
.Y(n_12436)
);

AOI21xp5_ASAP7_75t_L g12437 ( 
.A1(n_12356),
.A2(n_7436),
.B(n_7555),
.Y(n_12437)
);

O2A1O1Ixp5_ASAP7_75t_L g12438 ( 
.A1(n_12270),
.A2(n_7580),
.B(n_7589),
.C(n_7578),
.Y(n_12438)
);

AOI221x1_ASAP7_75t_L g12439 ( 
.A1(n_12320),
.A2(n_12326),
.B1(n_12313),
.B2(n_12311),
.C(n_12331),
.Y(n_12439)
);

OAI21xp33_ASAP7_75t_L g12440 ( 
.A1(n_12295),
.A2(n_7589),
.B(n_7580),
.Y(n_12440)
);

INVx1_ASAP7_75t_L g12441 ( 
.A(n_12369),
.Y(n_12441)
);

OAI22xp5_ASAP7_75t_L g12442 ( 
.A1(n_12324),
.A2(n_7598),
.B1(n_7600),
.B2(n_7595),
.Y(n_12442)
);

O2A1O1Ixp33_ASAP7_75t_L g12443 ( 
.A1(n_12354),
.A2(n_7600),
.B(n_7629),
.C(n_7598),
.Y(n_12443)
);

O2A1O1Ixp5_ASAP7_75t_L g12444 ( 
.A1(n_12367),
.A2(n_7338),
.B(n_7371),
.C(n_7275),
.Y(n_12444)
);

AOI221xp5_ASAP7_75t_L g12445 ( 
.A1(n_12298),
.A2(n_6529),
.B1(n_6545),
.B2(n_6537),
.C(n_6530),
.Y(n_12445)
);

AND2x2_ASAP7_75t_L g12446 ( 
.A(n_12352),
.B(n_6900),
.Y(n_12446)
);

NAND2xp5_ASAP7_75t_L g12447 ( 
.A(n_12326),
.B(n_6874),
.Y(n_12447)
);

NAND2xp5_ASAP7_75t_SL g12448 ( 
.A(n_12286),
.B(n_7480),
.Y(n_12448)
);

OAI221xp5_ASAP7_75t_L g12449 ( 
.A1(n_12252),
.A2(n_6995),
.B1(n_6969),
.B2(n_7227),
.C(n_7289),
.Y(n_12449)
);

AOI21xp5_ASAP7_75t_L g12450 ( 
.A1(n_12348),
.A2(n_6995),
.B(n_6969),
.Y(n_12450)
);

AOI221xp5_ASAP7_75t_L g12451 ( 
.A1(n_12359),
.A2(n_6529),
.B1(n_6567),
.B2(n_6545),
.C(n_6537),
.Y(n_12451)
);

NAND2xp5_ASAP7_75t_L g12452 ( 
.A(n_12259),
.B(n_6874),
.Y(n_12452)
);

OAI22xp5_ASAP7_75t_L g12453 ( 
.A1(n_12351),
.A2(n_6567),
.B1(n_6568),
.B2(n_6379),
.Y(n_12453)
);

NAND2xp5_ASAP7_75t_L g12454 ( 
.A(n_12342),
.B(n_6874),
.Y(n_12454)
);

OAI321xp33_ASAP7_75t_L g12455 ( 
.A1(n_12273),
.A2(n_7371),
.A3(n_7534),
.B1(n_7566),
.B2(n_7564),
.C(n_6197),
.Y(n_12455)
);

O2A1O1Ixp5_ASAP7_75t_SL g12456 ( 
.A1(n_12293),
.A2(n_6372),
.B(n_6383),
.C(n_6366),
.Y(n_12456)
);

INVx1_ASAP7_75t_L g12457 ( 
.A(n_12284),
.Y(n_12457)
);

OAI211xp5_ASAP7_75t_L g12458 ( 
.A1(n_12240),
.A2(n_7482),
.B(n_6969),
.C(n_6995),
.Y(n_12458)
);

INVx1_ASAP7_75t_L g12459 ( 
.A(n_12355),
.Y(n_12459)
);

AOI21xp5_ASAP7_75t_L g12460 ( 
.A1(n_12336),
.A2(n_6995),
.B(n_6969),
.Y(n_12460)
);

NAND2xp5_ASAP7_75t_L g12461 ( 
.A(n_12294),
.B(n_6874),
.Y(n_12461)
);

OAI21xp33_ASAP7_75t_SL g12462 ( 
.A1(n_12330),
.A2(n_7389),
.B(n_7379),
.Y(n_12462)
);

NOR2xp33_ASAP7_75t_L g12463 ( 
.A(n_12340),
.B(n_7289),
.Y(n_12463)
);

INVx1_ASAP7_75t_L g12464 ( 
.A(n_12376),
.Y(n_12464)
);

INVx1_ASAP7_75t_L g12465 ( 
.A(n_12337),
.Y(n_12465)
);

OAI21xp33_ASAP7_75t_L g12466 ( 
.A1(n_12303),
.A2(n_6361),
.B(n_6360),
.Y(n_12466)
);

OAI221xp5_ASAP7_75t_L g12467 ( 
.A1(n_12375),
.A2(n_7289),
.B1(n_7258),
.B2(n_7256),
.C(n_6367),
.Y(n_12467)
);

OAI22xp33_ASAP7_75t_SL g12468 ( 
.A1(n_12274),
.A2(n_6440),
.B1(n_6415),
.B2(n_6361),
.Y(n_12468)
);

AOI21xp5_ASAP7_75t_L g12469 ( 
.A1(n_12306),
.A2(n_7018),
.B(n_7010),
.Y(n_12469)
);

AOI21xp5_ASAP7_75t_L g12470 ( 
.A1(n_12332),
.A2(n_7018),
.B(n_7010),
.Y(n_12470)
);

INVx1_ASAP7_75t_L g12471 ( 
.A(n_12307),
.Y(n_12471)
);

OAI221xp5_ASAP7_75t_L g12472 ( 
.A1(n_12339),
.A2(n_7289),
.B1(n_7258),
.B2(n_7256),
.C(n_6367),
.Y(n_12472)
);

OAI22xp5_ASAP7_75t_L g12473 ( 
.A1(n_12304),
.A2(n_12276),
.B1(n_12373),
.B2(n_12366),
.Y(n_12473)
);

AO21x1_ASAP7_75t_L g12474 ( 
.A1(n_12362),
.A2(n_6361),
.B(n_6360),
.Y(n_12474)
);

AOI22xp5_ASAP7_75t_L g12475 ( 
.A1(n_12301),
.A2(n_12282),
.B1(n_12296),
.B2(n_12269),
.Y(n_12475)
);

AOI21xp5_ASAP7_75t_L g12476 ( 
.A1(n_12277),
.A2(n_12343),
.B(n_12297),
.Y(n_12476)
);

INVx2_ASAP7_75t_SL g12477 ( 
.A(n_12341),
.Y(n_12477)
);

AOI21xp33_ASAP7_75t_SL g12478 ( 
.A1(n_12364),
.A2(n_6884),
.B(n_7056),
.Y(n_12478)
);

OAI21xp5_ASAP7_75t_L g12479 ( 
.A1(n_12333),
.A2(n_7056),
.B(n_6884),
.Y(n_12479)
);

OAI221xp5_ASAP7_75t_SL g12480 ( 
.A1(n_12292),
.A2(n_6367),
.B1(n_6363),
.B2(n_6361),
.C(n_6360),
.Y(n_12480)
);

AOI21xp33_ASAP7_75t_L g12481 ( 
.A1(n_12368),
.A2(n_7258),
.B(n_7256),
.Y(n_12481)
);

AOI21xp33_ASAP7_75t_SL g12482 ( 
.A1(n_12291),
.A2(n_7294),
.B(n_7291),
.Y(n_12482)
);

NAND2xp33_ASAP7_75t_L g12483 ( 
.A(n_12372),
.B(n_6440),
.Y(n_12483)
);

OAI221xp5_ASAP7_75t_SL g12484 ( 
.A1(n_12347),
.A2(n_6367),
.B1(n_6379),
.B2(n_6363),
.C(n_6360),
.Y(n_12484)
);

NAND2xp5_ASAP7_75t_L g12485 ( 
.A(n_12363),
.B(n_6874),
.Y(n_12485)
);

OAI21xp5_ASAP7_75t_L g12486 ( 
.A1(n_12309),
.A2(n_7294),
.B(n_7291),
.Y(n_12486)
);

AOI322xp5_ASAP7_75t_L g12487 ( 
.A1(n_12334),
.A2(n_6440),
.A3(n_6379),
.B1(n_6384),
.B2(n_6363),
.C1(n_6172),
.C2(n_6162),
.Y(n_12487)
);

O2A1O1Ixp33_ASAP7_75t_L g12488 ( 
.A1(n_12361),
.A2(n_6440),
.B(n_6379),
.C(n_6384),
.Y(n_12488)
);

AOI221xp5_ASAP7_75t_L g12489 ( 
.A1(n_12345),
.A2(n_6363),
.B1(n_6384),
.B2(n_6383),
.C(n_6372),
.Y(n_12489)
);

OAI222xp33_ASAP7_75t_L g12490 ( 
.A1(n_12314),
.A2(n_6384),
.B1(n_6175),
.B2(n_6162),
.C1(n_6201),
.C2(n_6184),
.Y(n_12490)
);

NOR3xp33_ASAP7_75t_SL g12491 ( 
.A(n_12338),
.B(n_5765),
.C(n_5755),
.Y(n_12491)
);

NOR2xp33_ASAP7_75t_SL g12492 ( 
.A(n_12344),
.B(n_12323),
.Y(n_12492)
);

INVx3_ASAP7_75t_L g12493 ( 
.A(n_12327),
.Y(n_12493)
);

NAND2xp5_ASAP7_75t_SL g12494 ( 
.A(n_12323),
.B(n_7303),
.Y(n_12494)
);

AOI21xp5_ASAP7_75t_L g12495 ( 
.A1(n_12327),
.A2(n_6879),
.B(n_6875),
.Y(n_12495)
);

AOI211x1_ASAP7_75t_SL g12496 ( 
.A1(n_12322),
.A2(n_6172),
.B(n_6175),
.C(n_6162),
.Y(n_12496)
);

AOI22xp5_ASAP7_75t_L g12497 ( 
.A1(n_12365),
.A2(n_7258),
.B1(n_7256),
.B2(n_7168),
.Y(n_12497)
);

NAND2xp5_ASAP7_75t_L g12498 ( 
.A(n_12237),
.B(n_6874),
.Y(n_12498)
);

AOI221xp5_ASAP7_75t_L g12499 ( 
.A1(n_12253),
.A2(n_6390),
.B1(n_6401),
.B2(n_6383),
.C(n_6372),
.Y(n_12499)
);

AOI221xp5_ASAP7_75t_L g12500 ( 
.A1(n_12253),
.A2(n_6421),
.B1(n_6429),
.B2(n_6401),
.C(n_6390),
.Y(n_12500)
);

NAND2xp5_ASAP7_75t_L g12501 ( 
.A(n_12237),
.B(n_7567),
.Y(n_12501)
);

NAND2xp5_ASAP7_75t_L g12502 ( 
.A(n_12237),
.B(n_7567),
.Y(n_12502)
);

INVx1_ASAP7_75t_L g12503 ( 
.A(n_12290),
.Y(n_12503)
);

AND2x2_ASAP7_75t_L g12504 ( 
.A(n_12244),
.B(n_6900),
.Y(n_12504)
);

INVx1_ASAP7_75t_L g12505 ( 
.A(n_12290),
.Y(n_12505)
);

OAI22xp33_ASAP7_75t_SL g12506 ( 
.A1(n_12244),
.A2(n_6259),
.B1(n_6264),
.B2(n_6044),
.Y(n_12506)
);

INVx1_ASAP7_75t_L g12507 ( 
.A(n_12290),
.Y(n_12507)
);

OAI221xp5_ASAP7_75t_SL g12508 ( 
.A1(n_12289),
.A2(n_6175),
.B1(n_6184),
.B2(n_6172),
.C(n_6162),
.Y(n_12508)
);

AOI22xp5_ASAP7_75t_L g12509 ( 
.A1(n_12378),
.A2(n_7168),
.B1(n_7143),
.B2(n_6098),
.Y(n_12509)
);

AOI322xp5_ASAP7_75t_L g12510 ( 
.A1(n_12378),
.A2(n_6172),
.A3(n_6201),
.B1(n_6175),
.B2(n_6216),
.C1(n_6209),
.C2(n_6184),
.Y(n_12510)
);

NAND2xp33_ASAP7_75t_L g12511 ( 
.A(n_12237),
.B(n_5579),
.Y(n_12511)
);

AOI22xp5_ASAP7_75t_L g12512 ( 
.A1(n_12378),
.A2(n_7168),
.B1(n_7143),
.B2(n_6098),
.Y(n_12512)
);

NAND2x1_ASAP7_75t_L g12513 ( 
.A(n_12237),
.B(n_7606),
.Y(n_12513)
);

AOI22xp5_ASAP7_75t_L g12514 ( 
.A1(n_12378),
.A2(n_7168),
.B1(n_7143),
.B2(n_6098),
.Y(n_12514)
);

AOI22xp5_ASAP7_75t_L g12515 ( 
.A1(n_12378),
.A2(n_7143),
.B1(n_6098),
.B2(n_6135),
.Y(n_12515)
);

INVx1_ASAP7_75t_L g12516 ( 
.A(n_12290),
.Y(n_12516)
);

OAI211xp5_ASAP7_75t_L g12517 ( 
.A1(n_12253),
.A2(n_7303),
.B(n_7454),
.C(n_7439),
.Y(n_12517)
);

NAND2xp5_ASAP7_75t_L g12518 ( 
.A(n_12237),
.B(n_6900),
.Y(n_12518)
);

NAND2xp5_ASAP7_75t_L g12519 ( 
.A(n_12237),
.B(n_6900),
.Y(n_12519)
);

AOI21xp5_ASAP7_75t_L g12520 ( 
.A1(n_12237),
.A2(n_6879),
.B(n_6875),
.Y(n_12520)
);

OAI21xp33_ASAP7_75t_L g12521 ( 
.A1(n_12275),
.A2(n_5745),
.B(n_5618),
.Y(n_12521)
);

OAI221xp5_ASAP7_75t_L g12522 ( 
.A1(n_12420),
.A2(n_6271),
.B1(n_6412),
.B2(n_6264),
.C(n_6259),
.Y(n_12522)
);

OAI21xp33_ASAP7_75t_SL g12523 ( 
.A1(n_12389),
.A2(n_7454),
.B(n_7439),
.Y(n_12523)
);

OAI221xp5_ASAP7_75t_L g12524 ( 
.A1(n_12396),
.A2(n_6414),
.B1(n_6575),
.B2(n_6412),
.C(n_6271),
.Y(n_12524)
);

NOR3xp33_ASAP7_75t_L g12525 ( 
.A(n_12380),
.B(n_6644),
.C(n_7309),
.Y(n_12525)
);

AOI32xp33_ASAP7_75t_L g12526 ( 
.A1(n_12432),
.A2(n_12382),
.A3(n_12507),
.B1(n_12505),
.B2(n_12503),
.Y(n_12526)
);

NAND2xp5_ASAP7_75t_SL g12527 ( 
.A(n_12516),
.B(n_7462),
.Y(n_12527)
);

OAI22xp33_ASAP7_75t_L g12528 ( 
.A1(n_12461),
.A2(n_6201),
.B1(n_6209),
.B2(n_6184),
.Y(n_12528)
);

NAND3xp33_ASAP7_75t_L g12529 ( 
.A(n_12384),
.B(n_12439),
.C(n_12407),
.Y(n_12529)
);

INVx1_ASAP7_75t_L g12530 ( 
.A(n_12394),
.Y(n_12530)
);

OAI211xp5_ASAP7_75t_L g12531 ( 
.A1(n_12441),
.A2(n_7462),
.B(n_6830),
.C(n_6825),
.Y(n_12531)
);

OR3x1_ASAP7_75t_L g12532 ( 
.A(n_12457),
.B(n_6575),
.C(n_6414),
.Y(n_12532)
);

NOR2xp33_ASAP7_75t_L g12533 ( 
.A(n_12390),
.B(n_6825),
.Y(n_12533)
);

AOI21xp5_ASAP7_75t_L g12534 ( 
.A1(n_12419),
.A2(n_7031),
.B(n_6830),
.Y(n_12534)
);

INVx1_ASAP7_75t_L g12535 ( 
.A(n_12504),
.Y(n_12535)
);

AOI211xp5_ASAP7_75t_L g12536 ( 
.A1(n_12473),
.A2(n_7309),
.B(n_7342),
.C(n_7356),
.Y(n_12536)
);

AOI211xp5_ASAP7_75t_L g12537 ( 
.A1(n_12411),
.A2(n_7342),
.B(n_7356),
.C(n_7031),
.Y(n_12537)
);

HB1xp67_ASAP7_75t_L g12538 ( 
.A(n_12477),
.Y(n_12538)
);

OAI21xp33_ASAP7_75t_L g12539 ( 
.A1(n_12521),
.A2(n_5745),
.B(n_5618),
.Y(n_12539)
);

A2O1A1Ixp33_ASAP7_75t_L g12540 ( 
.A1(n_12385),
.A2(n_6962),
.B(n_6957),
.C(n_6989),
.Y(n_12540)
);

AOI22xp33_ASAP7_75t_L g12541 ( 
.A1(n_12390),
.A2(n_6098),
.B1(n_6135),
.B2(n_6106),
.Y(n_12541)
);

AOI222xp33_ASAP7_75t_L g12542 ( 
.A1(n_12462),
.A2(n_6909),
.B1(n_6910),
.B2(n_6989),
.C1(n_6962),
.C2(n_6957),
.Y(n_12542)
);

AND2x2_ASAP7_75t_L g12543 ( 
.A(n_12386),
.B(n_7481),
.Y(n_12543)
);

AOI21xp5_ASAP7_75t_L g12544 ( 
.A1(n_12393),
.A2(n_7026),
.B(n_7020),
.Y(n_12544)
);

NAND4xp25_ASAP7_75t_SL g12545 ( 
.A(n_12379),
.B(n_6216),
.C(n_6217),
.D(n_6201),
.Y(n_12545)
);

OAI31xp33_ASAP7_75t_L g12546 ( 
.A1(n_12458),
.A2(n_3017),
.A3(n_3023),
.B(n_2992),
.Y(n_12546)
);

NAND3xp33_ASAP7_75t_SL g12547 ( 
.A(n_12435),
.B(n_12464),
.C(n_12465),
.Y(n_12547)
);

AND4x1_ASAP7_75t_L g12548 ( 
.A(n_12459),
.B(n_6900),
.C(n_7036),
.D(n_7004),
.Y(n_12548)
);

OAI221xp5_ASAP7_75t_L g12549 ( 
.A1(n_12475),
.A2(n_6579),
.B1(n_6421),
.B2(n_6429),
.C(n_6401),
.Y(n_12549)
);

NAND4xp25_ASAP7_75t_L g12550 ( 
.A(n_12498),
.B(n_3017),
.C(n_3023),
.D(n_2992),
.Y(n_12550)
);

INVxp67_ASAP7_75t_L g12551 ( 
.A(n_12492),
.Y(n_12551)
);

AOI21xp5_ASAP7_75t_L g12552 ( 
.A1(n_12476),
.A2(n_7026),
.B(n_7020),
.Y(n_12552)
);

NAND2xp5_ASAP7_75t_L g12553 ( 
.A(n_12399),
.B(n_6900),
.Y(n_12553)
);

OAI211xp5_ASAP7_75t_L g12554 ( 
.A1(n_12429),
.A2(n_6910),
.B(n_6909),
.C(n_7606),
.Y(n_12554)
);

OAI22xp5_ASAP7_75t_L g12555 ( 
.A1(n_12518),
.A2(n_6216),
.B1(n_6217),
.B2(n_6209),
.Y(n_12555)
);

NAND3xp33_ASAP7_75t_L g12556 ( 
.A(n_12471),
.B(n_7606),
.C(n_7582),
.Y(n_12556)
);

AOI222xp33_ASAP7_75t_L g12557 ( 
.A1(n_12483),
.A2(n_6902),
.B1(n_6915),
.B2(n_6645),
.C1(n_6155),
.C2(n_6216),
.Y(n_12557)
);

NAND2xp33_ASAP7_75t_L g12558 ( 
.A(n_12519),
.B(n_5579),
.Y(n_12558)
);

OAI31xp33_ASAP7_75t_L g12559 ( 
.A1(n_12447),
.A2(n_3017),
.A3(n_3023),
.B(n_2992),
.Y(n_12559)
);

AOI21xp5_ASAP7_75t_L g12560 ( 
.A1(n_12423),
.A2(n_6349),
.B(n_7019),
.Y(n_12560)
);

NOR2x1_ASAP7_75t_L g12561 ( 
.A(n_12493),
.B(n_12425),
.Y(n_12561)
);

AOI321xp33_ASAP7_75t_L g12562 ( 
.A1(n_12446),
.A2(n_6217),
.A3(n_6222),
.B1(n_6258),
.B2(n_6251),
.C(n_6209),
.Y(n_12562)
);

AOI221xp5_ASAP7_75t_L g12563 ( 
.A1(n_12499),
.A2(n_6719),
.B1(n_6794),
.B2(n_6646),
.C(n_6563),
.Y(n_12563)
);

AOI221xp5_ASAP7_75t_L g12564 ( 
.A1(n_12500),
.A2(n_6719),
.B1(n_6794),
.B2(n_6646),
.C(n_6563),
.Y(n_12564)
);

NAND3xp33_ASAP7_75t_SL g12565 ( 
.A(n_12454),
.B(n_3072),
.C(n_6217),
.Y(n_12565)
);

O2A1O1Ixp33_ASAP7_75t_L g12566 ( 
.A1(n_12511),
.A2(n_6629),
.B(n_6490),
.C(n_6496),
.Y(n_12566)
);

AOI31xp33_ASAP7_75t_L g12567 ( 
.A1(n_12383),
.A2(n_5104),
.A3(n_5095),
.B(n_7004),
.Y(n_12567)
);

NAND4xp25_ASAP7_75t_SL g12568 ( 
.A(n_12388),
.B(n_6261),
.C(n_6258),
.D(n_6251),
.Y(n_12568)
);

AOI221xp5_ASAP7_75t_L g12569 ( 
.A1(n_12418),
.A2(n_12422),
.B1(n_12406),
.B2(n_12412),
.C(n_12400),
.Y(n_12569)
);

AOI211xp5_ASAP7_75t_L g12570 ( 
.A1(n_12501),
.A2(n_6861),
.B(n_6857),
.C(n_6645),
.Y(n_12570)
);

A2O1A1Ixp33_ASAP7_75t_L g12571 ( 
.A1(n_12463),
.A2(n_7609),
.B(n_6861),
.C(n_6857),
.Y(n_12571)
);

AOI221xp5_ASAP7_75t_L g12572 ( 
.A1(n_12502),
.A2(n_12448),
.B1(n_12442),
.B2(n_12416),
.C(n_12402),
.Y(n_12572)
);

NAND2xp5_ASAP7_75t_L g12573 ( 
.A(n_12491),
.B(n_7004),
.Y(n_12573)
);

AOI211xp5_ASAP7_75t_L g12574 ( 
.A1(n_12428),
.A2(n_6645),
.B(n_6373),
.C(n_7495),
.Y(n_12574)
);

OR2x2_ASAP7_75t_L g12575 ( 
.A(n_12452),
.B(n_12485),
.Y(n_12575)
);

O2A1O1Ixp5_ASAP7_75t_L g12576 ( 
.A1(n_12493),
.A2(n_6490),
.B(n_6496),
.C(n_6489),
.Y(n_12576)
);

OAI21xp33_ASAP7_75t_L g12577 ( 
.A1(n_12434),
.A2(n_5745),
.B(n_5618),
.Y(n_12577)
);

NAND4xp25_ASAP7_75t_SL g12578 ( 
.A(n_12417),
.B(n_12443),
.C(n_12456),
.D(n_12489),
.Y(n_12578)
);

AOI221x1_ASAP7_75t_L g12579 ( 
.A1(n_12437),
.A2(n_6258),
.B1(n_6261),
.B2(n_6251),
.C(n_6222),
.Y(n_12579)
);

AOI322xp5_ASAP7_75t_L g12580 ( 
.A1(n_12440),
.A2(n_6222),
.A3(n_6261),
.B1(n_6251),
.B2(n_6258),
.C1(n_7036),
.C2(n_7004),
.Y(n_12580)
);

O2A1O1Ixp33_ASAP7_75t_SL g12581 ( 
.A1(n_12387),
.A2(n_6490),
.B(n_6496),
.C(n_6489),
.Y(n_12581)
);

INVx1_ASAP7_75t_L g12582 ( 
.A(n_12392),
.Y(n_12582)
);

AOI221xp5_ASAP7_75t_SL g12583 ( 
.A1(n_12413),
.A2(n_6261),
.B1(n_6222),
.B2(n_6421),
.C(n_6390),
.Y(n_12583)
);

AOI222xp33_ASAP7_75t_L g12584 ( 
.A1(n_12408),
.A2(n_12494),
.B1(n_12479),
.B2(n_12405),
.C1(n_12517),
.C2(n_12466),
.Y(n_12584)
);

AOI211xp5_ASAP7_75t_L g12585 ( 
.A1(n_12395),
.A2(n_6373),
.B(n_7506),
.C(n_7495),
.Y(n_12585)
);

AOI21xp5_ASAP7_75t_SL g12586 ( 
.A1(n_12410),
.A2(n_3023),
.B(n_3017),
.Y(n_12586)
);

NOR3xp33_ASAP7_75t_L g12587 ( 
.A(n_12438),
.B(n_3072),
.C(n_7019),
.Y(n_12587)
);

OAI21xp33_ASAP7_75t_L g12588 ( 
.A1(n_12480),
.A2(n_5944),
.B(n_5801),
.Y(n_12588)
);

OAI211xp5_ASAP7_75t_L g12589 ( 
.A1(n_12409),
.A2(n_7606),
.B(n_6579),
.C(n_7582),
.Y(n_12589)
);

AOI21xp33_ASAP7_75t_L g12590 ( 
.A1(n_12414),
.A2(n_6349),
.B(n_6155),
.Y(n_12590)
);

AOI21xp5_ASAP7_75t_L g12591 ( 
.A1(n_12513),
.A2(n_6349),
.B(n_6902),
.Y(n_12591)
);

NAND3xp33_ASAP7_75t_SL g12592 ( 
.A(n_12397),
.B(n_3072),
.C(n_6489),
.Y(n_12592)
);

OAI221xp5_ASAP7_75t_L g12593 ( 
.A1(n_12433),
.A2(n_6433),
.B1(n_6443),
.B2(n_6438),
.C(n_6429),
.Y(n_12593)
);

AND2x2_ASAP7_75t_L g12594 ( 
.A(n_12486),
.B(n_7481),
.Y(n_12594)
);

HB1xp67_ASAP7_75t_L g12595 ( 
.A(n_12496),
.Y(n_12595)
);

O2A1O1Ixp33_ASAP7_75t_L g12596 ( 
.A1(n_12506),
.A2(n_6629),
.B(n_6496),
.C(n_6499),
.Y(n_12596)
);

OAI221xp5_ASAP7_75t_L g12597 ( 
.A1(n_12431),
.A2(n_6438),
.B1(n_6443),
.B2(n_6433),
.C(n_6430),
.Y(n_12597)
);

INVx1_ASAP7_75t_SL g12598 ( 
.A(n_12424),
.Y(n_12598)
);

OAI21xp33_ASAP7_75t_SL g12599 ( 
.A1(n_12430),
.A2(n_6915),
.B(n_7506),
.Y(n_12599)
);

AOI311xp33_ASAP7_75t_L g12600 ( 
.A1(n_12470),
.A2(n_6430),
.A3(n_6443),
.B(n_6438),
.C(n_6433),
.Y(n_12600)
);

INVx1_ASAP7_75t_L g12601 ( 
.A(n_12474),
.Y(n_12601)
);

NOR2xp33_ASAP7_75t_L g12602 ( 
.A(n_12401),
.B(n_6098),
.Y(n_12602)
);

AOI221xp5_ASAP7_75t_L g12603 ( 
.A1(n_12415),
.A2(n_6532),
.B1(n_6543),
.B2(n_6522),
.C(n_6468),
.Y(n_12603)
);

AOI21xp5_ASAP7_75t_L g12604 ( 
.A1(n_12520),
.A2(n_6155),
.B(n_7609),
.Y(n_12604)
);

NAND2xp5_ASAP7_75t_L g12605 ( 
.A(n_12478),
.B(n_7004),
.Y(n_12605)
);

NAND2xp5_ASAP7_75t_SL g12606 ( 
.A(n_12509),
.B(n_5579),
.Y(n_12606)
);

AOI221xp5_ASAP7_75t_L g12607 ( 
.A1(n_12508),
.A2(n_6636),
.B1(n_6688),
.B2(n_6547),
.C(n_6471),
.Y(n_12607)
);

NAND3xp33_ASAP7_75t_SL g12608 ( 
.A(n_12482),
.B(n_6499),
.C(n_6490),
.Y(n_12608)
);

O2A1O1Ixp33_ASAP7_75t_L g12609 ( 
.A1(n_12398),
.A2(n_6629),
.B(n_6499),
.C(n_6527),
.Y(n_12609)
);

AOI221xp5_ASAP7_75t_L g12610 ( 
.A1(n_12484),
.A2(n_6638),
.B1(n_6690),
.B2(n_6515),
.C(n_6471),
.Y(n_12610)
);

NAND4xp25_ASAP7_75t_L g12611 ( 
.A(n_12469),
.B(n_12514),
.C(n_12512),
.D(n_12391),
.Y(n_12611)
);

NOR2xp33_ASAP7_75t_L g12612 ( 
.A(n_12481),
.B(n_6106),
.Y(n_12612)
);

NAND2xp5_ASAP7_75t_L g12613 ( 
.A(n_12436),
.B(n_12450),
.Y(n_12613)
);

NOR2xp33_ASAP7_75t_L g12614 ( 
.A(n_12427),
.B(n_12421),
.Y(n_12614)
);

OAI211xp5_ASAP7_75t_L g12615 ( 
.A1(n_12515),
.A2(n_7582),
.B(n_6515),
.C(n_6638),
.Y(n_12615)
);

AOI221xp5_ASAP7_75t_L g12616 ( 
.A1(n_12468),
.A2(n_12453),
.B1(n_12455),
.B2(n_12444),
.C(n_12495),
.Y(n_12616)
);

AOI21xp5_ASAP7_75t_L g12617 ( 
.A1(n_12460),
.A2(n_6950),
.B(n_6927),
.Y(n_12617)
);

AOI221xp5_ASAP7_75t_SL g12618 ( 
.A1(n_12488),
.A2(n_6455),
.B1(n_6465),
.B2(n_6450),
.C(n_6430),
.Y(n_12618)
);

INVx1_ASAP7_75t_L g12619 ( 
.A(n_12404),
.Y(n_12619)
);

INVx1_ASAP7_75t_L g12620 ( 
.A(n_12497),
.Y(n_12620)
);

OAI21xp5_ASAP7_75t_L g12621 ( 
.A1(n_12449),
.A2(n_7561),
.B(n_7559),
.Y(n_12621)
);

OAI211xp5_ASAP7_75t_L g12622 ( 
.A1(n_12451),
.A2(n_7582),
.B(n_6516),
.C(n_6535),
.Y(n_12622)
);

INVx1_ASAP7_75t_L g12623 ( 
.A(n_12472),
.Y(n_12623)
);

OA21x2_ASAP7_75t_L g12624 ( 
.A1(n_12490),
.A2(n_6950),
.B(n_6927),
.Y(n_12624)
);

AOI221xp5_ASAP7_75t_SL g12625 ( 
.A1(n_12467),
.A2(n_6465),
.B1(n_6468),
.B2(n_6455),
.C(n_6450),
.Y(n_12625)
);

AOI21xp5_ASAP7_75t_L g12626 ( 
.A1(n_12426),
.A2(n_7561),
.B(n_7559),
.Y(n_12626)
);

NAND3xp33_ASAP7_75t_L g12627 ( 
.A(n_12510),
.B(n_7514),
.C(n_7471),
.Y(n_12627)
);

OAI22xp5_ASAP7_75t_L g12628 ( 
.A1(n_12445),
.A2(n_6106),
.B1(n_6135),
.B2(n_6047),
.Y(n_12628)
);

NAND3xp33_ASAP7_75t_SL g12629 ( 
.A(n_12381),
.B(n_6507),
.C(n_6499),
.Y(n_12629)
);

AND4x1_ASAP7_75t_L g12630 ( 
.A(n_12403),
.B(n_7036),
.C(n_7004),
.D(n_7210),
.Y(n_12630)
);

O2A1O1Ixp33_ASAP7_75t_L g12631 ( 
.A1(n_12487),
.A2(n_6629),
.B(n_6507),
.C(n_6527),
.Y(n_12631)
);

OAI21xp5_ASAP7_75t_L g12632 ( 
.A1(n_12389),
.A2(n_6633),
.B(n_7509),
.Y(n_12632)
);

AOI221xp5_ASAP7_75t_L g12633 ( 
.A1(n_12529),
.A2(n_12526),
.B1(n_12551),
.B2(n_12547),
.C(n_12522),
.Y(n_12633)
);

NOR2xp67_ASAP7_75t_L g12634 ( 
.A(n_12578),
.B(n_12582),
.Y(n_12634)
);

NOR3xp33_ASAP7_75t_L g12635 ( 
.A(n_12530),
.B(n_6633),
.C(n_7509),
.Y(n_12635)
);

NAND2xp5_ASAP7_75t_L g12636 ( 
.A(n_12538),
.B(n_7036),
.Y(n_12636)
);

OAI21xp5_ASAP7_75t_L g12637 ( 
.A1(n_12552),
.A2(n_6633),
.B(n_6194),
.Y(n_12637)
);

OAI22xp5_ASAP7_75t_L g12638 ( 
.A1(n_12573),
.A2(n_6106),
.B1(n_6135),
.B2(n_6047),
.Y(n_12638)
);

NOR3x1_ASAP7_75t_L g12639 ( 
.A(n_12620),
.B(n_6373),
.C(n_6194),
.Y(n_12639)
);

NAND4xp25_ASAP7_75t_L g12640 ( 
.A(n_12572),
.B(n_3051),
.C(n_3083),
.D(n_3023),
.Y(n_12640)
);

AOI21xp33_ASAP7_75t_L g12641 ( 
.A1(n_12598),
.A2(n_6629),
.B(n_7514),
.Y(n_12641)
);

AOI221xp5_ASAP7_75t_L g12642 ( 
.A1(n_12525),
.A2(n_6465),
.B1(n_6468),
.B2(n_6455),
.C(n_6450),
.Y(n_12642)
);

AOI211xp5_ASAP7_75t_L g12643 ( 
.A1(n_12623),
.A2(n_6194),
.B(n_7587),
.C(n_6385),
.Y(n_12643)
);

OAI21xp33_ASAP7_75t_SL g12644 ( 
.A1(n_12561),
.A2(n_7587),
.B(n_6385),
.Y(n_12644)
);

NOR3x1_ASAP7_75t_L g12645 ( 
.A(n_12535),
.B(n_6119),
.C(n_6118),
.Y(n_12645)
);

NAND3xp33_ASAP7_75t_L g12646 ( 
.A(n_12619),
.B(n_6135),
.C(n_6106),
.Y(n_12646)
);

INVx1_ASAP7_75t_L g12647 ( 
.A(n_12532),
.Y(n_12647)
);

NAND2xp5_ASAP7_75t_L g12648 ( 
.A(n_12595),
.B(n_7036),
.Y(n_12648)
);

AOI22xp5_ASAP7_75t_L g12649 ( 
.A1(n_12539),
.A2(n_6106),
.B1(n_6135),
.B2(n_6047),
.Y(n_12649)
);

OAI211xp5_ASAP7_75t_SL g12650 ( 
.A1(n_12569),
.A2(n_12575),
.B(n_12613),
.C(n_12616),
.Y(n_12650)
);

OAI321xp33_ASAP7_75t_L g12651 ( 
.A1(n_12611),
.A2(n_6197),
.A3(n_5824),
.B1(n_5956),
.B2(n_5805),
.C(n_6471),
.Y(n_12651)
);

O2A1O1Ixp33_ASAP7_75t_L g12652 ( 
.A1(n_12601),
.A2(n_6527),
.B(n_6507),
.C(n_3083),
.Y(n_12652)
);

AO21x1_ASAP7_75t_L g12653 ( 
.A1(n_12614),
.A2(n_6527),
.B(n_6507),
.Y(n_12653)
);

OAI22xp5_ASAP7_75t_L g12654 ( 
.A1(n_12605),
.A2(n_6047),
.B1(n_5824),
.B2(n_5956),
.Y(n_12654)
);

AOI222xp33_ASAP7_75t_L g12655 ( 
.A1(n_12608),
.A2(n_6501),
.B1(n_6506),
.B2(n_6515),
.C1(n_6511),
.C2(n_6480),
.Y(n_12655)
);

AOI21xp33_ASAP7_75t_L g12656 ( 
.A1(n_12584),
.A2(n_12577),
.B(n_12533),
.Y(n_12656)
);

OAI221xp5_ASAP7_75t_SL g12657 ( 
.A1(n_12559),
.A2(n_6501),
.B1(n_6511),
.B2(n_6506),
.C(n_6480),
.Y(n_12657)
);

NOR2xp33_ASAP7_75t_L g12658 ( 
.A(n_12550),
.B(n_6047),
.Y(n_12658)
);

AOI22xp33_ASAP7_75t_L g12659 ( 
.A1(n_12588),
.A2(n_6047),
.B1(n_7471),
.B2(n_7514),
.Y(n_12659)
);

INVx2_ASAP7_75t_SL g12660 ( 
.A(n_12543),
.Y(n_12660)
);

AOI22xp5_ASAP7_75t_L g12661 ( 
.A1(n_12612),
.A2(n_5805),
.B1(n_5598),
.B2(n_5685),
.Y(n_12661)
);

AOI221xp5_ASAP7_75t_L g12662 ( 
.A1(n_12558),
.A2(n_6506),
.B1(n_6511),
.B2(n_6501),
.C(n_6480),
.Y(n_12662)
);

AOI21xp5_ASAP7_75t_L g12663 ( 
.A1(n_12586),
.A2(n_7514),
.B(n_7520),
.Y(n_12663)
);

AOI22xp5_ASAP7_75t_L g12664 ( 
.A1(n_12553),
.A2(n_5598),
.B1(n_5685),
.B2(n_5579),
.Y(n_12664)
);

O2A1O1Ixp33_ASAP7_75t_L g12665 ( 
.A1(n_12565),
.A2(n_3083),
.B(n_3051),
.C(n_6572),
.Y(n_12665)
);

OAI211xp5_ASAP7_75t_L g12666 ( 
.A1(n_12546),
.A2(n_12592),
.B(n_12606),
.C(n_12600),
.Y(n_12666)
);

NAND2xp5_ASAP7_75t_SL g12667 ( 
.A(n_12528),
.B(n_5579),
.Y(n_12667)
);

AOI221x1_ASAP7_75t_L g12668 ( 
.A1(n_12587),
.A2(n_6522),
.B1(n_6532),
.B2(n_6517),
.C(n_6516),
.Y(n_12668)
);

NOR3xp33_ASAP7_75t_L g12669 ( 
.A(n_12625),
.B(n_6129),
.C(n_6124),
.Y(n_12669)
);

AO21x1_ASAP7_75t_L g12670 ( 
.A1(n_12631),
.A2(n_7526),
.B(n_7520),
.Y(n_12670)
);

AOI21xp5_ASAP7_75t_L g12671 ( 
.A1(n_12581),
.A2(n_7533),
.B(n_7526),
.Y(n_12671)
);

OAI21xp5_ASAP7_75t_L g12672 ( 
.A1(n_12594),
.A2(n_6329),
.B(n_6119),
.Y(n_12672)
);

AOI221xp5_ASAP7_75t_L g12673 ( 
.A1(n_12568),
.A2(n_6522),
.B1(n_6532),
.B2(n_6517),
.C(n_6516),
.Y(n_12673)
);

AND2x2_ASAP7_75t_L g12674 ( 
.A(n_12618),
.B(n_7481),
.Y(n_12674)
);

AOI221xp5_ASAP7_75t_L g12675 ( 
.A1(n_12549),
.A2(n_6543),
.B1(n_6547),
.B2(n_6535),
.C(n_6517),
.Y(n_12675)
);

NAND2xp5_ASAP7_75t_L g12676 ( 
.A(n_12536),
.B(n_7036),
.Y(n_12676)
);

OR2x2_ASAP7_75t_L g12677 ( 
.A(n_12629),
.B(n_7210),
.Y(n_12677)
);

AOI21xp5_ASAP7_75t_L g12678 ( 
.A1(n_12617),
.A2(n_7533),
.B(n_7535),
.Y(n_12678)
);

AND2x2_ASAP7_75t_L g12679 ( 
.A(n_12583),
.B(n_7481),
.Y(n_12679)
);

AOI31xp33_ASAP7_75t_L g12680 ( 
.A1(n_12557),
.A2(n_5104),
.A3(n_5095),
.B(n_5755),
.Y(n_12680)
);

OAI221xp5_ASAP7_75t_L g12681 ( 
.A1(n_12597),
.A2(n_6535),
.B1(n_6552),
.B2(n_6547),
.C(n_6543),
.Y(n_12681)
);

AOI221xp5_ASAP7_75t_L g12682 ( 
.A1(n_12545),
.A2(n_6804),
.B1(n_6563),
.B2(n_6570),
.C(n_6562),
.Y(n_12682)
);

O2A1O1Ixp33_ASAP7_75t_L g12683 ( 
.A1(n_12593),
.A2(n_12523),
.B(n_12576),
.C(n_12524),
.Y(n_12683)
);

NAND2xp5_ASAP7_75t_L g12684 ( 
.A(n_12602),
.B(n_7210),
.Y(n_12684)
);

OAI221xp5_ASAP7_75t_L g12685 ( 
.A1(n_12599),
.A2(n_6552),
.B1(n_6580),
.B2(n_6570),
.C(n_6562),
.Y(n_12685)
);

AOI211xp5_ASAP7_75t_SL g12686 ( 
.A1(n_12622),
.A2(n_6562),
.B(n_6570),
.C(n_6552),
.Y(n_12686)
);

AOI21xp5_ASAP7_75t_L g12687 ( 
.A1(n_12534),
.A2(n_12604),
.B(n_12596),
.Y(n_12687)
);

AOI221xp5_ASAP7_75t_L g12688 ( 
.A1(n_12615),
.A2(n_6804),
.B1(n_6586),
.B2(n_6617),
.C(n_6615),
.Y(n_12688)
);

AOI221x1_ASAP7_75t_L g12689 ( 
.A1(n_12544),
.A2(n_6586),
.B1(n_6617),
.B2(n_6615),
.C(n_6580),
.Y(n_12689)
);

AOI221xp5_ASAP7_75t_L g12690 ( 
.A1(n_12563),
.A2(n_6804),
.B1(n_6586),
.B2(n_6617),
.C(n_6615),
.Y(n_12690)
);

AOI221xp5_ASAP7_75t_L g12691 ( 
.A1(n_12564),
.A2(n_6638),
.B1(n_6646),
.B2(n_6636),
.C(n_6580),
.Y(n_12691)
);

NAND4xp25_ASAP7_75t_L g12692 ( 
.A(n_12570),
.B(n_3083),
.C(n_3051),
.D(n_5801),
.Y(n_12692)
);

AND2x2_ASAP7_75t_L g12693 ( 
.A(n_12632),
.B(n_7481),
.Y(n_12693)
);

NAND2xp5_ASAP7_75t_L g12694 ( 
.A(n_12589),
.B(n_7210),
.Y(n_12694)
);

AOI22xp5_ASAP7_75t_L g12695 ( 
.A1(n_12556),
.A2(n_5685),
.B1(n_5723),
.B2(n_5598),
.Y(n_12695)
);

AOI211xp5_ASAP7_75t_L g12696 ( 
.A1(n_12590),
.A2(n_6385),
.B(n_6118),
.C(n_6119),
.Y(n_12696)
);

AOI22xp5_ASAP7_75t_L g12697 ( 
.A1(n_12555),
.A2(n_5685),
.B1(n_5723),
.B2(n_5598),
.Y(n_12697)
);

OAI31xp33_ASAP7_75t_L g12698 ( 
.A1(n_12540),
.A2(n_3083),
.A3(n_3051),
.B(n_6636),
.Y(n_12698)
);

NOR2xp33_ASAP7_75t_L g12699 ( 
.A(n_12548),
.B(n_5801),
.Y(n_12699)
);

AND2x2_ASAP7_75t_L g12700 ( 
.A(n_12630),
.B(n_7518),
.Y(n_12700)
);

NOR3xp33_ASAP7_75t_L g12701 ( 
.A(n_12621),
.B(n_6129),
.C(n_6124),
.Y(n_12701)
);

AOI22xp5_ASAP7_75t_L g12702 ( 
.A1(n_12527),
.A2(n_5685),
.B1(n_5723),
.B2(n_5598),
.Y(n_12702)
);

AOI221xp5_ASAP7_75t_L g12703 ( 
.A1(n_12609),
.A2(n_6666),
.B1(n_6668),
.B2(n_6654),
.C(n_6649),
.Y(n_12703)
);

OAI21xp33_ASAP7_75t_L g12704 ( 
.A1(n_12567),
.A2(n_5962),
.B(n_5944),
.Y(n_12704)
);

NAND2xp5_ASAP7_75t_L g12705 ( 
.A(n_12560),
.B(n_7210),
.Y(n_12705)
);

AOI22xp5_ASAP7_75t_L g12706 ( 
.A1(n_12542),
.A2(n_5685),
.B1(n_5723),
.B2(n_5598),
.Y(n_12706)
);

OAI221xp5_ASAP7_75t_L g12707 ( 
.A1(n_12537),
.A2(n_6666),
.B1(n_6668),
.B2(n_6654),
.C(n_6649),
.Y(n_12707)
);

O2A1O1Ixp33_ASAP7_75t_L g12708 ( 
.A1(n_12566),
.A2(n_3051),
.B(n_6596),
.C(n_6572),
.Y(n_12708)
);

OAI221xp5_ASAP7_75t_L g12709 ( 
.A1(n_12571),
.A2(n_6666),
.B1(n_6668),
.B2(n_6654),
.C(n_6649),
.Y(n_12709)
);

NAND3xp33_ASAP7_75t_L g12710 ( 
.A(n_12585),
.B(n_6684),
.C(n_6681),
.Y(n_12710)
);

NOR3x1_ASAP7_75t_L g12711 ( 
.A(n_12627),
.B(n_6118),
.C(n_6705),
.Y(n_12711)
);

AOI21xp5_ASAP7_75t_L g12712 ( 
.A1(n_12626),
.A2(n_12591),
.B(n_12628),
.Y(n_12712)
);

OAI221xp5_ASAP7_75t_L g12713 ( 
.A1(n_12574),
.A2(n_6688),
.B1(n_6690),
.B2(n_6684),
.C(n_6681),
.Y(n_12713)
);

NAND2xp5_ASAP7_75t_L g12714 ( 
.A(n_12603),
.B(n_7210),
.Y(n_12714)
);

NAND4xp25_ASAP7_75t_L g12715 ( 
.A(n_12610),
.B(n_3147),
.C(n_3129),
.D(n_5944),
.Y(n_12715)
);

AOI211xp5_ASAP7_75t_L g12716 ( 
.A1(n_12531),
.A2(n_6129),
.B(n_6705),
.C(n_6764),
.Y(n_12716)
);

NOR3xp33_ASAP7_75t_L g12717 ( 
.A(n_12554),
.B(n_6329),
.C(n_6730),
.Y(n_12717)
);

AOI221xp5_ASAP7_75t_L g12718 ( 
.A1(n_12607),
.A2(n_6688),
.B1(n_6690),
.B2(n_6684),
.C(n_6681),
.Y(n_12718)
);

AOI221x1_ASAP7_75t_L g12719 ( 
.A1(n_12624),
.A2(n_6719),
.B1(n_6722),
.B2(n_6718),
.C(n_6714),
.Y(n_12719)
);

AOI21xp5_ASAP7_75t_L g12720 ( 
.A1(n_12624),
.A2(n_7535),
.B(n_7517),
.Y(n_12720)
);

AOI221xp5_ASAP7_75t_L g12721 ( 
.A1(n_12541),
.A2(n_6795),
.B1(n_6722),
.B2(n_6748),
.C(n_6718),
.Y(n_12721)
);

AOI221xp5_ASAP7_75t_L g12722 ( 
.A1(n_12562),
.A2(n_6795),
.B1(n_6722),
.B2(n_6748),
.C(n_6718),
.Y(n_12722)
);

OAI221xp5_ASAP7_75t_L g12723 ( 
.A1(n_12580),
.A2(n_6762),
.B1(n_6764),
.B2(n_6748),
.C(n_6714),
.Y(n_12723)
);

OAI21xp5_ASAP7_75t_L g12724 ( 
.A1(n_12579),
.A2(n_6329),
.B(n_6244),
.Y(n_12724)
);

NAND2xp5_ASAP7_75t_L g12725 ( 
.A(n_12526),
.B(n_7231),
.Y(n_12725)
);

OAI21xp5_ASAP7_75t_SL g12726 ( 
.A1(n_12526),
.A2(n_3021),
.B(n_3003),
.Y(n_12726)
);

AOI22xp5_ASAP7_75t_L g12727 ( 
.A1(n_12551),
.A2(n_5764),
.B1(n_5839),
.B2(n_5723),
.Y(n_12727)
);

NOR2xp33_ASAP7_75t_SL g12728 ( 
.A(n_12529),
.B(n_2876),
.Y(n_12728)
);

OAI21xp5_ASAP7_75t_L g12729 ( 
.A1(n_12529),
.A2(n_6244),
.B(n_6241),
.Y(n_12729)
);

NAND4xp25_ASAP7_75t_L g12730 ( 
.A(n_12526),
.B(n_6002),
.C(n_5962),
.D(n_3147),
.Y(n_12730)
);

INVxp33_ASAP7_75t_L g12731 ( 
.A(n_12538),
.Y(n_12731)
);

NAND3xp33_ASAP7_75t_SL g12732 ( 
.A(n_12526),
.B(n_6596),
.C(n_6572),
.Y(n_12732)
);

NAND3xp33_ASAP7_75t_SL g12733 ( 
.A(n_12526),
.B(n_6596),
.C(n_6572),
.Y(n_12733)
);

NAND3xp33_ASAP7_75t_L g12734 ( 
.A(n_12633),
.B(n_6762),
.C(n_6714),
.Y(n_12734)
);

NOR3x1_ASAP7_75t_L g12735 ( 
.A(n_12640),
.B(n_12726),
.C(n_12725),
.Y(n_12735)
);

NOR3xp33_ASAP7_75t_SL g12736 ( 
.A(n_12650),
.B(n_5787),
.C(n_5765),
.Y(n_12736)
);

NAND2xp5_ASAP7_75t_L g12737 ( 
.A(n_12634),
.B(n_7518),
.Y(n_12737)
);

INVx1_ASAP7_75t_L g12738 ( 
.A(n_12699),
.Y(n_12738)
);

NOR2x1_ASAP7_75t_L g12739 ( 
.A(n_12647),
.B(n_6762),
.Y(n_12739)
);

AOI211xp5_ASAP7_75t_L g12740 ( 
.A1(n_12731),
.A2(n_6765),
.B(n_6766),
.C(n_6764),
.Y(n_12740)
);

AOI311xp33_ASAP7_75t_L g12741 ( 
.A1(n_12656),
.A2(n_12712),
.A3(n_12666),
.B(n_12687),
.C(n_12685),
.Y(n_12741)
);

NOR3xp33_ASAP7_75t_SL g12742 ( 
.A(n_12733),
.B(n_5787),
.C(n_6765),
.Y(n_12742)
);

NOR2xp33_ASAP7_75t_L g12743 ( 
.A(n_12728),
.B(n_5962),
.Y(n_12743)
);

AOI21xp5_ASAP7_75t_L g12744 ( 
.A1(n_12683),
.A2(n_7517),
.B(n_6311),
.Y(n_12744)
);

AOI32xp33_ASAP7_75t_L g12745 ( 
.A1(n_12648),
.A2(n_6705),
.A3(n_6733),
.B1(n_6735),
.B2(n_6730),
.Y(n_12745)
);

OAI222xp33_ASAP7_75t_L g12746 ( 
.A1(n_12636),
.A2(n_6622),
.B1(n_6596),
.B2(n_6624),
.C1(n_6623),
.C2(n_6603),
.Y(n_12746)
);

AOI21xp33_ASAP7_75t_L g12747 ( 
.A1(n_12660),
.A2(n_7517),
.B(n_6225),
.Y(n_12747)
);

NAND2xp5_ASAP7_75t_L g12748 ( 
.A(n_12642),
.B(n_7518),
.Y(n_12748)
);

NAND2xp5_ASAP7_75t_L g12749 ( 
.A(n_12704),
.B(n_7518),
.Y(n_12749)
);

NAND4xp25_ASAP7_75t_L g12750 ( 
.A(n_12730),
.B(n_6002),
.C(n_3147),
.D(n_3129),
.Y(n_12750)
);

NAND3xp33_ASAP7_75t_L g12751 ( 
.A(n_12698),
.B(n_6795),
.C(n_6794),
.Y(n_12751)
);

NAND3xp33_ASAP7_75t_SL g12752 ( 
.A(n_12670),
.B(n_6622),
.C(n_6603),
.Y(n_12752)
);

OAI211xp5_ASAP7_75t_SL g12753 ( 
.A1(n_12661),
.A2(n_6766),
.B(n_6765),
.C(n_6622),
.Y(n_12753)
);

AND4x1_ASAP7_75t_L g12754 ( 
.A(n_12665),
.B(n_7231),
.C(n_6766),
.D(n_7518),
.Y(n_12754)
);

NOR2xp67_ASAP7_75t_SL g12755 ( 
.A(n_12677),
.B(n_12692),
.Y(n_12755)
);

NAND4xp25_ASAP7_75t_SL g12756 ( 
.A(n_12652),
.B(n_6622),
.C(n_6623),
.D(n_6603),
.Y(n_12756)
);

INVx1_ASAP7_75t_L g12757 ( 
.A(n_12732),
.Y(n_12757)
);

AOI21xp5_ASAP7_75t_L g12758 ( 
.A1(n_12708),
.A2(n_7517),
.B(n_6311),
.Y(n_12758)
);

NAND2xp5_ASAP7_75t_L g12759 ( 
.A(n_12674),
.B(n_7518),
.Y(n_12759)
);

OAI21xp33_ASAP7_75t_SL g12760 ( 
.A1(n_12700),
.A2(n_7616),
.B(n_6711),
.Y(n_12760)
);

OAI211xp5_ASAP7_75t_L g12761 ( 
.A1(n_12714),
.A2(n_6603),
.B(n_6624),
.C(n_6623),
.Y(n_12761)
);

OAI211xp5_ASAP7_75t_L g12762 ( 
.A1(n_12676),
.A2(n_6623),
.B(n_6648),
.C(n_6624),
.Y(n_12762)
);

NOR2x1_ASAP7_75t_L g12763 ( 
.A(n_12710),
.B(n_12715),
.Y(n_12763)
);

INVx1_ASAP7_75t_L g12764 ( 
.A(n_12679),
.Y(n_12764)
);

NAND2xp5_ASAP7_75t_L g12765 ( 
.A(n_12693),
.B(n_7231),
.Y(n_12765)
);

NAND2xp5_ASAP7_75t_L g12766 ( 
.A(n_12715),
.B(n_7231),
.Y(n_12766)
);

NAND2xp5_ASAP7_75t_L g12767 ( 
.A(n_12686),
.B(n_7231),
.Y(n_12767)
);

A2O1A1Ixp33_ASAP7_75t_L g12768 ( 
.A1(n_12644),
.A2(n_7616),
.B(n_6709),
.C(n_6711),
.Y(n_12768)
);

AOI211xp5_ASAP7_75t_L g12769 ( 
.A1(n_12657),
.A2(n_12654),
.B(n_12707),
.C(n_12667),
.Y(n_12769)
);

NAND4xp25_ASAP7_75t_L g12770 ( 
.A(n_12689),
.B(n_6002),
.C(n_3147),
.D(n_3129),
.Y(n_12770)
);

OAI211xp5_ASAP7_75t_L g12771 ( 
.A1(n_12729),
.A2(n_6624),
.B(n_6673),
.C(n_6648),
.Y(n_12771)
);

NAND4xp25_ASAP7_75t_L g12772 ( 
.A(n_12711),
.B(n_12668),
.C(n_12727),
.D(n_12719),
.Y(n_12772)
);

NAND4xp25_ASAP7_75t_L g12773 ( 
.A(n_12703),
.B(n_3147),
.C(n_3129),
.D(n_3177),
.Y(n_12773)
);

NOR3xp33_ASAP7_75t_L g12774 ( 
.A(n_12713),
.B(n_6244),
.C(n_6241),
.Y(n_12774)
);

NOR3xp33_ASAP7_75t_L g12775 ( 
.A(n_12684),
.B(n_6241),
.C(n_6730),
.Y(n_12775)
);

NAND2xp5_ASAP7_75t_L g12776 ( 
.A(n_12658),
.B(n_7231),
.Y(n_12776)
);

AND2x2_ASAP7_75t_L g12777 ( 
.A(n_12717),
.B(n_7334),
.Y(n_12777)
);

AOI221xp5_ASAP7_75t_SL g12778 ( 
.A1(n_12680),
.A2(n_6692),
.B1(n_6786),
.B2(n_6784),
.C(n_6673),
.Y(n_12778)
);

NAND3xp33_ASAP7_75t_L g12779 ( 
.A(n_12701),
.B(n_6225),
.C(n_6265),
.Y(n_12779)
);

NAND4xp25_ASAP7_75t_SL g12780 ( 
.A(n_12694),
.B(n_12653),
.C(n_12696),
.D(n_12705),
.Y(n_12780)
);

NOR3xp33_ASAP7_75t_L g12781 ( 
.A(n_12651),
.B(n_6735),
.C(n_6733),
.Y(n_12781)
);

OAI21xp5_ASAP7_75t_L g12782 ( 
.A1(n_12672),
.A2(n_6080),
.B(n_6077),
.Y(n_12782)
);

NOR2xp33_ASAP7_75t_L g12783 ( 
.A(n_12681),
.B(n_5723),
.Y(n_12783)
);

INVx1_ASAP7_75t_L g12784 ( 
.A(n_12709),
.Y(n_12784)
);

NAND2xp5_ASAP7_75t_L g12785 ( 
.A(n_12678),
.B(n_7334),
.Y(n_12785)
);

AOI221xp5_ASAP7_75t_L g12786 ( 
.A1(n_12723),
.A2(n_6797),
.B1(n_6789),
.B2(n_6786),
.C(n_6692),
.Y(n_12786)
);

NOR2x1_ASAP7_75t_L g12787 ( 
.A(n_12646),
.B(n_6648),
.Y(n_12787)
);

OAI21xp5_ASAP7_75t_SL g12788 ( 
.A1(n_12664),
.A2(n_12655),
.B(n_12662),
.Y(n_12788)
);

INVx1_ASAP7_75t_L g12789 ( 
.A(n_12637),
.Y(n_12789)
);

NAND2x1_ASAP7_75t_SL g12790 ( 
.A(n_12702),
.B(n_12706),
.Y(n_12790)
);

NAND2xp5_ASAP7_75t_L g12791 ( 
.A(n_12716),
.B(n_7334),
.Y(n_12791)
);

NAND3xp33_ASAP7_75t_L g12792 ( 
.A(n_12669),
.B(n_6225),
.C(n_6265),
.Y(n_12792)
);

NAND4xp25_ASAP7_75t_L g12793 ( 
.A(n_12718),
.B(n_3177),
.C(n_4483),
.D(n_4441),
.Y(n_12793)
);

INVx1_ASAP7_75t_L g12794 ( 
.A(n_12645),
.Y(n_12794)
);

AND4x1_ASAP7_75t_L g12795 ( 
.A(n_12639),
.B(n_6307),
.C(n_6592),
.D(n_6312),
.Y(n_12795)
);

AND4x1_ASAP7_75t_L g12796 ( 
.A(n_12643),
.B(n_12721),
.C(n_12691),
.D(n_12690),
.Y(n_12796)
);

OAI322xp33_ASAP7_75t_SL g12797 ( 
.A1(n_12663),
.A2(n_6789),
.A3(n_6797),
.B1(n_6786),
.B2(n_6740),
.C1(n_6648),
.C2(n_6692),
.Y(n_12797)
);

NAND4xp25_ASAP7_75t_L g12798 ( 
.A(n_12688),
.B(n_3177),
.C(n_4483),
.D(n_4441),
.Y(n_12798)
);

NOR4xp25_ASAP7_75t_L g12799 ( 
.A(n_12641),
.B(n_6692),
.C(n_6703),
.D(n_6673),
.Y(n_12799)
);

INVx1_ASAP7_75t_L g12800 ( 
.A(n_12695),
.Y(n_12800)
);

NAND2xp5_ASAP7_75t_SL g12801 ( 
.A(n_12697),
.B(n_5764),
.Y(n_12801)
);

NOR2x1_ASAP7_75t_L g12802 ( 
.A(n_12671),
.B(n_6673),
.Y(n_12802)
);

NOR2xp33_ASAP7_75t_SL g12803 ( 
.A(n_12638),
.B(n_3165),
.Y(n_12803)
);

INVx1_ASAP7_75t_L g12804 ( 
.A(n_12675),
.Y(n_12804)
);

NAND2xp5_ASAP7_75t_SL g12805 ( 
.A(n_12682),
.B(n_12720),
.Y(n_12805)
);

NOR2x1_ASAP7_75t_L g12806 ( 
.A(n_12724),
.B(n_6703),
.Y(n_12806)
);

NAND3xp33_ASAP7_75t_SL g12807 ( 
.A(n_12635),
.B(n_6740),
.C(n_6703),
.Y(n_12807)
);

NAND2xp5_ASAP7_75t_L g12808 ( 
.A(n_12673),
.B(n_7334),
.Y(n_12808)
);

NOR3x1_ASAP7_75t_L g12809 ( 
.A(n_12722),
.B(n_6735),
.C(n_6733),
.Y(n_12809)
);

INVx2_ASAP7_75t_SL g12810 ( 
.A(n_12649),
.Y(n_12810)
);

NOR2x1_ASAP7_75t_L g12811 ( 
.A(n_12659),
.B(n_6703),
.Y(n_12811)
);

NAND3xp33_ASAP7_75t_L g12812 ( 
.A(n_12633),
.B(n_6225),
.C(n_6265),
.Y(n_12812)
);

NOR4xp25_ASAP7_75t_L g12813 ( 
.A(n_12741),
.B(n_6741),
.C(n_6763),
.D(n_6740),
.Y(n_12813)
);

NOR3x1_ASAP7_75t_L g12814 ( 
.A(n_12810),
.B(n_6711),
.C(n_6709),
.Y(n_12814)
);

NAND2xp33_ASAP7_75t_SL g12815 ( 
.A(n_12736),
.B(n_12755),
.Y(n_12815)
);

NOR2xp33_ASAP7_75t_L g12816 ( 
.A(n_12738),
.B(n_12757),
.Y(n_12816)
);

NOR4xp75_ASAP7_75t_L g12817 ( 
.A(n_12790),
.B(n_4963),
.C(n_4991),
.D(n_4844),
.Y(n_12817)
);

INVx1_ASAP7_75t_L g12818 ( 
.A(n_12737),
.Y(n_12818)
);

NOR3xp33_ASAP7_75t_L g12819 ( 
.A(n_12764),
.B(n_6188),
.C(n_6709),
.Y(n_12819)
);

OAI211xp5_ASAP7_75t_L g12820 ( 
.A1(n_12794),
.A2(n_6740),
.B(n_6763),
.C(n_6741),
.Y(n_12820)
);

AOI211xp5_ASAP7_75t_L g12821 ( 
.A1(n_12780),
.A2(n_6080),
.B(n_6077),
.C(n_6069),
.Y(n_12821)
);

NOR2x1_ASAP7_75t_L g12822 ( 
.A(n_12739),
.B(n_6741),
.Y(n_12822)
);

AOI221xp5_ASAP7_75t_L g12823 ( 
.A1(n_12752),
.A2(n_6773),
.B1(n_6783),
.B2(n_6763),
.C(n_6741),
.Y(n_12823)
);

AOI211xp5_ASAP7_75t_L g12824 ( 
.A1(n_12804),
.A2(n_12805),
.B(n_12800),
.C(n_12788),
.Y(n_12824)
);

NOR3xp33_ASAP7_75t_L g12825 ( 
.A(n_12789),
.B(n_6188),
.C(n_6080),
.Y(n_12825)
);

NAND3xp33_ASAP7_75t_L g12826 ( 
.A(n_12784),
.B(n_12769),
.C(n_12763),
.Y(n_12826)
);

OAI22xp5_ASAP7_75t_L g12827 ( 
.A1(n_12734),
.A2(n_6773),
.B1(n_6783),
.B2(n_6763),
.Y(n_12827)
);

XOR2xp5_ASAP7_75t_L g12828 ( 
.A(n_12772),
.B(n_3003),
.Y(n_12828)
);

NAND4xp25_ASAP7_75t_L g12829 ( 
.A(n_12735),
.B(n_3177),
.C(n_4483),
.D(n_4441),
.Y(n_12829)
);

OAI211xp5_ASAP7_75t_L g12830 ( 
.A1(n_12761),
.A2(n_6784),
.B(n_6786),
.C(n_6783),
.Y(n_12830)
);

NOR2x1_ASAP7_75t_L g12831 ( 
.A(n_12807),
.B(n_6773),
.Y(n_12831)
);

INVxp67_ASAP7_75t_L g12832 ( 
.A(n_12743),
.Y(n_12832)
);

NAND2xp5_ASAP7_75t_SL g12833 ( 
.A(n_12796),
.B(n_5839),
.Y(n_12833)
);

NAND3xp33_ASAP7_75t_L g12834 ( 
.A(n_12803),
.B(n_3433),
.C(n_6773),
.Y(n_12834)
);

NAND5xp2_ASAP7_75t_L g12835 ( 
.A(n_12778),
.B(n_5104),
.C(n_5095),
.D(n_4727),
.E(n_4825),
.Y(n_12835)
);

AOI221xp5_ASAP7_75t_L g12836 ( 
.A1(n_12799),
.A2(n_6789),
.B1(n_6797),
.B2(n_6784),
.C(n_6783),
.Y(n_12836)
);

NAND2xp5_ASAP7_75t_L g12837 ( 
.A(n_12742),
.B(n_12783),
.Y(n_12837)
);

NOR2xp33_ASAP7_75t_L g12838 ( 
.A(n_12750),
.B(n_5764),
.Y(n_12838)
);

OAI21xp5_ASAP7_75t_L g12839 ( 
.A1(n_12759),
.A2(n_6077),
.B(n_6069),
.Y(n_12839)
);

NOR3xp33_ASAP7_75t_SL g12840 ( 
.A(n_12776),
.B(n_12798),
.C(n_12749),
.Y(n_12840)
);

NAND4xp75_ASAP7_75t_L g12841 ( 
.A(n_12802),
.B(n_12809),
.C(n_12806),
.D(n_12811),
.Y(n_12841)
);

OAI21xp5_ASAP7_75t_L g12842 ( 
.A1(n_12765),
.A2(n_6069),
.B(n_6093),
.Y(n_12842)
);

NOR2xp33_ASAP7_75t_L g12843 ( 
.A(n_12770),
.B(n_5764),
.Y(n_12843)
);

AND2x2_ASAP7_75t_L g12844 ( 
.A(n_12777),
.B(n_12808),
.Y(n_12844)
);

NAND3xp33_ASAP7_75t_L g12845 ( 
.A(n_12762),
.B(n_3433),
.C(n_6784),
.Y(n_12845)
);

AOI21xp33_ASAP7_75t_SL g12846 ( 
.A1(n_12785),
.A2(n_6169),
.B(n_7562),
.Y(n_12846)
);

NAND4xp25_ASAP7_75t_L g12847 ( 
.A(n_12793),
.B(n_3177),
.C(n_4483),
.D(n_4441),
.Y(n_12847)
);

INVx1_ASAP7_75t_L g12848 ( 
.A(n_12767),
.Y(n_12848)
);

AOI211xp5_ASAP7_75t_L g12849 ( 
.A1(n_12756),
.A2(n_3021),
.B(n_3036),
.C(n_3003),
.Y(n_12849)
);

NAND4xp25_ASAP7_75t_L g12850 ( 
.A(n_12773),
.B(n_4509),
.C(n_4531),
.D(n_4441),
.Y(n_12850)
);

NAND4xp25_ASAP7_75t_SL g12851 ( 
.A(n_12791),
.B(n_6797),
.C(n_6789),
.D(n_7334),
.Y(n_12851)
);

AOI33xp33_ASAP7_75t_L g12852 ( 
.A1(n_12740),
.A2(n_4991),
.A3(n_5060),
.B1(n_5129),
.B2(n_4963),
.B3(n_5107),
.Y(n_12852)
);

AND2x4_ASAP7_75t_L g12853 ( 
.A(n_12801),
.B(n_7334),
.Y(n_12853)
);

NOR2x1_ASAP7_75t_L g12854 ( 
.A(n_12773),
.B(n_3003),
.Y(n_12854)
);

INVx1_ASAP7_75t_L g12855 ( 
.A(n_12748),
.Y(n_12855)
);

NAND4xp75_ASAP7_75t_L g12856 ( 
.A(n_12787),
.B(n_6169),
.C(n_7562),
.D(n_6627),
.Y(n_12856)
);

NAND4xp25_ASAP7_75t_L g12857 ( 
.A(n_12812),
.B(n_4531),
.C(n_4560),
.D(n_4509),
.Y(n_12857)
);

NAND2xp5_ASAP7_75t_L g12858 ( 
.A(n_12766),
.B(n_6170),
.Y(n_12858)
);

NAND2xp5_ASAP7_75t_L g12859 ( 
.A(n_12744),
.B(n_6170),
.Y(n_12859)
);

NOR2x1_ASAP7_75t_L g12860 ( 
.A(n_12753),
.B(n_3003),
.Y(n_12860)
);

NAND2xp5_ASAP7_75t_L g12861 ( 
.A(n_12775),
.B(n_12758),
.Y(n_12861)
);

NOR3x1_ASAP7_75t_L g12862 ( 
.A(n_12792),
.B(n_6311),
.C(n_6188),
.Y(n_12862)
);

NOR3xp33_ASAP7_75t_L g12863 ( 
.A(n_12774),
.B(n_6154),
.C(n_6262),
.Y(n_12863)
);

NOR4xp25_ASAP7_75t_L g12864 ( 
.A(n_12760),
.B(n_5060),
.C(n_5129),
.D(n_4991),
.Y(n_12864)
);

NAND3xp33_ASAP7_75t_L g12865 ( 
.A(n_12754),
.B(n_3433),
.C(n_6169),
.Y(n_12865)
);

AOI211xp5_ASAP7_75t_L g12866 ( 
.A1(n_12747),
.A2(n_3021),
.B(n_3036),
.C(n_3003),
.Y(n_12866)
);

NOR3xp33_ASAP7_75t_L g12867 ( 
.A(n_12779),
.B(n_6154),
.C(n_6262),
.Y(n_12867)
);

OAI211xp5_ASAP7_75t_L g12868 ( 
.A1(n_12771),
.A2(n_6169),
.B(n_7562),
.C(n_6627),
.Y(n_12868)
);

OR2x2_ASAP7_75t_L g12869 ( 
.A(n_12751),
.B(n_6170),
.Y(n_12869)
);

OAI211xp5_ASAP7_75t_L g12870 ( 
.A1(n_12781),
.A2(n_6169),
.B(n_7562),
.C(n_6627),
.Y(n_12870)
);

NAND4xp25_ASAP7_75t_L g12871 ( 
.A(n_12782),
.B(n_4531),
.C(n_4560),
.D(n_4509),
.Y(n_12871)
);

OAI21xp33_ASAP7_75t_L g12872 ( 
.A1(n_12745),
.A2(n_5839),
.B(n_5764),
.Y(n_12872)
);

NAND4xp25_ASAP7_75t_L g12873 ( 
.A(n_12768),
.B(n_4531),
.C(n_4560),
.D(n_4509),
.Y(n_12873)
);

NAND4xp25_ASAP7_75t_SL g12874 ( 
.A(n_12786),
.B(n_12797),
.C(n_12795),
.D(n_12746),
.Y(n_12874)
);

AOI221xp5_ASAP7_75t_L g12875 ( 
.A1(n_12794),
.A2(n_5764),
.B1(n_5922),
.B2(n_5839),
.C(n_5129),
.Y(n_12875)
);

AOI211xp5_ASAP7_75t_L g12876 ( 
.A1(n_12780),
.A2(n_3036),
.B(n_3048),
.C(n_3021),
.Y(n_12876)
);

NOR4xp25_ASAP7_75t_L g12877 ( 
.A(n_12741),
.B(n_5060),
.C(n_4560),
.D(n_4705),
.Y(n_12877)
);

NOR4xp25_ASAP7_75t_L g12878 ( 
.A(n_12741),
.B(n_4560),
.C(n_4705),
.D(n_4531),
.Y(n_12878)
);

AOI221xp5_ASAP7_75t_L g12879 ( 
.A1(n_12794),
.A2(n_5922),
.B1(n_5839),
.B2(n_4718),
.C(n_4780),
.Y(n_12879)
);

NAND3xp33_ASAP7_75t_SL g12880 ( 
.A(n_12738),
.B(n_4727),
.C(n_4709),
.Y(n_12880)
);

NAND3xp33_ASAP7_75t_L g12881 ( 
.A(n_12741),
.B(n_3433),
.C(n_6169),
.Y(n_12881)
);

OAI21xp5_ASAP7_75t_L g12882 ( 
.A1(n_12736),
.A2(n_6097),
.B(n_6093),
.Y(n_12882)
);

NAND4xp25_ASAP7_75t_L g12883 ( 
.A(n_12741),
.B(n_4740),
.C(n_4854),
.D(n_4705),
.Y(n_12883)
);

INVx1_ASAP7_75t_L g12884 ( 
.A(n_12737),
.Y(n_12884)
);

INVx2_ASAP7_75t_L g12885 ( 
.A(n_12841),
.Y(n_12885)
);

NOR2x1_ASAP7_75t_L g12886 ( 
.A(n_12826),
.B(n_3021),
.Y(n_12886)
);

OAI22xp5_ASAP7_75t_L g12887 ( 
.A1(n_12881),
.A2(n_5839),
.B1(n_5922),
.B2(n_6609),
.Y(n_12887)
);

NOR2x1_ASAP7_75t_L g12888 ( 
.A(n_12818),
.B(n_3021),
.Y(n_12888)
);

AOI22xp5_ASAP7_75t_L g12889 ( 
.A1(n_12815),
.A2(n_5922),
.B1(n_6627),
.B2(n_6609),
.Y(n_12889)
);

AOI22x1_ASAP7_75t_SL g12890 ( 
.A1(n_12884),
.A2(n_2995),
.B1(n_3026),
.B2(n_2977),
.Y(n_12890)
);

INVx1_ASAP7_75t_L g12891 ( 
.A(n_12828),
.Y(n_12891)
);

INVxp67_ASAP7_75t_L g12892 ( 
.A(n_12816),
.Y(n_12892)
);

AND2x2_ASAP7_75t_L g12893 ( 
.A(n_12833),
.B(n_6170),
.Y(n_12893)
);

AND2x4_ASAP7_75t_L g12894 ( 
.A(n_12832),
.B(n_6531),
.Y(n_12894)
);

HB1xp67_ASAP7_75t_L g12895 ( 
.A(n_12837),
.Y(n_12895)
);

INVx1_ASAP7_75t_L g12896 ( 
.A(n_12861),
.Y(n_12896)
);

NOR2x1_ASAP7_75t_L g12897 ( 
.A(n_12848),
.B(n_3021),
.Y(n_12897)
);

AND2x2_ASAP7_75t_L g12898 ( 
.A(n_12824),
.B(n_6170),
.Y(n_12898)
);

INVxp67_ASAP7_75t_L g12899 ( 
.A(n_12844),
.Y(n_12899)
);

OR2x2_ASAP7_75t_L g12900 ( 
.A(n_12883),
.B(n_6170),
.Y(n_12900)
);

NOR2xp67_ASAP7_75t_L g12901 ( 
.A(n_12874),
.B(n_3021),
.Y(n_12901)
);

INVx1_ASAP7_75t_L g12902 ( 
.A(n_12855),
.Y(n_12902)
);

INVx1_ASAP7_75t_L g12903 ( 
.A(n_12876),
.Y(n_12903)
);

A2O1A1Ixp33_ASAP7_75t_SL g12904 ( 
.A1(n_12843),
.A2(n_2995),
.B(n_3026),
.C(n_2977),
.Y(n_12904)
);

INVx1_ASAP7_75t_L g12905 ( 
.A(n_12840),
.Y(n_12905)
);

INVx1_ASAP7_75t_SL g12906 ( 
.A(n_12822),
.Y(n_12906)
);

AO22x1_ASAP7_75t_L g12907 ( 
.A1(n_12854),
.A2(n_3108),
.B1(n_3021),
.B2(n_3048),
.Y(n_12907)
);

INVx1_ASAP7_75t_L g12908 ( 
.A(n_12860),
.Y(n_12908)
);

INVx1_ASAP7_75t_L g12909 ( 
.A(n_12813),
.Y(n_12909)
);

NAND2xp5_ASAP7_75t_L g12910 ( 
.A(n_12877),
.B(n_6170),
.Y(n_12910)
);

NOR2xp67_ASAP7_75t_L g12911 ( 
.A(n_12851),
.B(n_3021),
.Y(n_12911)
);

NOR2x1_ASAP7_75t_L g12912 ( 
.A(n_12865),
.B(n_3036),
.Y(n_12912)
);

INVx2_ASAP7_75t_L g12913 ( 
.A(n_12831),
.Y(n_12913)
);

INVxp33_ASAP7_75t_SL g12914 ( 
.A(n_12878),
.Y(n_12914)
);

INVx2_ASAP7_75t_L g12915 ( 
.A(n_12858),
.Y(n_12915)
);

INVx1_ASAP7_75t_L g12916 ( 
.A(n_12834),
.Y(n_12916)
);

NOR2x1_ASAP7_75t_L g12917 ( 
.A(n_12873),
.B(n_3036),
.Y(n_12917)
);

INVx1_ASAP7_75t_L g12918 ( 
.A(n_12838),
.Y(n_12918)
);

AND2x2_ASAP7_75t_L g12919 ( 
.A(n_12864),
.B(n_6170),
.Y(n_12919)
);

NOR2x1_ASAP7_75t_L g12920 ( 
.A(n_12845),
.B(n_3036),
.Y(n_12920)
);

AOI211xp5_ASAP7_75t_SL g12921 ( 
.A1(n_12872),
.A2(n_12849),
.B(n_12866),
.C(n_12821),
.Y(n_12921)
);

INVx2_ASAP7_75t_L g12922 ( 
.A(n_12869),
.Y(n_12922)
);

NAND2xp5_ASAP7_75t_L g12923 ( 
.A(n_12829),
.B(n_6207),
.Y(n_12923)
);

INVx2_ASAP7_75t_L g12924 ( 
.A(n_12862),
.Y(n_12924)
);

INVx1_ASAP7_75t_L g12925 ( 
.A(n_12817),
.Y(n_12925)
);

OR2x2_ASAP7_75t_L g12926 ( 
.A(n_12850),
.B(n_6207),
.Y(n_12926)
);

NOR2x1_ASAP7_75t_L g12927 ( 
.A(n_12857),
.B(n_3036),
.Y(n_12927)
);

INVx1_ASAP7_75t_L g12928 ( 
.A(n_12847),
.Y(n_12928)
);

AOI22xp5_ASAP7_75t_L g12929 ( 
.A1(n_12863),
.A2(n_5922),
.B1(n_6627),
.B2(n_6609),
.Y(n_12929)
);

INVx1_ASAP7_75t_L g12930 ( 
.A(n_12859),
.Y(n_12930)
);

AND3x4_ASAP7_75t_L g12931 ( 
.A(n_12867),
.B(n_3336),
.C(n_3326),
.Y(n_12931)
);

NOR2xp33_ASAP7_75t_L g12932 ( 
.A(n_12871),
.B(n_3165),
.Y(n_12932)
);

INVx2_ASAP7_75t_L g12933 ( 
.A(n_12853),
.Y(n_12933)
);

AOI22xp5_ASAP7_75t_L g12934 ( 
.A1(n_12820),
.A2(n_5922),
.B1(n_6627),
.B2(n_6609),
.Y(n_12934)
);

AOI22xp5_ASAP7_75t_L g12935 ( 
.A1(n_12870),
.A2(n_6609),
.B1(n_6696),
.B2(n_6679),
.Y(n_12935)
);

OR2x2_ASAP7_75t_L g12936 ( 
.A(n_12835),
.B(n_6207),
.Y(n_12936)
);

AND2x2_ASAP7_75t_L g12937 ( 
.A(n_12852),
.B(n_6531),
.Y(n_12937)
);

INVx2_ASAP7_75t_L g12938 ( 
.A(n_12853),
.Y(n_12938)
);

INVx1_ASAP7_75t_L g12939 ( 
.A(n_12846),
.Y(n_12939)
);

INVx2_ASAP7_75t_L g12940 ( 
.A(n_12842),
.Y(n_12940)
);

NAND4xp75_ASAP7_75t_L g12941 ( 
.A(n_12905),
.B(n_12875),
.C(n_12879),
.D(n_12839),
.Y(n_12941)
);

NAND3x2_ASAP7_75t_L g12942 ( 
.A(n_12909),
.B(n_12880),
.C(n_12868),
.Y(n_12942)
);

NAND4xp25_ASAP7_75t_L g12943 ( 
.A(n_12901),
.B(n_12882),
.C(n_12825),
.D(n_12814),
.Y(n_12943)
);

NOR3xp33_ASAP7_75t_L g12944 ( 
.A(n_12892),
.B(n_12830),
.C(n_12827),
.Y(n_12944)
);

INVx2_ASAP7_75t_L g12945 ( 
.A(n_12888),
.Y(n_12945)
);

INVx1_ASAP7_75t_L g12946 ( 
.A(n_12897),
.Y(n_12946)
);

NAND4xp25_ASAP7_75t_SL g12947 ( 
.A(n_12885),
.B(n_12823),
.C(n_12819),
.D(n_12836),
.Y(n_12947)
);

NAND4xp75_ASAP7_75t_L g12948 ( 
.A(n_12902),
.B(n_12856),
.C(n_6609),
.D(n_6225),
.Y(n_12948)
);

NAND3xp33_ASAP7_75t_SL g12949 ( 
.A(n_12906),
.B(n_4727),
.C(n_4709),
.Y(n_12949)
);

NOR3xp33_ASAP7_75t_L g12950 ( 
.A(n_12899),
.B(n_3026),
.C(n_2995),
.Y(n_12950)
);

NAND2xp5_ASAP7_75t_L g12951 ( 
.A(n_12898),
.B(n_6207),
.Y(n_12951)
);

NOR4xp25_ASAP7_75t_L g12952 ( 
.A(n_12924),
.B(n_4740),
.C(n_4854),
.D(n_4705),
.Y(n_12952)
);

NOR4xp25_ASAP7_75t_L g12953 ( 
.A(n_12896),
.B(n_4740),
.C(n_4854),
.D(n_4705),
.Y(n_12953)
);

NAND3xp33_ASAP7_75t_L g12954 ( 
.A(n_12895),
.B(n_3433),
.C(n_3048),
.Y(n_12954)
);

NOR2xp33_ASAP7_75t_SL g12955 ( 
.A(n_12891),
.B(n_3036),
.Y(n_12955)
);

NAND4xp25_ASAP7_75t_L g12956 ( 
.A(n_12886),
.B(n_12928),
.C(n_12921),
.D(n_12918),
.Y(n_12956)
);

NAND2xp5_ASAP7_75t_L g12957 ( 
.A(n_12914),
.B(n_6207),
.Y(n_12957)
);

NOR3xp33_ASAP7_75t_L g12958 ( 
.A(n_12922),
.B(n_3026),
.C(n_2995),
.Y(n_12958)
);

NOR2x1_ASAP7_75t_L g12959 ( 
.A(n_12913),
.B(n_3036),
.Y(n_12959)
);

NOR3xp33_ASAP7_75t_L g12960 ( 
.A(n_12930),
.B(n_3054),
.C(n_3026),
.Y(n_12960)
);

NOR2xp33_ASAP7_75t_L g12961 ( 
.A(n_12925),
.B(n_12903),
.Y(n_12961)
);

NAND4xp25_ASAP7_75t_L g12962 ( 
.A(n_12908),
.B(n_4854),
.C(n_4889),
.D(n_4740),
.Y(n_12962)
);

NOR2x1p5_ASAP7_75t_L g12963 ( 
.A(n_12940),
.B(n_3036),
.Y(n_12963)
);

NAND3xp33_ASAP7_75t_SL g12964 ( 
.A(n_12915),
.B(n_4727),
.C(n_4709),
.Y(n_12964)
);

NAND4xp75_ASAP7_75t_L g12965 ( 
.A(n_12933),
.B(n_6265),
.C(n_6696),
.D(n_6327),
.Y(n_12965)
);

NOR5xp2_ASAP7_75t_L g12966 ( 
.A(n_12939),
.B(n_6307),
.C(n_6592),
.D(n_6312),
.E(n_6034),
.Y(n_12966)
);

NAND5xp2_ASAP7_75t_L g12967 ( 
.A(n_12916),
.B(n_4825),
.C(n_4709),
.D(n_6207),
.E(n_3076),
.Y(n_12967)
);

INVx1_ASAP7_75t_L g12968 ( 
.A(n_12938),
.Y(n_12968)
);

NOR2x1_ASAP7_75t_L g12969 ( 
.A(n_12911),
.B(n_3048),
.Y(n_12969)
);

AND2x2_ASAP7_75t_L g12970 ( 
.A(n_12932),
.B(n_6531),
.Y(n_12970)
);

NOR3xp33_ASAP7_75t_L g12971 ( 
.A(n_12920),
.B(n_3058),
.C(n_3054),
.Y(n_12971)
);

NOR3xp33_ASAP7_75t_L g12972 ( 
.A(n_12912),
.B(n_3058),
.C(n_3054),
.Y(n_12972)
);

NOR2x1_ASAP7_75t_L g12973 ( 
.A(n_12917),
.B(n_3048),
.Y(n_12973)
);

NOR2x1p5_ASAP7_75t_L g12974 ( 
.A(n_12936),
.B(n_3048),
.Y(n_12974)
);

NAND2xp5_ASAP7_75t_SL g12975 ( 
.A(n_12927),
.B(n_3048),
.Y(n_12975)
);

NAND3x1_ASAP7_75t_SL g12976 ( 
.A(n_12893),
.B(n_6312),
.C(n_6307),
.Y(n_12976)
);

OR2x2_ASAP7_75t_L g12977 ( 
.A(n_12900),
.B(n_6207),
.Y(n_12977)
);

AND4x1_ASAP7_75t_L g12978 ( 
.A(n_12937),
.B(n_6312),
.C(n_6592),
.D(n_6307),
.Y(n_12978)
);

NAND4xp25_ASAP7_75t_L g12979 ( 
.A(n_12904),
.B(n_4854),
.C(n_4889),
.D(n_4740),
.Y(n_12979)
);

NOR4xp25_ASAP7_75t_L g12980 ( 
.A(n_12910),
.B(n_4948),
.C(n_5041),
.D(n_4889),
.Y(n_12980)
);

NOR3xp33_ASAP7_75t_L g12981 ( 
.A(n_12907),
.B(n_3058),
.C(n_3054),
.Y(n_12981)
);

NAND4xp25_ASAP7_75t_L g12982 ( 
.A(n_12923),
.B(n_4948),
.C(n_5041),
.D(n_4889),
.Y(n_12982)
);

INVx1_ASAP7_75t_L g12983 ( 
.A(n_12931),
.Y(n_12983)
);

INVx1_ASAP7_75t_L g12984 ( 
.A(n_12890),
.Y(n_12984)
);

NOR2x1_ASAP7_75t_L g12985 ( 
.A(n_12919),
.B(n_3048),
.Y(n_12985)
);

NAND2xp5_ASAP7_75t_L g12986 ( 
.A(n_12926),
.B(n_6207),
.Y(n_12986)
);

OR2x2_ASAP7_75t_L g12987 ( 
.A(n_12929),
.B(n_6531),
.Y(n_12987)
);

INVx2_ASAP7_75t_L g12988 ( 
.A(n_12887),
.Y(n_12988)
);

AOI21xp5_ASAP7_75t_L g12989 ( 
.A1(n_12968),
.A2(n_12934),
.B(n_12889),
.Y(n_12989)
);

NOR4xp75_ASAP7_75t_SL g12990 ( 
.A(n_12956),
.B(n_12935),
.C(n_12894),
.D(n_6312),
.Y(n_12990)
);

INVx2_ASAP7_75t_SL g12991 ( 
.A(n_12974),
.Y(n_12991)
);

NOR2xp33_ASAP7_75t_L g12992 ( 
.A(n_12943),
.B(n_12894),
.Y(n_12992)
);

INVx2_ASAP7_75t_L g12993 ( 
.A(n_12963),
.Y(n_12993)
);

NAND2xp5_ASAP7_75t_L g12994 ( 
.A(n_12955),
.B(n_6531),
.Y(n_12994)
);

NAND4xp25_ASAP7_75t_L g12995 ( 
.A(n_12961),
.B(n_3054),
.C(n_3079),
.D(n_3058),
.Y(n_12995)
);

NAND4xp75_ASAP7_75t_L g12996 ( 
.A(n_12946),
.B(n_6327),
.C(n_6381),
.D(n_6696),
.Y(n_12996)
);

NAND2xp5_ASAP7_75t_L g12997 ( 
.A(n_12944),
.B(n_6531),
.Y(n_12997)
);

OAI221xp5_ASAP7_75t_L g12998 ( 
.A1(n_12988),
.A2(n_3076),
.B1(n_3075),
.B2(n_3048),
.C(n_3407),
.Y(n_12998)
);

OAI22xp33_ASAP7_75t_L g12999 ( 
.A1(n_12957),
.A2(n_3075),
.B1(n_3076),
.B2(n_3048),
.Y(n_12999)
);

O2A1O1Ixp33_ASAP7_75t_L g13000 ( 
.A1(n_12945),
.A2(n_3058),
.B(n_3079),
.C(n_3054),
.Y(n_13000)
);

NAND3xp33_ASAP7_75t_SL g13001 ( 
.A(n_12984),
.B(n_4825),
.C(n_5687),
.Y(n_13001)
);

AND3x4_ASAP7_75t_L g13002 ( 
.A(n_12985),
.B(n_3336),
.C(n_3326),
.Y(n_13002)
);

NAND4xp25_ASAP7_75t_L g13003 ( 
.A(n_12983),
.B(n_3079),
.C(n_3096),
.D(n_3058),
.Y(n_13003)
);

INVx1_ASAP7_75t_L g13004 ( 
.A(n_12959),
.Y(n_13004)
);

OR2x2_ASAP7_75t_L g13005 ( 
.A(n_12942),
.B(n_6531),
.Y(n_13005)
);

AND2x2_ASAP7_75t_L g13006 ( 
.A(n_12969),
.B(n_6531),
.Y(n_13006)
);

NAND2xp5_ASAP7_75t_L g13007 ( 
.A(n_12973),
.B(n_6326),
.Y(n_13007)
);

AOI22xp33_ASAP7_75t_SL g13008 ( 
.A1(n_12954),
.A2(n_3076),
.B1(n_3075),
.B2(n_3407),
.Y(n_13008)
);

NAND2x1p5_ASAP7_75t_L g13009 ( 
.A(n_12975),
.B(n_3075),
.Y(n_13009)
);

NAND2xp5_ASAP7_75t_L g13010 ( 
.A(n_12941),
.B(n_6326),
.Y(n_13010)
);

NAND5xp2_ASAP7_75t_L g13011 ( 
.A(n_12960),
.B(n_4825),
.C(n_3076),
.D(n_3075),
.E(n_6630),
.Y(n_13011)
);

OAI211xp5_ASAP7_75t_SL g13012 ( 
.A1(n_12947),
.A2(n_3096),
.B(n_3107),
.C(n_3079),
.Y(n_13012)
);

OR2x2_ASAP7_75t_L g13013 ( 
.A(n_12982),
.B(n_6326),
.Y(n_13013)
);

INVx2_ASAP7_75t_L g13014 ( 
.A(n_12986),
.Y(n_13014)
);

INVx1_ASAP7_75t_L g13015 ( 
.A(n_12950),
.Y(n_13015)
);

OR2x6_ASAP7_75t_L g13016 ( 
.A(n_12951),
.B(n_3075),
.Y(n_13016)
);

AOI21xp5_ASAP7_75t_L g13017 ( 
.A1(n_12980),
.A2(n_6210),
.B(n_6441),
.Y(n_13017)
);

INVx1_ASAP7_75t_L g13018 ( 
.A(n_12958),
.Y(n_13018)
);

OR2x2_ASAP7_75t_L g13019 ( 
.A(n_12952),
.B(n_6326),
.Y(n_13019)
);

BUFx10_ASAP7_75t_L g13020 ( 
.A(n_12971),
.Y(n_13020)
);

NAND4xp25_ASAP7_75t_L g13021 ( 
.A(n_12972),
.B(n_3096),
.C(n_3107),
.D(n_3079),
.Y(n_13021)
);

INVx1_ASAP7_75t_SL g13022 ( 
.A(n_12970),
.Y(n_13022)
);

NOR2xp67_ASAP7_75t_L g13023 ( 
.A(n_12979),
.B(n_3075),
.Y(n_13023)
);

NAND2xp5_ASAP7_75t_L g13024 ( 
.A(n_12981),
.B(n_6326),
.Y(n_13024)
);

NOR2x1_ASAP7_75t_L g13025 ( 
.A(n_12948),
.B(n_3075),
.Y(n_13025)
);

AOI22xp5_ASAP7_75t_L g13026 ( 
.A1(n_12992),
.A2(n_12962),
.B1(n_12949),
.B2(n_12964),
.Y(n_13026)
);

NAND4xp25_ASAP7_75t_L g13027 ( 
.A(n_12989),
.B(n_12987),
.C(n_12977),
.D(n_12967),
.Y(n_13027)
);

INVx2_ASAP7_75t_L g13028 ( 
.A(n_13009),
.Y(n_13028)
);

NAND4xp25_ASAP7_75t_L g13029 ( 
.A(n_13022),
.B(n_12966),
.C(n_12953),
.D(n_12976),
.Y(n_13029)
);

NAND2x1p5_ASAP7_75t_L g13030 ( 
.A(n_13004),
.B(n_12978),
.Y(n_13030)
);

INVx1_ASAP7_75t_L g13031 ( 
.A(n_12993),
.Y(n_13031)
);

NAND2xp5_ASAP7_75t_SL g13032 ( 
.A(n_12990),
.B(n_12965),
.Y(n_13032)
);

HB1xp67_ASAP7_75t_L g13033 ( 
.A(n_13016),
.Y(n_13033)
);

NOR3xp33_ASAP7_75t_L g13034 ( 
.A(n_13014),
.B(n_3096),
.C(n_3079),
.Y(n_13034)
);

NAND4xp75_ASAP7_75t_L g13035 ( 
.A(n_12991),
.B(n_6327),
.C(n_6381),
.D(n_6607),
.Y(n_13035)
);

NAND4xp75_ASAP7_75t_L g13036 ( 
.A(n_13010),
.B(n_6327),
.C(n_6381),
.D(n_6607),
.Y(n_13036)
);

OR2x2_ASAP7_75t_L g13037 ( 
.A(n_13005),
.B(n_6326),
.Y(n_13037)
);

NOR2x1_ASAP7_75t_L g13038 ( 
.A(n_13016),
.B(n_3075),
.Y(n_13038)
);

INVx1_ASAP7_75t_L g13039 ( 
.A(n_13018),
.Y(n_13039)
);

INVx1_ASAP7_75t_SL g13040 ( 
.A(n_13020),
.Y(n_13040)
);

AND3x4_ASAP7_75t_L g13041 ( 
.A(n_13025),
.B(n_3336),
.C(n_3326),
.Y(n_13041)
);

HB1xp67_ASAP7_75t_L g13042 ( 
.A(n_13015),
.Y(n_13042)
);

NAND2xp5_ASAP7_75t_L g13043 ( 
.A(n_12997),
.B(n_6326),
.Y(n_13043)
);

BUFx4f_ASAP7_75t_SL g13044 ( 
.A(n_13002),
.Y(n_13044)
);

INVx1_ASAP7_75t_L g13045 ( 
.A(n_13023),
.Y(n_13045)
);

XOR2x1_ASAP7_75t_L g13046 ( 
.A(n_12999),
.B(n_13006),
.Y(n_13046)
);

NOR3xp33_ASAP7_75t_L g13047 ( 
.A(n_13012),
.B(n_3107),
.C(n_3096),
.Y(n_13047)
);

NAND2xp5_ASAP7_75t_L g13048 ( 
.A(n_13008),
.B(n_6326),
.Y(n_13048)
);

INVx2_ASAP7_75t_L g13049 ( 
.A(n_13013),
.Y(n_13049)
);

AND4x2_ASAP7_75t_L g13050 ( 
.A(n_12998),
.B(n_6307),
.C(n_6592),
.D(n_6312),
.Y(n_13050)
);

INVx1_ASAP7_75t_L g13051 ( 
.A(n_13007),
.Y(n_13051)
);

AND3x4_ASAP7_75t_L g13052 ( 
.A(n_13021),
.B(n_3336),
.C(n_3326),
.Y(n_13052)
);

NOR3xp33_ASAP7_75t_L g13053 ( 
.A(n_13001),
.B(n_3107),
.C(n_3096),
.Y(n_13053)
);

NOR3xp33_ASAP7_75t_L g13054 ( 
.A(n_13003),
.B(n_3107),
.C(n_3096),
.Y(n_13054)
);

NAND2x1p5_ASAP7_75t_L g13055 ( 
.A(n_13019),
.B(n_3076),
.Y(n_13055)
);

NOR3xp33_ASAP7_75t_L g13056 ( 
.A(n_12995),
.B(n_3131),
.C(n_3107),
.Y(n_13056)
);

NAND2x1p5_ASAP7_75t_L g13057 ( 
.A(n_12994),
.B(n_3076),
.Y(n_13057)
);

INVx2_ASAP7_75t_L g13058 ( 
.A(n_13024),
.Y(n_13058)
);

AND2x2_ASAP7_75t_L g13059 ( 
.A(n_13000),
.B(n_6307),
.Y(n_13059)
);

NOR2xp67_ASAP7_75t_L g13060 ( 
.A(n_13011),
.B(n_3076),
.Y(n_13060)
);

NOR2xp67_ASAP7_75t_SL g13061 ( 
.A(n_13017),
.B(n_12996),
.Y(n_13061)
);

NAND4xp25_ASAP7_75t_L g13062 ( 
.A(n_12992),
.B(n_3107),
.C(n_3140),
.D(n_3131),
.Y(n_13062)
);

AND2x4_ASAP7_75t_SL g13063 ( 
.A(n_13020),
.B(n_3076),
.Y(n_13063)
);

NOR2xp67_ASAP7_75t_SL g13064 ( 
.A(n_13014),
.B(n_3076),
.Y(n_13064)
);

NAND2xp5_ASAP7_75t_L g13065 ( 
.A(n_12993),
.B(n_6034),
.Y(n_13065)
);

INVx1_ASAP7_75t_L g13066 ( 
.A(n_13055),
.Y(n_13066)
);

BUFx3_ASAP7_75t_L g13067 ( 
.A(n_13030),
.Y(n_13067)
);

BUFx2_ASAP7_75t_L g13068 ( 
.A(n_13033),
.Y(n_13068)
);

INVx2_ASAP7_75t_L g13069 ( 
.A(n_13057),
.Y(n_13069)
);

INVx1_ASAP7_75t_L g13070 ( 
.A(n_13038),
.Y(n_13070)
);

HB1xp67_ASAP7_75t_L g13071 ( 
.A(n_13028),
.Y(n_13071)
);

AND3x1_ASAP7_75t_L g13072 ( 
.A(n_13031),
.B(n_3140),
.C(n_3131),
.Y(n_13072)
);

AND2x4_ASAP7_75t_L g13073 ( 
.A(n_13060),
.B(n_3407),
.Y(n_13073)
);

INVxp33_ASAP7_75t_SL g13074 ( 
.A(n_13042),
.Y(n_13074)
);

OR3x1_ASAP7_75t_L g13075 ( 
.A(n_13027),
.B(n_13029),
.C(n_13045),
.Y(n_13075)
);

AND2x4_ASAP7_75t_L g13076 ( 
.A(n_13063),
.B(n_3407),
.Y(n_13076)
);

AND2x4_ASAP7_75t_L g13077 ( 
.A(n_13039),
.B(n_3407),
.Y(n_13077)
);

AOI22xp5_ASAP7_75t_L g13078 ( 
.A1(n_13040),
.A2(n_6324),
.B1(n_6322),
.B2(n_3411),
.Y(n_13078)
);

INVx2_ASAP7_75t_L g13079 ( 
.A(n_13046),
.Y(n_13079)
);

INVx3_ASAP7_75t_SL g13080 ( 
.A(n_13049),
.Y(n_13080)
);

INVx1_ASAP7_75t_L g13081 ( 
.A(n_13032),
.Y(n_13081)
);

AND2x2_ASAP7_75t_L g13082 ( 
.A(n_13026),
.B(n_6307),
.Y(n_13082)
);

INVxp67_ASAP7_75t_SL g13083 ( 
.A(n_13058),
.Y(n_13083)
);

INVx1_ASAP7_75t_L g13084 ( 
.A(n_13061),
.Y(n_13084)
);

AOI22xp5_ASAP7_75t_L g13085 ( 
.A1(n_13044),
.A2(n_6324),
.B1(n_6322),
.B2(n_3411),
.Y(n_13085)
);

OA22x2_ASAP7_75t_L g13086 ( 
.A1(n_13051),
.A2(n_6749),
.B1(n_6048),
.B2(n_6045),
.Y(n_13086)
);

INVx1_ASAP7_75t_L g13087 ( 
.A(n_13064),
.Y(n_13087)
);

OR3x2_ASAP7_75t_L g13088 ( 
.A(n_13062),
.B(n_5447),
.C(n_5441),
.Y(n_13088)
);

INVx1_ASAP7_75t_L g13089 ( 
.A(n_13041),
.Y(n_13089)
);

INVxp67_ASAP7_75t_L g13090 ( 
.A(n_13065),
.Y(n_13090)
);

INVx2_ASAP7_75t_L g13091 ( 
.A(n_13043),
.Y(n_13091)
);

INVx1_ASAP7_75t_L g13092 ( 
.A(n_13052),
.Y(n_13092)
);

INVx1_ASAP7_75t_L g13093 ( 
.A(n_13053),
.Y(n_13093)
);

INVx1_ASAP7_75t_L g13094 ( 
.A(n_13034),
.Y(n_13094)
);

NAND2x1_ASAP7_75t_L g13095 ( 
.A(n_13068),
.B(n_13048),
.Y(n_13095)
);

AOI22xp33_ASAP7_75t_SL g13096 ( 
.A1(n_13074),
.A2(n_13059),
.B1(n_13037),
.B2(n_13047),
.Y(n_13096)
);

AOI21x1_ASAP7_75t_L g13097 ( 
.A1(n_13068),
.A2(n_13050),
.B(n_13054),
.Y(n_13097)
);

XNOR2xp5_ASAP7_75t_L g13098 ( 
.A(n_13075),
.B(n_13071),
.Y(n_13098)
);

INVx2_ASAP7_75t_L g13099 ( 
.A(n_13067),
.Y(n_13099)
);

HB1xp67_ASAP7_75t_L g13100 ( 
.A(n_13079),
.Y(n_13100)
);

INVx1_ASAP7_75t_L g13101 ( 
.A(n_13081),
.Y(n_13101)
);

AND2x4_ASAP7_75t_L g13102 ( 
.A(n_13077),
.B(n_13056),
.Y(n_13102)
);

INVx2_ASAP7_75t_L g13103 ( 
.A(n_13069),
.Y(n_13103)
);

AOI22xp5_ASAP7_75t_L g13104 ( 
.A1(n_13084),
.A2(n_13036),
.B1(n_13035),
.B2(n_3407),
.Y(n_13104)
);

INVx3_ASAP7_75t_L g13105 ( 
.A(n_13073),
.Y(n_13105)
);

BUFx6f_ASAP7_75t_L g13106 ( 
.A(n_13080),
.Y(n_13106)
);

INVx1_ASAP7_75t_L g13107 ( 
.A(n_13087),
.Y(n_13107)
);

XNOR2xp5_ASAP7_75t_L g13108 ( 
.A(n_13092),
.B(n_3326),
.Y(n_13108)
);

AND2x4_ASAP7_75t_L g13109 ( 
.A(n_13083),
.B(n_3407),
.Y(n_13109)
);

INVx2_ASAP7_75t_L g13110 ( 
.A(n_13070),
.Y(n_13110)
);

NAND2xp5_ASAP7_75t_L g13111 ( 
.A(n_13089),
.B(n_6034),
.Y(n_13111)
);

AND2x4_ASAP7_75t_L g13112 ( 
.A(n_13066),
.B(n_3407),
.Y(n_13112)
);

INVx2_ASAP7_75t_L g13113 ( 
.A(n_13091),
.Y(n_13113)
);

OAI22xp5_ASAP7_75t_L g13114 ( 
.A1(n_13090),
.A2(n_3421),
.B1(n_3411),
.B2(n_3333),
.Y(n_13114)
);

BUFx2_ASAP7_75t_L g13115 ( 
.A(n_13093),
.Y(n_13115)
);

INVx3_ASAP7_75t_L g13116 ( 
.A(n_13094),
.Y(n_13116)
);

INVx2_ASAP7_75t_L g13117 ( 
.A(n_13076),
.Y(n_13117)
);

NAND3xp33_ASAP7_75t_L g13118 ( 
.A(n_13072),
.B(n_3421),
.C(n_3411),
.Y(n_13118)
);

AND2x2_ASAP7_75t_L g13119 ( 
.A(n_13099),
.B(n_13082),
.Y(n_13119)
);

AOI22xp5_ASAP7_75t_L g13120 ( 
.A1(n_13101),
.A2(n_13088),
.B1(n_13078),
.B2(n_13085),
.Y(n_13120)
);

INVx2_ASAP7_75t_L g13121 ( 
.A(n_13109),
.Y(n_13121)
);

INVx1_ASAP7_75t_L g13122 ( 
.A(n_13100),
.Y(n_13122)
);

AOI22xp5_ASAP7_75t_L g13123 ( 
.A1(n_13098),
.A2(n_13086),
.B1(n_3411),
.B2(n_3421),
.Y(n_13123)
);

INVx1_ASAP7_75t_L g13124 ( 
.A(n_13106),
.Y(n_13124)
);

INVx2_ASAP7_75t_L g13125 ( 
.A(n_13106),
.Y(n_13125)
);

NAND2xp5_ASAP7_75t_L g13126 ( 
.A(n_13105),
.B(n_6034),
.Y(n_13126)
);

NOR2xp67_ASAP7_75t_L g13127 ( 
.A(n_13103),
.B(n_3411),
.Y(n_13127)
);

XOR2xp5_ASAP7_75t_L g13128 ( 
.A(n_13107),
.B(n_13115),
.Y(n_13128)
);

INVx1_ASAP7_75t_L g13129 ( 
.A(n_13095),
.Y(n_13129)
);

INVx2_ASAP7_75t_L g13130 ( 
.A(n_13110),
.Y(n_13130)
);

AND2x4_ASAP7_75t_L g13131 ( 
.A(n_13112),
.B(n_13113),
.Y(n_13131)
);

NAND2xp5_ASAP7_75t_L g13132 ( 
.A(n_13117),
.B(n_6034),
.Y(n_13132)
);

BUFx2_ASAP7_75t_L g13133 ( 
.A(n_13122),
.Y(n_13133)
);

AOI22xp5_ASAP7_75t_L g13134 ( 
.A1(n_13130),
.A2(n_13116),
.B1(n_13102),
.B2(n_13096),
.Y(n_13134)
);

OAI22xp5_ASAP7_75t_SL g13135 ( 
.A1(n_13128),
.A2(n_13104),
.B1(n_13108),
.B2(n_13097),
.Y(n_13135)
);

BUFx2_ASAP7_75t_L g13136 ( 
.A(n_13129),
.Y(n_13136)
);

OAI22xp5_ASAP7_75t_L g13137 ( 
.A1(n_13124),
.A2(n_13123),
.B1(n_13125),
.B2(n_13120),
.Y(n_13137)
);

NAND2x1_ASAP7_75t_L g13138 ( 
.A(n_13131),
.B(n_13111),
.Y(n_13138)
);

OAI22xp5_ASAP7_75t_L g13139 ( 
.A1(n_13127),
.A2(n_13118),
.B1(n_13114),
.B2(n_3421),
.Y(n_13139)
);

NAND2xp5_ASAP7_75t_L g13140 ( 
.A(n_13121),
.B(n_6034),
.Y(n_13140)
);

XNOR2xp5_ASAP7_75t_L g13141 ( 
.A(n_13119),
.B(n_3326),
.Y(n_13141)
);

OAI22xp5_ASAP7_75t_L g13142 ( 
.A1(n_13132),
.A2(n_3421),
.B1(n_3411),
.B2(n_3333),
.Y(n_13142)
);

OA22x2_ASAP7_75t_L g13143 ( 
.A1(n_13126),
.A2(n_6749),
.B1(n_6048),
.B2(n_6045),
.Y(n_13143)
);

OAI21xp5_ASAP7_75t_SL g13144 ( 
.A1(n_13134),
.A2(n_3421),
.B(n_3411),
.Y(n_13144)
);

AOI21xp5_ASAP7_75t_L g13145 ( 
.A1(n_13136),
.A2(n_3421),
.B(n_6210),
.Y(n_13145)
);

OAI21xp5_ASAP7_75t_L g13146 ( 
.A1(n_13133),
.A2(n_6154),
.B(n_6210),
.Y(n_13146)
);

OAI22x1_ASAP7_75t_L g13147 ( 
.A1(n_13141),
.A2(n_13135),
.B1(n_13138),
.B2(n_13137),
.Y(n_13147)
);

NAND4xp25_ASAP7_75t_L g13148 ( 
.A(n_13139),
.B(n_3131),
.C(n_3162),
.D(n_3140),
.Y(n_13148)
);

AO21x1_ASAP7_75t_L g13149 ( 
.A1(n_13140),
.A2(n_6749),
.B(n_3341),
.Y(n_13149)
);

AOI21x1_ASAP7_75t_L g13150 ( 
.A1(n_13142),
.A2(n_6687),
.B(n_6747),
.Y(n_13150)
);

OAI22xp5_ASAP7_75t_L g13151 ( 
.A1(n_13144),
.A2(n_13143),
.B1(n_3421),
.B2(n_3333),
.Y(n_13151)
);

INVx2_ASAP7_75t_L g13152 ( 
.A(n_13147),
.Y(n_13152)
);

NOR2x1_ASAP7_75t_L g13153 ( 
.A(n_13148),
.B(n_3421),
.Y(n_13153)
);

XNOR2xp5_ASAP7_75t_L g13154 ( 
.A(n_13152),
.B(n_13149),
.Y(n_13154)
);

HB1xp67_ASAP7_75t_L g13155 ( 
.A(n_13153),
.Y(n_13155)
);

OAI221xp5_ASAP7_75t_L g13156 ( 
.A1(n_13154),
.A2(n_13151),
.B1(n_13146),
.B2(n_13145),
.C(n_13150),
.Y(n_13156)
);

INVx1_ASAP7_75t_L g13157 ( 
.A(n_13156),
.Y(n_13157)
);

OAI21xp5_ASAP7_75t_L g13158 ( 
.A1(n_13157),
.A2(n_13155),
.B(n_6097),
.Y(n_13158)
);

INVx1_ASAP7_75t_L g13159 ( 
.A(n_13158),
.Y(n_13159)
);

NOR2x1p5_ASAP7_75t_SL g13160 ( 
.A(n_13159),
.B(n_5441),
.Y(n_13160)
);

OAI221xp5_ASAP7_75t_R g13161 ( 
.A1(n_13160),
.A2(n_6592),
.B1(n_6312),
.B2(n_6307),
.C(n_6034),
.Y(n_13161)
);

AOI21xp33_ASAP7_75t_SL g13162 ( 
.A1(n_13161),
.A2(n_6607),
.B(n_3140),
.Y(n_13162)
);

AOI211xp5_ASAP7_75t_L g13163 ( 
.A1(n_13162),
.A2(n_3421),
.B(n_3333),
.C(n_3338),
.Y(n_13163)
);


endmodule