module fake_aes_8607_n_791 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_791);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_791;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g103 ( .A(n_72), .Y(n_103) );
BUFx10_ASAP7_75t_L g104 ( .A(n_89), .Y(n_104) );
BUFx6f_ASAP7_75t_L g105 ( .A(n_70), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_2), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_66), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_43), .Y(n_108) );
INVx1_ASAP7_75t_SL g109 ( .A(n_68), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_59), .Y(n_110) );
BUFx6f_ASAP7_75t_L g111 ( .A(n_34), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_3), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_41), .Y(n_113) );
INVxp67_ASAP7_75t_L g114 ( .A(n_49), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_38), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_14), .Y(n_116) );
INVx2_ASAP7_75t_SL g117 ( .A(n_19), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_15), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_27), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_98), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_42), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_94), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_44), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_11), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_4), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_57), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_17), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_97), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_93), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_20), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_39), .Y(n_131) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_50), .Y(n_132) );
INVxp67_ASAP7_75t_L g133 ( .A(n_4), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_51), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_65), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_25), .Y(n_136) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_86), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_77), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_74), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_1), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_33), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_105), .Y(n_142) );
INVx5_ASAP7_75t_L g143 ( .A(n_105), .Y(n_143) );
BUFx8_ASAP7_75t_SL g144 ( .A(n_119), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_103), .Y(n_145) );
BUFx2_ASAP7_75t_L g146 ( .A(n_106), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_105), .Y(n_147) );
BUFx3_ASAP7_75t_L g148 ( .A(n_117), .Y(n_148) );
HB1xp67_ASAP7_75t_L g149 ( .A(n_133), .Y(n_149) );
BUFx12f_ASAP7_75t_L g150 ( .A(n_104), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_107), .Y(n_151) );
AOI22x1_ASAP7_75t_SL g152 ( .A1(n_119), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_152) );
HB1xp67_ASAP7_75t_L g153 ( .A(n_112), .Y(n_153) );
AND2x4_ASAP7_75t_L g154 ( .A(n_136), .B(n_118), .Y(n_154) );
HB1xp67_ASAP7_75t_L g155 ( .A(n_116), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_105), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_111), .Y(n_157) );
AND2x4_ASAP7_75t_L g158 ( .A(n_136), .B(n_0), .Y(n_158) );
AND2x4_ASAP7_75t_L g159 ( .A(n_125), .B(n_3), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_108), .Y(n_160) );
AND2x2_ASAP7_75t_L g161 ( .A(n_104), .B(n_5), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_110), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_123), .Y(n_163) );
INVx6_ASAP7_75t_L g164 ( .A(n_111), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_128), .Y(n_165) );
INVx3_ASAP7_75t_L g166 ( .A(n_111), .Y(n_166) );
BUFx3_ASAP7_75t_L g167 ( .A(n_130), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_111), .Y(n_168) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_144), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g170 ( .A(n_150), .Y(n_170) );
INVx1_ASAP7_75t_SL g171 ( .A(n_146), .Y(n_171) );
INVxp67_ASAP7_75t_L g172 ( .A(n_146), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_150), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_158), .Y(n_174) );
HB1xp67_ASAP7_75t_L g175 ( .A(n_153), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_166), .Y(n_176) );
CKINVDCx20_ASAP7_75t_R g177 ( .A(n_155), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_149), .Y(n_178) );
CKINVDCx20_ASAP7_75t_R g179 ( .A(n_161), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_158), .Y(n_180) );
CKINVDCx5p33_ASAP7_75t_R g181 ( .A(n_152), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_158), .Y(n_182) );
CKINVDCx5p33_ASAP7_75t_R g183 ( .A(n_152), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_158), .Y(n_184) );
CKINVDCx5p33_ASAP7_75t_R g185 ( .A(n_148), .Y(n_185) );
CKINVDCx5p33_ASAP7_75t_R g186 ( .A(n_148), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_159), .Y(n_187) );
BUFx10_ASAP7_75t_L g188 ( .A(n_154), .Y(n_188) );
CKINVDCx20_ASAP7_75t_R g189 ( .A(n_167), .Y(n_189) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_147), .Y(n_190) );
INVx3_ASAP7_75t_L g191 ( .A(n_159), .Y(n_191) );
CKINVDCx20_ASAP7_75t_R g192 ( .A(n_167), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_166), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_166), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_159), .Y(n_195) );
CKINVDCx5p33_ASAP7_75t_R g196 ( .A(n_167), .Y(n_196) );
CKINVDCx11_ASAP7_75t_R g197 ( .A(n_159), .Y(n_197) );
CKINVDCx5p33_ASAP7_75t_R g198 ( .A(n_154), .Y(n_198) );
CKINVDCx5p33_ASAP7_75t_R g199 ( .A(n_154), .Y(n_199) );
CKINVDCx20_ASAP7_75t_R g200 ( .A(n_145), .Y(n_200) );
INVx3_ASAP7_75t_L g201 ( .A(n_160), .Y(n_201) );
CKINVDCx5p33_ASAP7_75t_R g202 ( .A(n_145), .Y(n_202) );
INVx3_ASAP7_75t_L g203 ( .A(n_160), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_151), .B(n_124), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_162), .Y(n_205) );
CKINVDCx20_ASAP7_75t_R g206 ( .A(n_151), .Y(n_206) );
CKINVDCx5p33_ASAP7_75t_R g207 ( .A(n_163), .Y(n_207) );
CKINVDCx5p33_ASAP7_75t_R g208 ( .A(n_163), .Y(n_208) );
BUFx16f_ASAP7_75t_R g209 ( .A(n_162), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_166), .Y(n_210) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_165), .Y(n_211) );
AOI21x1_ASAP7_75t_L g212 ( .A1(n_165), .A2(n_131), .B(n_138), .Y(n_212) );
CKINVDCx20_ASAP7_75t_R g213 ( .A(n_164), .Y(n_213) );
CKINVDCx20_ASAP7_75t_R g214 ( .A(n_164), .Y(n_214) );
CKINVDCx5p33_ASAP7_75t_R g215 ( .A(n_143), .Y(n_215) );
CKINVDCx5p33_ASAP7_75t_R g216 ( .A(n_143), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_142), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_142), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_164), .Y(n_219) );
BUFx3_ASAP7_75t_L g220 ( .A(n_143), .Y(n_220) );
CKINVDCx8_ASAP7_75t_R g221 ( .A(n_143), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_142), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_185), .B(n_114), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_188), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_188), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_188), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_196), .B(n_202), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_207), .B(n_113), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_208), .B(n_115), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_211), .B(n_120), .Y(n_230) );
INVx8_ASAP7_75t_L g231 ( .A(n_189), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_186), .B(n_109), .Y(n_232) );
NOR2xp33_ASAP7_75t_SL g233 ( .A(n_171), .B(n_121), .Y(n_233) );
BUFx4_ASAP7_75t_L g234 ( .A(n_209), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_204), .B(n_122), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_205), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_198), .B(n_126), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_199), .B(n_129), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_187), .B(n_132), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_172), .B(n_134), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_201), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_195), .B(n_135), .Y(n_242) );
INVxp67_ASAP7_75t_L g243 ( .A(n_175), .Y(n_243) );
NAND2x1p5_ASAP7_75t_L g244 ( .A(n_191), .B(n_140), .Y(n_244) );
INVx4_ASAP7_75t_L g245 ( .A(n_197), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_197), .B(n_139), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_174), .B(n_180), .Y(n_247) );
INVx8_ASAP7_75t_L g248 ( .A(n_192), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_201), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g250 ( .A(n_191), .B(n_141), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_182), .B(n_127), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_203), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_184), .B(n_137), .Y(n_253) );
INVxp33_ASAP7_75t_L g254 ( .A(n_178), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_203), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_212), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_219), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_217), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_217), .Y(n_259) );
CKINVDCx5p33_ASAP7_75t_R g260 ( .A(n_169), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g261 ( .A(n_179), .B(n_137), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_206), .B(n_137), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_206), .B(n_156), .Y(n_263) );
INVx2_ASAP7_75t_SL g264 ( .A(n_177), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_213), .Y(n_265) );
INVxp67_ASAP7_75t_L g266 ( .A(n_170), .Y(n_266) );
INVx2_ASAP7_75t_SL g267 ( .A(n_200), .Y(n_267) );
INVx3_ASAP7_75t_L g268 ( .A(n_221), .Y(n_268) );
AO221x1_ASAP7_75t_L g269 ( .A1(n_181), .A2(n_183), .B1(n_173), .B2(n_214), .C(n_147), .Y(n_269) );
AO221x1_ASAP7_75t_L g270 ( .A1(n_176), .A2(n_147), .B1(n_157), .B2(n_7), .C(n_8), .Y(n_270) );
NAND3xp33_ASAP7_75t_L g271 ( .A(n_215), .B(n_157), .C(n_147), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_220), .B(n_156), .Y(n_272) );
NAND2xp5_ASAP7_75t_SL g273 ( .A(n_216), .B(n_147), .Y(n_273) );
AND2x2_ASAP7_75t_L g274 ( .A(n_176), .B(n_5), .Y(n_274) );
OAI21xp33_ASAP7_75t_L g275 ( .A1(n_193), .A2(n_168), .B(n_156), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_193), .B(n_168), .Y(n_276) );
INVx3_ASAP7_75t_L g277 ( .A(n_194), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_218), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_194), .B(n_168), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_278), .Y(n_280) );
NOR2xp67_ASAP7_75t_L g281 ( .A(n_245), .B(n_18), .Y(n_281) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_244), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_236), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_244), .B(n_6), .Y(n_284) );
BUFx8_ASAP7_75t_L g285 ( .A(n_264), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_258), .Y(n_286) );
XNOR2xp5_ASAP7_75t_L g287 ( .A(n_267), .B(n_6), .Y(n_287) );
BUFx3_ASAP7_75t_L g288 ( .A(n_245), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_247), .Y(n_289) );
NAND2x1p5_ASAP7_75t_L g290 ( .A(n_224), .B(n_210), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_259), .Y(n_291) );
NOR2xp33_ASAP7_75t_L g292 ( .A(n_243), .B(n_7), .Y(n_292) );
BUFx3_ASAP7_75t_L g293 ( .A(n_268), .Y(n_293) );
NAND2x1p5_ASAP7_75t_L g294 ( .A(n_225), .B(n_210), .Y(n_294) );
NOR2xp33_ASAP7_75t_L g295 ( .A(n_254), .B(n_8), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_277), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_276), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_276), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_279), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_241), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_228), .B(n_9), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_249), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_279), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_233), .B(n_9), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_256), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_228), .B(n_10), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_252), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_255), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_272), .Y(n_309) );
NAND2xp5_ASAP7_75t_SL g310 ( .A(n_226), .B(n_218), .Y(n_310) );
CKINVDCx5p33_ASAP7_75t_R g311 ( .A(n_260), .Y(n_311) );
BUFx2_ASAP7_75t_L g312 ( .A(n_231), .Y(n_312) );
BUFx3_ASAP7_75t_L g313 ( .A(n_268), .Y(n_313) );
INVx4_ASAP7_75t_L g314 ( .A(n_274), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_257), .Y(n_315) );
NOR2x2_ASAP7_75t_L g316 ( .A(n_231), .B(n_10), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_272), .Y(n_317) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_239), .A2(n_222), .B(n_190), .Y(n_318) );
INVx5_ASAP7_75t_L g319 ( .A(n_270), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_251), .Y(n_320) );
OAI21xp5_ASAP7_75t_L g321 ( .A1(n_239), .A2(n_222), .B(n_157), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_242), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_271), .Y(n_323) );
OAI22xp5_ASAP7_75t_L g324 ( .A1(n_242), .A2(n_147), .B1(n_157), .B2(n_13), .Y(n_324) );
OAI22xp5_ASAP7_75t_L g325 ( .A1(n_289), .A2(n_263), .B1(n_227), .B2(n_232), .Y(n_325) );
OAI21xp5_ASAP7_75t_L g326 ( .A1(n_322), .A2(n_235), .B(n_253), .Y(n_326) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_282), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_283), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_289), .B(n_240), .Y(n_329) );
INVx3_ASAP7_75t_L g330 ( .A(n_282), .Y(n_330) );
AOI22xp33_ASAP7_75t_SL g331 ( .A1(n_304), .A2(n_248), .B1(n_269), .B2(n_261), .Y(n_331) );
OAI22xp5_ASAP7_75t_L g332 ( .A1(n_314), .A2(n_230), .B1(n_229), .B2(n_262), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_322), .B(n_223), .Y(n_333) );
OR2x6_ASAP7_75t_L g334 ( .A(n_312), .B(n_248), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_320), .B(n_265), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_297), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_320), .B(n_237), .Y(n_337) );
OR2x6_ASAP7_75t_SL g338 ( .A(n_311), .B(n_248), .Y(n_338) );
O2A1O1Ixp33_ASAP7_75t_L g339 ( .A1(n_301), .A2(n_250), .B(n_266), .C(n_238), .Y(n_339) );
NAND2x1p5_ASAP7_75t_L g340 ( .A(n_282), .B(n_246), .Y(n_340) );
NOR3xp33_ASAP7_75t_SL g341 ( .A(n_311), .B(n_234), .C(n_273), .Y(n_341) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_282), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_297), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_283), .Y(n_344) );
INVxp67_ASAP7_75t_L g345 ( .A(n_282), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_298), .Y(n_346) );
A2O1A1Ixp33_ASAP7_75t_L g347 ( .A1(n_306), .A2(n_275), .B(n_157), .C(n_190), .Y(n_347) );
CKINVDCx20_ASAP7_75t_R g348 ( .A(n_285), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_298), .B(n_11), .Y(n_349) );
AOI21xp5_ASAP7_75t_L g350 ( .A1(n_305), .A2(n_190), .B(n_157), .Y(n_350) );
AOI21xp5_ASAP7_75t_L g351 ( .A1(n_347), .A2(n_318), .B(n_321), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_335), .B(n_292), .Y(n_352) );
AOI22x1_ASAP7_75t_L g353 ( .A1(n_336), .A2(n_323), .B1(n_280), .B2(n_305), .Y(n_353) );
OR2x2_ASAP7_75t_L g354 ( .A(n_343), .B(n_299), .Y(n_354) );
INVx8_ASAP7_75t_L g355 ( .A(n_348), .Y(n_355) );
AOI21xp5_ASAP7_75t_L g356 ( .A1(n_332), .A2(n_280), .B(n_323), .Y(n_356) );
BUFx2_ASAP7_75t_SL g357 ( .A(n_327), .Y(n_357) );
OR2x2_ASAP7_75t_L g358 ( .A(n_346), .B(n_299), .Y(n_358) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_334), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_328), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_344), .B(n_303), .Y(n_361) );
CKINVDCx11_ASAP7_75t_R g362 ( .A(n_338), .Y(n_362) );
AO21x2_ASAP7_75t_L g363 ( .A1(n_349), .A2(n_324), .B(n_284), .Y(n_363) );
INVx1_ASAP7_75t_SL g364 ( .A(n_334), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_327), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_337), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_342), .Y(n_367) );
NAND2x1p5_ASAP7_75t_L g368 ( .A(n_327), .B(n_303), .Y(n_368) );
OAI21xp5_ASAP7_75t_L g369 ( .A1(n_329), .A2(n_317), .B(n_315), .Y(n_369) );
NAND2x1p5_ASAP7_75t_L g370 ( .A(n_327), .B(n_309), .Y(n_370) );
AOI21x1_ASAP7_75t_L g371 ( .A1(n_350), .A2(n_315), .B(n_281), .Y(n_371) );
AND2x4_ASAP7_75t_L g372 ( .A(n_330), .B(n_300), .Y(n_372) );
OAI21xp5_ASAP7_75t_L g373 ( .A1(n_333), .A2(n_317), .B(n_302), .Y(n_373) );
BUFx12f_ASAP7_75t_L g374 ( .A(n_334), .Y(n_374) );
OAI21x1_ASAP7_75t_L g375 ( .A1(n_330), .A2(n_290), .B(n_294), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_337), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_342), .B(n_309), .Y(n_377) );
INVx5_ASAP7_75t_L g378 ( .A(n_345), .Y(n_378) );
OAI21x1_ASAP7_75t_L g379 ( .A1(n_340), .A2(n_294), .B(n_290), .Y(n_379) );
OAI21x1_ASAP7_75t_L g380 ( .A1(n_326), .A2(n_294), .B(n_290), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_345), .Y(n_381) );
BUFx12f_ASAP7_75t_L g382 ( .A(n_362), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_360), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_367), .Y(n_384) );
BUFx3_ASAP7_75t_L g385 ( .A(n_379), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_353), .Y(n_386) );
AOI22xp33_ASAP7_75t_SL g387 ( .A1(n_374), .A2(n_319), .B1(n_285), .B2(n_288), .Y(n_387) );
CKINVDCx5p33_ASAP7_75t_R g388 ( .A(n_362), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_353), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_361), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_361), .Y(n_391) );
OAI22xp5_ASAP7_75t_L g392 ( .A1(n_369), .A2(n_331), .B1(n_319), .B2(n_287), .Y(n_392) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_379), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_354), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_354), .Y(n_395) );
BUFx12f_ASAP7_75t_L g396 ( .A(n_355), .Y(n_396) );
CKINVDCx6p67_ASAP7_75t_R g397 ( .A(n_355), .Y(n_397) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_373), .A2(n_331), .B1(n_319), .B2(n_325), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_358), .Y(n_399) );
INVx3_ASAP7_75t_L g400 ( .A(n_375), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_377), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_377), .Y(n_402) );
BUFx2_ASAP7_75t_L g403 ( .A(n_368), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_381), .Y(n_404) );
CKINVDCx20_ASAP7_75t_R g405 ( .A(n_355), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_381), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_368), .Y(n_407) );
OAI21x1_ASAP7_75t_L g408 ( .A1(n_371), .A2(n_281), .B(n_307), .Y(n_408) );
OAI21x1_ASAP7_75t_L g409 ( .A1(n_351), .A2(n_307), .B(n_286), .Y(n_409) );
OAI21xp5_ASAP7_75t_L g410 ( .A1(n_352), .A2(n_339), .B(n_295), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_368), .Y(n_411) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_359), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_370), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_365), .Y(n_414) );
BUFx2_ASAP7_75t_R g415 ( .A(n_357), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_370), .Y(n_416) );
INVx3_ASAP7_75t_L g417 ( .A(n_375), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_370), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_366), .B(n_300), .Y(n_419) );
INVx3_ASAP7_75t_L g420 ( .A(n_380), .Y(n_420) );
OAI21x1_ASAP7_75t_L g421 ( .A1(n_380), .A2(n_286), .B(n_291), .Y(n_421) );
INVx3_ASAP7_75t_L g422 ( .A(n_378), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_372), .Y(n_423) );
HB1xp67_ASAP7_75t_L g424 ( .A(n_355), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_376), .B(n_302), .Y(n_425) );
OAI21x1_ASAP7_75t_SL g426 ( .A1(n_356), .A2(n_291), .B(n_296), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_372), .B(n_308), .Y(n_427) );
BUFx2_ASAP7_75t_L g428 ( .A(n_378), .Y(n_428) );
BUFx12f_ASAP7_75t_L g429 ( .A(n_382), .Y(n_429) );
CKINVDCx5p33_ASAP7_75t_R g430 ( .A(n_382), .Y(n_430) );
NOR2xp33_ASAP7_75t_R g431 ( .A(n_397), .B(n_364), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_392), .A2(n_363), .B1(n_378), .B2(n_313), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_383), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g434 ( .A1(n_398), .A2(n_363), .B1(n_341), .B2(n_378), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_401), .B(n_378), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g436 ( .A1(n_419), .A2(n_363), .B1(n_341), .B2(n_293), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_427), .B(n_12), .Y(n_437) );
NAND2xp33_ASAP7_75t_R g438 ( .A(n_388), .B(n_316), .Y(n_438) );
NAND2xp33_ASAP7_75t_R g439 ( .A(n_428), .B(n_13), .Y(n_439) );
OR2x6_ASAP7_75t_L g440 ( .A(n_428), .B(n_357), .Y(n_440) );
CKINVDCx5p33_ASAP7_75t_R g441 ( .A(n_396), .Y(n_441) );
NAND2xp33_ASAP7_75t_R g442 ( .A(n_422), .B(n_14), .Y(n_442) );
OR2x2_ASAP7_75t_SL g443 ( .A(n_424), .B(n_15), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_384), .Y(n_444) );
CKINVDCx5p33_ASAP7_75t_R g445 ( .A(n_396), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_427), .B(n_16), .Y(n_446) );
NAND2xp33_ASAP7_75t_R g447 ( .A(n_422), .B(n_17), .Y(n_447) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_394), .Y(n_448) );
CKINVDCx5p33_ASAP7_75t_R g449 ( .A(n_405), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_401), .B(n_296), .Y(n_450) );
BUFx2_ASAP7_75t_SL g451 ( .A(n_422), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_402), .B(n_21), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_404), .Y(n_453) );
CKINVDCx16_ASAP7_75t_R g454 ( .A(n_412), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_404), .Y(n_455) );
BUFx12f_ASAP7_75t_L g456 ( .A(n_419), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_406), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_390), .B(n_310), .Y(n_458) );
INVx3_ASAP7_75t_L g459 ( .A(n_385), .Y(n_459) );
NAND2xp33_ASAP7_75t_R g460 ( .A(n_403), .B(n_22), .Y(n_460) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_406), .Y(n_461) );
CKINVDCx16_ASAP7_75t_R g462 ( .A(n_385), .Y(n_462) );
INVx3_ASAP7_75t_L g463 ( .A(n_385), .Y(n_463) );
NAND3xp33_ASAP7_75t_SL g464 ( .A(n_387), .B(n_23), .C(n_24), .Y(n_464) );
CKINVDCx5p33_ASAP7_75t_R g465 ( .A(n_415), .Y(n_465) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_395), .Y(n_466) );
AO31x2_ASAP7_75t_L g467 ( .A1(n_386), .A2(n_26), .A3(n_28), .B(n_29), .Y(n_467) );
NOR3xp33_ASAP7_75t_SL g468 ( .A(n_410), .B(n_30), .C(n_31), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_391), .Y(n_469) );
AND2x4_ASAP7_75t_L g470 ( .A(n_423), .B(n_32), .Y(n_470) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_399), .Y(n_471) );
NOR3xp33_ASAP7_75t_SL g472 ( .A(n_425), .B(n_35), .C(n_36), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_399), .B(n_37), .Y(n_473) );
BUFx6f_ASAP7_75t_L g474 ( .A(n_393), .Y(n_474) );
BUFx4f_ASAP7_75t_SL g475 ( .A(n_403), .Y(n_475) );
INVx3_ASAP7_75t_L g476 ( .A(n_400), .Y(n_476) );
OAI21x1_ASAP7_75t_L g477 ( .A1(n_408), .A2(n_190), .B(n_40), .Y(n_477) );
CKINVDCx5p33_ASAP7_75t_R g478 ( .A(n_407), .Y(n_478) );
INVx8_ASAP7_75t_L g479 ( .A(n_400), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_407), .A2(n_45), .B1(n_46), .B2(n_47), .Y(n_480) );
AO32x2_ASAP7_75t_L g481 ( .A1(n_400), .A2(n_48), .A3(n_52), .B1(n_53), .B2(n_54), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g482 ( .A1(n_411), .A2(n_55), .B1(n_56), .B2(n_58), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_411), .Y(n_483) );
NOR2xp33_ASAP7_75t_R g484 ( .A(n_413), .B(n_418), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_414), .B(n_102), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g486 ( .A1(n_413), .A2(n_60), .B1(n_61), .B2(n_62), .Y(n_486) );
OAI21xp5_ASAP7_75t_SL g487 ( .A1(n_417), .A2(n_63), .B(n_64), .Y(n_487) );
CKINVDCx5p33_ASAP7_75t_R g488 ( .A(n_393), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_416), .B(n_67), .Y(n_489) );
CKINVDCx16_ASAP7_75t_R g490 ( .A(n_393), .Y(n_490) );
OAI22xp5_ASAP7_75t_L g491 ( .A1(n_417), .A2(n_69), .B1(n_71), .B2(n_73), .Y(n_491) );
BUFx6f_ASAP7_75t_L g492 ( .A(n_393), .Y(n_492) );
OAI22xp5_ASAP7_75t_L g493 ( .A1(n_417), .A2(n_75), .B1(n_76), .B2(n_78), .Y(n_493) );
OAI22xp5_ASAP7_75t_SL g494 ( .A1(n_417), .A2(n_79), .B1(n_80), .B2(n_81), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_409), .Y(n_495) );
NOR2xp33_ASAP7_75t_R g496 ( .A(n_393), .B(n_82), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_416), .B(n_83), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_466), .B(n_416), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_433), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_484), .B(n_483), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_453), .Y(n_501) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_461), .Y(n_502) );
INVxp33_ASAP7_75t_L g503 ( .A(n_496), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_454), .B(n_420), .Y(n_504) );
AOI32xp33_ASAP7_75t_L g505 ( .A1(n_437), .A2(n_420), .A3(n_408), .B1(n_389), .B2(n_386), .Y(n_505) );
AOI22xp33_ASAP7_75t_SL g506 ( .A1(n_475), .A2(n_426), .B1(n_389), .B2(n_421), .Y(n_506) );
INVx3_ASAP7_75t_L g507 ( .A(n_440), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_444), .Y(n_508) );
NAND2x1p5_ASAP7_75t_L g509 ( .A(n_470), .B(n_421), .Y(n_509) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_448), .Y(n_510) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_443), .B(n_409), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_446), .B(n_84), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_469), .B(n_85), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_455), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_457), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_451), .B(n_87), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_435), .B(n_88), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_440), .B(n_90), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_450), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_436), .B(n_432), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_450), .Y(n_521) );
OAI22xp33_ASAP7_75t_L g522 ( .A1(n_439), .A2(n_91), .B1(n_92), .B2(n_95), .Y(n_522) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_490), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_436), .Y(n_524) );
AO21x2_ASAP7_75t_L g525 ( .A1(n_434), .A2(n_96), .B(n_99), .Y(n_525) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_459), .Y(n_526) );
HB1xp67_ASAP7_75t_L g527 ( .A(n_459), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_458), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_462), .B(n_100), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_489), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_473), .B(n_101), .Y(n_531) );
HB1xp67_ASAP7_75t_L g532 ( .A(n_463), .Y(n_532) );
BUFx6f_ASAP7_75t_L g533 ( .A(n_474), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_489), .Y(n_534) );
INVx1_ASAP7_75t_SL g535 ( .A(n_431), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_452), .Y(n_536) );
BUFx3_ASAP7_75t_L g537 ( .A(n_441), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_479), .Y(n_538) );
AND2x4_ASAP7_75t_L g539 ( .A(n_488), .B(n_476), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_497), .Y(n_540) );
AND2x4_ASAP7_75t_L g541 ( .A(n_476), .B(n_492), .Y(n_541) );
INVx5_ASAP7_75t_L g542 ( .A(n_474), .Y(n_542) );
NOR2x1_ASAP7_75t_L g543 ( .A(n_487), .B(n_464), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_465), .B(n_449), .Y(n_544) );
OAI332xp33_ASAP7_75t_L g545 ( .A1(n_438), .A2(n_494), .A3(n_493), .B1(n_491), .B2(n_442), .B3(n_447), .C1(n_429), .C2(n_460), .Y(n_545) );
OR2x6_ASAP7_75t_L g546 ( .A(n_487), .B(n_494), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_472), .B(n_445), .Y(n_547) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_492), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_485), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_481), .Y(n_550) );
INVxp67_ASAP7_75t_L g551 ( .A(n_491), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_481), .Y(n_552) );
AND2x4_ASAP7_75t_L g553 ( .A(n_468), .B(n_467), .Y(n_553) );
OR2x6_ASAP7_75t_L g554 ( .A(n_493), .B(n_477), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_481), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_467), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_467), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_430), .Y(n_558) );
AO31x2_ASAP7_75t_L g559 ( .A1(n_486), .A2(n_386), .A3(n_389), .B(n_495), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_480), .B(n_482), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_456), .B(n_478), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_456), .A2(n_392), .B1(n_410), .B2(n_382), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_454), .B(n_461), .Y(n_563) );
BUFx2_ASAP7_75t_L g564 ( .A(n_484), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_456), .A2(n_392), .B1(n_410), .B2(n_382), .Y(n_565) );
BUFx6f_ASAP7_75t_L g566 ( .A(n_440), .Y(n_566) );
BUFx2_ASAP7_75t_L g567 ( .A(n_484), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_456), .B(n_478), .Y(n_568) );
INVx4_ASAP7_75t_L g569 ( .A(n_440), .Y(n_569) );
OAI21x1_ASAP7_75t_L g570 ( .A1(n_477), .A2(n_408), .B(n_426), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_456), .B(n_478), .Y(n_571) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_461), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_456), .B(n_478), .Y(n_573) );
NOR2x1_ASAP7_75t_L g574 ( .A(n_487), .B(n_483), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_456), .B(n_478), .Y(n_575) );
INVx6_ASAP7_75t_L g576 ( .A(n_456), .Y(n_576) );
CKINVDCx5p33_ASAP7_75t_R g577 ( .A(n_429), .Y(n_577) );
NOR2xp67_ASAP7_75t_L g578 ( .A(n_487), .B(n_382), .Y(n_578) );
INVx2_ASAP7_75t_SL g579 ( .A(n_431), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_466), .B(n_471), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_454), .B(n_461), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_466), .B(n_471), .Y(n_582) );
AND2x4_ASAP7_75t_L g583 ( .A(n_539), .B(n_504), .Y(n_583) );
NOR2x1_ASAP7_75t_SL g584 ( .A(n_546), .B(n_500), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_523), .B(n_563), .Y(n_585) );
NOR2x1_ASAP7_75t_L g586 ( .A(n_578), .B(n_535), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_523), .B(n_581), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_580), .Y(n_588) );
OR2x2_ASAP7_75t_L g589 ( .A(n_580), .B(n_582), .Y(n_589) );
OR2x2_ASAP7_75t_L g590 ( .A(n_582), .B(n_510), .Y(n_590) );
HB1xp67_ASAP7_75t_L g591 ( .A(n_572), .Y(n_591) );
AND2x4_ASAP7_75t_SL g592 ( .A(n_569), .B(n_546), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_499), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_564), .B(n_567), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_501), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_528), .B(n_519), .Y(n_596) );
INVx3_ASAP7_75t_L g597 ( .A(n_569), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_521), .B(n_508), .Y(n_598) );
OR2x2_ASAP7_75t_L g599 ( .A(n_498), .B(n_514), .Y(n_599) );
NAND2x1_ASAP7_75t_L g600 ( .A(n_574), .B(n_576), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_515), .B(n_524), .Y(n_601) );
BUFx2_ASAP7_75t_L g602 ( .A(n_535), .Y(n_602) );
BUFx2_ASAP7_75t_L g603 ( .A(n_579), .Y(n_603) );
AOI221xp5_ASAP7_75t_L g604 ( .A1(n_545), .A2(n_565), .B1(n_562), .B2(n_522), .C(n_551), .Y(n_604) );
AND2x4_ASAP7_75t_L g605 ( .A(n_507), .B(n_566), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_520), .B(n_530), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_526), .B(n_532), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_527), .B(n_532), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_534), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_538), .B(n_507), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_520), .B(n_550), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_540), .B(n_561), .Y(n_612) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_548), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_568), .B(n_571), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_573), .B(n_575), .Y(n_615) );
AND2x4_ASAP7_75t_SL g616 ( .A(n_546), .B(n_566), .Y(n_616) );
AND2x4_ASAP7_75t_L g617 ( .A(n_566), .B(n_541), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_536), .B(n_529), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_552), .B(n_555), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_551), .B(n_511), .Y(n_620) );
OR2x2_ASAP7_75t_L g621 ( .A(n_549), .B(n_517), .Y(n_621) );
INVxp67_ASAP7_75t_L g622 ( .A(n_511), .Y(n_622) );
AND2x4_ASAP7_75t_L g623 ( .A(n_541), .B(n_542), .Y(n_623) );
OR2x2_ASAP7_75t_L g624 ( .A(n_509), .B(n_503), .Y(n_624) );
AND2x4_ASAP7_75t_L g625 ( .A(n_542), .B(n_533), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_576), .B(n_565), .Y(n_626) );
INVx3_ASAP7_75t_L g627 ( .A(n_576), .Y(n_627) );
OAI22xp5_ASAP7_75t_L g628 ( .A1(n_562), .A2(n_543), .B1(n_503), .B2(n_554), .Y(n_628) );
OR2x2_ASAP7_75t_L g629 ( .A(n_509), .B(n_558), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_518), .B(n_512), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_513), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_505), .B(n_557), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_556), .B(n_506), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_547), .B(n_554), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_533), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_554), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_542), .B(n_533), .Y(n_637) );
OR2x2_ASAP7_75t_L g638 ( .A(n_537), .B(n_544), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_542), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_506), .B(n_516), .Y(n_640) );
INVxp67_ASAP7_75t_L g641 ( .A(n_525), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_545), .B(n_553), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_525), .Y(n_643) );
OR2x2_ASAP7_75t_L g644 ( .A(n_559), .B(n_560), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g645 ( .A(n_522), .B(n_553), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_570), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_531), .B(n_577), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_559), .B(n_504), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_559), .B(n_504), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_559), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_580), .Y(n_651) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_502), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_510), .B(n_528), .Y(n_653) );
AND2x4_ASAP7_75t_SL g654 ( .A(n_500), .B(n_483), .Y(n_654) );
AND2x4_ASAP7_75t_L g655 ( .A(n_539), .B(n_504), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_653), .Y(n_656) );
INVx1_ASAP7_75t_SL g657 ( .A(n_654), .Y(n_657) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_591), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_653), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_611), .B(n_606), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_604), .A2(n_642), .B1(n_645), .B2(n_592), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_611), .B(n_606), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_588), .B(n_651), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_591), .Y(n_664) );
AND2x2_ASAP7_75t_L g665 ( .A(n_648), .B(n_649), .Y(n_665) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_652), .Y(n_666) );
AND2x2_ASAP7_75t_L g667 ( .A(n_622), .B(n_636), .Y(n_667) );
AND2x2_ASAP7_75t_L g668 ( .A(n_622), .B(n_620), .Y(n_668) );
INVx2_ASAP7_75t_L g669 ( .A(n_595), .Y(n_669) );
AND2x2_ASAP7_75t_L g670 ( .A(n_620), .B(n_634), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_652), .Y(n_671) );
BUFx3_ASAP7_75t_L g672 ( .A(n_627), .Y(n_672) );
INVx2_ASAP7_75t_SL g673 ( .A(n_607), .Y(n_673) );
INVxp67_ASAP7_75t_SL g674 ( .A(n_613), .Y(n_674) );
OR2x2_ASAP7_75t_L g675 ( .A(n_589), .B(n_590), .Y(n_675) );
OR2x2_ASAP7_75t_SL g676 ( .A(n_642), .B(n_584), .Y(n_676) );
NAND2xp5_ASAP7_75t_SL g677 ( .A(n_586), .B(n_628), .Y(n_677) );
NAND4xp25_ASAP7_75t_L g678 ( .A(n_604), .B(n_628), .C(n_645), .D(n_626), .Y(n_678) );
HB1xp67_ASAP7_75t_L g679 ( .A(n_613), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_599), .Y(n_680) );
AND2x2_ASAP7_75t_L g681 ( .A(n_608), .B(n_587), .Y(n_681) );
INVx3_ASAP7_75t_L g682 ( .A(n_592), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_585), .B(n_583), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_583), .B(n_655), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_619), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_619), .Y(n_686) );
AND2x2_ASAP7_75t_L g687 ( .A(n_655), .B(n_609), .Y(n_687) );
AND2x2_ASAP7_75t_L g688 ( .A(n_644), .B(n_593), .Y(n_688) );
HB1xp67_ASAP7_75t_L g689 ( .A(n_602), .Y(n_689) );
OR2x2_ASAP7_75t_L g690 ( .A(n_596), .B(n_601), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_598), .Y(n_691) );
AND2x2_ASAP7_75t_L g692 ( .A(n_633), .B(n_632), .Y(n_692) );
NAND4xp25_ASAP7_75t_L g693 ( .A(n_632), .B(n_640), .C(n_594), .D(n_633), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_598), .Y(n_694) );
AND2x2_ASAP7_75t_L g695 ( .A(n_650), .B(n_610), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_596), .Y(n_696) );
NAND2x1_ASAP7_75t_L g697 ( .A(n_597), .B(n_627), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_612), .B(n_601), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_691), .Y(n_699) );
NAND5xp2_ASAP7_75t_L g700 ( .A(n_661), .B(n_647), .C(n_603), .D(n_641), .E(n_643), .Y(n_700) );
INVx2_ASAP7_75t_L g701 ( .A(n_679), .Y(n_701) );
OAI31xp33_ASAP7_75t_L g702 ( .A1(n_677), .A2(n_654), .A3(n_616), .B(n_630), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_691), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_694), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_694), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_670), .B(n_616), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_696), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_692), .B(n_641), .Y(n_708) );
AOI32xp33_ASAP7_75t_L g709 ( .A1(n_692), .A2(n_597), .A3(n_647), .B1(n_614), .B2(n_615), .Y(n_709) );
INVx2_ASAP7_75t_L g710 ( .A(n_669), .Y(n_710) );
NAND2xp5_ASAP7_75t_SL g711 ( .A(n_682), .B(n_639), .Y(n_711) );
AOI32xp33_ASAP7_75t_L g712 ( .A1(n_682), .A2(n_618), .A3(n_638), .B1(n_623), .B2(n_639), .Y(n_712) );
NAND4xp75_ASAP7_75t_L g713 ( .A(n_668), .B(n_637), .C(n_600), .D(n_631), .Y(n_713) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_676), .A2(n_624), .B1(n_621), .B2(n_629), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g715 ( .A1(n_678), .A2(n_605), .B1(n_617), .B2(n_623), .Y(n_715) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_657), .B(n_617), .Y(n_716) );
INVxp33_ASAP7_75t_L g717 ( .A(n_689), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_685), .B(n_646), .Y(n_718) );
OR2x2_ASAP7_75t_L g719 ( .A(n_675), .B(n_605), .Y(n_719) );
OAI22xp33_ASAP7_75t_L g720 ( .A1(n_682), .A2(n_625), .B1(n_635), .B2(n_693), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_688), .Y(n_721) );
NAND2xp5_ASAP7_75t_SL g722 ( .A(n_672), .B(n_625), .Y(n_722) );
AND2x4_ASAP7_75t_L g723 ( .A(n_667), .B(n_635), .Y(n_723) );
INVx2_ASAP7_75t_L g724 ( .A(n_658), .Y(n_724) );
NAND2x2_ASAP7_75t_L g725 ( .A(n_676), .B(n_697), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_688), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_685), .B(n_686), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_656), .Y(n_728) );
AND2x2_ASAP7_75t_L g729 ( .A(n_670), .B(n_683), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_656), .Y(n_730) );
INVx2_ASAP7_75t_SL g731 ( .A(n_684), .Y(n_731) );
OAI22xp33_ASAP7_75t_R g732 ( .A1(n_716), .A2(n_675), .B1(n_674), .B2(n_673), .Y(n_732) );
INVx1_ASAP7_75t_L g733 ( .A(n_727), .Y(n_733) );
INVxp67_ASAP7_75t_SL g734 ( .A(n_718), .Y(n_734) );
INVx1_ASAP7_75t_SL g735 ( .A(n_717), .Y(n_735) );
OAI211xp5_ASAP7_75t_L g736 ( .A1(n_702), .A2(n_709), .B(n_715), .C(n_712), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_727), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_699), .Y(n_738) );
XNOR2x1_ASAP7_75t_L g739 ( .A(n_714), .B(n_684), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g740 ( .A1(n_700), .A2(n_668), .B1(n_667), .B2(n_665), .Y(n_740) );
INVx2_ASAP7_75t_L g741 ( .A(n_710), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_703), .Y(n_742) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_718), .Y(n_743) );
NAND3xp33_ASAP7_75t_L g744 ( .A(n_702), .B(n_664), .C(n_671), .Y(n_744) );
INVx1_ASAP7_75t_SL g745 ( .A(n_711), .Y(n_745) );
AOI211xp5_ASAP7_75t_L g746 ( .A1(n_720), .A2(n_672), .B(n_662), .C(n_660), .Y(n_746) );
AOI22xp5_ASAP7_75t_L g747 ( .A1(n_714), .A2(n_665), .B1(n_687), .B2(n_680), .Y(n_747) );
OAI21xp33_ASAP7_75t_L g748 ( .A1(n_700), .A2(n_659), .B(n_695), .Y(n_748) );
OAI21xp33_ASAP7_75t_L g749 ( .A1(n_708), .A2(n_659), .B(n_695), .Y(n_749) );
XNOR2xp5_ASAP7_75t_L g750 ( .A(n_713), .B(n_683), .Y(n_750) );
AOI22xp5_ASAP7_75t_L g751 ( .A1(n_725), .A2(n_687), .B1(n_680), .B2(n_698), .Y(n_751) );
OAI31xp33_ASAP7_75t_L g752 ( .A1(n_708), .A2(n_666), .A3(n_673), .B(n_690), .Y(n_752) );
INVxp67_ASAP7_75t_L g753 ( .A(n_735), .Y(n_753) );
INVx2_ASAP7_75t_L g754 ( .A(n_741), .Y(n_754) );
OAI32xp33_ASAP7_75t_L g755 ( .A1(n_745), .A2(n_722), .A3(n_719), .B1(n_721), .B2(n_726), .Y(n_755) );
INVx2_ASAP7_75t_L g756 ( .A(n_741), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_738), .Y(n_757) );
AOI21xp5_ASAP7_75t_L g758 ( .A1(n_732), .A2(n_697), .B(n_663), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_742), .Y(n_759) );
AOI222xp33_ASAP7_75t_L g760 ( .A1(n_736), .A2(n_724), .B1(n_701), .B2(n_730), .C1(n_728), .C2(n_707), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_733), .B(n_698), .Y(n_761) );
OAI21xp33_ASAP7_75t_SL g762 ( .A1(n_752), .A2(n_731), .B(n_729), .Y(n_762) );
OAI22xp33_ASAP7_75t_SL g763 ( .A1(n_747), .A2(n_664), .B1(n_671), .B2(n_705), .Y(n_763) );
NOR2xp33_ASAP7_75t_L g764 ( .A(n_739), .B(n_690), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_753), .B(n_737), .Y(n_765) );
INVx1_ASAP7_75t_L g766 ( .A(n_761), .Y(n_766) );
AOI221xp5_ASAP7_75t_L g767 ( .A1(n_762), .A2(n_763), .B1(n_755), .B2(n_764), .C(n_744), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_757), .Y(n_768) );
OAI21xp33_ASAP7_75t_L g769 ( .A1(n_760), .A2(n_748), .B(n_740), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_759), .Y(n_770) );
INVxp33_ASAP7_75t_SL g771 ( .A(n_765), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_766), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_768), .Y(n_773) );
INVx1_ASAP7_75t_L g774 ( .A(n_770), .Y(n_774) );
NAND2xp5_ASAP7_75t_L g775 ( .A(n_771), .B(n_769), .Y(n_775) );
NOR3xp33_ASAP7_75t_L g776 ( .A(n_772), .B(n_767), .C(n_763), .Y(n_776) );
AOI311xp33_ASAP7_75t_L g777 ( .A1(n_773), .A2(n_746), .A3(n_758), .B(n_734), .C(n_704), .Y(n_777) );
AO22x1_ASAP7_75t_L g778 ( .A1(n_776), .A2(n_774), .B1(n_734), .B2(n_754), .Y(n_778) );
AOI22xp5_ASAP7_75t_SL g779 ( .A1(n_775), .A2(n_750), .B1(n_777), .B2(n_743), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_778), .Y(n_780) );
INVx2_ASAP7_75t_L g781 ( .A(n_779), .Y(n_781) );
CKINVDCx5p33_ASAP7_75t_R g782 ( .A(n_781), .Y(n_782) );
CKINVDCx20_ASAP7_75t_R g783 ( .A(n_780), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_783), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_784), .Y(n_785) );
CKINVDCx20_ASAP7_75t_R g786 ( .A(n_785), .Y(n_786) );
AOI21xp5_ASAP7_75t_L g787 ( .A1(n_786), .A2(n_782), .B(n_743), .Y(n_787) );
AOI21xp33_ASAP7_75t_L g788 ( .A1(n_787), .A2(n_756), .B(n_751), .Y(n_788) );
AOI22xp33_ASAP7_75t_SL g789 ( .A1(n_788), .A2(n_706), .B1(n_681), .B2(n_723), .Y(n_789) );
OR2x6_ASAP7_75t_L g790 ( .A(n_789), .B(n_723), .Y(n_790) );
AOI22xp5_ASAP7_75t_L g791 ( .A1(n_790), .A2(n_749), .B1(n_740), .B2(n_681), .Y(n_791) );
endmodule