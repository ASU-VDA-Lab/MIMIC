module real_jpeg_28450_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_68;
wire n_78;
wire n_83;
wire n_64;
wire n_11;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_9;
wire n_72;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_85;
wire n_89;
wire n_16;

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_0),
.A2(n_15),
.B1(n_16),
.B2(n_26),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_0),
.A2(n_20),
.B1(n_21),
.B2(n_26),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_0),
.B(n_36),
.Y(n_35)
);

AOI21xp33_ASAP7_75t_SL g42 ( 
.A1(n_0),
.A2(n_16),
.B(n_43),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_0),
.A2(n_26),
.B1(n_44),
.B2(n_45),
.Y(n_57)
);

AOI21xp33_ASAP7_75t_L g71 ( 
.A1(n_0),
.A2(n_4),
.B(n_21),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_4),
.A2(n_18),
.B1(n_20),
.B2(n_21),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_5),
.A2(n_15),
.B1(n_16),
.B2(n_24),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_5),
.A2(n_20),
.B1(n_21),
.B2(n_24),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_5),
.A2(n_24),
.B1(n_44),
.B2(n_45),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_6),
.A2(n_15),
.B1(n_16),
.B2(n_37),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_7),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_67),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_65),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_38),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_11),
.B(n_38),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_27),
.C(n_34),
.Y(n_11)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_12),
.A2(n_34),
.B1(n_35),
.B2(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_12),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g12 ( 
.A1(n_13),
.A2(n_19),
.B1(n_23),
.B2(n_25),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_13),
.B(n_25),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_19),
.Y(n_13)
);

OAI22xp33_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_16),
.Y(n_15)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_16),
.A2(n_18),
.B(n_26),
.C(n_71),
.Y(n_70)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_19),
.B(n_26),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_20),
.B(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_21),
.B(n_30),
.Y(n_29)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_26),
.A2(n_41),
.B(n_42),
.C(n_44),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_26),
.B(n_89),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_27),
.A2(n_73),
.B1(n_75),
.B2(n_76),
.Y(n_72)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_27),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_27),
.B(n_92),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_28),
.A2(n_33),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_29),
.B(n_30),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_59),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_37),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_51),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_46),
.B1(n_47),
.B2(n_50),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_40),
.Y(n_50)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_48),
.B(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_60),
.B2(n_61),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B(n_56),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_58),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_60),
.A2(n_61),
.B1(n_70),
.B2(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_61),
.B(n_70),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_63),
.B(n_64),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_77),
.B(n_95),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_72),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_70),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_73),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_85),
.B(n_94),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_83),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_79),
.B(n_83),
.Y(n_94)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_80),
.B(n_87),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_91),
.B(n_93),
.Y(n_85)
);

INVx5_ASAP7_75t_SL g89 ( 
.A(n_90),
.Y(n_89)
);


endmodule