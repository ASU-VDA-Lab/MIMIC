module fake_jpeg_24257_n_284 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_284);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_284;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_155;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_36),
.B(n_40),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

CKINVDCx9p33_ASAP7_75t_R g49 ( 
.A(n_37),
.Y(n_49)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

AOI21xp33_ASAP7_75t_L g42 ( 
.A1(n_37),
.A2(n_20),
.B(n_1),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_42),
.A2(n_46),
.B(n_20),
.C(n_31),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_36),
.B(n_18),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_55),
.Y(n_79)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_34),
.A2(n_27),
.B1(n_33),
.B2(n_29),
.Y(n_46)
);

CKINVDCx12_ASAP7_75t_R g48 ( 
.A(n_37),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_48),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_33),
.B1(n_27),
.B2(n_17),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_50),
.A2(n_24),
.B1(n_22),
.B2(n_18),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_27),
.B1(n_33),
.B2(n_22),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_52),
.A2(n_23),
.B(n_19),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_22),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_54),
.B(n_24),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_20),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_58),
.B(n_60),
.Y(n_91)
);

CKINVDCx5p33_ASAP7_75t_R g60 ( 
.A(n_48),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_61),
.A2(n_64),
.B1(n_72),
.B2(n_80),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_53),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_62),
.B(n_65),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_63),
.A2(n_0),
.B(n_2),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_42),
.A2(n_41),
.B1(n_40),
.B2(n_35),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_53),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_46),
.A2(n_29),
.B1(n_18),
.B2(n_30),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_66),
.A2(n_77),
.B1(n_81),
.B2(n_52),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_L g67 ( 
.A1(n_55),
.A2(n_56),
.B1(n_35),
.B2(n_46),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_67),
.A2(n_51),
.B1(n_31),
.B2(n_28),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_68),
.Y(n_94)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_69),
.A2(n_75),
.B1(n_0),
.B2(n_2),
.Y(n_109)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_70),
.B(n_74),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_47),
.Y(n_71)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_50),
.A2(n_17),
.B1(n_19),
.B2(n_23),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_45),
.A2(n_30),
.B1(n_29),
.B2(n_24),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_45),
.A2(n_30),
.B1(n_21),
.B2(n_17),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_57),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_76),
.B(n_78),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_43),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_50),
.A2(n_23),
.B1(n_19),
.B2(n_16),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_51),
.A2(n_21),
.B1(n_32),
.B2(n_25),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_82),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_20),
.C(n_32),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_64),
.C(n_77),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_47),
.B(n_26),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_84),
.Y(n_97)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_3),
.Y(n_114)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_89),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_90),
.B(n_80),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_108),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_55),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_93),
.B(n_102),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_63),
.A2(n_51),
.B1(n_45),
.B2(n_56),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_101),
.A2(n_105),
.B1(n_115),
.B2(n_89),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_20),
.Y(n_102)
);

NAND3xp33_ASAP7_75t_SL g103 ( 
.A(n_78),
.B(n_25),
.C(n_49),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_117),
.Y(n_124)
);

A2O1A1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_62),
.A2(n_16),
.B(n_28),
.C(n_31),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_104),
.A2(n_107),
.B(n_59),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_58),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_106),
.Y(n_128)
);

OA21x2_ASAP7_75t_L g107 ( 
.A1(n_67),
.A2(n_31),
.B(n_28),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_65),
.B(n_26),
.C(n_1),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_111),
.A2(n_85),
.B(n_12),
.Y(n_138)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_114),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_69),
.A2(n_9),
.B1(n_14),
.B2(n_5),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_61),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_106),
.B(n_83),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_118),
.B(n_122),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_119),
.A2(n_136),
.B1(n_6),
.B2(n_7),
.Y(n_169)
);

OA22x2_ASAP7_75t_L g121 ( 
.A1(n_107),
.A2(n_76),
.B1(n_72),
.B2(n_87),
.Y(n_121)
);

OA22x2_ASAP7_75t_L g164 ( 
.A1(n_121),
.A2(n_98),
.B1(n_95),
.B2(n_4),
.Y(n_164)
);

A2O1A1Ixp33_ASAP7_75t_L g122 ( 
.A1(n_100),
.A2(n_60),
.B(n_85),
.C(n_68),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_3),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_139),
.Y(n_155)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_96),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_130),
.Y(n_150)
);

NAND2x1p5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_68),
.Y(n_127)
);

AO22x1_ASAP7_75t_SL g152 ( 
.A1(n_127),
.A2(n_104),
.B1(n_107),
.B2(n_91),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_100),
.A2(n_59),
.B1(n_86),
.B2(n_87),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_129),
.A2(n_131),
.B1(n_141),
.B2(n_105),
.Y(n_147)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_74),
.Y(n_132)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_116),
.Y(n_134)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_134),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_135),
.B(n_94),
.Y(n_154)
);

FAx1_ASAP7_75t_SL g146 ( 
.A(n_138),
.B(n_108),
.CI(n_114),
.CON(n_146),
.SN(n_146)
);

INVx2_ASAP7_75t_R g139 ( 
.A(n_91),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_70),
.Y(n_140)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_140),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_117),
.A2(n_88),
.B1(n_82),
.B2(n_3),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_3),
.Y(n_142)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_142),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_99),
.A2(n_4),
.B(n_5),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_12),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_93),
.B(n_102),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_144),
.B(n_145),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_82),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_146),
.B(n_147),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_134),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_149),
.B(n_173),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_127),
.A2(n_107),
.B1(n_90),
.B2(n_101),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_151),
.Y(n_197)
);

A2O1A1Ixp33_ASAP7_75t_SL g186 ( 
.A1(n_152),
.A2(n_175),
.B(n_138),
.C(n_143),
.Y(n_186)
);

AND2x6_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_97),
.Y(n_153)
);

NAND3xp33_ASAP7_75t_L g189 ( 
.A(n_153),
.B(n_171),
.C(n_126),
.Y(n_189)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_154),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_144),
.B(n_97),
.C(n_113),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_157),
.B(n_165),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_130),
.B(n_113),
.Y(n_159)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_159),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_104),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_167),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_119),
.A2(n_98),
.B1(n_95),
.B2(n_4),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_161),
.A2(n_133),
.B1(n_122),
.B2(n_136),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_162),
.B(n_172),
.Y(n_198)
);

OA21x2_ASAP7_75t_L g177 ( 
.A1(n_164),
.A2(n_135),
.B(n_139),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_6),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_6),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_168),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_169),
.A2(n_118),
.B1(n_124),
.B2(n_139),
.Y(n_185)
);

AND2x6_ASAP7_75t_L g171 ( 
.A(n_120),
.B(n_7),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_127),
.B(n_8),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_132),
.Y(n_173)
);

INVxp33_ASAP7_75t_L g174 ( 
.A(n_135),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_174),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_129),
.B(n_8),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_150),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_176),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_177),
.B(n_181),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_149),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_178),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_174),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_180),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_147),
.A2(n_124),
.B1(n_131),
.B2(n_121),
.Y(n_184)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_184),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_185),
.B(n_195),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_186),
.A2(n_189),
.B1(n_200),
.B2(n_158),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_152),
.A2(n_121),
.B1(n_141),
.B2(n_128),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_196),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_165),
.B(n_120),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_193),
.B(n_199),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_161),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_153),
.A2(n_121),
.B1(n_137),
.B2(n_128),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_157),
.B(n_123),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_152),
.A2(n_121),
.B1(n_123),
.B2(n_125),
.Y(n_200)
);

INVxp33_ASAP7_75t_SL g202 ( 
.A(n_191),
.Y(n_202)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_202),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_177),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_204),
.B(n_214),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_206),
.A2(n_209),
.B1(n_200),
.B2(n_188),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_148),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_207),
.B(n_212),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_197),
.A2(n_172),
.B1(n_156),
.B2(n_163),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_187),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_210),
.A2(n_218),
.B1(n_125),
.B2(n_164),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_183),
.B(n_148),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_185),
.B(n_142),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_190),
.B(n_166),
.Y(n_216)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_216),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_177),
.A2(n_170),
.B(n_164),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_217),
.A2(n_179),
.B(n_192),
.Y(n_224)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_194),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_207),
.B(n_212),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_222),
.B(n_229),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_224),
.A2(n_232),
.B1(n_235),
.B2(n_204),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_182),
.C(n_199),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_228),
.C(n_219),
.Y(n_237)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_208),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_227),
.B(n_230),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_182),
.C(n_196),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_206),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_205),
.Y(n_230)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_231),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_215),
.A2(n_197),
.B1(n_184),
.B2(n_181),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_192),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_233),
.B(n_229),
.Y(n_242)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_209),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_172),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_215),
.A2(n_171),
.B1(n_186),
.B2(n_164),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_236),
.A2(n_186),
.B1(n_146),
.B2(n_198),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_249),
.C(n_228),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_233),
.B(n_203),
.Y(n_238)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_238),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_241),
.B(n_247),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_242),
.B(n_243),
.Y(n_256)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_226),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_244),
.A2(n_245),
.B(n_246),
.Y(n_253)
);

A2O1A1Ixp33_ASAP7_75t_SL g245 ( 
.A1(n_236),
.A2(n_211),
.B(n_213),
.C(n_232),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_218),
.Y(n_246)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_231),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_250),
.B(n_252),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_225),
.C(n_223),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_245),
.Y(n_254)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_254),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_223),
.C(n_220),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_257),
.B(n_258),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_162),
.C(n_222),
.Y(n_258)
);

AOI21x1_ASAP7_75t_L g259 ( 
.A1(n_245),
.A2(n_186),
.B(n_155),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_259),
.A2(n_239),
.B(n_247),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_261),
.A2(n_265),
.B(n_267),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_253),
.Y(n_264)
);

OA21x2_ASAP7_75t_L g269 ( 
.A1(n_264),
.A2(n_198),
.B(n_155),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_259),
.A2(n_240),
.B(n_245),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_251),
.B(n_242),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_266),
.B(n_155),
.C(n_146),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_255),
.A2(n_210),
.B(n_198),
.Y(n_267)
);

OR2x2_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_256),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_268),
.B(n_273),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_269),
.B(n_272),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_271),
.A2(n_10),
.B(n_12),
.Y(n_276)
);

NOR3xp33_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_175),
.C(n_11),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_266),
.B(n_175),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_270),
.B(n_263),
.Y(n_275)
);

INVxp33_ASAP7_75t_L g279 ( 
.A(n_275),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_276),
.A2(n_10),
.B1(n_13),
.B2(n_14),
.Y(n_278)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_278),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_279),
.A2(n_274),
.B(n_277),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_280),
.A2(n_15),
.B(n_10),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_282),
.B(n_281),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_13),
.Y(n_284)
);


endmodule