module fake_netlist_6_2323_n_1744 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1744);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1744;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_719;
wire n_228;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_110),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_21),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_39),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_153),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_96),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_119),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_59),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_67),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_95),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_76),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_117),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_98),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_145),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_28),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_23),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_149),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_27),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_80),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_122),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_61),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_48),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_154),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_130),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_53),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_34),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_144),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_123),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_129),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_45),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_114),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_150),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_5),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_60),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_88),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_127),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_103),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_147),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_31),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_65),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_63),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_126),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_120),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_121),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_93),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_91),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_27),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_7),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_29),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_72),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_38),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_125),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_11),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_143),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_68),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_75),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_69),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_112),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_4),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_87),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_1),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_18),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_151),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_32),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_44),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_36),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_22),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_13),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_43),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_58),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_128),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_140),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_2),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_50),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_47),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_16),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_77),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_0),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_5),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_10),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_13),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_42),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_21),
.Y(n_237)
);

BUFx5_ASAP7_75t_L g238 ( 
.A(n_31),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_139),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_101),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_90),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_8),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_25),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_102),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_23),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_24),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_71),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_104),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_85),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_100),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_64),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_42),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_17),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_89),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_39),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_70),
.Y(n_256)
);

BUFx10_ASAP7_75t_L g257 ( 
.A(n_131),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_74),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_48),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_92),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_51),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_137),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_148),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_105),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_84),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_45),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_29),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_78),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_58),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_142),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_6),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_6),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g273 ( 
.A(n_11),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_136),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_44),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_83),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_22),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_135),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_46),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_9),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_30),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_81),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_12),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_116),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_46),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_26),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_20),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_52),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_0),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_107),
.Y(n_290)
);

INVx4_ASAP7_75t_R g291 ( 
.A(n_124),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_17),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_152),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_111),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_25),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_55),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_30),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_38),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_133),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_50),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_106),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_20),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_8),
.Y(n_303)
);

BUFx10_ASAP7_75t_L g304 ( 
.A(n_62),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_34),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_16),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_24),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_18),
.Y(n_308)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_73),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_141),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_159),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_238),
.B(n_1),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_243),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_156),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_243),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_192),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_273),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_160),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_238),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_161),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_238),
.Y(n_321)
);

BUFx6f_ASAP7_75t_SL g322 ( 
.A(n_257),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_163),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_238),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_194),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_238),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_165),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_310),
.Y(n_328)
);

INVxp33_ASAP7_75t_SL g329 ( 
.A(n_172),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_273),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_204),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_238),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_238),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_200),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_238),
.B(n_2),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_226),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_238),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_205),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_241),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_166),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_157),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_244),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_248),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_254),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_222),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_167),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_262),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_282),
.Y(n_348)
);

INVxp67_ASAP7_75t_SL g349 ( 
.A(n_157),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_232),
.B(n_3),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_205),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_205),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_173),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_182),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_183),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_205),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_205),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_170),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_193),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_185),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_257),
.Y(n_361)
);

INVxp33_ASAP7_75t_L g362 ( 
.A(n_158),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_193),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_197),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_206),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_222),
.B(n_3),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_158),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_237),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_276),
.B(n_4),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_162),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_237),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_208),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_242),
.Y(n_373)
);

INVxp67_ASAP7_75t_SL g374 ( 
.A(n_162),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_210),
.Y(n_375)
);

NOR2xp67_ASAP7_75t_L g376 ( 
.A(n_309),
.B(n_7),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_211),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_242),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_212),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_267),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_267),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_319),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_319),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_338),
.Y(n_384)
);

INVx4_ASAP7_75t_L g385 ( 
.A(n_331),
.Y(n_385)
);

AND2x4_ASAP7_75t_L g386 ( 
.A(n_376),
.B(n_309),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_338),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_321),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_321),
.B(n_309),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_324),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_350),
.B(n_276),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_324),
.B(n_171),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_326),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_326),
.B(n_171),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_350),
.B(n_164),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_369),
.B(n_175),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_332),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_351),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_332),
.B(n_174),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_329),
.B(n_164),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_351),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_333),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_333),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_352),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_331),
.B(n_168),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_358),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_330),
.Y(n_407)
);

INVx6_ASAP7_75t_L g408 ( 
.A(n_331),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_352),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_337),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_341),
.B(n_168),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_356),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_356),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_337),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_357),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_341),
.B(n_177),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_357),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_312),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_312),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_335),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_359),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_335),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_359),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_363),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_363),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_368),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_368),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_371),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_376),
.B(n_174),
.Y(n_429)
);

NOR2x1_ASAP7_75t_L g430 ( 
.A(n_371),
.B(n_177),
.Y(n_430)
);

BUFx2_ASAP7_75t_L g431 ( 
.A(n_315),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_373),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_373),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_378),
.B(n_178),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_378),
.Y(n_435)
);

AND3x2_ASAP7_75t_L g436 ( 
.A(n_315),
.B(n_303),
.C(n_287),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_380),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_349),
.B(n_178),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_380),
.Y(n_439)
);

NAND2xp33_ASAP7_75t_L g440 ( 
.A(n_366),
.B(n_189),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_381),
.Y(n_441)
);

INVx4_ASAP7_75t_L g442 ( 
.A(n_381),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_349),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_374),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_374),
.Y(n_445)
);

BUFx8_ASAP7_75t_L g446 ( 
.A(n_322),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_420),
.B(n_311),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_420),
.B(n_318),
.Y(n_448)
);

INVx4_ASAP7_75t_L g449 ( 
.A(n_418),
.Y(n_449)
);

BUFx4f_ASAP7_75t_L g450 ( 
.A(n_418),
.Y(n_450)
);

AND3x2_ASAP7_75t_L g451 ( 
.A(n_407),
.B(n_345),
.C(n_317),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_390),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_420),
.B(n_320),
.Y(n_453)
);

BUFx10_ASAP7_75t_L g454 ( 
.A(n_396),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_383),
.Y(n_455)
);

AND2x4_ASAP7_75t_L g456 ( 
.A(n_405),
.B(n_181),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_383),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_390),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_390),
.Y(n_459)
);

BUFx8_ASAP7_75t_SL g460 ( 
.A(n_431),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_383),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_407),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_390),
.Y(n_463)
);

OR2x6_ASAP7_75t_L g464 ( 
.A(n_422),
.B(n_366),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_383),
.Y(n_465)
);

BUFx4f_ASAP7_75t_L g466 ( 
.A(n_418),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_390),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_396),
.B(n_323),
.Y(n_468)
);

AND2x4_ASAP7_75t_L g469 ( 
.A(n_405),
.B(n_181),
.Y(n_469)
);

INVxp33_ASAP7_75t_L g470 ( 
.A(n_431),
.Y(n_470)
);

BUFx3_ASAP7_75t_L g471 ( 
.A(n_408),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_383),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_400),
.B(n_361),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_422),
.B(n_419),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_410),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_410),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_410),
.Y(n_477)
);

NAND3xp33_ASAP7_75t_L g478 ( 
.A(n_400),
.B(n_340),
.C(n_327),
.Y(n_478)
);

INVxp67_ASAP7_75t_SL g479 ( 
.A(n_418),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_410),
.Y(n_480)
);

OR2x6_ASAP7_75t_L g481 ( 
.A(n_422),
.B(n_367),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_406),
.B(n_361),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_390),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_443),
.B(n_346),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_443),
.B(n_353),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_406),
.B(n_328),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_419),
.B(n_354),
.Y(n_487)
);

AND2x4_ASAP7_75t_L g488 ( 
.A(n_405),
.B(n_186),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_388),
.Y(n_489)
);

INVx5_ASAP7_75t_L g490 ( 
.A(n_382),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_443),
.B(n_328),
.Y(n_491)
);

OR2x6_ASAP7_75t_L g492 ( 
.A(n_391),
.B(n_419),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_388),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_388),
.Y(n_494)
);

INVx1_ASAP7_75t_SL g495 ( 
.A(n_431),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_388),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_410),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_408),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_397),
.Y(n_499)
);

AOI22xp33_ASAP7_75t_L g500 ( 
.A1(n_419),
.A2(n_330),
.B1(n_313),
.B2(n_281),
.Y(n_500)
);

NAND2xp33_ASAP7_75t_L g501 ( 
.A(n_418),
.B(n_189),
.Y(n_501)
);

INVx2_ASAP7_75t_SL g502 ( 
.A(n_419),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_397),
.Y(n_503)
);

AND2x6_ASAP7_75t_L g504 ( 
.A(n_418),
.B(n_186),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_414),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_397),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_382),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_414),
.Y(n_508)
);

INVx4_ASAP7_75t_L g509 ( 
.A(n_418),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_382),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_397),
.Y(n_511)
);

BUFx3_ASAP7_75t_L g512 ( 
.A(n_408),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_385),
.B(n_355),
.Y(n_513)
);

AOI21x1_ASAP7_75t_L g514 ( 
.A1(n_389),
.A2(n_191),
.B(n_190),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_384),
.Y(n_515)
);

INVx1_ASAP7_75t_SL g516 ( 
.A(n_391),
.Y(n_516)
);

AOI22xp33_ASAP7_75t_L g517 ( 
.A1(n_418),
.A2(n_281),
.B1(n_246),
.B2(n_233),
.Y(n_517)
);

AND2x6_ASAP7_75t_L g518 ( 
.A(n_418),
.B(n_190),
.Y(n_518)
);

AND2x6_ASAP7_75t_L g519 ( 
.A(n_418),
.B(n_191),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_414),
.Y(n_520)
);

AOI22xp33_ASAP7_75t_L g521 ( 
.A1(n_391),
.A2(n_246),
.B1(n_233),
.B2(n_232),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_414),
.Y(n_522)
);

AOI22xp33_ASAP7_75t_SL g523 ( 
.A1(n_391),
.A2(n_322),
.B1(n_188),
.B2(n_229),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_384),
.Y(n_524)
);

NAND2xp33_ASAP7_75t_L g525 ( 
.A(n_411),
.B(n_189),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_382),
.Y(n_526)
);

AOI22xp33_ASAP7_75t_L g527 ( 
.A1(n_395),
.A2(n_416),
.B1(n_438),
.B2(n_411),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_414),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_408),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_382),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_444),
.B(n_360),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_384),
.Y(n_532)
);

OR2x2_ASAP7_75t_L g533 ( 
.A(n_444),
.B(n_345),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_387),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_387),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_387),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_398),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_398),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_444),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_398),
.Y(n_540)
);

OR2x6_ASAP7_75t_L g541 ( 
.A(n_445),
.B(n_411),
.Y(n_541)
);

NAND2xp33_ASAP7_75t_SL g542 ( 
.A(n_411),
.B(n_221),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_401),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_382),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_385),
.B(n_364),
.Y(n_545)
);

INVx8_ASAP7_75t_L g546 ( 
.A(n_395),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_401),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_401),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_404),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_445),
.B(n_372),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_404),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_404),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_409),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_409),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_409),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_395),
.A2(n_236),
.B1(n_227),
.B2(n_253),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_412),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_445),
.A2(n_379),
.B1(n_377),
.B2(n_365),
.Y(n_558)
);

OAI22xp33_ASAP7_75t_L g559 ( 
.A1(n_416),
.A2(n_234),
.B1(n_235),
.B2(n_184),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_416),
.A2(n_375),
.B1(n_322),
.B2(n_347),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_416),
.B(n_322),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_412),
.Y(n_562)
);

NAND2xp33_ASAP7_75t_L g563 ( 
.A(n_438),
.B(n_189),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_412),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_413),
.Y(n_565)
);

NAND2xp33_ASAP7_75t_L g566 ( 
.A(n_438),
.B(n_189),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_L g567 ( 
.A1(n_395),
.A2(n_438),
.B1(n_429),
.B2(n_440),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_382),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_L g569 ( 
.A1(n_429),
.A2(n_169),
.B1(n_180),
.B2(n_187),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_446),
.B(n_257),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_385),
.B(n_217),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_413),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_413),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_415),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_385),
.B(n_362),
.Y(n_575)
);

AND3x2_ASAP7_75t_L g576 ( 
.A(n_429),
.B(n_370),
.C(n_367),
.Y(n_576)
);

INVxp67_ASAP7_75t_L g577 ( 
.A(n_405),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_382),
.Y(n_578)
);

BUFx6f_ASAP7_75t_L g579 ( 
.A(n_382),
.Y(n_579)
);

INVx4_ASAP7_75t_L g580 ( 
.A(n_382),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_446),
.B(n_385),
.Y(n_581)
);

OR2x2_ASAP7_75t_L g582 ( 
.A(n_429),
.B(n_370),
.Y(n_582)
);

INVx5_ASAP7_75t_L g583 ( 
.A(n_393),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_415),
.Y(n_584)
);

INVx1_ASAP7_75t_SL g585 ( 
.A(n_436),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_385),
.B(n_348),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_415),
.Y(n_587)
);

CKINVDCx20_ASAP7_75t_R g588 ( 
.A(n_446),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_385),
.B(n_314),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_417),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_SL g591 ( 
.A(n_446),
.B(n_316),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_417),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_429),
.B(n_225),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_549),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_534),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_549),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_450),
.B(n_466),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_546),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_555),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_555),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_534),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_447),
.B(n_436),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_536),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_450),
.B(n_429),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_516),
.B(n_325),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_L g606 ( 
.A1(n_502),
.A2(n_429),
.B1(n_386),
.B2(n_440),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_527),
.B(n_446),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_450),
.B(n_386),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_466),
.B(n_386),
.Y(n_609)
);

BUFx3_ASAP7_75t_L g610 ( 
.A(n_546),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_462),
.B(n_334),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_502),
.B(n_386),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_479),
.B(n_386),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_448),
.B(n_245),
.Y(n_614)
);

HB1xp67_ASAP7_75t_L g615 ( 
.A(n_495),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_567),
.B(n_386),
.Y(n_616)
);

INVxp67_ASAP7_75t_L g617 ( 
.A(n_468),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_575),
.B(n_386),
.Y(n_618)
);

NAND2x1p5_ASAP7_75t_L g619 ( 
.A(n_449),
.B(n_430),
.Y(n_619)
);

OAI22xp33_ASAP7_75t_L g620 ( 
.A1(n_492),
.A2(n_260),
.B1(n_293),
.B2(n_299),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_466),
.B(n_446),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_484),
.B(n_408),
.Y(n_622)
);

OR2x2_ASAP7_75t_SL g623 ( 
.A(n_478),
.B(n_169),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_577),
.B(n_430),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_453),
.B(n_280),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_470),
.B(n_336),
.Y(n_626)
);

OR2x6_ASAP7_75t_L g627 ( 
.A(n_492),
.B(n_180),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_485),
.B(n_408),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_449),
.B(n_446),
.Y(n_629)
);

NAND2xp33_ASAP7_75t_L g630 ( 
.A(n_546),
.B(n_231),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_487),
.B(n_292),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_536),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_531),
.B(n_442),
.Y(n_633)
);

INVx8_ASAP7_75t_L g634 ( 
.A(n_546),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_550),
.B(n_442),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_449),
.B(n_393),
.Y(n_636)
);

NAND3xp33_ASAP7_75t_L g637 ( 
.A(n_539),
.B(n_491),
.C(n_542),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_537),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_470),
.B(n_339),
.Y(n_639)
);

NOR2x1p5_ASAP7_75t_L g640 ( 
.A(n_533),
.B(n_176),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_474),
.B(n_408),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_561),
.B(n_408),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_557),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_537),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_571),
.A2(n_389),
.B(n_392),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_509),
.B(n_492),
.Y(n_646)
);

OR2x2_ASAP7_75t_L g647 ( 
.A(n_533),
.B(n_434),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_509),
.B(n_393),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_492),
.B(n_393),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_541),
.B(n_393),
.Y(n_650)
);

INVxp67_ASAP7_75t_L g651 ( 
.A(n_482),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_541),
.B(n_393),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_539),
.B(n_442),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_454),
.B(n_393),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_454),
.B(n_393),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_557),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_454),
.B(n_442),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_562),
.Y(n_658)
);

OAI22xp5_ASAP7_75t_L g659 ( 
.A1(n_541),
.A2(n_342),
.B1(n_343),
.B2(n_344),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_473),
.B(n_442),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_541),
.B(n_393),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_576),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_481),
.B(n_442),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_538),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_562),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_481),
.B(n_430),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_464),
.B(n_393),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_538),
.Y(n_668)
);

OAI22xp5_ASAP7_75t_SL g669 ( 
.A1(n_523),
.A2(n_272),
.B1(n_277),
.B2(n_255),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_SL g670 ( 
.A(n_588),
.B(n_304),
.Y(n_670)
);

AOI22xp5_ASAP7_75t_L g671 ( 
.A1(n_464),
.A2(n_239),
.B1(n_240),
.B2(n_247),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_481),
.B(n_442),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_481),
.B(n_464),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_565),
.Y(n_674)
);

OR2x2_ASAP7_75t_L g675 ( 
.A(n_464),
.B(n_434),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_565),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_582),
.B(n_179),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_573),
.Y(n_678)
);

HB1xp67_ASAP7_75t_L g679 ( 
.A(n_582),
.Y(n_679)
);

NAND2xp33_ASAP7_75t_SL g680 ( 
.A(n_588),
.B(n_201),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_551),
.Y(n_681)
);

INVxp67_ASAP7_75t_L g682 ( 
.A(n_486),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_463),
.B(n_467),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_463),
.B(n_402),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_500),
.B(n_434),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_551),
.Y(n_686)
);

AND2x2_ASAP7_75t_SL g687 ( 
.A(n_525),
.B(n_563),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_467),
.B(n_402),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_586),
.A2(n_265),
.B1(n_263),
.B2(n_278),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_456),
.A2(n_389),
.B1(n_392),
.B2(n_394),
.Y(n_690)
);

BUFx6f_ASAP7_75t_L g691 ( 
.A(n_507),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_456),
.B(n_402),
.Y(n_692)
);

O2A1O1Ixp5_ASAP7_75t_L g693 ( 
.A1(n_456),
.A2(n_399),
.B(n_392),
.C(n_394),
.Y(n_693)
);

A2O1A1Ixp33_ASAP7_75t_L g694 ( 
.A1(n_469),
.A2(n_394),
.B(n_399),
.C(n_195),
.Y(n_694)
);

OAI22xp5_ASAP7_75t_L g695 ( 
.A1(n_581),
.A2(n_264),
.B1(n_199),
.B2(n_198),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_573),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_469),
.B(n_402),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_560),
.B(n_249),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_574),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_469),
.B(n_402),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_488),
.B(n_402),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_488),
.B(n_402),
.Y(n_702)
);

AOI22xp33_ASAP7_75t_L g703 ( 
.A1(n_488),
.A2(n_399),
.B1(n_198),
.B2(n_260),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_525),
.B(n_402),
.Y(n_704)
);

AOI221xp5_ASAP7_75t_L g705 ( 
.A1(n_559),
.A2(n_227),
.B1(n_215),
.B2(n_213),
.C(n_187),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_574),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_513),
.B(n_402),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_592),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_592),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_545),
.B(n_402),
.Y(n_710)
);

INVxp67_ASAP7_75t_L g711 ( 
.A(n_460),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_552),
.Y(n_712)
);

OR2x2_ASAP7_75t_L g713 ( 
.A(n_542),
.B(n_202),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_552),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_558),
.B(n_432),
.Y(n_715)
);

INVx3_ASAP7_75t_L g716 ( 
.A(n_553),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_553),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_563),
.B(n_566),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_566),
.B(n_403),
.Y(n_719)
);

INVx2_ASAP7_75t_SL g720 ( 
.A(n_451),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_564),
.Y(n_721)
);

OAI22xp5_ASAP7_75t_L g722 ( 
.A1(n_589),
.A2(n_264),
.B1(n_196),
.B2(n_299),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_507),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_515),
.B(n_403),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_564),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_593),
.B(n_452),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_572),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_524),
.B(n_403),
.Y(n_728)
);

INVx2_ASAP7_75t_SL g729 ( 
.A(n_585),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_572),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_532),
.B(n_403),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_458),
.B(n_403),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_535),
.B(n_403),
.Y(n_733)
);

NOR3xp33_ASAP7_75t_L g734 ( 
.A(n_570),
.B(n_223),
.C(n_218),
.Y(n_734)
);

BUFx6f_ASAP7_75t_L g735 ( 
.A(n_507),
.Y(n_735)
);

AND2x6_ASAP7_75t_SL g736 ( 
.A(n_460),
.B(n_213),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_459),
.B(n_403),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_540),
.B(n_403),
.Y(n_738)
);

AND2x6_ASAP7_75t_SL g739 ( 
.A(n_591),
.B(n_215),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_483),
.B(n_403),
.Y(n_740)
);

AO22x2_ASAP7_75t_L g741 ( 
.A1(n_543),
.A2(n_270),
.B1(n_293),
.B2(n_256),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_584),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_521),
.B(n_432),
.Y(n_743)
);

OAI22xp33_ASAP7_75t_L g744 ( 
.A1(n_547),
.A2(n_214),
.B1(n_209),
.B2(n_199),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_584),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_548),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_554),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_587),
.B(n_203),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_556),
.B(n_432),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_590),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_504),
.A2(n_519),
.B1(n_518),
.B2(n_501),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_510),
.B(n_441),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_503),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_503),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_510),
.B(n_441),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_510),
.B(n_441),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_506),
.Y(n_757)
);

OR2x2_ASAP7_75t_L g758 ( 
.A(n_517),
.B(n_207),
.Y(n_758)
);

O2A1O1Ixp33_ASAP7_75t_L g759 ( 
.A1(n_501),
.A2(n_285),
.B(n_236),
.C(n_253),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_530),
.B(n_544),
.Y(n_760)
);

OR2x6_ASAP7_75t_L g761 ( 
.A(n_514),
.B(n_269),
.Y(n_761)
);

NOR2xp67_ASAP7_75t_L g762 ( 
.A(n_514),
.B(n_439),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_530),
.B(n_441),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_633),
.B(n_504),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_633),
.B(n_504),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_659),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_604),
.A2(n_613),
.B(n_597),
.Y(n_767)
);

OAI22xp5_ASAP7_75t_L g768 ( 
.A1(n_616),
.A2(n_617),
.B1(n_635),
.B2(n_606),
.Y(n_768)
);

O2A1O1Ixp33_ASAP7_75t_L g769 ( 
.A1(n_722),
.A2(n_511),
.B(n_506),
.C(n_569),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_624),
.B(n_507),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_635),
.B(n_504),
.Y(n_771)
);

INVx3_ASAP7_75t_L g772 ( 
.A(n_716),
.Y(n_772)
);

OAI22xp5_ASAP7_75t_L g773 ( 
.A1(n_687),
.A2(n_471),
.B1(n_498),
.B2(n_512),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_594),
.Y(n_774)
);

OAI21xp5_ASAP7_75t_L g775 ( 
.A1(n_693),
.A2(n_511),
.B(n_504),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_624),
.B(n_598),
.Y(n_776)
);

BUFx6f_ASAP7_75t_L g777 ( 
.A(n_598),
.Y(n_777)
);

OAI321xp33_ASAP7_75t_L g778 ( 
.A1(n_705),
.A2(n_283),
.A3(n_285),
.B1(n_275),
.B2(n_271),
.C(n_269),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_596),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_631),
.B(n_504),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_631),
.B(n_518),
.Y(n_781)
);

AOI21xp33_ASAP7_75t_L g782 ( 
.A1(n_614),
.A2(n_196),
.B(n_195),
.Y(n_782)
);

AOI21xp5_ASAP7_75t_L g783 ( 
.A1(n_604),
.A2(n_498),
.B(n_471),
.Y(n_783)
);

A2O1A1Ixp33_ASAP7_75t_L g784 ( 
.A1(n_614),
.A2(n_270),
.B(n_256),
.C(n_258),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_625),
.B(n_518),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_625),
.B(n_580),
.Y(n_786)
);

INVxp67_ASAP7_75t_L g787 ( 
.A(n_615),
.Y(n_787)
);

A2O1A1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_660),
.A2(n_284),
.B(n_258),
.C(n_268),
.Y(n_788)
);

INVxp67_ASAP7_75t_L g789 ( 
.A(n_605),
.Y(n_789)
);

OAI21xp33_ASAP7_75t_L g790 ( 
.A1(n_647),
.A2(n_219),
.B(n_216),
.Y(n_790)
);

AOI21xp5_ASAP7_75t_L g791 ( 
.A1(n_612),
.A2(n_609),
.B(n_608),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_624),
.B(n_518),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_679),
.B(n_580),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_608),
.A2(n_609),
.B(n_618),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_599),
.Y(n_795)
);

OAI21xp5_ASAP7_75t_L g796 ( 
.A1(n_645),
.A2(n_518),
.B(n_519),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_598),
.B(n_507),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_685),
.B(n_439),
.Y(n_798)
);

INVxp67_ASAP7_75t_L g799 ( 
.A(n_729),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_598),
.B(n_526),
.Y(n_800)
);

AOI21xp5_ASAP7_75t_L g801 ( 
.A1(n_622),
.A2(n_529),
.B(n_580),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_600),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_628),
.A2(n_544),
.B(n_530),
.Y(n_803)
);

HB1xp67_ASAP7_75t_L g804 ( 
.A(n_627),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_641),
.A2(n_544),
.B(n_579),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_619),
.A2(n_526),
.B(n_579),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_619),
.A2(n_526),
.B(n_579),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_653),
.B(n_518),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_707),
.A2(n_579),
.B(n_578),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_595),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_666),
.B(n_646),
.Y(n_811)
);

NAND2x1p5_ASAP7_75t_L g812 ( 
.A(n_610),
.B(n_526),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_707),
.A2(n_568),
.B(n_578),
.Y(n_813)
);

INVx2_ASAP7_75t_SL g814 ( 
.A(n_626),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_710),
.A2(n_636),
.B(n_648),
.Y(n_815)
);

CKINVDCx8_ASAP7_75t_R g816 ( 
.A(n_736),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_710),
.A2(n_568),
.B(n_578),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_653),
.B(n_519),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_643),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_690),
.B(n_519),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_682),
.B(n_637),
.Y(n_821)
);

AO21x2_ASAP7_75t_L g822 ( 
.A1(n_621),
.A2(n_209),
.B(n_214),
.Y(n_822)
);

NAND2xp33_ASAP7_75t_L g823 ( 
.A(n_634),
.B(n_519),
.Y(n_823)
);

OAI21x1_ASAP7_75t_L g824 ( 
.A1(n_760),
.A2(n_636),
.B(n_697),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_726),
.A2(n_578),
.B(n_568),
.Y(n_825)
);

AOI21xp5_ASAP7_75t_L g826 ( 
.A1(n_726),
.A2(n_578),
.B(n_568),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_SL g827 ( 
.A(n_611),
.B(n_304),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_687),
.B(n_677),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_677),
.B(n_519),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_642),
.A2(n_568),
.B(n_583),
.Y(n_830)
);

INVx2_ASAP7_75t_SL g831 ( 
.A(n_639),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_656),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_675),
.B(n_489),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_651),
.B(n_493),
.Y(n_834)
);

O2A1O1Ixp33_ASAP7_75t_L g835 ( 
.A1(n_694),
.A2(n_655),
.B(n_654),
.C(n_620),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_715),
.B(n_439),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_602),
.B(n_673),
.Y(n_837)
);

INVx11_ASAP7_75t_L g838 ( 
.A(n_623),
.Y(n_838)
);

A2O1A1Ixp33_ASAP7_75t_L g839 ( 
.A1(n_673),
.A2(n_271),
.B(n_288),
.C(n_286),
.Y(n_839)
);

O2A1O1Ixp33_ASAP7_75t_L g840 ( 
.A1(n_654),
.A2(n_655),
.B(n_667),
.C(n_744),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_692),
.A2(n_583),
.B(n_490),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_658),
.Y(n_842)
);

BUFx6f_ASAP7_75t_L g843 ( 
.A(n_610),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_660),
.B(n_494),
.Y(n_844)
);

HB1xp67_ASAP7_75t_L g845 ( 
.A(n_627),
.Y(n_845)
);

OAI22xp5_ASAP7_75t_L g846 ( 
.A1(n_718),
.A2(n_268),
.B1(n_274),
.B2(n_284),
.Y(n_846)
);

A2O1A1Ixp33_ASAP7_75t_L g847 ( 
.A1(n_749),
.A2(n_286),
.B(n_289),
.C(n_288),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_692),
.A2(n_583),
.B(n_490),
.Y(n_848)
);

OAI22xp5_ASAP7_75t_L g849 ( 
.A1(n_607),
.A2(n_650),
.B1(n_661),
.B2(n_652),
.Y(n_849)
);

O2A1O1Ixp5_ASAP7_75t_L g850 ( 
.A1(n_695),
.A2(n_461),
.B(n_528),
.C(n_522),
.Y(n_850)
);

HB1xp67_ASAP7_75t_L g851 ( 
.A(n_627),
.Y(n_851)
);

NOR2xp67_ASAP7_75t_L g852 ( 
.A(n_711),
.B(n_496),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_L g853 ( 
.A1(n_702),
.A2(n_499),
.B(n_528),
.Y(n_853)
);

A2O1A1Ixp33_ASAP7_75t_L g854 ( 
.A1(n_663),
.A2(n_274),
.B(n_522),
.C(n_520),
.Y(n_854)
);

AOI21xp33_ASAP7_75t_L g855 ( 
.A1(n_713),
.A2(n_300),
.B(n_224),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_700),
.A2(n_583),
.B(n_490),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_700),
.A2(n_583),
.B(n_490),
.Y(n_857)
);

INVx2_ASAP7_75t_SL g858 ( 
.A(n_640),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_701),
.A2(n_649),
.B(n_704),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_701),
.A2(n_490),
.B(n_508),
.Y(n_860)
);

A2O1A1Ixp33_ASAP7_75t_L g861 ( 
.A1(n_663),
.A2(n_465),
.B(n_508),
.C(n_505),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_SL g862 ( 
.A(n_670),
.B(n_669),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_719),
.A2(n_520),
.B(n_505),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_672),
.A2(n_250),
.B1(n_251),
.B2(n_290),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_665),
.B(n_455),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_674),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_691),
.A2(n_497),
.B(n_480),
.Y(n_867)
);

AO21x1_ASAP7_75t_L g868 ( 
.A1(n_621),
.A2(n_275),
.B(n_283),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_676),
.B(n_678),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_691),
.A2(n_497),
.B(n_480),
.Y(n_870)
);

AOI22xp5_ASAP7_75t_L g871 ( 
.A1(n_602),
.A2(n_294),
.B1(n_301),
.B2(n_475),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_696),
.Y(n_872)
);

OAI21xp5_ASAP7_75t_L g873 ( 
.A1(n_683),
.A2(n_477),
.B(n_476),
.Y(n_873)
);

OR2x2_ASAP7_75t_L g874 ( 
.A(n_680),
.B(n_220),
.Y(n_874)
);

AO21x1_ASAP7_75t_L g875 ( 
.A1(n_629),
.A2(n_289),
.B(n_307),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_699),
.B(n_455),
.Y(n_876)
);

O2A1O1Ixp5_ASAP7_75t_L g877 ( 
.A1(n_629),
.A2(n_477),
.B(n_476),
.C(n_475),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_657),
.B(n_457),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_706),
.B(n_457),
.Y(n_879)
);

AOI22xp5_ASAP7_75t_L g880 ( 
.A1(n_672),
.A2(n_472),
.B1(n_465),
.B2(n_461),
.Y(n_880)
);

O2A1O1Ixp33_ASAP7_75t_L g881 ( 
.A1(n_708),
.A2(n_472),
.B(n_307),
.C(n_441),
.Y(n_881)
);

AOI21x1_ASAP7_75t_L g882 ( 
.A1(n_684),
.A2(n_737),
.B(n_732),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_709),
.B(n_441),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_595),
.Y(n_884)
);

NOR2xp67_ASAP7_75t_L g885 ( 
.A(n_689),
.B(n_66),
.Y(n_885)
);

OAI22xp5_ASAP7_75t_L g886 ( 
.A1(n_703),
.A2(n_228),
.B1(n_230),
.B2(n_252),
.Y(n_886)
);

OAI21xp5_ASAP7_75t_L g887 ( 
.A1(n_724),
.A2(n_437),
.B(n_435),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_747),
.B(n_421),
.Y(n_888)
);

OAI21x1_ASAP7_75t_L g889 ( 
.A1(n_752),
.A2(n_437),
.B(n_435),
.Y(n_889)
);

INVx1_ASAP7_75t_SL g890 ( 
.A(n_720),
.Y(n_890)
);

NOR3xp33_ASAP7_75t_L g891 ( 
.A(n_698),
.B(n_259),
.C(n_261),
.Y(n_891)
);

OAI21xp5_ASAP7_75t_L g892 ( 
.A1(n_728),
.A2(n_437),
.B(n_435),
.Y(n_892)
);

INVxp67_ASAP7_75t_L g893 ( 
.A(n_748),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_746),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_657),
.B(n_421),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_739),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_743),
.B(n_746),
.Y(n_897)
);

AND2x4_ASAP7_75t_L g898 ( 
.A(n_662),
.B(n_421),
.Y(n_898)
);

OAI22xp5_ASAP7_75t_L g899 ( 
.A1(n_750),
.A2(n_306),
.B1(n_279),
.B2(n_295),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_750),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_748),
.B(n_266),
.Y(n_901)
);

O2A1O1Ixp33_ASAP7_75t_L g902 ( 
.A1(n_758),
.A2(n_426),
.B(n_423),
.C(n_433),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_601),
.Y(n_903)
);

BUFx6f_ASAP7_75t_L g904 ( 
.A(n_691),
.Y(n_904)
);

OAI21xp5_ASAP7_75t_L g905 ( 
.A1(n_731),
.A2(n_437),
.B(n_435),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_716),
.B(n_423),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_671),
.B(n_296),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_SL g908 ( 
.A(n_691),
.B(n_428),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_723),
.A2(n_437),
.B(n_435),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_601),
.Y(n_910)
);

OAI21xp5_ASAP7_75t_L g911 ( 
.A1(n_733),
.A2(n_433),
.B(n_421),
.Y(n_911)
);

BUFx4f_ASAP7_75t_L g912 ( 
.A(n_761),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_603),
.B(n_433),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_723),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_723),
.A2(n_433),
.B(n_423),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_603),
.B(n_427),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_632),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_723),
.A2(n_427),
.B(n_426),
.Y(n_918)
);

OAI21xp5_ASAP7_75t_L g919 ( 
.A1(n_738),
.A2(n_423),
.B(n_427),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_632),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_638),
.Y(n_921)
);

O2A1O1Ixp33_ASAP7_75t_L g922 ( 
.A1(n_759),
.A2(n_754),
.B(n_753),
.C(n_757),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_638),
.B(n_426),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_644),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_644),
.B(n_425),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_735),
.A2(n_425),
.B(n_291),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_734),
.B(n_305),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_735),
.A2(n_425),
.B(n_428),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_735),
.A2(n_763),
.B(n_756),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_755),
.A2(n_425),
.B(n_428),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_634),
.A2(n_428),
.B(n_424),
.Y(n_931)
);

O2A1O1Ixp33_ASAP7_75t_SL g932 ( 
.A1(n_688),
.A2(n_304),
.B(n_10),
.C(n_12),
.Y(n_932)
);

O2A1O1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_717),
.A2(n_308),
.B(n_302),
.C(n_298),
.Y(n_933)
);

CKINVDCx20_ASAP7_75t_R g934 ( 
.A(n_634),
.Y(n_934)
);

NOR2x2_ASAP7_75t_L g935 ( 
.A(n_761),
.B(n_297),
.Y(n_935)
);

OAI21xp5_ASAP7_75t_L g936 ( 
.A1(n_762),
.A2(n_428),
.B(n_424),
.Y(n_936)
);

OAI22xp5_ASAP7_75t_L g937 ( 
.A1(n_751),
.A2(n_428),
.B1(n_424),
.B2(n_155),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_630),
.A2(n_684),
.B(n_732),
.Y(n_938)
);

OAI21xp5_ASAP7_75t_L g939 ( 
.A1(n_664),
.A2(n_428),
.B(n_424),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_664),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_668),
.B(n_428),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_668),
.B(n_428),
.Y(n_942)
);

NAND2x1p5_ASAP7_75t_L g943 ( 
.A(n_721),
.B(n_424),
.Y(n_943)
);

AOI21x1_ASAP7_75t_L g944 ( 
.A1(n_737),
.A2(n_424),
.B(n_146),
.Y(n_944)
);

BUFx2_ASAP7_75t_L g945 ( 
.A(n_741),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_740),
.A2(n_424),
.B(n_138),
.Y(n_946)
);

INVx3_ASAP7_75t_L g947 ( 
.A(n_681),
.Y(n_947)
);

AOI22xp5_ASAP7_75t_L g948 ( 
.A1(n_725),
.A2(n_424),
.B1(n_134),
.B2(n_132),
.Y(n_948)
);

CKINVDCx16_ASAP7_75t_R g949 ( 
.A(n_934),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_866),
.Y(n_950)
);

O2A1O1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_782),
.A2(n_730),
.B(n_745),
.C(n_742),
.Y(n_951)
);

A2O1A1Ixp33_ASAP7_75t_SL g952 ( 
.A1(n_901),
.A2(n_714),
.B(n_686),
.C(n_712),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_794),
.A2(n_714),
.B(n_681),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_866),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_791),
.A2(n_712),
.B(n_686),
.Y(n_955)
);

INVx1_ASAP7_75t_SL g956 ( 
.A(n_890),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_L g957 ( 
.A1(n_901),
.A2(n_727),
.B1(n_740),
.B2(n_741),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_843),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_836),
.B(n_741),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_893),
.B(n_761),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_837),
.B(n_424),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_767),
.A2(n_118),
.B(n_115),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_837),
.B(n_113),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_862),
.B(n_821),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_947),
.Y(n_965)
);

OR2x2_ASAP7_75t_L g966 ( 
.A(n_787),
.B(n_789),
.Y(n_966)
);

O2A1O1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_855),
.A2(n_9),
.B(n_14),
.C(n_15),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_798),
.B(n_14),
.Y(n_968)
);

NAND3xp33_ASAP7_75t_SL g969 ( 
.A(n_827),
.B(n_15),
.C(n_19),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_R g970 ( 
.A(n_766),
.B(n_896),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_786),
.B(n_19),
.Y(n_971)
);

OR2x6_ASAP7_75t_L g972 ( 
.A(n_804),
.B(n_109),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_774),
.Y(n_973)
);

INVx5_ASAP7_75t_L g974 ( 
.A(n_777),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_786),
.B(n_26),
.Y(n_975)
);

BUFx2_ASAP7_75t_SL g976 ( 
.A(n_777),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_814),
.B(n_28),
.Y(n_977)
);

INVxp67_ASAP7_75t_L g978 ( 
.A(n_821),
.Y(n_978)
);

NAND2xp33_ASAP7_75t_SL g979 ( 
.A(n_843),
.B(n_32),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_SL g980 ( 
.A(n_816),
.B(n_799),
.Y(n_980)
);

OR2x2_ASAP7_75t_SL g981 ( 
.A(n_874),
.B(n_33),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_897),
.B(n_33),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_828),
.B(n_108),
.Y(n_983)
);

BUFx2_ASAP7_75t_L g984 ( 
.A(n_804),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_L g985 ( 
.A(n_831),
.B(n_35),
.Y(n_985)
);

OAI22xp5_ASAP7_75t_L g986 ( 
.A1(n_768),
.A2(n_99),
.B1(n_97),
.B2(n_94),
.Y(n_986)
);

INVx3_ASAP7_75t_L g987 ( 
.A(n_777),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_834),
.B(n_779),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_777),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_796),
.A2(n_86),
.B(n_82),
.Y(n_990)
);

OAI22xp5_ASAP7_75t_L g991 ( 
.A1(n_849),
.A2(n_79),
.B1(n_36),
.B2(n_37),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_907),
.B(n_35),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_834),
.B(n_37),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_838),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_904),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_844),
.A2(n_40),
.B(n_41),
.Y(n_996)
);

INVx4_ASAP7_75t_L g997 ( 
.A(n_843),
.Y(n_997)
);

A2O1A1Ixp33_ASAP7_75t_L g998 ( 
.A1(n_907),
.A2(n_40),
.B(n_41),
.C(n_43),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_764),
.A2(n_47),
.B(n_49),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_765),
.A2(n_49),
.B(n_51),
.Y(n_1000)
);

NOR3xp33_ASAP7_75t_L g1001 ( 
.A(n_790),
.B(n_52),
.C(n_53),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_771),
.A2(n_54),
.B(n_55),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_947),
.Y(n_1003)
);

OR2x2_ASAP7_75t_L g1004 ( 
.A(n_845),
.B(n_54),
.Y(n_1004)
);

OAI22x1_ASAP7_75t_L g1005 ( 
.A1(n_945),
.A2(n_56),
.B1(n_57),
.B2(n_59),
.Y(n_1005)
);

OR2x6_ASAP7_75t_L g1006 ( 
.A(n_845),
.B(n_56),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_815),
.A2(n_57),
.B(n_60),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_795),
.B(n_802),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_840),
.A2(n_835),
.B(n_785),
.C(n_859),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_912),
.B(n_843),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_895),
.A2(n_829),
.B(n_938),
.Y(n_1011)
);

OAI22x1_ASAP7_75t_L g1012 ( 
.A1(n_851),
.A2(n_927),
.B1(n_858),
.B2(n_832),
.Y(n_1012)
);

XOR2xp5_ASAP7_75t_L g1013 ( 
.A(n_811),
.B(n_851),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_811),
.B(n_819),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_842),
.Y(n_1015)
);

O2A1O1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_784),
.A2(n_839),
.B(n_847),
.C(n_788),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_878),
.A2(n_801),
.B(n_783),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_878),
.A2(n_773),
.B(n_818),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_R g1019 ( 
.A(n_912),
.B(n_882),
.Y(n_1019)
);

NOR2x1_ASAP7_75t_L g1020 ( 
.A(n_885),
.B(n_776),
.Y(n_1020)
);

HB1xp67_ASAP7_75t_L g1021 ( 
.A(n_898),
.Y(n_1021)
);

AOI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_891),
.A2(n_776),
.B1(n_792),
.B2(n_871),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_SL g1023 ( 
.A(n_891),
.B(n_869),
.Y(n_1023)
);

HB1xp67_ASAP7_75t_L g1024 ( 
.A(n_898),
.Y(n_1024)
);

BUFx3_ASAP7_75t_L g1025 ( 
.A(n_872),
.Y(n_1025)
);

AND2x2_ASAP7_75t_L g1026 ( 
.A(n_852),
.B(n_899),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_833),
.B(n_793),
.Y(n_1027)
);

OAI22x1_ASAP7_75t_L g1028 ( 
.A1(n_935),
.A2(n_793),
.B1(n_894),
.B2(n_900),
.Y(n_1028)
);

OR2x2_ASAP7_75t_L g1029 ( 
.A(n_886),
.B(n_864),
.Y(n_1029)
);

OAI21x1_ASAP7_75t_L g1030 ( 
.A1(n_889),
.A2(n_805),
.B(n_807),
.Y(n_1030)
);

AOI33xp33_ASAP7_75t_L g1031 ( 
.A1(n_932),
.A2(n_933),
.A3(n_940),
.B1(n_920),
.B2(n_921),
.B3(n_778),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_780),
.B(n_781),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_810),
.Y(n_1033)
);

BUFx2_ASAP7_75t_L g1034 ( 
.A(n_839),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_847),
.B(n_884),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_806),
.A2(n_770),
.B(n_823),
.Y(n_1036)
);

A2O1A1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_820),
.A2(n_769),
.B(n_922),
.C(n_808),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_770),
.B(n_772),
.Y(n_1038)
);

BUFx8_ASAP7_75t_SL g1039 ( 
.A(n_904),
.Y(n_1039)
);

AOI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_875),
.A2(n_868),
.B1(n_772),
.B2(n_888),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_903),
.B(n_910),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_917),
.B(n_924),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_812),
.A2(n_797),
.B1(n_800),
.B2(n_904),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_904),
.B(n_914),
.Y(n_1044)
);

OAI21xp33_ASAP7_75t_L g1045 ( 
.A1(n_846),
.A2(n_879),
.B(n_876),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_865),
.B(n_929),
.Y(n_1046)
);

NAND2x1p5_ASAP7_75t_L g1047 ( 
.A(n_914),
.B(n_797),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_883),
.B(n_923),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_830),
.A2(n_853),
.B(n_809),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_914),
.B(n_812),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_SL g1051 ( 
.A(n_914),
.B(n_880),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_913),
.Y(n_1052)
);

INVx6_ASAP7_75t_L g1053 ( 
.A(n_932),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_822),
.B(n_824),
.Y(n_1054)
);

NAND3xp33_ASAP7_75t_L g1055 ( 
.A(n_854),
.B(n_948),
.C(n_937),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_926),
.Y(n_1056)
);

AND2x4_ASAP7_75t_L g1057 ( 
.A(n_861),
.B(n_908),
.Y(n_1057)
);

INVx4_ASAP7_75t_L g1058 ( 
.A(n_943),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_813),
.A2(n_817),
.B(n_803),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_936),
.A2(n_775),
.B(n_825),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_822),
.B(n_942),
.Y(n_1061)
);

HB1xp67_ASAP7_75t_L g1062 ( 
.A(n_906),
.Y(n_1062)
);

BUFx2_ASAP7_75t_L g1063 ( 
.A(n_943),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_908),
.B(n_916),
.Y(n_1064)
);

O2A1O1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_881),
.A2(n_902),
.B(n_942),
.C(n_925),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_873),
.A2(n_826),
.B(n_919),
.Y(n_1066)
);

AOI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_941),
.A2(n_860),
.B1(n_911),
.B2(n_946),
.Y(n_1067)
);

INVx3_ASAP7_75t_L g1068 ( 
.A(n_944),
.Y(n_1068)
);

BUFx12f_ASAP7_75t_L g1069 ( 
.A(n_850),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_887),
.B(n_905),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_892),
.A2(n_863),
.B(n_877),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_939),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_909),
.Y(n_1073)
);

INVx5_ASAP7_75t_L g1074 ( 
.A(n_931),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_867),
.A2(n_870),
.B(n_930),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_915),
.B(n_918),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_928),
.B(n_841),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_848),
.A2(n_856),
.B(n_857),
.Y(n_1078)
);

A2O1A1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_901),
.A2(n_614),
.B(n_625),
.C(n_828),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_893),
.B(n_617),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_947),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_947),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_794),
.A2(n_466),
.B(n_450),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_794),
.A2(n_466),
.B(n_450),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_893),
.B(n_617),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_893),
.B(n_617),
.Y(n_1086)
);

NAND3xp33_ASAP7_75t_SL g1087 ( 
.A(n_862),
.B(n_827),
.C(n_901),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_836),
.B(n_617),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_893),
.B(n_617),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_794),
.A2(n_466),
.B(n_450),
.Y(n_1090)
);

AOI22x1_ASAP7_75t_L g1091 ( 
.A1(n_767),
.A2(n_794),
.B1(n_938),
.B2(n_791),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_836),
.B(n_407),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_794),
.A2(n_466),
.B(n_450),
.Y(n_1093)
);

AND2x4_ASAP7_75t_L g1094 ( 
.A(n_1025),
.B(n_1010),
.Y(n_1094)
);

OA21x2_ASAP7_75t_L g1095 ( 
.A1(n_1009),
.A2(n_1018),
.B(n_1011),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_1030),
.A2(n_955),
.B(n_953),
.Y(n_1096)
);

AOI31xp67_ASAP7_75t_L g1097 ( 
.A1(n_1067),
.A2(n_1040),
.A3(n_961),
.B(n_1022),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_1046),
.A2(n_1011),
.B(n_1066),
.Y(n_1098)
);

AO32x2_ASAP7_75t_L g1099 ( 
.A1(n_991),
.A2(n_986),
.A3(n_1043),
.B1(n_1058),
.B2(n_1053),
.Y(n_1099)
);

O2A1O1Ixp33_ASAP7_75t_SL g1100 ( 
.A1(n_1079),
.A2(n_1087),
.B(n_964),
.C(n_992),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_973),
.Y(n_1101)
);

INVx4_ASAP7_75t_L g1102 ( 
.A(n_974),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1015),
.Y(n_1103)
);

INVx2_ASAP7_75t_SL g1104 ( 
.A(n_956),
.Y(n_1104)
);

AO32x2_ASAP7_75t_L g1105 ( 
.A1(n_1058),
.A2(n_1053),
.A3(n_1031),
.B1(n_1069),
.B2(n_1034),
.Y(n_1105)
);

AOI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_1092),
.A2(n_1086),
.B1(n_1080),
.B2(n_978),
.Y(n_1106)
);

INVx8_ASAP7_75t_L g1107 ( 
.A(n_974),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_955),
.A2(n_953),
.B(n_1036),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1027),
.B(n_988),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1088),
.B(n_1014),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1066),
.A2(n_1093),
.B(n_1090),
.Y(n_1111)
);

AOI22xp33_ASAP7_75t_SL g1112 ( 
.A1(n_1029),
.A2(n_970),
.B1(n_1006),
.B2(n_985),
.Y(n_1112)
);

OAI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1037),
.A2(n_1018),
.B(n_1032),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_1083),
.A2(n_1093),
.B(n_1084),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1052),
.B(n_1062),
.Y(n_1115)
);

BUFx6f_ASAP7_75t_L g1116 ( 
.A(n_1039),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_SL g1117 ( 
.A(n_994),
.B(n_969),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_1021),
.B(n_1024),
.Y(n_1118)
);

O2A1O1Ixp5_ASAP7_75t_SL g1119 ( 
.A1(n_1023),
.A2(n_1068),
.B(n_1076),
.C(n_983),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1070),
.B(n_1035),
.Y(n_1120)
);

CKINVDCx20_ASAP7_75t_R g1121 ( 
.A(n_949),
.Y(n_1121)
);

AND2x4_ASAP7_75t_L g1122 ( 
.A(n_984),
.B(n_950),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_1085),
.Y(n_1123)
);

INVx3_ASAP7_75t_L g1124 ( 
.A(n_958),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_1078),
.A2(n_1075),
.B(n_1059),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1083),
.A2(n_1090),
.B(n_1084),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1017),
.A2(n_1049),
.B(n_1060),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_977),
.B(n_1013),
.Y(n_1128)
);

O2A1O1Ixp33_ASAP7_75t_SL g1129 ( 
.A1(n_963),
.A2(n_971),
.B(n_975),
.C(n_998),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1008),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1041),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_959),
.B(n_1038),
.Y(n_1132)
);

O2A1O1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_1089),
.A2(n_993),
.B(n_1001),
.C(n_967),
.Y(n_1133)
);

BUFx3_ASAP7_75t_L g1134 ( 
.A(n_958),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_1033),
.Y(n_1135)
);

O2A1O1Ixp33_ASAP7_75t_SL g1136 ( 
.A1(n_1051),
.A2(n_952),
.B(n_1050),
.C(n_990),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1017),
.A2(n_1074),
.B(n_1071),
.Y(n_1137)
);

AOI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_1026),
.A2(n_1028),
.B1(n_980),
.B2(n_1012),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1074),
.A2(n_1071),
.B(n_1045),
.Y(n_1139)
);

HB1xp67_ASAP7_75t_L g1140 ( 
.A(n_954),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1091),
.A2(n_1074),
.B(n_1077),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_1064),
.B(n_1042),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_965),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_966),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_968),
.B(n_982),
.Y(n_1145)
);

AO31x2_ASAP7_75t_L g1146 ( 
.A1(n_990),
.A2(n_1007),
.A3(n_962),
.B(n_1000),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1003),
.B(n_1082),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1074),
.A2(n_1048),
.B(n_1020),
.Y(n_1148)
);

OAI21xp33_ASAP7_75t_L g1149 ( 
.A1(n_960),
.A2(n_1004),
.B(n_1005),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_1081),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_957),
.B(n_1057),
.Y(n_1151)
);

O2A1O1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_996),
.A2(n_1007),
.B(n_1000),
.C(n_1002),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_962),
.A2(n_1054),
.B(n_1065),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_1047),
.A2(n_951),
.B(n_1061),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_995),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1055),
.A2(n_1057),
.B(n_1056),
.Y(n_1156)
);

OA21x2_ASAP7_75t_L g1157 ( 
.A1(n_999),
.A2(n_1002),
.B(n_996),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_L g1158 ( 
.A1(n_1047),
.A2(n_1016),
.B(n_1044),
.Y(n_1158)
);

BUFx2_ASAP7_75t_L g1159 ( 
.A(n_958),
.Y(n_1159)
);

AO31x2_ASAP7_75t_L g1160 ( 
.A1(n_999),
.A2(n_1072),
.A3(n_1063),
.B(n_1053),
.Y(n_1160)
);

NOR2xp33_ASAP7_75t_L g1161 ( 
.A(n_981),
.B(n_1006),
.Y(n_1161)
);

AO32x2_ASAP7_75t_L g1162 ( 
.A1(n_997),
.A2(n_1019),
.A3(n_979),
.B1(n_1006),
.B2(n_972),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_995),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_987),
.B(n_989),
.Y(n_1164)
);

OR2x2_ASAP7_75t_L g1165 ( 
.A(n_997),
.B(n_972),
.Y(n_1165)
);

A2O1A1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_1073),
.A2(n_987),
.B(n_989),
.C(n_976),
.Y(n_1166)
);

OA21x2_ASAP7_75t_L g1167 ( 
.A1(n_1073),
.A2(n_974),
.B(n_972),
.Y(n_1167)
);

NAND3xp33_ASAP7_75t_L g1168 ( 
.A(n_1073),
.B(n_1079),
.C(n_992),
.Y(n_1168)
);

A2O1A1Ixp33_ASAP7_75t_L g1169 ( 
.A1(n_974),
.A2(n_1079),
.B(n_992),
.C(n_901),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_992),
.A2(n_1079),
.B1(n_527),
.B2(n_988),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_973),
.Y(n_1171)
);

INVx3_ASAP7_75t_L g1172 ( 
.A(n_958),
.Y(n_1172)
);

AOI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_1046),
.A2(n_466),
.B(n_450),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_1030),
.A2(n_889),
.B(n_955),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_973),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1046),
.A2(n_466),
.B(n_450),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1079),
.B(n_798),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1030),
.A2(n_889),
.B(n_955),
.Y(n_1178)
);

AND2x2_ASAP7_75t_L g1179 ( 
.A(n_1092),
.B(n_1088),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1079),
.B(n_798),
.Y(n_1180)
);

A2O1A1Ixp33_ASAP7_75t_L g1181 ( 
.A1(n_1079),
.A2(n_992),
.B(n_901),
.C(n_617),
.Y(n_1181)
);

AO31x2_ASAP7_75t_L g1182 ( 
.A1(n_1009),
.A2(n_1032),
.A3(n_1066),
.B(n_1071),
.Y(n_1182)
);

INVx5_ASAP7_75t_L g1183 ( 
.A(n_974),
.Y(n_1183)
);

AO31x2_ASAP7_75t_L g1184 ( 
.A1(n_1009),
.A2(n_1032),
.A3(n_1066),
.B(n_1071),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1011),
.A2(n_466),
.B(n_450),
.Y(n_1185)
);

OAI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1079),
.A2(n_1009),
.B(n_1037),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1030),
.A2(n_889),
.B(n_955),
.Y(n_1187)
);

A2O1A1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_1079),
.A2(n_992),
.B(n_901),
.C(n_617),
.Y(n_1188)
);

O2A1O1Ixp33_ASAP7_75t_SL g1189 ( 
.A1(n_1079),
.A2(n_828),
.B(n_1087),
.C(n_782),
.Y(n_1189)
);

AO31x2_ASAP7_75t_L g1190 ( 
.A1(n_1009),
.A2(n_1032),
.A3(n_1066),
.B(n_1071),
.Y(n_1190)
);

AND2x2_ASAP7_75t_L g1191 ( 
.A(n_1092),
.B(n_1088),
.Y(n_1191)
);

A2O1A1Ixp33_ASAP7_75t_L g1192 ( 
.A1(n_1079),
.A2(n_992),
.B(n_901),
.C(n_617),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_973),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_1030),
.A2(n_889),
.B(n_955),
.Y(n_1194)
);

O2A1O1Ixp33_ASAP7_75t_L g1195 ( 
.A1(n_1079),
.A2(n_992),
.B(n_617),
.C(n_1087),
.Y(n_1195)
);

OA21x2_ASAP7_75t_L g1196 ( 
.A1(n_1009),
.A2(n_1018),
.B(n_1011),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1046),
.A2(n_466),
.B(n_450),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_973),
.Y(n_1198)
);

INVx3_ASAP7_75t_L g1199 ( 
.A(n_958),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1046),
.A2(n_466),
.B(n_450),
.Y(n_1200)
);

AOI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1083),
.A2(n_1090),
.B(n_1084),
.Y(n_1201)
);

INVx3_ASAP7_75t_L g1202 ( 
.A(n_958),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1079),
.B(n_798),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1030),
.A2(n_889),
.B(n_955),
.Y(n_1204)
);

OAI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1079),
.A2(n_1009),
.B(n_1037),
.Y(n_1205)
);

AO31x2_ASAP7_75t_L g1206 ( 
.A1(n_1009),
.A2(n_1032),
.A3(n_1066),
.B(n_1071),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_973),
.Y(n_1207)
);

NAND3xp33_ASAP7_75t_SL g1208 ( 
.A(n_992),
.B(n_1079),
.C(n_827),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_973),
.Y(n_1209)
);

O2A1O1Ixp33_ASAP7_75t_SL g1210 ( 
.A1(n_1079),
.A2(n_828),
.B(n_1087),
.C(n_782),
.Y(n_1210)
);

BUFx6f_ASAP7_75t_L g1211 ( 
.A(n_1039),
.Y(n_1211)
);

INVxp67_ASAP7_75t_SL g1212 ( 
.A(n_950),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1079),
.B(n_798),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1030),
.A2(n_889),
.B(n_955),
.Y(n_1214)
);

BUFx10_ASAP7_75t_L g1215 ( 
.A(n_992),
.Y(n_1215)
);

INVx3_ASAP7_75t_L g1216 ( 
.A(n_958),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_992),
.A2(n_1087),
.B1(n_964),
.B2(n_901),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1046),
.A2(n_466),
.B(n_450),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1011),
.A2(n_466),
.B(n_450),
.Y(n_1219)
);

O2A1O1Ixp33_ASAP7_75t_SL g1220 ( 
.A1(n_1079),
.A2(n_828),
.B(n_1087),
.C(n_782),
.Y(n_1220)
);

AO31x2_ASAP7_75t_L g1221 ( 
.A1(n_1009),
.A2(n_1032),
.A3(n_1066),
.B(n_1071),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1079),
.B(n_798),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1046),
.A2(n_466),
.B(n_450),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_973),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1079),
.B(n_798),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_973),
.Y(n_1226)
);

OAI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1079),
.A2(n_1009),
.B(n_1037),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1046),
.A2(n_466),
.B(n_450),
.Y(n_1228)
);

A2O1A1Ixp33_ASAP7_75t_L g1229 ( 
.A1(n_1079),
.A2(n_992),
.B(n_901),
.C(n_617),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_973),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1030),
.A2(n_889),
.B(n_955),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1079),
.B(n_798),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1046),
.A2(n_466),
.B(n_450),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1011),
.A2(n_466),
.B(n_450),
.Y(n_1234)
);

O2A1O1Ixp33_ASAP7_75t_SL g1235 ( 
.A1(n_1079),
.A2(n_828),
.B(n_1087),
.C(n_782),
.Y(n_1235)
);

CKINVDCx11_ASAP7_75t_R g1236 ( 
.A(n_1121),
.Y(n_1236)
);

INVx2_ASAP7_75t_SL g1237 ( 
.A(n_1107),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1208),
.A2(n_1217),
.B1(n_1170),
.B2(n_1168),
.Y(n_1238)
);

INVx3_ASAP7_75t_L g1239 ( 
.A(n_1183),
.Y(n_1239)
);

INVx3_ASAP7_75t_L g1240 ( 
.A(n_1183),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_SL g1241 ( 
.A1(n_1215),
.A2(n_1117),
.B1(n_1161),
.B2(n_1170),
.Y(n_1241)
);

BUFx3_ASAP7_75t_L g1242 ( 
.A(n_1107),
.Y(n_1242)
);

BUFx6f_ASAP7_75t_L g1243 ( 
.A(n_1183),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1106),
.A2(n_1188),
.B1(n_1181),
.B2(n_1192),
.Y(n_1244)
);

CKINVDCx11_ASAP7_75t_R g1245 ( 
.A(n_1116),
.Y(n_1245)
);

AOI22xp33_ASAP7_75t_L g1246 ( 
.A1(n_1168),
.A2(n_1215),
.B1(n_1112),
.B2(n_1205),
.Y(n_1246)
);

CKINVDCx11_ASAP7_75t_R g1247 ( 
.A(n_1116),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1186),
.A2(n_1205),
.B1(n_1227),
.B2(n_1149),
.Y(n_1248)
);

INVx8_ASAP7_75t_L g1249 ( 
.A(n_1107),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1207),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1186),
.A2(n_1227),
.B1(n_1156),
.B2(n_1117),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1128),
.A2(n_1151),
.B1(n_1191),
.B2(n_1179),
.Y(n_1252)
);

BUFx3_ASAP7_75t_L g1253 ( 
.A(n_1104),
.Y(n_1253)
);

BUFx12f_ASAP7_75t_L g1254 ( 
.A(n_1116),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1151),
.A2(n_1145),
.B1(n_1113),
.B2(n_1138),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1110),
.B(n_1109),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1145),
.A2(n_1113),
.B1(n_1123),
.B2(n_1142),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_1211),
.Y(n_1258)
);

OAI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1229),
.A2(n_1109),
.B1(n_1169),
.B2(n_1110),
.Y(n_1259)
);

OAI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1144),
.A2(n_1142),
.B1(n_1130),
.B2(n_1120),
.Y(n_1260)
);

INVx6_ASAP7_75t_L g1261 ( 
.A(n_1183),
.Y(n_1261)
);

BUFx3_ASAP7_75t_L g1262 ( 
.A(n_1122),
.Y(n_1262)
);

BUFx10_ASAP7_75t_L g1263 ( 
.A(n_1211),
.Y(n_1263)
);

AOI22xp33_ASAP7_75t_L g1264 ( 
.A1(n_1120),
.A2(n_1132),
.B1(n_1232),
.B2(n_1225),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1101),
.Y(n_1265)
);

BUFx2_ASAP7_75t_L g1266 ( 
.A(n_1122),
.Y(n_1266)
);

OAI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1115),
.A2(n_1132),
.B1(n_1165),
.B2(n_1203),
.Y(n_1267)
);

AOI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1177),
.A2(n_1222),
.B1(n_1225),
.B2(n_1180),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1103),
.Y(n_1269)
);

INVx6_ASAP7_75t_L g1270 ( 
.A(n_1102),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_SL g1271 ( 
.A1(n_1167),
.A2(n_1232),
.B(n_1222),
.Y(n_1271)
);

OAI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1195),
.A2(n_1115),
.B1(n_1094),
.B2(n_1212),
.Y(n_1272)
);

INVx1_ASAP7_75t_SL g1273 ( 
.A(n_1140),
.Y(n_1273)
);

AOI22xp5_ASAP7_75t_SL g1274 ( 
.A1(n_1094),
.A2(n_1167),
.B1(n_1118),
.B2(n_1131),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1177),
.A2(n_1180),
.B1(n_1203),
.B2(n_1213),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1175),
.Y(n_1276)
);

AOI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1100),
.A2(n_1129),
.B1(n_1213),
.B2(n_1189),
.Y(n_1277)
);

CKINVDCx11_ASAP7_75t_R g1278 ( 
.A(n_1211),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1193),
.Y(n_1279)
);

BUFx3_ASAP7_75t_L g1280 ( 
.A(n_1134),
.Y(n_1280)
);

BUFx12f_ASAP7_75t_L g1281 ( 
.A(n_1159),
.Y(n_1281)
);

INVx1_ASAP7_75t_SL g1282 ( 
.A(n_1164),
.Y(n_1282)
);

BUFx10_ASAP7_75t_L g1283 ( 
.A(n_1198),
.Y(n_1283)
);

BUFx3_ASAP7_75t_L g1284 ( 
.A(n_1124),
.Y(n_1284)
);

BUFx12f_ASAP7_75t_L g1285 ( 
.A(n_1102),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1209),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1224),
.Y(n_1287)
);

AOI22xp33_ASAP7_75t_SL g1288 ( 
.A1(n_1157),
.A2(n_1095),
.B1(n_1196),
.B2(n_1226),
.Y(n_1288)
);

OAI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1133),
.A2(n_1230),
.B1(n_1166),
.B2(n_1148),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1157),
.A2(n_1135),
.B1(n_1150),
.B2(n_1143),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1095),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_1124),
.Y(n_1292)
);

CKINVDCx6p67_ASAP7_75t_R g1293 ( 
.A(n_1164),
.Y(n_1293)
);

BUFx2_ASAP7_75t_SL g1294 ( 
.A(n_1172),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1158),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1154),
.A2(n_1163),
.B1(n_1139),
.B2(n_1155),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_SL g1297 ( 
.A1(n_1162),
.A2(n_1153),
.B1(n_1210),
.B2(n_1235),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_SL g1298 ( 
.A1(n_1152),
.A2(n_1127),
.B(n_1111),
.Y(n_1298)
);

OAI21xp5_ASAP7_75t_SL g1299 ( 
.A1(n_1098),
.A2(n_1137),
.B(n_1126),
.Y(n_1299)
);

INVx2_ASAP7_75t_SL g1300 ( 
.A(n_1172),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1147),
.Y(n_1301)
);

INVx6_ASAP7_75t_L g1302 ( 
.A(n_1162),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1147),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1141),
.A2(n_1197),
.B1(n_1233),
.B2(n_1228),
.Y(n_1304)
);

INVx1_ASAP7_75t_SL g1305 ( 
.A(n_1199),
.Y(n_1305)
);

OAI22xp33_ASAP7_75t_SL g1306 ( 
.A1(n_1220),
.A2(n_1162),
.B1(n_1199),
.B2(n_1216),
.Y(n_1306)
);

BUFx6f_ASAP7_75t_L g1307 ( 
.A(n_1202),
.Y(n_1307)
);

BUFx10_ASAP7_75t_L g1308 ( 
.A(n_1119),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1141),
.A2(n_1176),
.B1(n_1223),
.B2(n_1173),
.Y(n_1309)
);

BUFx2_ASAP7_75t_L g1310 ( 
.A(n_1202),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_SL g1311 ( 
.A1(n_1114),
.A2(n_1185),
.B1(n_1219),
.B2(n_1234),
.Y(n_1311)
);

BUFx3_ASAP7_75t_L g1312 ( 
.A(n_1216),
.Y(n_1312)
);

INVx4_ASAP7_75t_L g1313 ( 
.A(n_1099),
.Y(n_1313)
);

CKINVDCx20_ASAP7_75t_R g1314 ( 
.A(n_1200),
.Y(n_1314)
);

OAI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1218),
.A2(n_1234),
.B1(n_1219),
.B2(n_1185),
.Y(n_1315)
);

BUFx4_ASAP7_75t_R g1316 ( 
.A(n_1105),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_SL g1317 ( 
.A1(n_1097),
.A2(n_1099),
.B1(n_1105),
.B2(n_1125),
.Y(n_1317)
);

CKINVDCx11_ASAP7_75t_R g1318 ( 
.A(n_1105),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1108),
.A2(n_1096),
.B1(n_1187),
.B2(n_1231),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1201),
.A2(n_1099),
.B1(n_1136),
.B2(n_1184),
.Y(n_1320)
);

AOI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1174),
.A2(n_1178),
.B1(n_1214),
.B2(n_1204),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1182),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1184),
.Y(n_1323)
);

AOI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1194),
.A2(n_1146),
.B1(n_1190),
.B2(n_1206),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1190),
.A2(n_1206),
.B1(n_1221),
.B2(n_1146),
.Y(n_1325)
);

CKINVDCx11_ASAP7_75t_R g1326 ( 
.A(n_1190),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1221),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1221),
.A2(n_1217),
.B1(n_617),
.B2(n_992),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1171),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1208),
.A2(n_992),
.B1(n_1087),
.B2(n_1217),
.Y(n_1330)
);

OAI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1181),
.A2(n_1079),
.B(n_1188),
.Y(n_1331)
);

CKINVDCx14_ASAP7_75t_R g1332 ( 
.A(n_1121),
.Y(n_1332)
);

OAI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1217),
.A2(n_617),
.B1(n_992),
.B2(n_1106),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_1121),
.Y(n_1334)
);

INVx4_ASAP7_75t_L g1335 ( 
.A(n_1183),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1208),
.A2(n_992),
.B1(n_1087),
.B2(n_1217),
.Y(n_1336)
);

OAI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1217),
.A2(n_617),
.B1(n_992),
.B2(n_1106),
.Y(n_1337)
);

OAI22xp33_ASAP7_75t_L g1338 ( 
.A1(n_1117),
.A2(n_862),
.B1(n_670),
.B2(n_827),
.Y(n_1338)
);

NAND2x1p5_ASAP7_75t_L g1339 ( 
.A(n_1183),
.B(n_1167),
.Y(n_1339)
);

CKINVDCx6p67_ASAP7_75t_R g1340 ( 
.A(n_1116),
.Y(n_1340)
);

INVx3_ASAP7_75t_L g1341 ( 
.A(n_1183),
.Y(n_1341)
);

BUFx2_ASAP7_75t_L g1342 ( 
.A(n_1160),
.Y(n_1342)
);

BUFx2_ASAP7_75t_L g1343 ( 
.A(n_1144),
.Y(n_1343)
);

BUFx3_ASAP7_75t_L g1344 ( 
.A(n_1107),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1104),
.Y(n_1345)
);

BUFx8_ASAP7_75t_SL g1346 ( 
.A(n_1116),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1171),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1208),
.A2(n_992),
.B1(n_1087),
.B2(n_1217),
.Y(n_1348)
);

CKINVDCx20_ASAP7_75t_R g1349 ( 
.A(n_1121),
.Y(n_1349)
);

BUFx4f_ASAP7_75t_SL g1350 ( 
.A(n_1121),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1171),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1208),
.A2(n_992),
.B1(n_1087),
.B2(n_1217),
.Y(n_1352)
);

OAI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1251),
.A2(n_1248),
.B1(n_1257),
.B2(n_1330),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1291),
.Y(n_1354)
);

BUFx2_ASAP7_75t_R g1355 ( 
.A(n_1346),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1322),
.Y(n_1356)
);

AND2x4_ASAP7_75t_L g1357 ( 
.A(n_1274),
.B(n_1295),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1264),
.B(n_1255),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1323),
.Y(n_1359)
);

BUFx2_ASAP7_75t_L g1360 ( 
.A(n_1342),
.Y(n_1360)
);

OA21x2_ASAP7_75t_L g1361 ( 
.A1(n_1298),
.A2(n_1299),
.B(n_1304),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1327),
.Y(n_1362)
);

HB1xp67_ASAP7_75t_L g1363 ( 
.A(n_1342),
.Y(n_1363)
);

AO21x1_ASAP7_75t_SL g1364 ( 
.A1(n_1277),
.A2(n_1331),
.B(n_1238),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1313),
.B(n_1302),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1315),
.A2(n_1309),
.B(n_1319),
.Y(n_1366)
);

OAI21xp33_ASAP7_75t_SL g1367 ( 
.A1(n_1313),
.A2(n_1352),
.B(n_1336),
.Y(n_1367)
);

AO21x2_ASAP7_75t_L g1368 ( 
.A1(n_1324),
.A2(n_1321),
.B(n_1320),
.Y(n_1368)
);

AO21x2_ASAP7_75t_L g1369 ( 
.A1(n_1325),
.A2(n_1271),
.B(n_1295),
.Y(n_1369)
);

BUFx3_ASAP7_75t_L g1370 ( 
.A(n_1293),
.Y(n_1370)
);

INVx2_ASAP7_75t_SL g1371 ( 
.A(n_1339),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1276),
.Y(n_1372)
);

INVx2_ASAP7_75t_SL g1373 ( 
.A(n_1339),
.Y(n_1373)
);

HB1xp67_ASAP7_75t_L g1374 ( 
.A(n_1289),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1256),
.B(n_1267),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_L g1376 ( 
.A(n_1343),
.B(n_1333),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1326),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1326),
.Y(n_1378)
);

INVxp67_ASAP7_75t_L g1379 ( 
.A(n_1265),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1288),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1269),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1279),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1318),
.B(n_1282),
.Y(n_1383)
);

NAND2x1_ASAP7_75t_L g1384 ( 
.A(n_1271),
.B(n_1261),
.Y(n_1384)
);

AND2x4_ASAP7_75t_L g1385 ( 
.A(n_1314),
.B(n_1296),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1290),
.A2(n_1259),
.B(n_1244),
.Y(n_1386)
);

A2O1A1Ixp33_ASAP7_75t_L g1387 ( 
.A1(n_1348),
.A2(n_1337),
.B(n_1246),
.C(n_1241),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1268),
.B(n_1275),
.Y(n_1388)
);

HB1xp67_ASAP7_75t_L g1389 ( 
.A(n_1306),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1286),
.Y(n_1390)
);

AO21x2_ASAP7_75t_L g1391 ( 
.A1(n_1328),
.A2(n_1260),
.B(n_1287),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1272),
.A2(n_1341),
.B(n_1240),
.Y(n_1392)
);

OR2x2_ASAP7_75t_L g1393 ( 
.A(n_1252),
.B(n_1273),
.Y(n_1393)
);

AND2x4_ASAP7_75t_L g1394 ( 
.A(n_1314),
.B(n_1329),
.Y(n_1394)
);

INVx2_ASAP7_75t_SL g1395 ( 
.A(n_1283),
.Y(n_1395)
);

INVx3_ASAP7_75t_L g1396 ( 
.A(n_1308),
.Y(n_1396)
);

HB1xp67_ASAP7_75t_L g1397 ( 
.A(n_1316),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1338),
.A2(n_1266),
.B1(n_1332),
.B2(n_1262),
.Y(n_1398)
);

INVx1_ASAP7_75t_SL g1399 ( 
.A(n_1293),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1347),
.Y(n_1400)
);

OAI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1297),
.A2(n_1311),
.B(n_1317),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1308),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1301),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1303),
.Y(n_1404)
);

BUFx4f_ASAP7_75t_SL g1405 ( 
.A(n_1254),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1250),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_1346),
.Y(n_1407)
);

INVx2_ASAP7_75t_SL g1408 ( 
.A(n_1261),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1239),
.A2(n_1341),
.B(n_1240),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1308),
.B(n_1351),
.Y(n_1410)
);

INVx2_ASAP7_75t_SL g1411 ( 
.A(n_1261),
.Y(n_1411)
);

BUFx2_ASAP7_75t_R g1412 ( 
.A(n_1334),
.Y(n_1412)
);

CKINVDCx20_ASAP7_75t_R g1413 ( 
.A(n_1350),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1310),
.B(n_1262),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1261),
.Y(n_1415)
);

BUFx2_ASAP7_75t_SL g1416 ( 
.A(n_1243),
.Y(n_1416)
);

OR2x2_ASAP7_75t_L g1417 ( 
.A(n_1393),
.B(n_1345),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1365),
.B(n_1307),
.Y(n_1418)
);

OA21x2_ASAP7_75t_L g1419 ( 
.A1(n_1401),
.A2(n_1300),
.B(n_1305),
.Y(n_1419)
);

AOI22xp5_ASAP7_75t_L g1420 ( 
.A1(n_1353),
.A2(n_1332),
.B1(n_1349),
.B2(n_1334),
.Y(n_1420)
);

OAI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1387),
.A2(n_1349),
.B(n_1253),
.Y(n_1421)
);

A2O1A1Ixp33_ASAP7_75t_L g1422 ( 
.A1(n_1374),
.A2(n_1249),
.B(n_1242),
.C(n_1344),
.Y(n_1422)
);

OAI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1353),
.A2(n_1253),
.B(n_1237),
.Y(n_1423)
);

INVxp67_ASAP7_75t_SL g1424 ( 
.A(n_1400),
.Y(n_1424)
);

OAI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1374),
.A2(n_1386),
.B(n_1367),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1372),
.Y(n_1426)
);

A2O1A1Ixp33_ASAP7_75t_L g1427 ( 
.A1(n_1367),
.A2(n_1249),
.B(n_1242),
.C(n_1243),
.Y(n_1427)
);

NOR2xp33_ASAP7_75t_SL g1428 ( 
.A(n_1355),
.B(n_1254),
.Y(n_1428)
);

A2O1A1Ixp33_ASAP7_75t_L g1429 ( 
.A1(n_1386),
.A2(n_1249),
.B(n_1243),
.C(n_1237),
.Y(n_1429)
);

BUFx2_ASAP7_75t_L g1430 ( 
.A(n_1370),
.Y(n_1430)
);

CKINVDCx16_ASAP7_75t_R g1431 ( 
.A(n_1413),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1372),
.Y(n_1432)
);

AOI21xp5_ASAP7_75t_L g1433 ( 
.A1(n_1361),
.A2(n_1335),
.B(n_1249),
.Y(n_1433)
);

AOI221x1_ASAP7_75t_SL g1434 ( 
.A1(n_1376),
.A2(n_1236),
.B1(n_1340),
.B2(n_1247),
.C(n_1245),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1412),
.B(n_1236),
.Y(n_1435)
);

A2O1A1Ixp33_ASAP7_75t_L g1436 ( 
.A1(n_1386),
.A2(n_1292),
.B(n_1294),
.C(n_1312),
.Y(n_1436)
);

AO21x2_ASAP7_75t_L g1437 ( 
.A1(n_1401),
.A2(n_1270),
.B(n_1285),
.Y(n_1437)
);

NOR2x1_ASAP7_75t_L g1438 ( 
.A(n_1370),
.B(n_1280),
.Y(n_1438)
);

OAI221xp5_ASAP7_75t_SL g1439 ( 
.A1(n_1398),
.A2(n_1340),
.B1(n_1280),
.B2(n_1312),
.C(n_1284),
.Y(n_1439)
);

NOR2xp33_ASAP7_75t_L g1440 ( 
.A(n_1412),
.B(n_1393),
.Y(n_1440)
);

AOI221xp5_ASAP7_75t_L g1441 ( 
.A1(n_1358),
.A2(n_1258),
.B1(n_1281),
.B2(n_1263),
.C(n_1245),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1402),
.B(n_1258),
.Y(n_1442)
);

OA21x2_ASAP7_75t_L g1443 ( 
.A1(n_1366),
.A2(n_1270),
.B(n_1285),
.Y(n_1443)
);

INVx3_ASAP7_75t_L g1444 ( 
.A(n_1409),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1397),
.B(n_1263),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1361),
.A2(n_1384),
.B(n_1375),
.Y(n_1446)
);

OR2x2_ASAP7_75t_L g1447 ( 
.A(n_1402),
.B(n_1281),
.Y(n_1447)
);

OR2x2_ASAP7_75t_L g1448 ( 
.A(n_1402),
.B(n_1247),
.Y(n_1448)
);

AOI221xp5_ASAP7_75t_L g1449 ( 
.A1(n_1358),
.A2(n_1278),
.B1(n_1375),
.B2(n_1388),
.C(n_1389),
.Y(n_1449)
);

INVx1_ASAP7_75t_SL g1450 ( 
.A(n_1355),
.Y(n_1450)
);

AO21x2_ASAP7_75t_L g1451 ( 
.A1(n_1366),
.A2(n_1278),
.B(n_1369),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1366),
.A2(n_1392),
.B(n_1384),
.Y(n_1452)
);

AO32x2_ASAP7_75t_L g1453 ( 
.A1(n_1371),
.A2(n_1373),
.A3(n_1395),
.B1(n_1411),
.B2(n_1408),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1410),
.B(n_1381),
.Y(n_1454)
);

OA21x2_ASAP7_75t_L g1455 ( 
.A1(n_1392),
.A2(n_1380),
.B(n_1362),
.Y(n_1455)
);

OAI21xp5_ASAP7_75t_L g1456 ( 
.A1(n_1388),
.A2(n_1361),
.B(n_1385),
.Y(n_1456)
);

OR2x2_ASAP7_75t_L g1457 ( 
.A(n_1377),
.B(n_1378),
.Y(n_1457)
);

NOR2x1_ASAP7_75t_SL g1458 ( 
.A(n_1364),
.B(n_1391),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1377),
.B(n_1378),
.Y(n_1459)
);

OA21x2_ASAP7_75t_L g1460 ( 
.A1(n_1392),
.A2(n_1359),
.B(n_1356),
.Y(n_1460)
);

NOR2xp33_ASAP7_75t_L g1461 ( 
.A(n_1394),
.B(n_1399),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1382),
.B(n_1390),
.Y(n_1462)
);

BUFx3_ASAP7_75t_L g1463 ( 
.A(n_1370),
.Y(n_1463)
);

OAI22xp5_ASAP7_75t_SL g1464 ( 
.A1(n_1405),
.A2(n_1407),
.B1(n_1399),
.B2(n_1385),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1394),
.B(n_1383),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1379),
.Y(n_1466)
);

AND2x4_ASAP7_75t_L g1467 ( 
.A(n_1371),
.B(n_1373),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1379),
.Y(n_1468)
);

O2A1O1Ixp33_ASAP7_75t_L g1469 ( 
.A1(n_1389),
.A2(n_1391),
.B(n_1385),
.C(n_1414),
.Y(n_1469)
);

AO32x2_ASAP7_75t_L g1470 ( 
.A1(n_1373),
.A2(n_1395),
.A3(n_1411),
.B1(n_1408),
.B2(n_1363),
.Y(n_1470)
);

BUFx2_ASAP7_75t_L g1471 ( 
.A(n_1453),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1460),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1455),
.B(n_1368),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1444),
.B(n_1368),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1466),
.B(n_1391),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1460),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1444),
.B(n_1369),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1451),
.B(n_1454),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1470),
.B(n_1369),
.Y(n_1479)
);

AOI221xp5_ASAP7_75t_L g1480 ( 
.A1(n_1469),
.A2(n_1385),
.B1(n_1391),
.B2(n_1383),
.C(n_1406),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1462),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1470),
.B(n_1361),
.Y(n_1482)
);

INVxp67_ASAP7_75t_SL g1483 ( 
.A(n_1424),
.Y(n_1483)
);

BUFx2_ASAP7_75t_L g1484 ( 
.A(n_1453),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1462),
.Y(n_1485)
);

NAND2x1p5_ASAP7_75t_L g1486 ( 
.A(n_1419),
.B(n_1357),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1451),
.B(n_1360),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1470),
.B(n_1354),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1470),
.B(n_1354),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1426),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1432),
.Y(n_1491)
);

BUFx2_ASAP7_75t_L g1492 ( 
.A(n_1453),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1453),
.B(n_1354),
.Y(n_1493)
);

BUFx2_ASAP7_75t_L g1494 ( 
.A(n_1467),
.Y(n_1494)
);

BUFx3_ASAP7_75t_L g1495 ( 
.A(n_1463),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1449),
.A2(n_1357),
.B1(n_1415),
.B2(n_1396),
.Y(n_1496)
);

NOR2xp33_ASAP7_75t_L g1497 ( 
.A(n_1431),
.B(n_1415),
.Y(n_1497)
);

HB1xp67_ASAP7_75t_L g1498 ( 
.A(n_1468),
.Y(n_1498)
);

OR2x2_ASAP7_75t_L g1499 ( 
.A(n_1446),
.B(n_1362),
.Y(n_1499)
);

AOI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1420),
.A2(n_1357),
.B1(n_1403),
.B2(n_1404),
.Y(n_1500)
);

HB1xp67_ASAP7_75t_L g1501 ( 
.A(n_1493),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1498),
.B(n_1456),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_1497),
.Y(n_1503)
);

BUFx2_ASAP7_75t_L g1504 ( 
.A(n_1486),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1471),
.B(n_1443),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1471),
.B(n_1443),
.Y(n_1506)
);

NAND3xp33_ASAP7_75t_L g1507 ( 
.A(n_1480),
.B(n_1421),
.C(n_1425),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1484),
.B(n_1443),
.Y(n_1508)
);

INVx1_ASAP7_75t_SL g1509 ( 
.A(n_1494),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1482),
.B(n_1452),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1484),
.B(n_1492),
.Y(n_1511)
);

INVx1_ASAP7_75t_SL g1512 ( 
.A(n_1494),
.Y(n_1512)
);

INVx3_ASAP7_75t_L g1513 ( 
.A(n_1472),
.Y(n_1513)
);

AO221x2_ASAP7_75t_L g1514 ( 
.A1(n_1480),
.A2(n_1464),
.B1(n_1423),
.B2(n_1465),
.C(n_1434),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1472),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1490),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1498),
.B(n_1458),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1475),
.B(n_1467),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1492),
.B(n_1452),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1490),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1496),
.A2(n_1437),
.B1(n_1419),
.B2(n_1440),
.Y(n_1521)
);

BUFx2_ASAP7_75t_L g1522 ( 
.A(n_1486),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1491),
.Y(n_1523)
);

OAI31xp33_ASAP7_75t_L g1524 ( 
.A1(n_1486),
.A2(n_1427),
.A3(n_1436),
.B(n_1439),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1482),
.B(n_1418),
.Y(n_1525)
);

OAI21xp5_ASAP7_75t_L g1526 ( 
.A1(n_1500),
.A2(n_1436),
.B(n_1427),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1476),
.Y(n_1527)
);

AND2x2_ASAP7_75t_L g1528 ( 
.A(n_1479),
.B(n_1493),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1478),
.B(n_1419),
.Y(n_1529)
);

CKINVDCx5p33_ASAP7_75t_R g1530 ( 
.A(n_1495),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1479),
.B(n_1467),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1475),
.B(n_1483),
.Y(n_1532)
);

INVx5_ASAP7_75t_L g1533 ( 
.A(n_1473),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1478),
.B(n_1457),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1534),
.B(n_1478),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1528),
.B(n_1479),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1532),
.B(n_1502),
.Y(n_1537)
);

BUFx2_ASAP7_75t_L g1538 ( 
.A(n_1504),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1513),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1528),
.B(n_1493),
.Y(n_1540)
);

NAND2xp5_ASAP7_75t_L g1541 ( 
.A(n_1532),
.B(n_1488),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1502),
.B(n_1488),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1528),
.B(n_1488),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1501),
.B(n_1489),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_1503),
.Y(n_1545)
);

AOI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1514),
.A2(n_1437),
.B1(n_1500),
.B2(n_1441),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1534),
.B(n_1499),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1534),
.B(n_1518),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1501),
.B(n_1489),
.Y(n_1549)
);

INVx1_ASAP7_75t_SL g1550 ( 
.A(n_1509),
.Y(n_1550)
);

BUFx2_ASAP7_75t_L g1551 ( 
.A(n_1504),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1518),
.B(n_1489),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1516),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1516),
.B(n_1481),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1516),
.B(n_1481),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1511),
.B(n_1474),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1520),
.Y(n_1557)
);

AND2x4_ASAP7_75t_L g1558 ( 
.A(n_1504),
.B(n_1477),
.Y(n_1558)
);

INVx2_ASAP7_75t_SL g1559 ( 
.A(n_1533),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1513),
.Y(n_1560)
);

INVx2_ASAP7_75t_SL g1561 ( 
.A(n_1533),
.Y(n_1561)
);

AND2x4_ASAP7_75t_L g1562 ( 
.A(n_1522),
.B(n_1477),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1520),
.B(n_1485),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1520),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1511),
.B(n_1533),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1513),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1529),
.B(n_1499),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1511),
.B(n_1474),
.Y(n_1568)
);

HB1xp67_ASAP7_75t_L g1569 ( 
.A(n_1523),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1523),
.Y(n_1570)
);

OR2x6_ASAP7_75t_L g1571 ( 
.A(n_1526),
.B(n_1433),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1569),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1569),
.Y(n_1573)
);

NAND4xp75_ASAP7_75t_L g1574 ( 
.A(n_1546),
.B(n_1524),
.C(n_1526),
.D(n_1438),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1553),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1553),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1557),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1537),
.B(n_1514),
.Y(n_1578)
);

INVx1_ASAP7_75t_SL g1579 ( 
.A(n_1545),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1537),
.B(n_1514),
.Y(n_1580)
);

HB1xp67_ASAP7_75t_L g1581 ( 
.A(n_1550),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1557),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1565),
.B(n_1531),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1565),
.B(n_1531),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1550),
.B(n_1514),
.Y(n_1585)
);

A2O1A1Ixp33_ASAP7_75t_L g1586 ( 
.A1(n_1546),
.A2(n_1507),
.B(n_1524),
.C(n_1435),
.Y(n_1586)
);

INVx1_ASAP7_75t_SL g1587 ( 
.A(n_1565),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1564),
.Y(n_1588)
);

INVx2_ASAP7_75t_L g1589 ( 
.A(n_1564),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1548),
.B(n_1514),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1570),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1548),
.B(n_1514),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1570),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1554),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1554),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1540),
.B(n_1531),
.Y(n_1596)
);

NOR2x1p5_ASAP7_75t_SL g1597 ( 
.A(n_1539),
.B(n_1515),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1547),
.B(n_1529),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1555),
.Y(n_1599)
);

AO221x1_ASAP7_75t_L g1600 ( 
.A1(n_1538),
.A2(n_1514),
.B1(n_1522),
.B2(n_1430),
.C(n_1507),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1555),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1547),
.B(n_1529),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1563),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1542),
.B(n_1507),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1563),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1540),
.B(n_1531),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1538),
.Y(n_1607)
);

A2O1A1Ixp33_ASAP7_75t_L g1608 ( 
.A1(n_1542),
.A2(n_1521),
.B(n_1508),
.C(n_1505),
.Y(n_1608)
);

NAND2x1_ASAP7_75t_L g1609 ( 
.A(n_1559),
.B(n_1522),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1541),
.B(n_1517),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1567),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1540),
.B(n_1505),
.Y(n_1612)
);

INVxp67_ASAP7_75t_L g1613 ( 
.A(n_1551),
.Y(n_1613)
);

NOR3xp33_ASAP7_75t_L g1614 ( 
.A(n_1586),
.B(n_1561),
.C(n_1559),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1578),
.B(n_1517),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1607),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1581),
.B(n_1567),
.Y(n_1617)
);

INVxp67_ASAP7_75t_SL g1618 ( 
.A(n_1585),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1580),
.B(n_1552),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1582),
.Y(n_1620)
);

INVx1_ASAP7_75t_SL g1621 ( 
.A(n_1607),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1596),
.B(n_1571),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1604),
.B(n_1543),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1611),
.B(n_1541),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1590),
.B(n_1543),
.Y(n_1625)
);

AOI22xp33_ASAP7_75t_L g1626 ( 
.A1(n_1600),
.A2(n_1571),
.B1(n_1437),
.B2(n_1521),
.Y(n_1626)
);

NOR3xp33_ASAP7_75t_L g1627 ( 
.A(n_1574),
.B(n_1561),
.C(n_1559),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1592),
.B(n_1552),
.Y(n_1628)
);

INVx3_ASAP7_75t_L g1629 ( 
.A(n_1609),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1596),
.B(n_1571),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1611),
.B(n_1535),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1582),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1589),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1574),
.B(n_1525),
.Y(n_1634)
);

NAND2x1_ASAP7_75t_L g1635 ( 
.A(n_1600),
.B(n_1561),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1594),
.B(n_1601),
.Y(n_1636)
);

NAND2xp33_ASAP7_75t_L g1637 ( 
.A(n_1579),
.B(n_1503),
.Y(n_1637)
);

INVx2_ASAP7_75t_SL g1638 ( 
.A(n_1609),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1588),
.Y(n_1639)
);

AOI22xp5_ASAP7_75t_L g1640 ( 
.A1(n_1608),
.A2(n_1571),
.B1(n_1428),
.B2(n_1461),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1606),
.B(n_1571),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1606),
.B(n_1571),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1613),
.B(n_1525),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1583),
.B(n_1543),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1588),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1583),
.B(n_1536),
.Y(n_1646)
);

HB1xp67_ASAP7_75t_L g1647 ( 
.A(n_1572),
.Y(n_1647)
);

INVxp67_ASAP7_75t_L g1648 ( 
.A(n_1573),
.Y(n_1648)
);

AOI32xp33_ASAP7_75t_L g1649 ( 
.A1(n_1627),
.A2(n_1587),
.A3(n_1584),
.B1(n_1508),
.B2(n_1506),
.Y(n_1649)
);

OAI221xp5_ASAP7_75t_SL g1650 ( 
.A1(n_1640),
.A2(n_1598),
.B1(n_1602),
.B2(n_1610),
.C(n_1448),
.Y(n_1650)
);

INVxp67_ASAP7_75t_L g1651 ( 
.A(n_1637),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1620),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1644),
.B(n_1584),
.Y(n_1653)
);

NOR2xp33_ASAP7_75t_L g1654 ( 
.A(n_1648),
.B(n_1450),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1618),
.B(n_1595),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1621),
.B(n_1595),
.Y(n_1656)
);

AOI221xp5_ASAP7_75t_L g1657 ( 
.A1(n_1614),
.A2(n_1605),
.B1(n_1603),
.B2(n_1599),
.C(n_1572),
.Y(n_1657)
);

OAI221xp5_ASAP7_75t_SL g1658 ( 
.A1(n_1640),
.A2(n_1602),
.B1(n_1598),
.B2(n_1448),
.C(n_1551),
.Y(n_1658)
);

AOI22xp33_ASAP7_75t_L g1659 ( 
.A1(n_1634),
.A2(n_1533),
.B1(n_1605),
.B2(n_1603),
.Y(n_1659)
);

OAI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1635),
.A2(n_1626),
.B1(n_1621),
.B2(n_1615),
.Y(n_1660)
);

AOI21xp5_ASAP7_75t_L g1661 ( 
.A1(n_1635),
.A2(n_1576),
.B(n_1575),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1620),
.Y(n_1662)
);

OAI21xp33_ASAP7_75t_SL g1663 ( 
.A1(n_1638),
.A2(n_1612),
.B(n_1599),
.Y(n_1663)
);

AOI211x1_ASAP7_75t_L g1664 ( 
.A1(n_1619),
.A2(n_1544),
.B(n_1549),
.C(n_1612),
.Y(n_1664)
);

AOI222xp33_ASAP7_75t_L g1665 ( 
.A1(n_1628),
.A2(n_1508),
.B1(n_1505),
.B2(n_1506),
.C1(n_1473),
.C2(n_1597),
.Y(n_1665)
);

AOI21xp5_ASAP7_75t_L g1666 ( 
.A1(n_1636),
.A2(n_1647),
.B(n_1638),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1623),
.B(n_1535),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1644),
.B(n_1556),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1616),
.B(n_1577),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1623),
.B(n_1591),
.Y(n_1670)
);

AOI22xp5_ASAP7_75t_L g1671 ( 
.A1(n_1625),
.A2(n_1473),
.B1(n_1530),
.B2(n_1506),
.Y(n_1671)
);

NOR2xp33_ASAP7_75t_L g1672 ( 
.A(n_1617),
.B(n_1625),
.Y(n_1672)
);

AOI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1636),
.A2(n_1593),
.B(n_1589),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1652),
.Y(n_1674)
);

AOI22xp5_ASAP7_75t_L g1675 ( 
.A1(n_1660),
.A2(n_1643),
.B1(n_1641),
.B2(n_1622),
.Y(n_1675)
);

AOI21xp5_ASAP7_75t_L g1676 ( 
.A1(n_1666),
.A2(n_1616),
.B(n_1629),
.Y(n_1676)
);

INVxp67_ASAP7_75t_L g1677 ( 
.A(n_1654),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1662),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1669),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1669),
.Y(n_1680)
);

OAI221xp5_ASAP7_75t_L g1681 ( 
.A1(n_1658),
.A2(n_1617),
.B1(n_1629),
.B2(n_1616),
.C(n_1631),
.Y(n_1681)
);

INVxp67_ASAP7_75t_L g1682 ( 
.A(n_1672),
.Y(n_1682)
);

NOR2xp33_ASAP7_75t_L g1683 ( 
.A(n_1651),
.B(n_1631),
.Y(n_1683)
);

INVx1_ASAP7_75t_SL g1684 ( 
.A(n_1655),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1656),
.Y(n_1685)
);

AOI22xp33_ASAP7_75t_L g1686 ( 
.A1(n_1657),
.A2(n_1622),
.B1(n_1642),
.B2(n_1641),
.Y(n_1686)
);

INVx1_ASAP7_75t_SL g1687 ( 
.A(n_1656),
.Y(n_1687)
);

OAI21xp5_ASAP7_75t_L g1688 ( 
.A1(n_1661),
.A2(n_1629),
.B(n_1630),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_L g1689 ( 
.A(n_1650),
.B(n_1630),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1670),
.Y(n_1690)
);

NAND2x1p5_ASAP7_75t_L g1691 ( 
.A(n_1653),
.B(n_1629),
.Y(n_1691)
);

AOI221xp5_ASAP7_75t_L g1692 ( 
.A1(n_1649),
.A2(n_1645),
.B1(n_1639),
.B2(n_1632),
.C(n_1642),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1674),
.Y(n_1693)
);

AOI211xp5_ASAP7_75t_L g1694 ( 
.A1(n_1681),
.A2(n_1663),
.B(n_1671),
.C(n_1673),
.Y(n_1694)
);

O2A1O1Ixp33_ASAP7_75t_L g1695 ( 
.A1(n_1687),
.A2(n_1665),
.B(n_1659),
.C(n_1639),
.Y(n_1695)
);

INVxp67_ASAP7_75t_L g1696 ( 
.A(n_1683),
.Y(n_1696)
);

NAND3xp33_ASAP7_75t_L g1697 ( 
.A(n_1675),
.B(n_1664),
.C(n_1645),
.Y(n_1697)
);

AOI21xp33_ASAP7_75t_L g1698 ( 
.A1(n_1677),
.A2(n_1667),
.B(n_1633),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1678),
.Y(n_1699)
);

NOR2xp33_ASAP7_75t_L g1700 ( 
.A(n_1682),
.B(n_1624),
.Y(n_1700)
);

AOI32xp33_ASAP7_75t_L g1701 ( 
.A1(n_1689),
.A2(n_1668),
.A3(n_1646),
.B1(n_1632),
.B2(n_1519),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1684),
.B(n_1646),
.Y(n_1702)
);

INVx1_ASAP7_75t_SL g1703 ( 
.A(n_1691),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1702),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1703),
.B(n_1690),
.Y(n_1705)
);

NOR3xp33_ASAP7_75t_L g1706 ( 
.A(n_1696),
.B(n_1685),
.C(n_1688),
.Y(n_1706)
);

NOR3x1_ASAP7_75t_L g1707 ( 
.A(n_1697),
.B(n_1680),
.C(n_1679),
.Y(n_1707)
);

INVx1_ASAP7_75t_SL g1708 ( 
.A(n_1698),
.Y(n_1708)
);

OAI21xp5_ASAP7_75t_SL g1709 ( 
.A1(n_1701),
.A2(n_1686),
.B(n_1692),
.Y(n_1709)
);

NOR4xp25_ASAP7_75t_L g1710 ( 
.A(n_1693),
.B(n_1633),
.C(n_1676),
.D(n_1624),
.Y(n_1710)
);

AOI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1694),
.A2(n_1691),
.B1(n_1676),
.B2(n_1633),
.Y(n_1711)
);

AOI211xp5_ASAP7_75t_L g1712 ( 
.A1(n_1695),
.A2(n_1459),
.B(n_1422),
.C(n_1519),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1700),
.B(n_1536),
.Y(n_1713)
);

OAI211xp5_ASAP7_75t_L g1714 ( 
.A1(n_1699),
.A2(n_1533),
.B(n_1519),
.C(n_1544),
.Y(n_1714)
);

OAI211xp5_ASAP7_75t_L g1715 ( 
.A1(n_1711),
.A2(n_1533),
.B(n_1530),
.C(n_1422),
.Y(n_1715)
);

AOI222xp33_ASAP7_75t_L g1716 ( 
.A1(n_1709),
.A2(n_1597),
.B1(n_1533),
.B2(n_1544),
.C1(n_1549),
.C2(n_1510),
.Y(n_1716)
);

OAI321xp33_ASAP7_75t_L g1717 ( 
.A1(n_1705),
.A2(n_1447),
.A3(n_1486),
.B1(n_1442),
.B2(n_1593),
.C(n_1487),
.Y(n_1717)
);

AOI211x1_ASAP7_75t_L g1718 ( 
.A1(n_1704),
.A2(n_1549),
.B(n_1556),
.C(n_1568),
.Y(n_1718)
);

AOI221xp5_ASAP7_75t_SL g1719 ( 
.A1(n_1708),
.A2(n_1509),
.B1(n_1512),
.B2(n_1568),
.C(n_1556),
.Y(n_1719)
);

HB1xp67_ASAP7_75t_L g1720 ( 
.A(n_1715),
.Y(n_1720)
);

AOI221xp5_ASAP7_75t_L g1721 ( 
.A1(n_1718),
.A2(n_1710),
.B1(n_1706),
.B2(n_1712),
.C(n_1707),
.Y(n_1721)
);

OAI211xp5_ASAP7_75t_L g1722 ( 
.A1(n_1716),
.A2(n_1714),
.B(n_1713),
.C(n_1533),
.Y(n_1722)
);

OAI221xp5_ASAP7_75t_L g1723 ( 
.A1(n_1719),
.A2(n_1714),
.B1(n_1533),
.B2(n_1447),
.C(n_1417),
.Y(n_1723)
);

OAI211xp5_ASAP7_75t_L g1724 ( 
.A1(n_1717),
.A2(n_1533),
.B(n_1512),
.C(n_1463),
.Y(n_1724)
);

NAND3xp33_ASAP7_75t_SL g1725 ( 
.A(n_1715),
.B(n_1442),
.C(n_1429),
.Y(n_1725)
);

NOR2xp33_ASAP7_75t_L g1726 ( 
.A(n_1720),
.B(n_1558),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1722),
.Y(n_1727)
);

XNOR2xp5_ASAP7_75t_L g1728 ( 
.A(n_1721),
.B(n_1445),
.Y(n_1728)
);

INVx2_ASAP7_75t_SL g1729 ( 
.A(n_1725),
.Y(n_1729)
);

NOR2xp67_ASAP7_75t_L g1730 ( 
.A(n_1724),
.B(n_1539),
.Y(n_1730)
);

INVx1_ASAP7_75t_SL g1731 ( 
.A(n_1729),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1727),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1728),
.Y(n_1733)
);

NAND2xp5_ASAP7_75t_L g1734 ( 
.A(n_1731),
.B(n_1726),
.Y(n_1734)
);

OAI22x1_ASAP7_75t_L g1735 ( 
.A1(n_1734),
.A2(n_1733),
.B1(n_1732),
.B2(n_1730),
.Y(n_1735)
);

AO22x2_ASAP7_75t_L g1736 ( 
.A1(n_1735),
.A2(n_1723),
.B1(n_1560),
.B2(n_1566),
.Y(n_1736)
);

INVx1_ASAP7_75t_SL g1737 ( 
.A(n_1736),
.Y(n_1737)
);

AOI21xp5_ASAP7_75t_L g1738 ( 
.A1(n_1737),
.A2(n_1566),
.B(n_1560),
.Y(n_1738)
);

OAI221xp5_ASAP7_75t_L g1739 ( 
.A1(n_1738),
.A2(n_1566),
.B1(n_1560),
.B2(n_1539),
.C(n_1515),
.Y(n_1739)
);

OAI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1739),
.A2(n_1568),
.B(n_1536),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1740),
.Y(n_1741)
);

AOI22x1_ASAP7_75t_L g1742 ( 
.A1(n_1740),
.A2(n_1416),
.B1(n_1408),
.B2(n_1411),
.Y(n_1742)
);

AOI221xp5_ASAP7_75t_L g1743 ( 
.A1(n_1741),
.A2(n_1562),
.B1(n_1558),
.B2(n_1527),
.C(n_1515),
.Y(n_1743)
);

AOI211xp5_ASAP7_75t_L g1744 ( 
.A1(n_1743),
.A2(n_1742),
.B(n_1562),
.C(n_1558),
.Y(n_1744)
);


endmodule