module fake_jpeg_4089_n_91 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_91);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_91;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_0),
.B(n_1),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_2),
.B(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx6_ASAP7_75t_SL g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

A2O1A1Ixp33_ASAP7_75t_L g23 ( 
.A1(n_18),
.A2(n_6),
.B(n_1),
.C(n_4),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_23),
.B(n_22),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g24 ( 
.A(n_21),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_18),
.B(n_0),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_22),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_14),
.A2(n_5),
.B1(n_8),
.B2(n_9),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_28),
.A2(n_15),
.B1(n_19),
.B2(n_12),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_15),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_24),
.A2(n_13),
.B(n_20),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_31),
.B(n_32),
.C(n_35),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_29),
.A2(n_17),
.B(n_14),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_33),
.B(n_38),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_34),
.B(n_36),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_29),
.A2(n_20),
.B(n_16),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_28),
.B(n_16),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_44),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_40),
.A2(n_43),
.B1(n_46),
.B2(n_47),
.Y(n_59)
);

NOR2x1_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_24),
.B(n_19),
.Y(n_42)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_25),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_26),
.B(n_5),
.Y(n_45)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_30),
.A2(n_19),
.B1(n_10),
.B2(n_11),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_46),
.A2(n_11),
.B1(n_41),
.B2(n_36),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_24),
.B(n_8),
.Y(n_47)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_48),
.A2(n_59),
.B1(n_34),
.B2(n_47),
.Y(n_66)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_35),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_51),
.B(n_53),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_39),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_57),
.B(n_33),
.Y(n_63)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_33),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_SL g76 ( 
.A(n_64),
.B(n_58),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_66),
.A2(n_68),
.B1(n_54),
.B2(n_49),
.Y(n_72)
);

XOR2xp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_31),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_69),
.C(n_70),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_50),
.A2(n_40),
.B1(n_43),
.B2(n_32),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_55),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_37),
.C(n_39),
.Y(n_78)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_54),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_58),
.Y(n_83)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_78),
.B(n_67),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_76),
.A2(n_61),
.B(n_74),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_79),
.A2(n_77),
.B(n_65),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_82),
.B(n_83),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

OAI21x1_ASAP7_75t_L g85 ( 
.A1(n_80),
.A2(n_68),
.B(n_73),
.Y(n_85)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_85),
.B(n_81),
.Y(n_87)
);

AOI21x1_ASAP7_75t_L g89 ( 
.A1(n_87),
.A2(n_86),
.B(n_79),
.Y(n_89)
);

MAJx2_ASAP7_75t_L g91 ( 
.A(n_89),
.B(n_90),
.C(n_71),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_88),
.A2(n_56),
.B(n_62),
.Y(n_90)
);


endmodule