module fake_jpeg_932_n_77 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_77);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_77;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_44;
wire n_24;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_61;
wire n_45;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_0),
.Y(n_28)
);

OAI21xp33_ASAP7_75t_L g34 ( 
.A1(n_28),
.A2(n_31),
.B(n_1),
.Y(n_34)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_32),
.Y(n_37)
);

AOI21xp33_ASAP7_75t_L g31 ( 
.A1(n_22),
.A2(n_19),
.B(n_18),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_38),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_22),
.C(n_28),
.Y(n_35)
);

AND2x2_ASAP7_75t_SL g43 ( 
.A(n_35),
.B(n_26),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_30),
.A2(n_27),
.B1(n_23),
.B2(n_25),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_36),
.A2(n_29),
.B1(n_32),
.B2(n_27),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_25),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_32),
.Y(n_48)
);

AND2x6_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_31),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_24),
.B(n_17),
.C(n_14),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_45),
.A2(n_37),
.B1(n_32),
.B2(n_33),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_50),
.C(n_2),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_49),
.A2(n_41),
.B1(n_43),
.B2(n_21),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_1),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_13),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_55),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_41),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_54),
.B(n_56),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_52),
.B(n_47),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_21),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_57),
.B(n_58),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_46),
.A2(n_2),
.B(n_3),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_4),
.C(n_5),
.Y(n_62)
);

XNOR2x2_ASAP7_75t_SL g60 ( 
.A(n_56),
.B(n_3),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_63),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_46),
.C(n_6),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_65),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_68)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_68),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_61),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g70 ( 
.A1(n_69),
.A2(n_64),
.B(n_9),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_66),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_66),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_73),
.A2(n_67),
.B(n_71),
.C(n_11),
.Y(n_74)
);

BUFx24_ASAP7_75t_SL g75 ( 
.A(n_74),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_8),
.Y(n_76)
);

FAx1_ASAP7_75t_SL g77 ( 
.A(n_76),
.B(n_10),
.CI(n_11),
.CON(n_77),
.SN(n_77)
);


endmodule