module fake_jpeg_5517_n_284 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_284);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_284;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

HB1xp67_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_5),
.B(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_5),
.B(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_SL g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_39),
.B(n_43),
.Y(n_93)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_42),
.Y(n_56)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_15),
.B(n_8),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_16),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_19),
.B(n_7),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_46),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_7),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_18),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_51),
.Y(n_72)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_52),
.B(n_53),
.Y(n_77)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_26),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_27),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_55),
.B(n_61),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_39),
.A2(n_18),
.B1(n_15),
.B2(n_32),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g100 ( 
.A1(n_58),
.A2(n_64),
.B(n_78),
.C(n_21),
.Y(n_100)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_27),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_62),
.A2(n_6),
.B(n_10),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVxp33_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_48),
.A2(n_16),
.B1(n_22),
.B2(n_34),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_53),
.A2(n_22),
.B1(n_16),
.B2(n_36),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_67),
.A2(n_88),
.B1(n_90),
.B2(n_92),
.Y(n_107)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

INVx3_ASAP7_75t_SL g70 ( 
.A(n_45),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_41),
.A2(n_22),
.B1(n_36),
.B2(n_29),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_73),
.A2(n_98),
.B1(n_23),
.B2(n_9),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_74),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_30),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_75),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_30),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_76),
.B(n_95),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_38),
.A2(n_35),
.B1(n_34),
.B2(n_29),
.Y(n_78)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_80),
.Y(n_113)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_35),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_82),
.B(n_83),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_44),
.B(n_20),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_39),
.A2(n_20),
.B1(n_28),
.B2(n_19),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_85),
.A2(n_91),
.B1(n_31),
.B2(n_23),
.Y(n_111)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_50),
.A2(n_24),
.B1(n_21),
.B2(n_23),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_39),
.A2(n_28),
.B1(n_31),
.B2(n_24),
.Y(n_91)
);

OA22x2_ASAP7_75t_L g92 ( 
.A1(n_48),
.A2(n_24),
.B1(n_31),
.B2(n_23),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_44),
.B(n_24),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_52),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_97),
.B(n_74),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_39),
.A2(n_31),
.B1(n_24),
.B2(n_21),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_100),
.B(n_111),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_92),
.A2(n_23),
.B(n_21),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_101),
.B(n_123),
.Y(n_132)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_114),
.B(n_13),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_55),
.B(n_0),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_93),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_92),
.A2(n_0),
.B(n_1),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_92),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_124),
.A2(n_125),
.B1(n_66),
.B2(n_94),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_93),
.A2(n_66),
.B1(n_61),
.B2(n_62),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_76),
.A2(n_2),
.B(n_3),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_126),
.A2(n_127),
.B(n_100),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_100),
.A2(n_58),
.B1(n_78),
.B2(n_64),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_128),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_75),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_129),
.B(n_153),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_96),
.Y(n_130)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_130),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_131),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_109),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_134),
.B(n_137),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_136),
.B(n_152),
.Y(n_183)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

AO22x1_ASAP7_75t_L g138 ( 
.A1(n_101),
.A2(n_70),
.B1(n_84),
.B2(n_57),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_138),
.A2(n_117),
.B(n_106),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_102),
.B(n_68),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_139),
.B(n_143),
.Y(n_171)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_141),
.Y(n_166)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_103),
.Y(n_141)
);

NAND3xp33_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_70),
.C(n_56),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_142),
.B(n_146),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_103),
.B(n_65),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_105),
.B(n_96),
.Y(n_144)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_144),
.Y(n_163)
);

NOR2x1_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_125),
.Y(n_145)
);

NOR2x1_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_127),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_105),
.B(n_77),
.Y(n_147)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_81),
.Y(n_148)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_148),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_149),
.A2(n_154),
.B1(n_110),
.B2(n_106),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_86),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_150),
.B(n_4),
.Y(n_187)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_156),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_107),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_97),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_113),
.B(n_60),
.Y(n_155)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_116),
.B(n_88),
.Y(n_157)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_157),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_116),
.B(n_120),
.Y(n_158)
);

INVxp33_ASAP7_75t_L g173 ( 
.A(n_158),
.Y(n_173)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_110),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_120),
.Y(n_169)
);

INVx5_ASAP7_75t_SL g160 ( 
.A(n_121),
.Y(n_160)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_160),
.Y(n_164)
);

AOI32xp33_ASAP7_75t_L g161 ( 
.A1(n_111),
.A2(n_84),
.A3(n_72),
.B1(n_69),
.B2(n_94),
.Y(n_161)
);

AOI32xp33_ASAP7_75t_L g184 ( 
.A1(n_161),
.A2(n_108),
.A3(n_74),
.B1(n_71),
.B2(n_87),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_165),
.A2(n_180),
.B(n_138),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_167),
.A2(n_193),
.B(n_160),
.Y(n_210)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_169),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_134),
.Y(n_170)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_170),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_128),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_150),
.A2(n_79),
.B(n_87),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_132),
.B(n_112),
.C(n_99),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_181),
.B(n_189),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_184),
.B(n_187),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_135),
.B(n_143),
.Y(n_186)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_186),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_136),
.B(n_112),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_192),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_132),
.B(n_135),
.C(n_139),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_151),
.A2(n_59),
.B1(n_99),
.B2(n_115),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_191),
.A2(n_149),
.B1(n_156),
.B2(n_160),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_145),
.B(n_141),
.C(n_133),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_145),
.B(n_74),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_166),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_196),
.Y(n_223)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_195),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_178),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_193),
.A2(n_133),
.B1(n_152),
.B2(n_153),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_197),
.A2(n_217),
.B1(n_183),
.B2(n_187),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_175),
.A2(n_146),
.B1(n_138),
.B2(n_154),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_198),
.A2(n_174),
.B1(n_201),
.B2(n_209),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_199),
.B(n_208),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_180),
.A2(n_153),
.B(n_161),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_201),
.Y(n_230)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_205),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_178),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_206),
.B(n_209),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_175),
.A2(n_159),
.B(n_129),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_179),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_165),
.A2(n_129),
.B(n_137),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_188),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_210),
.B(n_211),
.Y(n_225)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_171),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_168),
.Y(n_212)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_212),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_171),
.B(n_104),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_215),
.B(n_216),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_173),
.B(n_63),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_193),
.A2(n_192),
.B1(n_182),
.B2(n_167),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_189),
.C(n_181),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_221),
.C(n_232),
.Y(n_244)
);

AOI322xp5_ASAP7_75t_L g221 ( 
.A1(n_198),
.A2(n_174),
.A3(n_167),
.B1(n_183),
.B2(n_182),
.C1(n_184),
.C2(n_176),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_233),
.Y(n_240)
);

OA22x2_ASAP7_75t_L g226 ( 
.A1(n_199),
.A2(n_191),
.B1(n_182),
.B2(n_164),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_226),
.A2(n_227),
.B1(n_234),
.B2(n_237),
.Y(n_242)
);

NAND3xp33_ASAP7_75t_L g231 ( 
.A(n_196),
.B(n_172),
.C(n_190),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_231),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_190),
.C(n_172),
.Y(n_232)
);

NAND2x1_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_164),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_211),
.A2(n_179),
.B1(n_185),
.B2(n_163),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_207),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_214),
.A2(n_185),
.B1(n_163),
.B2(n_162),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_220),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_250),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_218),
.A2(n_195),
.B1(n_208),
.B2(n_206),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_239),
.A2(n_241),
.B1(n_247),
.B2(n_240),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_230),
.A2(n_197),
.B1(n_212),
.B2(n_217),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_225),
.B(n_215),
.Y(n_243)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_243),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_230),
.A2(n_226),
.B1(n_233),
.B2(n_222),
.Y(n_245)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_245),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_214),
.C(n_204),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_237),
.C(n_234),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_226),
.A2(n_203),
.B1(n_202),
.B2(n_194),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_233),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_249),
.Y(n_262)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_223),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_251),
.B(n_236),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_243),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_248),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_245),
.A2(n_226),
.B(n_225),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_255),
.A2(n_240),
.B(n_248),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_256),
.A2(n_259),
.B1(n_229),
.B2(n_244),
.Y(n_269)
);

AOI321xp33_ASAP7_75t_L g257 ( 
.A1(n_251),
.A2(n_224),
.A3(n_236),
.B1(n_227),
.B2(n_235),
.C(n_204),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_257),
.B(n_242),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_240),
.A2(n_232),
.B1(n_203),
.B2(n_202),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_242),
.C(n_244),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_263),
.A2(n_266),
.B(n_267),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_252),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_254),
.B(n_228),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_200),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_268),
.A2(n_261),
.B(n_200),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_269),
.B(n_260),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_270),
.B(n_272),
.C(n_275),
.Y(n_277)
);

NAND3xp33_ASAP7_75t_SL g271 ( 
.A(n_263),
.B(n_258),
.C(n_256),
.Y(n_271)
);

A2O1A1Ixp33_ASAP7_75t_SL g278 ( 
.A1(n_271),
.A2(n_276),
.B(n_259),
.C(n_265),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_264),
.A2(n_255),
.B(n_262),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_274),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_177),
.Y(n_276)
);

O2A1O1Ixp33_ASAP7_75t_L g281 ( 
.A1(n_278),
.A2(n_279),
.B(n_13),
.C(n_10),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_277),
.B(n_177),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_280),
.B(n_79),
.Y(n_283)
);

A2O1A1O1Ixp25_ASAP7_75t_L g282 ( 
.A1(n_281),
.A2(n_278),
.B(n_11),
.C(n_12),
.D(n_14),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_282),
.B(n_283),
.Y(n_284)
);


endmodule