module real_aes_556_n_222 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_222);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_222;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_578;
wire n_528;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_281;
wire n_496;
wire n_468;
wire n_234;
wire n_284;
wire n_656;
wire n_316;
wire n_532;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_504;
wire n_310;
wire n_455;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_430;
wire n_269;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_622;
wire n_470;
wire n_494;
wire n_377;
wire n_273;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_291;
wire n_498;
wire n_481;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_243;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_681;
wire n_456;
wire n_359;
wire n_312;
wire n_266;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_541;
wire n_224;
wire n_546;
wire n_587;
wire n_639;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_646;
wire n_650;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
XNOR2x1_ASAP7_75t_L g450 ( .A(n_0), .B(n_451), .Y(n_450) );
AOI22xp33_ASAP7_75t_L g279 ( .A1(n_1), .A2(n_202), .B1(n_280), .B2(n_281), .Y(n_279) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_2), .A2(n_210), .B1(n_289), .B2(n_348), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g453 ( .A1(n_3), .A2(n_122), .B1(n_454), .B2(n_456), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_4), .A2(n_134), .B1(n_387), .B2(n_388), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g613 ( .A1(n_5), .A2(n_118), .B1(n_280), .B2(n_281), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_6), .A2(n_106), .B1(n_671), .B2(n_672), .Y(n_670) );
AO22x2_ASAP7_75t_L g246 ( .A1(n_7), .A2(n_154), .B1(n_243), .B2(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g628 ( .A(n_7), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_8), .A2(n_155), .B1(n_265), .B2(n_402), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_9), .A2(n_204), .B1(n_268), .B2(n_591), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_10), .A2(n_94), .B1(n_349), .B2(n_408), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_11), .A2(n_172), .B1(n_507), .B2(n_509), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_12), .B(n_363), .Y(n_362) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_13), .Y(n_496) );
CKINVDCx20_ASAP7_75t_R g644 ( .A(n_14), .Y(n_644) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_15), .A2(n_146), .B1(n_408), .B2(n_474), .Y(n_473) );
AO22x2_ASAP7_75t_L g242 ( .A1(n_16), .A2(n_56), .B1(n_243), .B2(n_244), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g626 ( .A(n_16), .B(n_627), .Y(n_626) );
AOI22xp5_ASAP7_75t_L g564 ( .A1(n_17), .A2(n_184), .B1(n_465), .B2(n_509), .Y(n_564) );
AOI22xp33_ASAP7_75t_SL g588 ( .A1(n_18), .A2(n_72), .B1(n_271), .B2(n_589), .Y(n_588) );
CKINVDCx20_ASAP7_75t_R g604 ( .A(n_19), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_20), .A2(n_221), .B1(n_468), .B2(n_669), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_21), .A2(n_180), .B1(n_285), .B2(n_615), .Y(n_653) );
AO222x2_ASAP7_75t_SL g239 ( .A1(n_22), .A2(n_40), .B1(n_127), .B2(n_240), .C1(n_256), .C2(n_259), .Y(n_239) );
AO22x2_ASAP7_75t_L g416 ( .A1(n_23), .A2(n_417), .B1(n_447), .B2(n_448), .Y(n_416) );
INVx1_ASAP7_75t_L g448 ( .A(n_23), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g411 ( .A(n_24), .Y(n_411) );
AOI22xp5_ASAP7_75t_L g291 ( .A1(n_25), .A2(n_130), .B1(n_292), .B2(n_293), .Y(n_291) );
AOI22xp33_ASAP7_75t_L g264 ( .A1(n_26), .A2(n_123), .B1(n_265), .B2(n_268), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_27), .A2(n_162), .B1(n_442), .B2(n_443), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_28), .A2(n_168), .B1(n_383), .B2(n_424), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_29), .A2(n_201), .B1(n_382), .B2(n_384), .Y(n_381) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_30), .A2(n_197), .B1(n_271), .B2(n_274), .Y(n_610) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_31), .A2(n_632), .B1(n_655), .B2(n_656), .Y(n_631) );
CKINVDCx20_ASAP7_75t_R g655 ( .A(n_31), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_32), .A2(n_124), .B1(n_289), .B2(n_290), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_33), .A2(n_174), .B1(n_365), .B2(n_555), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_34), .A2(n_109), .B1(n_471), .B2(n_472), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g321 ( .A1(n_35), .A2(n_150), .B1(n_322), .B2(n_324), .Y(n_321) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_36), .A2(n_133), .B1(n_427), .B2(n_428), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_37), .A2(n_147), .B1(n_427), .B2(n_428), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_38), .A2(n_112), .B1(n_285), .B2(n_615), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_39), .A2(n_97), .B1(n_495), .B2(n_552), .Y(n_551) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_41), .Y(n_498) );
AOI22xp5_ASAP7_75t_L g503 ( .A1(n_42), .A2(n_205), .B1(n_504), .B2(n_505), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g350 ( .A1(n_43), .A2(n_152), .B1(n_351), .B2(n_354), .Y(n_350) );
AOI22xp5_ASAP7_75t_L g379 ( .A1(n_44), .A2(n_209), .B1(n_305), .B2(n_380), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_45), .A2(n_63), .B1(n_281), .B2(n_406), .Y(n_405) );
AOI22xp5_ASAP7_75t_L g368 ( .A1(n_46), .A2(n_95), .B1(n_369), .B2(n_370), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_47), .A2(n_76), .B1(n_271), .B2(n_274), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_48), .A2(n_93), .B1(n_265), .B2(n_402), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g674 ( .A1(n_49), .A2(n_213), .B1(n_437), .B2(n_460), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g567 ( .A1(n_50), .A2(n_208), .B1(n_334), .B2(n_408), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_51), .A2(n_136), .B1(n_284), .B2(n_285), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_52), .A2(n_104), .B1(n_271), .B2(n_274), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_53), .A2(n_148), .B1(n_434), .B2(n_435), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_54), .A2(n_121), .B1(n_240), .B2(n_256), .Y(n_637) );
AOI222xp33_ASAP7_75t_L g676 ( .A1(n_55), .A2(n_58), .B1(n_212), .B2(n_572), .C1(n_575), .C2(n_677), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_57), .A2(n_163), .B1(n_240), .B2(n_256), .Y(n_586) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_59), .Y(n_544) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_60), .A2(n_181), .B1(n_387), .B2(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g487 ( .A(n_61), .B(n_488), .Y(n_487) );
INVx3_ASAP7_75t_L g243 ( .A(n_62), .Y(n_243) );
AOI22xp33_ASAP7_75t_L g283 ( .A1(n_64), .A2(n_116), .B1(n_284), .B2(n_285), .Y(n_283) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_65), .A2(n_173), .B1(n_340), .B2(n_430), .Y(n_429) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_66), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_67), .A2(n_189), .B1(n_240), .B2(n_256), .Y(n_400) );
CKINVDCx20_ASAP7_75t_R g548 ( .A(n_68), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_69), .A2(n_211), .B1(n_240), .B2(n_256), .Y(n_608) );
OA22x2_ASAP7_75t_L g660 ( .A1(n_70), .A2(n_661), .B1(n_662), .B2(n_678), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_70), .Y(n_661) );
AOI222xp33_ASAP7_75t_L g571 ( .A1(n_71), .A2(n_84), .B1(n_156), .B2(n_572), .C1(n_573), .C2(n_575), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_73), .A2(n_200), .B1(n_280), .B2(n_281), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_74), .A2(n_107), .B1(n_367), .B2(n_460), .Y(n_459) );
INVx1_ASAP7_75t_SL g251 ( .A(n_75), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_75), .B(n_105), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_77), .A2(n_206), .B1(n_336), .B2(n_340), .Y(n_335) );
AOI22xp5_ASAP7_75t_SL g377 ( .A1(n_78), .A2(n_170), .B1(n_354), .B2(n_378), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_79), .A2(n_219), .B1(n_430), .B2(n_468), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g457 ( .A1(n_80), .A2(n_144), .B1(n_434), .B2(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g230 ( .A(n_81), .Y(n_230) );
AO22x1_ASAP7_75t_L g490 ( .A1(n_82), .A2(n_131), .B1(n_385), .B2(n_491), .Y(n_490) );
XOR2x2_ASAP7_75t_L g298 ( .A(n_83), .B(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_85), .B(n_462), .Y(n_607) );
CKINVDCx20_ASAP7_75t_R g518 ( .A(n_86), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g642 ( .A(n_87), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_88), .A2(n_115), .B1(n_347), .B2(n_351), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_89), .A2(n_100), .B1(n_330), .B2(n_369), .Y(n_512) );
CKINVDCx20_ASAP7_75t_R g522 ( .A(n_90), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g540 ( .A(n_91), .Y(n_540) );
AOI22xp33_ASAP7_75t_SL g594 ( .A1(n_92), .A2(n_149), .B1(n_280), .B2(n_281), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g570 ( .A1(n_96), .A2(n_198), .B1(n_367), .B2(n_495), .Y(n_570) );
INVx1_ASAP7_75t_L g482 ( .A(n_98), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_99), .A2(n_157), .B1(n_289), .B2(n_290), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g329 ( .A1(n_101), .A2(n_214), .B1(n_330), .B2(n_333), .Y(n_329) );
AOI22xp5_ASAP7_75t_L g313 ( .A1(n_102), .A2(n_215), .B1(n_314), .B2(n_317), .Y(n_313) );
AOI22xp33_ASAP7_75t_L g342 ( .A1(n_103), .A2(n_159), .B1(n_343), .B2(n_347), .Y(n_342) );
AO22x2_ASAP7_75t_L g254 ( .A1(n_105), .A2(n_165), .B1(n_243), .B2(n_255), .Y(n_254) );
CKINVDCx20_ASAP7_75t_R g533 ( .A(n_108), .Y(n_533) );
CKINVDCx20_ASAP7_75t_R g556 ( .A(n_110), .Y(n_556) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_111), .Y(n_537) );
AOI22xp5_ASAP7_75t_L g436 ( .A1(n_113), .A2(n_194), .B1(n_437), .B2(n_438), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g288 ( .A1(n_114), .A2(n_178), .B1(n_289), .B2(n_290), .Y(n_288) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_117), .A2(n_129), .B1(n_268), .B2(n_591), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_119), .A2(n_132), .B1(n_408), .B2(n_666), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_120), .A2(n_220), .B1(n_374), .B2(n_468), .Y(n_563) );
INVx1_ASAP7_75t_L g252 ( .A(n_125), .Y(n_252) );
CKINVDCx20_ASAP7_75t_R g640 ( .A(n_126), .Y(n_640) );
CKINVDCx20_ASAP7_75t_R g294 ( .A(n_128), .Y(n_294) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_135), .A2(n_179), .B1(n_389), .B2(n_427), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_137), .A2(n_207), .B1(n_465), .B2(n_466), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g301 ( .A1(n_138), .A2(n_182), .B1(n_302), .B2(n_305), .Y(n_301) );
INVx1_ASAP7_75t_L g359 ( .A(n_139), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_140), .A2(n_143), .B1(n_284), .B2(n_285), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_141), .A2(n_153), .B1(n_372), .B2(n_375), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_142), .B(n_310), .Y(n_403) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_145), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_151), .A2(n_196), .B1(n_292), .B2(n_293), .Y(n_598) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_158), .A2(n_176), .B1(n_402), .B2(n_591), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_160), .A2(n_193), .B1(n_289), .B2(n_290), .Y(n_595) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_161), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_164), .B(n_462), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_166), .A2(n_188), .B1(n_365), .B2(n_366), .Y(n_364) );
AOI211xp5_ASAP7_75t_L g222 ( .A1(n_167), .A2(n_223), .B(n_231), .C(n_630), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_169), .B(n_309), .Y(n_308) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_171), .A2(n_217), .B1(n_290), .B2(n_408), .Y(n_407) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_175), .B(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g624 ( .A(n_175), .Y(n_624) );
CKINVDCx20_ASAP7_75t_R g585 ( .A(n_177), .Y(n_585) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_183), .A2(n_187), .B1(n_348), .B2(n_408), .Y(n_616) );
INVx1_ASAP7_75t_L g226 ( .A(n_185), .Y(n_226) );
AND2x2_ASAP7_75t_R g658 ( .A(n_185), .B(n_624), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_186), .B(n_572), .Y(n_638) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_190), .Y(n_541) );
CKINVDCx20_ASAP7_75t_R g422 ( .A(n_191), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_192), .B(n_524), .Y(n_523) );
INVxp67_ASAP7_75t_L g228 ( .A(n_195), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g646 ( .A(n_199), .Y(n_646) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_203), .Y(n_500) );
AO21x2_ASAP7_75t_L g560 ( .A1(n_216), .A2(n_561), .B(n_576), .Y(n_560) );
INVx1_ASAP7_75t_L g578 ( .A(n_216), .Y(n_578) );
OA22x2_ASAP7_75t_L g599 ( .A1(n_216), .A2(n_561), .B1(n_578), .B2(n_600), .Y(n_599) );
XNOR2xp5_ASAP7_75t_L g580 ( .A(n_218), .B(n_581), .Y(n_580) );
AND2x4_ASAP7_75t_SL g223 ( .A(n_224), .B(n_227), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
OR2x2_ASAP7_75t_L g684 ( .A(n_225), .B(n_227), .Y(n_684) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g623 ( .A(n_226), .B(n_624), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_228), .B(n_229), .Y(n_227) );
AOI221xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_476), .B1(n_619), .B2(n_620), .C(n_621), .Y(n_231) );
INVx1_ASAP7_75t_L g620 ( .A(n_232), .Y(n_620) );
XOR2xp5_ASAP7_75t_L g232 ( .A(n_233), .B(n_393), .Y(n_232) );
AOI22xp5_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_295), .B1(n_296), .B2(n_392), .Y(n_233) );
INVx1_ASAP7_75t_L g392 ( .A(n_234), .Y(n_392) );
HB1xp67_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
XOR2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_294), .Y(n_236) );
NAND2x1_ASAP7_75t_L g237 ( .A(n_238), .B(n_277), .Y(n_237) );
NOR2x1_ASAP7_75t_L g238 ( .A(n_239), .B(n_263), .Y(n_238) );
INVx1_ASAP7_75t_SL g574 ( .A(n_240), .Y(n_574) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_240), .Y(n_677) );
AND2x4_ASAP7_75t_L g240 ( .A(n_241), .B(n_248), .Y(n_240) );
AND2x2_ASAP7_75t_L g265 ( .A(n_241), .B(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g293 ( .A(n_241), .B(n_286), .Y(n_293) );
AND2x4_ASAP7_75t_L g304 ( .A(n_241), .B(n_266), .Y(n_304) );
AND2x2_ASAP7_75t_L g316 ( .A(n_241), .B(n_248), .Y(n_316) );
AND2x4_ASAP7_75t_L g349 ( .A(n_241), .B(n_286), .Y(n_349) );
AND2x2_ASAP7_75t_L g591 ( .A(n_241), .B(n_266), .Y(n_591) );
AND2x4_ASAP7_75t_L g241 ( .A(n_242), .B(n_245), .Y(n_241) );
AND2x2_ASAP7_75t_L g258 ( .A(n_242), .B(n_246), .Y(n_258) );
INVx1_ASAP7_75t_L g262 ( .A(n_242), .Y(n_262) );
INVx1_ASAP7_75t_L g273 ( .A(n_242), .Y(n_273) );
INVx2_ASAP7_75t_L g244 ( .A(n_243), .Y(n_244) );
INVx1_ASAP7_75t_L g247 ( .A(n_243), .Y(n_247) );
OAI22x1_ASAP7_75t_L g249 ( .A1(n_243), .A2(n_250), .B1(n_251), .B2(n_252), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_243), .Y(n_250) );
INVx1_ASAP7_75t_L g255 ( .A(n_243), .Y(n_255) );
AND2x4_ASAP7_75t_L g261 ( .A(n_245), .B(n_262), .Y(n_261) );
INVxp67_ASAP7_75t_L g269 ( .A(n_245), .Y(n_269) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g272 ( .A(n_246), .B(n_273), .Y(n_272) );
AND2x4_ASAP7_75t_L g271 ( .A(n_248), .B(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g284 ( .A(n_248), .B(n_261), .Y(n_284) );
AND2x2_ASAP7_75t_L g323 ( .A(n_248), .B(n_272), .Y(n_323) );
AND2x4_ASAP7_75t_L g332 ( .A(n_248), .B(n_261), .Y(n_332) );
AND2x2_ASAP7_75t_L g615 ( .A(n_248), .B(n_261), .Y(n_615) );
AND2x2_ASAP7_75t_L g248 ( .A(n_249), .B(n_253), .Y(n_248) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_249), .Y(n_257) );
AND2x2_ASAP7_75t_L g260 ( .A(n_249), .B(n_254), .Y(n_260) );
INVx2_ASAP7_75t_L g267 ( .A(n_249), .Y(n_267) );
AND2x4_ASAP7_75t_L g286 ( .A(n_253), .B(n_267), .Y(n_286) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g266 ( .A(n_254), .B(n_267), .Y(n_266) );
BUFx2_ASAP7_75t_L g282 ( .A(n_254), .Y(n_282) );
AND2x2_ASAP7_75t_SL g256 ( .A(n_257), .B(n_258), .Y(n_256) );
AND2x2_ASAP7_75t_L g320 ( .A(n_257), .B(n_258), .Y(n_320) );
AND2x2_ASAP7_75t_SL g575 ( .A(n_257), .B(n_258), .Y(n_575) );
AND2x4_ASAP7_75t_L g281 ( .A(n_258), .B(n_282), .Y(n_281) );
AND2x4_ASAP7_75t_L g285 ( .A(n_258), .B(n_286), .Y(n_285) );
AND2x4_ASAP7_75t_L g334 ( .A(n_258), .B(n_286), .Y(n_334) );
AND2x4_ASAP7_75t_L g341 ( .A(n_258), .B(n_282), .Y(n_341) );
BUFx2_ASAP7_75t_L g572 ( .A(n_259), .Y(n_572) );
INVx2_ASAP7_75t_SL g584 ( .A(n_259), .Y(n_584) );
AND2x4_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
AND2x2_ASAP7_75t_L g268 ( .A(n_260), .B(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g274 ( .A(n_260), .B(n_275), .Y(n_274) );
AND2x4_ASAP7_75t_L g307 ( .A(n_260), .B(n_269), .Y(n_307) );
AND2x2_ASAP7_75t_L g312 ( .A(n_260), .B(n_261), .Y(n_312) );
AND2x4_ASAP7_75t_L g327 ( .A(n_260), .B(n_275), .Y(n_327) );
AND2x2_ASAP7_75t_L g402 ( .A(n_260), .B(n_269), .Y(n_402) );
AND2x2_ASAP7_75t_L g589 ( .A(n_260), .B(n_275), .Y(n_589) );
AND2x6_ASAP7_75t_L g289 ( .A(n_261), .B(n_266), .Y(n_289) );
AND2x2_ASAP7_75t_L g292 ( .A(n_261), .B(n_286), .Y(n_292) );
AND2x4_ASAP7_75t_L g346 ( .A(n_261), .B(n_286), .Y(n_346) );
AND2x2_ASAP7_75t_L g353 ( .A(n_261), .B(n_266), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_270), .Y(n_263) );
INVxp67_ASAP7_75t_L g645 ( .A(n_265), .Y(n_645) );
AND2x2_ASAP7_75t_SL g280 ( .A(n_266), .B(n_272), .Y(n_280) );
AND2x2_ASAP7_75t_L g339 ( .A(n_266), .B(n_272), .Y(n_339) );
AND2x2_ASAP7_75t_L g406 ( .A(n_266), .B(n_272), .Y(n_406) );
INVxp67_ASAP7_75t_L g647 ( .A(n_268), .Y(n_647) );
AND2x6_ASAP7_75t_L g290 ( .A(n_272), .B(n_286), .Y(n_290) );
AND2x4_ASAP7_75t_L g356 ( .A(n_272), .B(n_286), .Y(n_356) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_273), .Y(n_276) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NOR2x1_ASAP7_75t_L g277 ( .A(n_278), .B(n_287), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_283), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_291), .Y(n_287) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
OAI22xp5_ASAP7_75t_SL g296 ( .A1(n_297), .A2(n_357), .B1(n_358), .B2(n_391), .Y(n_296) );
INVx3_ASAP7_75t_L g391 ( .A(n_297), .Y(n_391) );
INVx5_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NOR2x1_ASAP7_75t_L g299 ( .A(n_300), .B(n_328), .Y(n_299) );
NAND4xp25_ASAP7_75t_L g300 ( .A(n_301), .B(n_308), .C(n_313), .D(n_321), .Y(n_300) );
BUFx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
BUFx2_ASAP7_75t_L g365 ( .A(n_303), .Y(n_365) );
INVx1_ASAP7_75t_L g499 ( .A(n_303), .Y(n_499) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
BUFx3_ASAP7_75t_L g434 ( .A(n_304), .Y(n_434) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx2_ASAP7_75t_SL g435 ( .A(n_306), .Y(n_435) );
INVx2_ASAP7_75t_L g458 ( .A(n_306), .Y(n_458) );
OAI22xp5_ASAP7_75t_L g497 ( .A1(n_306), .A2(n_498), .B1(n_499), .B2(n_500), .Y(n_497) );
INVx2_ASAP7_75t_L g555 ( .A(n_306), .Y(n_555) );
INVx6_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
BUFx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx4_ASAP7_75t_SL g310 ( .A(n_311), .Y(n_310) );
INVx3_ASAP7_75t_L g363 ( .A(n_311), .Y(n_363) );
INVx3_ASAP7_75t_SL g421 ( .A(n_311), .Y(n_421) );
INVx4_ASAP7_75t_SL g462 ( .A(n_311), .Y(n_462) );
BUFx2_ASAP7_75t_L g489 ( .A(n_311), .Y(n_489) );
INVx6_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
BUFx6f_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
BUFx3_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
BUFx3_ASAP7_75t_L g383 ( .A(n_316), .Y(n_383) );
INVx2_ASAP7_75t_L g455 ( .A(n_316), .Y(n_455) );
BUFx6f_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx3_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx2_ASAP7_75t_L g424 ( .A(n_319), .Y(n_424) );
INVx2_ASAP7_75t_L g456 ( .A(n_319), .Y(n_456) );
INVx3_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
BUFx12f_ASAP7_75t_L g385 ( .A(n_320), .Y(n_385) );
BUFx6f_ASAP7_75t_SL g380 ( .A(n_322), .Y(n_380) );
INVx1_ASAP7_75t_L g641 ( .A(n_322), .Y(n_641) );
BUFx6f_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx3_ASAP7_75t_L g439 ( .A(n_323), .Y(n_439) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_323), .Y(n_460) );
INVx3_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_325), .A2(n_493), .B1(n_494), .B2(n_496), .Y(n_492) );
BUFx2_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
BUFx3_ASAP7_75t_L g367 ( .A(n_327), .Y(n_367) );
BUFx6f_ASAP7_75t_SL g437 ( .A(n_327), .Y(n_437) );
INVx1_ASAP7_75t_L g553 ( .A(n_327), .Y(n_553) );
NAND4xp25_ASAP7_75t_L g328 ( .A(n_329), .B(n_335), .C(n_342), .D(n_350), .Y(n_328) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx2_ASAP7_75t_L g370 ( .A(n_331), .Y(n_370) );
INVx3_ASAP7_75t_L g471 ( .A(n_331), .Y(n_471) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_331), .A2(n_540), .B1(n_541), .B2(n_542), .Y(n_539) );
INVx6_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
BUFx3_ASAP7_75t_L g427 ( .A(n_332), .Y(n_427) );
BUFx2_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
BUFx2_ASAP7_75t_SL g369 ( .A(n_334), .Y(n_369) );
INVx2_ASAP7_75t_L g444 ( .A(n_334), .Y(n_444) );
BUFx3_ASAP7_75t_L g474 ( .A(n_334), .Y(n_474) );
BUFx3_ASAP7_75t_L g666 ( .A(n_334), .Y(n_666) );
BUFx6f_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g374 ( .A(n_338), .Y(n_374) );
INVx1_ASAP7_75t_L g669 ( .A(n_338), .Y(n_669) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
BUFx6f_ASAP7_75t_L g430 ( .A(n_339), .Y(n_430) );
BUFx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
BUFx3_ASAP7_75t_L g375 ( .A(n_341), .Y(n_375) );
INVx5_ASAP7_75t_SL g469 ( .A(n_341), .Y(n_469) );
BUFx6f_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g508 ( .A(n_344), .Y(n_508) );
INVx4_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx2_ASAP7_75t_L g378 ( .A(n_345), .Y(n_378) );
INVx3_ASAP7_75t_L g408 ( .A(n_345), .Y(n_408) );
INVx2_ASAP7_75t_SL g442 ( .A(n_345), .Y(n_442) );
INVx2_ASAP7_75t_SL g547 ( .A(n_345), .Y(n_547) );
INVx8_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
BUFx6f_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx2_ASAP7_75t_L g549 ( .A(n_348), .Y(n_549) );
BUFx6f_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g390 ( .A(n_349), .Y(n_390) );
BUFx3_ASAP7_75t_L g428 ( .A(n_349), .Y(n_428) );
BUFx6f_ASAP7_75t_L g472 ( .A(n_349), .Y(n_472) );
INVx2_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
INVx3_ASAP7_75t_L g465 ( .A(n_352), .Y(n_465) );
INVx2_ASAP7_75t_L g536 ( .A(n_352), .Y(n_536) );
INVx3_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
BUFx2_ASAP7_75t_L g387 ( .A(n_353), .Y(n_387) );
BUFx2_ASAP7_75t_L g671 ( .A(n_353), .Y(n_671) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g446 ( .A(n_355), .Y(n_446) );
INVx2_ASAP7_75t_L g466 ( .A(n_355), .Y(n_466) );
INVx2_ASAP7_75t_L g509 ( .A(n_355), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_355), .A2(n_533), .B1(n_534), .B2(n_537), .Y(n_532) );
INVx2_ASAP7_75t_L g672 ( .A(n_355), .Y(n_672) );
INVx8_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
XNOR2xp5_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
NOR2x1_ASAP7_75t_L g360 ( .A(n_361), .B(n_376), .Y(n_360) );
NAND4xp25_ASAP7_75t_L g361 ( .A(n_362), .B(n_364), .C(n_368), .D(n_371), .Y(n_361) );
BUFx6f_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g542 ( .A(n_369), .Y(n_542) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g504 ( .A(n_373), .Y(n_504) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
NAND4xp25_ASAP7_75t_L g376 ( .A(n_377), .B(n_379), .C(n_381), .D(n_386), .Y(n_376) );
INVx1_ASAP7_75t_SL g521 ( .A(n_382), .Y(n_521) );
BUFx6f_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
BUFx3_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx2_ASAP7_75t_L g525 ( .A(n_385), .Y(n_525) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AOI22xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_395), .B1(n_412), .B2(n_413), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
XNOR2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_411), .Y(n_396) );
NOR2x1_ASAP7_75t_L g397 ( .A(n_398), .B(n_404), .Y(n_397) );
NAND4xp25_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .C(n_401), .D(n_403), .Y(n_398) );
NAND4xp25_ASAP7_75t_L g404 ( .A(n_405), .B(n_407), .C(n_409), .D(n_410), .Y(n_404) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
OAI22xp33_ASAP7_75t_SL g413 ( .A1(n_414), .A2(n_415), .B1(n_449), .B2(n_475), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx3_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_SL g447 ( .A(n_417), .Y(n_447) );
AND2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_431), .Y(n_417) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_419), .B(n_425), .Y(n_418) );
OAI21xp33_ASAP7_75t_SL g419 ( .A1(n_420), .A2(n_422), .B(n_423), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
BUFx6f_ASAP7_75t_L g520 ( .A(n_421), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_426), .B(n_429), .Y(n_425) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_430), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g431 ( .A(n_432), .B(n_440), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_433), .B(n_436), .Y(n_432) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx4_ASAP7_75t_L g495 ( .A(n_439), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_441), .B(n_445), .Y(n_440) );
INVx2_ASAP7_75t_SL g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g475 ( .A(n_449), .Y(n_475) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
OR2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_463), .Y(n_451) );
NAND4xp25_ASAP7_75t_L g452 ( .A(n_453), .B(n_457), .C(n_459), .D(n_461), .Y(n_452) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g491 ( .A(n_455), .Y(n_491) );
NAND4xp25_ASAP7_75t_L g463 ( .A(n_464), .B(n_467), .C(n_470), .D(n_473), .Y(n_463) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g505 ( .A(n_469), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g527 ( .A1(n_469), .A2(n_528), .B1(n_529), .B2(n_531), .Y(n_527) );
INVx1_ASAP7_75t_L g619 ( .A(n_476), .Y(n_619) );
AOI22xp5_ASAP7_75t_SL g476 ( .A1(n_477), .A2(n_602), .B1(n_617), .B2(n_618), .Y(n_476) );
INVx1_ASAP7_75t_L g618 ( .A(n_477), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_479), .B1(n_557), .B2(n_558), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
XNOR2xp5_ASAP7_75t_L g480 ( .A(n_481), .B(n_514), .Y(n_480) );
OAI21x1_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_483), .B(n_513), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_482), .B(n_485), .Y(n_513) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_486), .B(n_501), .Y(n_485) );
NOR4xp75_ASAP7_75t_L g486 ( .A(n_487), .B(n_490), .C(n_492), .D(n_497), .Y(n_486) );
INVx2_ASAP7_75t_SL g488 ( .A(n_489), .Y(n_488) );
INVx2_ASAP7_75t_SL g494 ( .A(n_495), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_502), .B(n_510), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_503), .B(n_506), .Y(n_502) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_512), .Y(n_510) );
XNOR2x1_ASAP7_75t_L g514 ( .A(n_515), .B(n_556), .Y(n_514) );
NAND4xp75_ASAP7_75t_L g515 ( .A(n_516), .B(n_526), .C(n_538), .D(n_550), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
OAI221xp5_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_519), .B1(n_521), .B2(n_522), .C(n_523), .Y(n_517) );
INVx3_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
NOR2x1_ASAP7_75t_L g526 ( .A(n_527), .B(n_532), .Y(n_526) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
BUFx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
NOR2x1_ASAP7_75t_L g538 ( .A(n_539), .B(n_543), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g543 ( .A1(n_544), .A2(n_545), .B1(n_548), .B2(n_549), .Y(n_543) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
BUFx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AND2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_554), .Y(n_550) );
INVx2_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g639 ( .A1(n_553), .A2(n_640), .B1(n_641), .B2(n_642), .Y(n_639) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
OAI22xp33_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_579), .B1(n_599), .B2(n_601), .Y(n_558) );
INVx3_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
NOR2x1_ASAP7_75t_SL g576 ( .A(n_561), .B(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g600 ( .A(n_561), .Y(n_600) );
NAND4xp75_ASAP7_75t_L g561 ( .A(n_562), .B(n_565), .C(n_568), .D(n_571), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
AND2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
CKINVDCx20_ASAP7_75t_R g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g601 ( .A(n_579), .Y(n_601) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_SL g581 ( .A(n_582), .B(n_592), .Y(n_581) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_583), .B(n_587), .Y(n_582) );
OAI21xp5_ASAP7_75t_SL g583 ( .A1(n_584), .A2(n_585), .B(n_586), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_588), .B(n_590), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_593), .B(n_596), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
INVx2_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_603), .Y(n_617) );
XNOR2x1_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
NOR2x1_ASAP7_75t_L g605 ( .A(n_606), .B(n_611), .Y(n_605) );
NAND4xp25_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .C(n_609), .D(n_610), .Y(n_606) );
NAND4xp25_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .C(n_614), .D(n_616), .Y(n_611) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_623), .B(n_625), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_623), .B(n_626), .Y(n_681) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
OAI222xp33_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_657), .B1(n_659), .B2(n_661), .C1(n_679), .C2(n_682), .Y(n_630) );
CKINVDCx20_ASAP7_75t_R g656 ( .A(n_632), .Y(n_656) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_635), .B(n_648), .Y(n_634) );
NOR3xp33_ASAP7_75t_L g635 ( .A(n_636), .B(n_639), .C(n_643), .Y(n_635) );
NAND2xp5_ASAP7_75t_SL g636 ( .A(n_637), .B(n_638), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_645), .B1(n_646), .B2(n_647), .Y(n_643) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_649), .B(n_652), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
INVx1_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
BUFx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx2_ASAP7_75t_L g678 ( .A(n_662), .Y(n_678) );
NAND4xp75_ASAP7_75t_L g662 ( .A(n_663), .B(n_667), .C(n_673), .D(n_676), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
AND2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_670), .Y(n_667) );
AND2x2_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
CKINVDCx20_ASAP7_75t_R g679 ( .A(n_680), .Y(n_679) );
CKINVDCx6p67_ASAP7_75t_R g680 ( .A(n_681), .Y(n_680) );
CKINVDCx20_ASAP7_75t_R g682 ( .A(n_683), .Y(n_682) );
CKINVDCx20_ASAP7_75t_R g683 ( .A(n_684), .Y(n_683) );
endmodule