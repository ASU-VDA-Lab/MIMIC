module real_aes_18221_n_102 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_856, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_102);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_856;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_102;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_545;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_626;
wire n_400;
wire n_539;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_728;
wire n_713;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g846 ( .A(n_0), .B(n_847), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_1), .A2(n_34), .B1(n_144), .B2(n_181), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g555 ( .A1(n_2), .A2(n_10), .B1(n_507), .B2(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g847 ( .A(n_3), .Y(n_847) );
CKINVDCx5p33_ASAP7_75t_R g519 ( .A(n_4), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_5), .B(n_810), .Y(n_809) );
AOI22xp5_ASAP7_75t_L g542 ( .A1(n_6), .A2(n_11), .B1(n_543), .B2(n_544), .Y(n_542) );
OR2x2_ASAP7_75t_L g808 ( .A(n_7), .B(n_31), .Y(n_808) );
BUFx2_ASAP7_75t_L g852 ( .A(n_7), .Y(n_852) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_8), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g559 ( .A(n_9), .Y(n_559) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_12), .B(n_165), .Y(n_164) );
AOI22xp5_ASAP7_75t_L g506 ( .A1(n_13), .A2(n_99), .B1(n_237), .B2(n_507), .Y(n_506) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_14), .A2(n_30), .B1(n_524), .B2(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_15), .B(n_165), .Y(n_521) );
OAI21x1_ASAP7_75t_L g121 ( .A1(n_16), .A2(n_45), .B(n_122), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_17), .B(n_212), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g512 ( .A(n_18), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g833 ( .A1(n_19), .A2(n_87), .B1(n_483), .B2(n_834), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_19), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g533 ( .A1(n_20), .A2(n_38), .B1(n_143), .B2(n_242), .Y(n_533) );
CKINVDCx5p33_ASAP7_75t_R g132 ( .A(n_21), .Y(n_132) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_22), .A2(n_43), .B1(n_143), .B2(n_507), .Y(n_604) );
CKINVDCx5p33_ASAP7_75t_R g570 ( .A(n_23), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_24), .B(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_25), .B(n_175), .Y(n_210) );
CKINVDCx5p33_ASAP7_75t_R g587 ( .A(n_26), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_27), .B(n_152), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_28), .Y(n_236) );
CKINVDCx20_ASAP7_75t_R g841 ( .A(n_29), .Y(n_841) );
HB1xp67_ASAP7_75t_L g850 ( .A(n_31), .Y(n_850) );
AOI22xp5_ASAP7_75t_L g564 ( .A1(n_32), .A2(n_82), .B1(n_144), .B2(n_565), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_33), .A2(n_37), .B1(n_144), .B2(n_520), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_35), .A2(n_48), .B1(n_507), .B2(n_509), .Y(n_508) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_36), .Y(n_142) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_39), .B(n_165), .Y(n_196) );
INVx2_ASAP7_75t_L g803 ( .A(n_40), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_41), .B(n_200), .Y(n_207) );
BUFx3_ASAP7_75t_L g806 ( .A(n_42), .Y(n_806) );
INVx1_ASAP7_75t_L g830 ( .A(n_42), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_44), .B(n_147), .Y(n_215) );
AND2x2_ASAP7_75t_L g146 ( .A(n_46), .B(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_47), .B(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_49), .B(n_175), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_50), .B(n_242), .Y(n_241) );
AOI22xp5_ASAP7_75t_L g490 ( .A1(n_51), .A2(n_88), .B1(n_491), .B2(n_492), .Y(n_490) );
CKINVDCx5p33_ASAP7_75t_R g492 ( .A(n_51), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_52), .A2(n_70), .B1(n_242), .B2(n_509), .Y(n_603) );
AOI22xp33_ASAP7_75t_SL g102 ( .A1(n_53), .A2(n_103), .B1(n_842), .B2(n_853), .Y(n_102) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_54), .A2(n_73), .B1(n_144), .B2(n_520), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_55), .B(n_180), .Y(n_179) );
A2O1A1Ixp33_ASAP7_75t_L g128 ( .A1(n_56), .A2(n_129), .B(n_131), .C(n_134), .Y(n_128) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_57), .A2(n_96), .B1(n_507), .B2(n_544), .Y(n_584) );
AND2x4_ASAP7_75t_L g125 ( .A(n_58), .B(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g122 ( .A(n_59), .Y(n_122) );
AOI22xp33_ASAP7_75t_L g222 ( .A1(n_60), .A2(n_61), .B1(n_143), .B2(n_223), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_62), .B(n_152), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_63), .B(n_147), .Y(n_270) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_64), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_65), .B(n_143), .Y(n_199) );
INVx1_ASAP7_75t_L g126 ( .A(n_66), .Y(n_126) );
OAI22xp5_ASAP7_75t_L g832 ( .A1(n_67), .A2(n_833), .B1(n_835), .B2(n_836), .Y(n_832) );
CKINVDCx14_ASAP7_75t_R g835 ( .A(n_67), .Y(n_835) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_68), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_69), .B(n_152), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_71), .B(n_144), .Y(n_173) );
NAND3xp33_ASAP7_75t_L g208 ( .A(n_72), .B(n_181), .C(n_200), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_74), .B(n_144), .Y(n_156) );
INVx2_ASAP7_75t_L g136 ( .A(n_75), .Y(n_136) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_76), .B(n_165), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g264 ( .A(n_77), .B(n_214), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_78), .B(n_161), .Y(n_160) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_79), .A2(n_95), .B1(n_129), .B2(n_143), .Y(n_566) );
CKINVDCx5p33_ASAP7_75t_R g606 ( .A(n_80), .Y(n_606) );
CKINVDCx5p33_ASAP7_75t_R g536 ( .A(n_81), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g219 ( .A1(n_83), .A2(n_90), .B1(n_175), .B2(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_84), .B(n_165), .Y(n_238) );
NAND2xp33_ASAP7_75t_SL g269 ( .A(n_85), .B(n_158), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_86), .B(n_195), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_87), .B(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g483 ( .A(n_87), .Y(n_483) );
CKINVDCx5p33_ASAP7_75t_R g491 ( .A(n_88), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_89), .B(n_152), .Y(n_528) );
CKINVDCx5p33_ASAP7_75t_R g549 ( .A(n_91), .Y(n_549) );
INVx1_ASAP7_75t_L g488 ( .A(n_92), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g828 ( .A(n_92), .B(n_829), .Y(n_828) );
NAND2xp33_ASAP7_75t_L g525 ( .A(n_93), .B(n_165), .Y(n_525) );
NAND2xp33_ASAP7_75t_L g157 ( .A(n_94), .B(n_158), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_97), .B(n_147), .Y(n_183) );
NAND3xp33_ASAP7_75t_L g265 ( .A(n_98), .B(n_158), .C(n_214), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_100), .B(n_144), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_101), .B(n_175), .Y(n_178) );
OAI21x1_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_817), .B(n_821), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
A2O1A1Ixp33_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_489), .B(n_800), .C(n_809), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_107), .B(n_482), .Y(n_106) );
NAND2xp5_ASAP7_75t_SL g820 ( .A(n_107), .B(n_482), .Y(n_820) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_109), .A2(n_483), .B(n_484), .Y(n_482) );
XNOR2xp5_ASAP7_75t_L g831 ( .A(n_109), .B(n_832), .Y(n_831) );
AND2x4_ASAP7_75t_L g109 ( .A(n_110), .B(n_370), .Y(n_109) );
NOR4xp75_ASAP7_75t_L g110 ( .A(n_111), .B(n_309), .C(n_333), .D(n_352), .Y(n_110) );
NAND3x1_ASAP7_75t_L g111 ( .A(n_112), .B(n_249), .C(n_300), .Y(n_111) );
AOI22xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_184), .B1(n_227), .B2(n_245), .Y(n_112) );
AND2x2_ASAP7_75t_L g431 ( .A(n_113), .B(n_306), .Y(n_431) );
AND2x2_ASAP7_75t_L g113 ( .A(n_114), .B(n_149), .Y(n_113) );
AND2x2_ASAP7_75t_L g381 ( .A(n_114), .B(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_114), .B(n_386), .Y(n_385) );
INVx2_ASAP7_75t_L g408 ( .A(n_114), .Y(n_408) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g253 ( .A(n_115), .Y(n_253) );
INVx2_ASAP7_75t_L g275 ( .A(n_115), .Y(n_275) );
AND2x2_ASAP7_75t_L g369 ( .A(n_115), .B(n_332), .Y(n_369) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g248 ( .A(n_116), .Y(n_248) );
AND2x2_ASAP7_75t_L g348 ( .A(n_116), .B(n_260), .Y(n_348) );
AOI21x1_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_127), .B(n_146), .Y(n_116) );
NOR2xp67_ASAP7_75t_SL g117 ( .A(n_118), .B(n_123), .Y(n_117) );
INVx2_ASAP7_75t_L g510 ( .A(n_118), .Y(n_510) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AO31x2_ASAP7_75t_L g217 ( .A1(n_119), .A2(n_124), .A3(n_218), .B(n_224), .Y(n_217) );
NOR2xp33_ASAP7_75t_SL g548 ( .A(n_119), .B(n_549), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_119), .B(n_570), .Y(n_569) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g148 ( .A(n_120), .Y(n_148) );
INVx2_ASAP7_75t_L g226 ( .A(n_120), .Y(n_226) );
INVx2_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_121), .Y(n_153) );
INVx1_ASAP7_75t_L g504 ( .A(n_123), .Y(n_504) );
INVx2_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AO31x2_ASAP7_75t_L g530 ( .A1(n_124), .A2(n_531), .A3(n_534), .B(n_535), .Y(n_530) );
AO31x2_ASAP7_75t_L g540 ( .A1(n_124), .A2(n_541), .A3(n_547), .B(n_548), .Y(n_540) );
AO31x2_ASAP7_75t_L g551 ( .A1(n_124), .A2(n_552), .A3(n_557), .B(n_558), .Y(n_551) );
BUFx10_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
BUFx10_ASAP7_75t_L g167 ( .A(n_125), .Y(n_167) );
INVx1_ASAP7_75t_L g527 ( .A(n_125), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_137), .Y(n_127) );
INVx1_ASAP7_75t_L g163 ( .A(n_129), .Y(n_163) );
INVx1_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g133 ( .A(n_130), .Y(n_133) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_130), .Y(n_143) );
INVx3_ASAP7_75t_L g144 ( .A(n_130), .Y(n_144) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_130), .Y(n_158) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_130), .Y(n_165) );
INVx1_ASAP7_75t_L g176 ( .A(n_130), .Y(n_176) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_130), .Y(n_181) );
INVx1_ASAP7_75t_L g195 ( .A(n_130), .Y(n_195) );
INVx1_ASAP7_75t_L g223 ( .A(n_130), .Y(n_223) );
INVx1_ASAP7_75t_L g268 ( .A(n_130), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
INVx2_ASAP7_75t_SL g565 ( .A(n_133), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_134), .A2(n_156), .B(n_157), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_134), .A2(n_173), .B(n_174), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_134), .A2(n_194), .B(n_196), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_134), .A2(n_267), .B(n_269), .Y(n_266) );
BUFx4f_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g140 ( .A(n_136), .Y(n_140) );
BUFx8_ASAP7_75t_L g200 ( .A(n_136), .Y(n_200) );
INVx1_ASAP7_75t_L g214 ( .A(n_136), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_141), .Y(n_137) );
OAI22xp5_ASAP7_75t_L g218 ( .A1(n_138), .A2(n_219), .B1(n_221), .B2(n_222), .Y(n_218) );
OAI22xp5_ASAP7_75t_L g505 ( .A1(n_138), .A2(n_221), .B1(n_506), .B2(n_508), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g531 ( .A1(n_138), .A2(n_221), .B1(n_532), .B2(n_533), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_138), .A2(n_221), .B1(n_553), .B2(n_555), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g602 ( .A1(n_138), .A2(n_221), .B1(n_603), .B2(n_604), .Y(n_602) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g182 ( .A(n_139), .Y(n_182) );
BUFx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g162 ( .A(n_140), .Y(n_162) );
OAI22xp33_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_143), .B1(n_144), .B2(n_145), .Y(n_141) );
OAI21xp5_ASAP7_75t_L g206 ( .A1(n_143), .A2(n_207), .B(n_208), .Y(n_206) );
INVx2_ASAP7_75t_L g220 ( .A(n_143), .Y(n_220) );
INVx1_ASAP7_75t_L g509 ( .A(n_144), .Y(n_509) );
INVx4_ASAP7_75t_L g520 ( .A(n_144), .Y(n_520) );
INVx1_ASAP7_75t_L g544 ( .A(n_144), .Y(n_544) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g170 ( .A(n_148), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_148), .B(n_512), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_148), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g301 ( .A(n_149), .B(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g416 ( .A(n_149), .Y(n_416) );
AND2x2_ASAP7_75t_L g422 ( .A(n_149), .B(n_286), .Y(n_422) );
AND2x2_ASAP7_75t_L g149 ( .A(n_150), .B(n_168), .Y(n_149) );
INVx1_ASAP7_75t_L g258 ( .A(n_150), .Y(n_258) );
INVx4_ASAP7_75t_L g279 ( .A(n_150), .Y(n_279) );
OR2x2_ASAP7_75t_L g328 ( .A(n_150), .B(n_308), .Y(n_328) );
BUFx2_ASAP7_75t_L g397 ( .A(n_150), .Y(n_397) );
AND2x4_ASAP7_75t_L g150 ( .A(n_151), .B(n_154), .Y(n_150) );
INVx2_ASAP7_75t_L g534 ( .A(n_152), .Y(n_534) );
INVx4_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
AND2x4_ASAP7_75t_SL g166 ( .A(n_153), .B(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g191 ( .A(n_153), .Y(n_191) );
INVx1_ASAP7_75t_SL g261 ( .A(n_153), .Y(n_261) );
INVx2_ASAP7_75t_SL g516 ( .A(n_153), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_153), .B(n_536), .Y(n_535) );
BUFx3_ASAP7_75t_L g557 ( .A(n_153), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_153), .B(n_559), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_153), .B(n_587), .Y(n_586) );
OAI21x1_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_159), .B(n_166), .Y(n_154) );
INVx2_ASAP7_75t_L g242 ( .A(n_158), .Y(n_242) );
INVx1_ASAP7_75t_L g524 ( .A(n_158), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_162), .B1(n_163), .B2(n_164), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_161), .A2(n_240), .B(n_241), .Y(n_239) );
INVx2_ASAP7_75t_SL g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g212 ( .A(n_165), .Y(n_212) );
OAI21xp5_ASAP7_75t_L g263 ( .A1(n_165), .A2(n_264), .B(n_265), .Y(n_263) );
INVx3_ASAP7_75t_L g507 ( .A(n_165), .Y(n_507) );
OAI21x1_ASAP7_75t_L g171 ( .A1(n_167), .A2(n_172), .B(n_177), .Y(n_171) );
OAI21x1_ASAP7_75t_L g192 ( .A1(n_167), .A2(n_193), .B(n_197), .Y(n_192) );
OAI21x1_ASAP7_75t_L g205 ( .A1(n_167), .A2(n_206), .B(n_209), .Y(n_205) );
OAI21x1_ASAP7_75t_L g234 ( .A1(n_167), .A2(n_235), .B(n_239), .Y(n_234) );
OAI21x1_ASAP7_75t_L g262 ( .A1(n_167), .A2(n_263), .B(n_266), .Y(n_262) );
AND2x2_ASAP7_75t_L g247 ( .A(n_168), .B(n_248), .Y(n_247) );
INVx2_ASAP7_75t_L g350 ( .A(n_168), .Y(n_350) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g274 ( .A(n_169), .Y(n_274) );
OAI21x1_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_171), .B(n_183), .Y(n_169) );
OAI21xp5_ASAP7_75t_L g233 ( .A1(n_170), .A2(n_234), .B(n_243), .Y(n_233) );
OAI21xp33_ASAP7_75t_SL g288 ( .A1(n_170), .A2(n_171), .B(n_183), .Y(n_288) );
OAI21x1_ASAP7_75t_L g299 ( .A1(n_170), .A2(n_234), .B(n_243), .Y(n_299) );
INVx1_ASAP7_75t_L g543 ( .A(n_175), .Y(n_543) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_179), .B(n_182), .Y(n_177) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
NAND2x1_ASAP7_75t_L g419 ( .A(n_186), .B(n_359), .Y(n_419) );
AND2x4_ASAP7_75t_L g186 ( .A(n_187), .B(n_202), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
OR2x2_ASAP7_75t_L g304 ( .A(n_188), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g324 ( .A(n_188), .B(n_325), .Y(n_324) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_188), .Y(n_358) );
INVx3_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AND2x2_ASAP7_75t_L g314 ( .A(n_189), .B(n_204), .Y(n_314) );
NOR2xp67_ASAP7_75t_L g469 ( .A(n_189), .B(n_203), .Y(n_469) );
BUFx3_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx1_ASAP7_75t_L g391 ( .A(n_190), .Y(n_391) );
OAI21x1_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .B(n_201), .Y(n_190) );
OAI21x1_ASAP7_75t_L g204 ( .A1(n_191), .A2(n_205), .B(n_215), .Y(n_204) );
OAI21x1_ASAP7_75t_L g231 ( .A1(n_191), .A2(n_192), .B(n_201), .Y(n_231) );
OA21x2_ASAP7_75t_L g244 ( .A1(n_191), .A2(n_205), .B(n_215), .Y(n_244) );
INVx2_ASAP7_75t_L g237 ( .A(n_195), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_199), .B(n_200), .Y(n_197) );
INVx6_ASAP7_75t_L g221 ( .A(n_200), .Y(n_221) );
O2A1O1Ixp5_ASAP7_75t_L g235 ( .A1(n_200), .A2(n_236), .B(n_237), .C(n_238), .Y(n_235) );
O2A1O1Ixp5_ASAP7_75t_L g518 ( .A1(n_200), .A2(n_519), .B(n_520), .C(n_521), .Y(n_518) );
INVx2_ASAP7_75t_L g412 ( .A(n_202), .Y(n_412) );
AND2x4_ASAP7_75t_L g450 ( .A(n_202), .B(n_389), .Y(n_450) );
AND2x4_ASAP7_75t_L g202 ( .A(n_203), .B(n_216), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g290 ( .A(n_204), .Y(n_290) );
AND2x2_ASAP7_75t_L g325 ( .A(n_204), .B(n_217), .Y(n_325) );
AND2x2_ASAP7_75t_L g448 ( .A(n_204), .B(n_298), .Y(n_448) );
AND2x2_ASAP7_75t_L g459 ( .A(n_204), .B(n_233), .Y(n_459) );
AOI21x1_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B(n_213), .Y(n_209) );
INVx1_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx1_ASAP7_75t_SL g546 ( .A(n_214), .Y(n_546) );
INVx1_ASAP7_75t_L g567 ( .A(n_214), .Y(n_567) );
AND2x2_ASAP7_75t_L g317 ( .A(n_216), .B(n_231), .Y(n_317) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
OR2x2_ASAP7_75t_L g230 ( .A(n_217), .B(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g291 ( .A(n_217), .B(n_231), .Y(n_291) );
OR2x2_ASAP7_75t_L g305 ( .A(n_217), .B(n_244), .Y(n_305) );
AND2x2_ASAP7_75t_L g390 ( .A(n_217), .B(n_391), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_217), .B(n_244), .Y(n_401) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_217), .Y(n_443) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_221), .A2(n_523), .B(n_525), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g541 ( .A1(n_221), .A2(n_542), .B1(n_545), .B2(n_546), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_221), .A2(n_564), .B1(n_566), .B2(n_567), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g583 ( .A1(n_221), .A2(n_546), .B1(n_584), .B2(n_585), .Y(n_583) );
INVx1_ASAP7_75t_L g556 ( .A(n_223), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_225), .B(n_226), .Y(n_224) );
BUFx2_ASAP7_75t_L g547 ( .A(n_226), .Y(n_547) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_229), .B(n_232), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
INVx1_ASAP7_75t_L g339 ( .A(n_230), .Y(n_339) );
NAND3xp33_ASAP7_75t_L g446 ( .A(n_230), .B(n_447), .C(n_449), .Y(n_446) );
INVx1_ASAP7_75t_L g283 ( .A(n_231), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_232), .B(n_291), .Y(n_413) );
AND2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_244), .Y(n_232) );
INVx1_ASAP7_75t_L g256 ( .A(n_233), .Y(n_256) );
AND2x2_ASAP7_75t_L g462 ( .A(n_244), .B(n_298), .Y(n_462) );
INVx1_ASAP7_75t_L g465 ( .A(n_245), .Y(n_465) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
OR2x2_ASAP7_75t_L g444 ( .A(n_246), .B(n_277), .Y(n_444) );
OR2x2_ASAP7_75t_L g455 ( .A(n_246), .B(n_328), .Y(n_455) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g331 ( .A(n_247), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g479 ( .A(n_247), .B(n_257), .Y(n_479) );
AND2x2_ASAP7_75t_L g287 ( .A(n_248), .B(n_288), .Y(n_287) );
A2O1A1O1Ixp25_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_254), .B(n_271), .C(n_280), .D(n_284), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g365 ( .A(n_252), .B(n_366), .Y(n_365) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g302 ( .A(n_253), .Y(n_302) );
INVx1_ASAP7_75t_L g337 ( .A(n_254), .Y(n_337) );
AND2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_257), .Y(n_254) );
AND2x2_ASAP7_75t_L g316 ( .A(n_255), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
OR2x2_ASAP7_75t_L g307 ( .A(n_256), .B(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g336 ( .A(n_257), .Y(n_336) );
AND2x2_ASAP7_75t_L g407 ( .A(n_257), .B(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g453 ( .A(n_257), .B(n_287), .Y(n_453) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
INVx1_ASAP7_75t_L g278 ( .A(n_259), .Y(n_278) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_259), .Y(n_286) );
INVx2_ASAP7_75t_L g332 ( .A(n_259), .Y(n_332) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g308 ( .A(n_260), .Y(n_308) );
OAI21x1_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_262), .B(n_270), .Y(n_260) );
INVx1_ASAP7_75t_L g554 ( .A(n_268), .Y(n_554) );
INVx1_ASAP7_75t_L g403 ( .A(n_271), .Y(n_403) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_276), .Y(n_271) );
OAI21xp33_ASAP7_75t_L g327 ( .A1(n_272), .A2(n_277), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
AND2x2_ASAP7_75t_L g293 ( .A(n_273), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g398 ( .A(n_273), .B(n_348), .Y(n_398) );
INVx2_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AND2x2_ASAP7_75t_L g330 ( .A(n_274), .B(n_308), .Y(n_330) );
AND2x2_ASAP7_75t_L g354 ( .A(n_275), .B(n_279), .Y(n_354) );
NAND2xp5_ASAP7_75t_SL g438 ( .A(n_275), .B(n_294), .Y(n_438) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx1_ASAP7_75t_SL g382 ( .A(n_277), .Y(n_382) );
OR2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
INVx2_ASAP7_75t_L g294 ( .A(n_279), .Y(n_294) );
NAND2x1_ASAP7_75t_L g349 ( .A(n_279), .B(n_350), .Y(n_349) );
OAI32xp33_ASAP7_75t_L g470 ( .A1(n_280), .A2(n_346), .A3(n_454), .B1(n_471), .B2(n_472), .Y(n_470) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g344 ( .A(n_282), .Y(n_344) );
AND2x2_ASAP7_75t_L g367 ( .A(n_282), .B(n_325), .Y(n_367) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g364 ( .A(n_283), .B(n_298), .Y(n_364) );
OAI22xp33_ASAP7_75t_SL g284 ( .A1(n_285), .A2(n_289), .B1(n_292), .B2(n_295), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
AND2x2_ASAP7_75t_L g321 ( .A(n_287), .B(n_322), .Y(n_321) );
BUFx2_ASAP7_75t_L g340 ( .A(n_288), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
INVx2_ASAP7_75t_L g454 ( .A(n_290), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_291), .B(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g433 ( .A(n_291), .Y(n_433) );
AND2x2_ASAP7_75t_L g461 ( .A(n_291), .B(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x4_ASAP7_75t_L g368 ( .A(n_293), .B(n_369), .Y(n_368) );
O2A1O1Ixp33_ASAP7_75t_L g417 ( .A1(n_293), .A2(n_348), .B(n_418), .C(n_420), .Y(n_417) );
INVx1_ASAP7_75t_L g322 ( .A(n_294), .Y(n_322) );
AND2x2_ASAP7_75t_L g366 ( .A(n_294), .B(n_332), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_296), .B(n_317), .Y(n_335) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVxp67_ASAP7_75t_SL g313 ( .A(n_298), .Y(n_313) );
INVxp67_ASAP7_75t_SL g360 ( .A(n_298), .Y(n_360) );
INVx1_ASAP7_75t_L g389 ( .A(n_298), .Y(n_389) );
BUFx3_ASAP7_75t_L g402 ( .A(n_298), .Y(n_402) );
INVx3_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND3xp33_ASAP7_75t_L g300 ( .A(n_301), .B(n_303), .C(n_306), .Y(n_300) );
INVx1_ASAP7_75t_L g424 ( .A(n_301), .Y(n_424) );
OR2x2_ASAP7_75t_L g351 ( .A(n_302), .B(n_336), .Y(n_351) );
OR2x2_ASAP7_75t_L g315 ( .A(n_303), .B(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OAI22xp33_ASAP7_75t_L g341 ( .A1(n_304), .A2(n_342), .B1(n_346), .B2(n_351), .Y(n_341) );
INVx2_ASAP7_75t_L g345 ( .A(n_305), .Y(n_345) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_305), .Y(n_357) );
INVx1_ASAP7_75t_L g376 ( .A(n_305), .Y(n_376) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVxp67_ASAP7_75t_L g320 ( .A(n_308), .Y(n_320) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_308), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_318), .B1(n_323), .B2(n_326), .Y(n_309) );
NOR2x1_ASAP7_75t_L g310 ( .A(n_311), .B(n_315), .Y(n_310) );
BUFx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x4_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_317), .Y(n_395) );
NAND2x1p5_ASAP7_75t_L g318 ( .A(n_319), .B(n_321), .Y(n_318) );
INVx1_ASAP7_75t_L g386 ( .A(n_319), .Y(n_386) );
BUFx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AOI221x1_ASAP7_75t_L g372 ( .A1(n_321), .A2(n_373), .B1(n_377), .B2(n_379), .C(n_383), .Y(n_372) );
BUFx2_ASAP7_75t_L g475 ( .A(n_322), .Y(n_475) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_325), .B(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_325), .B(n_402), .Y(n_427) );
AND2x2_ASAP7_75t_L g481 ( .A(n_325), .B(n_360), .Y(n_481) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_329), .B(n_331), .Y(n_326) );
AOI211xp5_ASAP7_75t_L g463 ( .A1(n_328), .A2(n_464), .B(n_470), .C(n_473), .Y(n_463) );
OAI222xp33_ASAP7_75t_L g451 ( .A1(n_329), .A2(n_452), .B1(n_454), .B2(n_455), .C1(n_456), .C2(n_460), .Y(n_451) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
AO21x1_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_340), .B(n_341), .Y(n_333) );
OAI22xp5_ASAP7_75t_L g334 ( .A1(n_335), .A2(n_336), .B1(n_337), .B2(n_338), .Y(n_334) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g477 ( .A(n_340), .Y(n_477) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x4_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
AND2x2_ASAP7_75t_L g378 ( .A(n_345), .B(n_364), .Y(n_378) );
INVx1_ASAP7_75t_L g404 ( .A(n_345), .Y(n_404) );
OAI22xp5_ASAP7_75t_L g399 ( .A1(n_346), .A2(n_400), .B1(n_403), .B2(n_404), .Y(n_399) );
INVx1_ASAP7_75t_L g430 ( .A(n_346), .Y(n_430) );
OR2x6_ASAP7_75t_L g346 ( .A(n_347), .B(n_349), .Y(n_346) );
INVx1_ASAP7_75t_L g476 ( .A(n_347), .Y(n_476) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_SL g437 ( .A(n_350), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_350), .B(n_366), .Y(n_471) );
OAI21xp33_ASAP7_75t_SL g352 ( .A1(n_353), .A2(n_355), .B(n_361), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NOR3x1_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .C(n_359), .Y(n_356) );
BUFx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
AOI22xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_365), .B1(n_367), .B2(n_368), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_364), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g449 ( .A(n_364), .Y(n_449) );
INVx2_ASAP7_75t_L g423 ( .A(n_367), .Y(n_423) );
INVx3_ASAP7_75t_L g384 ( .A(n_368), .Y(n_384) );
NOR2x1_ASAP7_75t_L g370 ( .A(n_371), .B(n_428), .Y(n_370) );
NAND3xp33_ASAP7_75t_L g371 ( .A(n_372), .B(n_392), .C(n_417), .Y(n_371) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AOI21xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_385), .B(n_387), .Y(n_383) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
INVx1_ASAP7_75t_L g440 ( .A(n_389), .Y(n_440) );
BUFx2_ASAP7_75t_L g411 ( .A(n_391), .Y(n_411) );
AOI211xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_396), .B(n_399), .C(n_405), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AND2x4_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
OR2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_402), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_402), .B(n_469), .Y(n_468) );
OAI22xp33_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_409), .B1(n_413), .B2(n_414), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OR2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_412), .Y(n_409) );
AND2x2_ASAP7_75t_L g457 ( .A(n_410), .B(n_448), .Y(n_457) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g458 ( .A(n_411), .B(n_459), .Y(n_458) );
OR2x2_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_423), .B1(n_424), .B2(n_425), .Y(n_420) );
INVx3_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVxp67_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
NAND3xp33_ASAP7_75t_L g428 ( .A(n_429), .B(n_434), .C(n_463), .Y(n_428) );
OAI21xp33_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_431), .B(n_432), .Y(n_429) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_435), .B(n_451), .Y(n_434) );
OAI22xp33_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_439), .B1(n_444), .B2(n_445), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_438), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NOR2xp67_ASAP7_75t_L g445 ( .A(n_446), .B(n_450), .Y(n_445) );
INVx2_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NOR2xp33_ASAP7_75t_SL g456 ( .A(n_457), .B(n_458), .Y(n_456) );
INVx2_ASAP7_75t_L g472 ( .A(n_458), .Y(n_472) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
AOI21xp33_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_478), .B(n_480), .Y(n_473) );
NAND3x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .C(n_477), .Y(n_474) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVxp67_ASAP7_75t_SL g480 ( .A(n_481), .Y(n_480) );
INVx4_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
BUFx12f_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
CKINVDCx5p33_ASAP7_75t_R g486 ( .A(n_487), .Y(n_486) );
BUFx8_ASAP7_75t_SL g799 ( .A(n_487), .Y(n_799) );
AND2x2_ASAP7_75t_L g815 ( .A(n_487), .B(n_816), .Y(n_815) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx2_ASAP7_75t_L g848 ( .A(n_488), .Y(n_848) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_490), .B(n_493), .Y(n_489) );
NAND2xp5_ASAP7_75t_SL g818 ( .A(n_490), .B(n_809), .Y(n_818) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g819 ( .A(n_494), .B(n_820), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_495), .B(n_799), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_702), .Y(n_495) );
NAND4xp25_ASAP7_75t_L g496 ( .A(n_497), .B(n_626), .C(n_657), .D(n_686), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_498), .B(n_593), .Y(n_497) );
OAI322xp33_ASAP7_75t_L g498 ( .A1(n_499), .A2(n_537), .A3(n_560), .B1(n_571), .B2(n_579), .C1(n_588), .C2(n_590), .Y(n_498) );
INVxp67_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_500), .B(n_783), .Y(n_782) );
AND2x2_ASAP7_75t_L g500 ( .A(n_501), .B(n_513), .Y(n_500) );
AND2x2_ASAP7_75t_L g623 ( .A(n_501), .B(n_624), .Y(n_623) );
INVx4_ASAP7_75t_L g659 ( .A(n_501), .Y(n_659) );
INVx3_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AND2x2_ASAP7_75t_L g634 ( .A(n_502), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g637 ( .A(n_502), .B(n_539), .Y(n_637) );
AND2x2_ASAP7_75t_L g654 ( .A(n_502), .B(n_551), .Y(n_654) );
AND2x2_ASAP7_75t_L g752 ( .A(n_502), .B(n_753), .Y(n_752) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx2_ASAP7_75t_L g575 ( .A(n_503), .Y(n_575) );
AND2x4_ASAP7_75t_L g758 ( .A(n_503), .B(n_753), .Y(n_758) );
AO31x2_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_505), .A3(n_510), .B(n_511), .Y(n_503) );
AO31x2_ASAP7_75t_L g582 ( .A1(n_504), .A2(n_547), .A3(n_583), .B(n_586), .Y(n_582) );
AO31x2_ASAP7_75t_L g601 ( .A1(n_510), .A2(n_568), .A3(n_602), .B(n_605), .Y(n_601) );
AND2x4_ASAP7_75t_L g763 ( .A(n_513), .B(n_664), .Y(n_763) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g592 ( .A(n_514), .Y(n_592) );
INVxp67_ASAP7_75t_SL g750 ( .A(n_514), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_515), .B(n_529), .Y(n_514) );
AND2x2_ASAP7_75t_L g580 ( .A(n_515), .B(n_530), .Y(n_580) );
INVx1_ASAP7_75t_L g621 ( .A(n_515), .Y(n_621) );
OAI21x1_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_517), .B(n_528), .Y(n_515) );
OAI21x1_ASAP7_75t_L g616 ( .A1(n_516), .A2(n_517), .B(n_528), .Y(n_616) );
OAI21x1_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_522), .B(n_526), .Y(n_517) );
INVx2_ASAP7_75t_SL g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_SL g568 ( .A(n_527), .Y(n_568) );
INVx2_ASAP7_75t_L g612 ( .A(n_529), .Y(n_612) );
AND2x2_ASAP7_75t_L g676 ( .A(n_529), .B(n_615), .Y(n_676) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g630 ( .A(n_530), .Y(n_630) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_530), .Y(n_683) );
OR2x2_ASAP7_75t_L g754 ( .A(n_530), .B(n_562), .Y(n_754) );
NAND4xp25_ASAP7_75t_L g632 ( .A(n_537), .B(n_633), .C(n_636), .D(n_638), .Y(n_632) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_L g770 ( .A(n_538), .B(n_758), .Y(n_770) );
AND2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_550), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_539), .B(n_599), .Y(n_598) );
AND2x4_ASAP7_75t_L g624 ( .A(n_539), .B(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g644 ( .A(n_539), .Y(n_644) );
INVx1_ASAP7_75t_L g661 ( .A(n_539), .Y(n_661) );
INVx1_ASAP7_75t_L g669 ( .A(n_539), .Y(n_669) );
HB1xp67_ASAP7_75t_L g783 ( .A(n_539), .Y(n_783) );
INVx4_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_540), .B(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g701 ( .A(n_540), .B(n_601), .Y(n_701) );
AND2x2_ASAP7_75t_L g709 ( .A(n_540), .B(n_551), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_540), .B(n_732), .Y(n_731) );
BUFx2_ASAP7_75t_L g774 ( .A(n_540), .Y(n_774) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g578 ( .A(n_551), .Y(n_578) );
OR2x2_ASAP7_75t_L g639 ( .A(n_551), .B(n_601), .Y(n_639) );
INVx2_ASAP7_75t_L g646 ( .A(n_551), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_551), .B(n_599), .Y(n_670) );
HB1xp67_ASAP7_75t_L g757 ( .A(n_551), .Y(n_757) );
AO31x2_ASAP7_75t_L g562 ( .A1(n_557), .A2(n_563), .A3(n_568), .B(n_569), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g728 ( .A(n_560), .B(n_729), .Y(n_728) );
BUFx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g581 ( .A(n_562), .B(n_582), .Y(n_581) );
BUFx2_ASAP7_75t_L g591 ( .A(n_562), .Y(n_591) );
INVx2_ASAP7_75t_L g609 ( .A(n_562), .Y(n_609) );
AND2x4_ASAP7_75t_L g641 ( .A(n_562), .B(n_613), .Y(n_641) );
OR2x2_ASAP7_75t_L g721 ( .A(n_562), .B(n_621), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_576), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_573), .B(n_589), .Y(n_588) );
OR2x2_ASAP7_75t_L g638 ( .A(n_573), .B(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_573), .B(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_574), .B(n_644), .Y(n_652) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx2_ASAP7_75t_L g597 ( .A(n_575), .Y(n_597) );
OR2x2_ASAP7_75t_L g690 ( .A(n_575), .B(n_600), .Y(n_690) );
INVx1_ASAP7_75t_L g617 ( .A(n_576), .Y(n_617) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g589 ( .A(n_577), .Y(n_589) );
INVx1_ASAP7_75t_L g625 ( .A(n_578), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
OAI322xp33_ASAP7_75t_L g593 ( .A1(n_580), .A2(n_594), .A3(n_607), .B1(n_610), .B2(n_617), .C1(n_618), .C2(n_622), .Y(n_593) );
AND2x4_ASAP7_75t_L g640 ( .A(n_580), .B(n_641), .Y(n_640) );
AOI211xp5_ASAP7_75t_SL g671 ( .A1(n_580), .A2(n_672), .B(n_673), .C(n_677), .Y(n_671) );
AND2x2_ASAP7_75t_L g691 ( .A(n_580), .B(n_581), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_580), .B(n_608), .Y(n_697) );
AND2x4_ASAP7_75t_SL g619 ( .A(n_581), .B(n_620), .Y(n_619) );
NAND3xp33_ASAP7_75t_L g710 ( .A(n_581), .B(n_637), .C(n_665), .Y(n_710) );
AND2x2_ASAP7_75t_L g741 ( .A(n_581), .B(n_742), .Y(n_741) );
AND2x2_ASAP7_75t_L g608 ( .A(n_582), .B(n_609), .Y(n_608) );
INVx3_ASAP7_75t_L g613 ( .A(n_582), .Y(n_613) );
BUFx2_ASAP7_75t_L g681 ( .A(n_582), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_591), .B(n_615), .Y(n_614) );
NAND2x1_ASAP7_75t_L g655 ( .A(n_591), .B(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g674 ( .A(n_591), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_592), .B(n_608), .Y(n_739) );
OR2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_598), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx3_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g682 ( .A(n_597), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_601), .Y(n_635) );
AND2x4_ASAP7_75t_L g645 ( .A(n_601), .B(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g732 ( .A(n_601), .Y(n_732) );
INVx2_ASAP7_75t_L g753 ( .A(n_601), .Y(n_753) );
OAI22xp33_ASAP7_75t_L g765 ( .A1(n_607), .A2(n_766), .B1(n_768), .B2(n_769), .Y(n_765) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AND2x2_ASAP7_75t_L g677 ( .A(n_608), .B(n_678), .Y(n_677) );
AND2x4_ASAP7_75t_L g631 ( .A(n_609), .B(n_615), .Y(n_631) );
OR2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_614), .Y(n_610) );
INVx1_ASAP7_75t_L g650 ( .A(n_611), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
AND2x4_ASAP7_75t_L g620 ( .A(n_612), .B(n_621), .Y(n_620) );
INVx1_ASAP7_75t_L g742 ( .A(n_612), .Y(n_742) );
INVx2_ASAP7_75t_L g628 ( .A(n_613), .Y(n_628) );
AND2x2_ASAP7_75t_L g656 ( .A(n_613), .B(n_615), .Y(n_656) );
INVx3_ASAP7_75t_L g664 ( .A(n_613), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_613), .B(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g649 ( .A(n_614), .Y(n_649) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
BUFx2_ASAP7_75t_L g665 ( .A(n_616), .Y(n_665) );
OAI222xp33_ASAP7_75t_L g788 ( .A1(n_618), .A2(n_778), .B1(n_789), .B2(n_792), .C1(n_794), .C2(n_796), .Y(n_788) );
INVx3_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g729 ( .A(n_620), .Y(n_729) );
AND2x2_ASAP7_75t_L g793 ( .A(n_620), .B(n_663), .Y(n_793) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_623), .B(n_714), .Y(n_713) );
AOI221xp5_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_632), .B1(n_640), .B2(n_642), .C(n_647), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_628), .B(n_629), .Y(n_627) );
INVx1_ASAP7_75t_L g715 ( .A(n_628), .Y(n_715) );
INVx2_ASAP7_75t_L g777 ( .A(n_629), .Y(n_777) );
AND2x4_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
INVx2_ASAP7_75t_L g678 ( .A(n_630), .Y(n_678) );
AND2x2_ASAP7_75t_L g714 ( .A(n_630), .B(n_715), .Y(n_714) );
AND2x4_ASAP7_75t_L g680 ( .A(n_631), .B(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g706 ( .A(n_631), .B(n_707), .Y(n_706) );
INVx1_ASAP7_75t_L g795 ( .A(n_631), .Y(n_795) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g744 ( .A(n_635), .Y(n_744) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g767 ( .A(n_637), .B(n_645), .Y(n_767) );
AND2x2_ASAP7_75t_L g790 ( .A(n_637), .B(n_791), .Y(n_790) );
OR2x2_ASAP7_75t_L g651 ( .A(n_639), .B(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g786 ( .A(n_639), .Y(n_786) );
AOI22xp5_ASAP7_75t_L g727 ( .A1(n_640), .A2(n_694), .B1(n_728), .B2(n_730), .Y(n_727) );
OAI21xp5_ASAP7_75t_L g755 ( .A1(n_640), .A2(n_756), .B(n_759), .Y(n_755) );
INVxp67_ASAP7_75t_L g672 ( .A(n_641), .Y(n_672) );
INVx2_ASAP7_75t_SL g776 ( .A(n_641), .Y(n_776) );
AND2x4_ASAP7_75t_L g642 ( .A(n_643), .B(n_645), .Y(n_642) );
OR2x2_ASAP7_75t_L g689 ( .A(n_643), .B(n_690), .Y(n_689) );
AND2x2_ASAP7_75t_L g787 ( .A(n_643), .B(n_786), .Y(n_787) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g660 ( .A(n_645), .B(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_645), .B(n_669), .Y(n_685) );
INVx2_ASAP7_75t_L g712 ( .A(n_645), .Y(n_712) );
OAI22xp33_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_651), .B1(n_653), .B2(n_655), .Y(n_647) );
NOR2xp33_ASAP7_75t_SL g648 ( .A(n_649), .B(n_650), .Y(n_648) );
AOI22xp5_ASAP7_75t_L g735 ( .A1(n_649), .A2(n_723), .B1(n_736), .B2(n_738), .Y(n_735) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g745 ( .A(n_654), .B(n_746), .Y(n_745) );
AOI21xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_662), .B(n_666), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
INVx1_ASAP7_75t_L g726 ( .A(n_659), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_659), .B(n_709), .Y(n_737) );
INVx1_ASAP7_75t_L g695 ( .A(n_661), .Y(n_695) );
AND2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_665), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_663), .B(n_676), .Y(n_768) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
OAI21xp33_ASAP7_75t_L g781 ( .A1(n_664), .A2(n_782), .B(n_784), .Y(n_781) );
OAI21xp5_ASAP7_75t_SL g666 ( .A1(n_667), .A2(n_671), .B(n_679), .Y(n_666) );
BUFx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
OR2x2_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
INVx1_ASAP7_75t_L g725 ( .A(n_670), .Y(n_725) );
INVx1_ASAP7_75t_L g791 ( .A(n_670), .Y(n_791) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
INVx1_ASAP7_75t_L g764 ( .A(n_674), .Y(n_764) );
OR2x2_ASAP7_75t_L g775 ( .A(n_675), .B(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
NAND3xp33_ASAP7_75t_L g679 ( .A(n_680), .B(n_682), .C(n_684), .Y(n_679) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_680), .A2(n_741), .B1(n_743), .B2(n_745), .Y(n_740) );
INVx1_ASAP7_75t_L g707 ( .A(n_681), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_682), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g720 ( .A(n_683), .Y(n_720) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_685), .B(n_689), .Y(n_688) );
OAI221xp5_ASAP7_75t_L g747 ( .A1(n_685), .A2(n_748), .B1(n_751), .B2(n_754), .C(n_755), .Y(n_747) );
AOI21xp5_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_691), .B(n_692), .Y(n_686) );
HB1xp67_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx2_ASAP7_75t_L g696 ( .A(n_690), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_697), .B1(n_698), .B2(n_856), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AND2x4_ASAP7_75t_L g694 ( .A(n_695), .B(n_696), .Y(n_694) );
INVxp67_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx2_ASAP7_75t_SL g699 ( .A(n_700), .Y(n_699) );
AND2x4_ASAP7_75t_L g779 ( .A(n_701), .B(n_757), .Y(n_779) );
NAND4xp25_ASAP7_75t_L g702 ( .A(n_703), .B(n_733), .C(n_760), .D(n_780), .Y(n_702) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_704), .B(n_716), .Y(n_703) );
OAI221xp5_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_708), .B1(n_710), .B2(n_711), .C(n_713), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_706), .A2(n_763), .B1(n_785), .B2(n_787), .Y(n_784) );
INVx1_ASAP7_75t_L g759 ( .A(n_708), .Y(n_759) );
INVx2_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
AND2x2_ASAP7_75t_L g743 ( .A(n_709), .B(n_744), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_709), .B(n_752), .Y(n_751) );
NAND2x1_ASAP7_75t_L g796 ( .A(n_709), .B(n_797), .Y(n_796) );
NOR2xp33_ASAP7_75t_L g772 ( .A(n_711), .B(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g718 ( .A(n_715), .B(n_719), .Y(n_718) );
OAI21xp33_ASAP7_75t_SL g716 ( .A1(n_717), .A2(n_722), .B(n_727), .Y(n_716) );
INVx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
NOR2x1_ASAP7_75t_L g719 ( .A(n_720), .B(n_721), .Y(n_719) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g746 ( .A(n_732), .Y(n_746) );
AOI211xp5_ASAP7_75t_L g760 ( .A1(n_732), .A2(n_761), .B(n_765), .C(n_771), .Y(n_760) );
NOR2xp33_ASAP7_75t_L g733 ( .A(n_734), .B(n_747), .Y(n_733) );
NAND2xp5_ASAP7_75t_SL g734 ( .A(n_735), .B(n_740), .Y(n_734) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
OR2x2_ASAP7_75t_L g794 ( .A(n_742), .B(n_795), .Y(n_794) );
HB1xp67_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
AND2x4_ASAP7_75t_L g756 ( .A(n_757), .B(n_758), .Y(n_756) );
INVx3_ASAP7_75t_L g798 ( .A(n_758), .Y(n_798) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
NAND2x1p5_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .Y(n_762) );
INVx2_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
OAI22xp33_ASAP7_75t_R g771 ( .A1(n_772), .A2(n_775), .B1(n_777), .B2(n_778), .Y(n_771) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
AND2x4_ASAP7_75t_L g785 ( .A(n_774), .B(n_786), .Y(n_785) );
INVx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
NOR2xp33_ASAP7_75t_L g780 ( .A(n_781), .B(n_788), .Y(n_780) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx2_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx6_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
AND2x6_ASAP7_75t_SL g801 ( .A(n_802), .B(n_804), .Y(n_801) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
NOR2xp33_ASAP7_75t_L g813 ( .A(n_803), .B(n_814), .Y(n_813) );
INVx3_ASAP7_75t_L g823 ( .A(n_803), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_805), .B(n_807), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
NOR2x1_ASAP7_75t_L g816 ( .A(n_806), .B(n_808), .Y(n_816) );
NOR3x1_ASAP7_75t_L g844 ( .A(n_806), .B(n_845), .C(n_848), .Y(n_844) );
AND2x6_ASAP7_75t_SL g827 ( .A(n_807), .B(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
INVx3_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx6_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
BUFx10_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
NOR2xp67_ASAP7_75t_L g817 ( .A(n_818), .B(n_819), .Y(n_817) );
OA21x2_ASAP7_75t_L g821 ( .A1(n_822), .A2(n_824), .B(n_837), .Y(n_821) );
BUFx6f_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
AND2x2_ASAP7_75t_L g825 ( .A(n_826), .B(n_831), .Y(n_825) );
CKINVDCx5p33_ASAP7_75t_R g826 ( .A(n_827), .Y(n_826) );
INVx5_ASAP7_75t_L g840 ( .A(n_827), .Y(n_840) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g836 ( .A(n_833), .Y(n_836) );
INVxp67_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
NOR2xp67_ASAP7_75t_SL g838 ( .A(n_839), .B(n_841), .Y(n_838) );
BUFx3_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
BUFx2_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
AND2x4_ASAP7_75t_L g843 ( .A(n_844), .B(n_849), .Y(n_843) );
AND2x2_ASAP7_75t_SL g854 ( .A(n_844), .B(n_849), .Y(n_854) );
INVx2_ASAP7_75t_SL g845 ( .A(n_846), .Y(n_845) );
NOR2x1p5_ASAP7_75t_L g849 ( .A(n_850), .B(n_851), .Y(n_849) );
INVx1_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
INVx6_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
endmodule