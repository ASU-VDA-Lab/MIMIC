module fake_jpeg_18355_n_109 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_109);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_109;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_31),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_54),
.Y(n_71)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_55),
.B(n_56),
.Y(n_62)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_57),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_44),
.B(n_0),
.Y(n_58)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_1),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_59),
.A2(n_42),
.B1(n_39),
.B2(n_38),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_53),
.A2(n_41),
.B1(n_48),
.B2(n_47),
.Y(n_61)
);

OAI22x1_ASAP7_75t_L g83 ( 
.A1(n_61),
.A2(n_63),
.B1(n_66),
.B2(n_18),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_54),
.A2(n_49),
.B1(n_45),
.B2(n_43),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_16),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_52),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_59),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_L g77 ( 
.A1(n_68),
.A2(n_37),
.B1(n_11),
.B2(n_12),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_7),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_77),
.Y(n_86)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_73),
.Y(n_87)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_71),
.Y(n_76)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_9),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_79),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_14),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

OA22x2_ASAP7_75t_SL g88 ( 
.A1(n_82),
.A2(n_83),
.B1(n_19),
.B2(n_20),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_79),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_92),
.A2(n_94),
.B1(n_96),
.B2(n_95),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_84),
.B(n_72),
.Y(n_93)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_93),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_89),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_74),
.C(n_25),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_95),
.B(n_91),
.Y(n_97)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_97),
.B(n_98),
.Y(n_101)
);

OAI322xp33_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_88),
.A3(n_90),
.B1(n_28),
.B2(n_29),
.C1(n_30),
.C2(n_32),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_100),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_101),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_87),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_105),
.Y(n_106)
);

OAI21x1_ASAP7_75t_L g107 ( 
.A1(n_106),
.A2(n_23),
.B(n_26),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_107),
.B(n_33),
.C(n_35),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_108),
.B(n_36),
.Y(n_109)
);


endmodule