module fake_jpeg_21591_n_103 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_103);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_103;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

AND2x2_ASAP7_75t_L g12 ( 
.A(n_7),
.B(n_1),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

OR2x2_ASAP7_75t_L g14 ( 
.A(n_6),
.B(n_11),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx4f_ASAP7_75t_SL g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx9p33_ASAP7_75t_R g24 ( 
.A(n_19),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_12),
.B(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_27),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_12),
.B(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_20),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_31),
.Y(n_34)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_22),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_30),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_22),
.A2(n_2),
.B1(n_5),
.B2(n_7),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_19),
.Y(n_35)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_14),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_42),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_14),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_26),
.B(n_12),
.Y(n_43)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_29),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_44),
.A2(n_45),
.B1(n_25),
.B2(n_40),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_17),
.B(n_20),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_33),
.B(n_18),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_47),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_33),
.B(n_18),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_13),
.Y(n_48)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_28),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_50),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_28),
.Y(n_50)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_60),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_37),
.A2(n_30),
.B1(n_31),
.B2(n_28),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_52),
.A2(n_32),
.B1(n_21),
.B2(n_13),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_38),
.A2(n_29),
.B1(n_25),
.B2(n_32),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g59 ( 
.A1(n_36),
.A2(n_25),
.B1(n_32),
.B2(n_17),
.Y(n_59)
);

OA21x2_ASAP7_75t_L g71 ( 
.A1(n_59),
.A2(n_50),
.B(n_49),
.Y(n_71)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_61),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_69),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_68),
.A2(n_71),
.B1(n_44),
.B2(n_59),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_56),
.B(n_19),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_23),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_72),
.B(n_59),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_44),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_64),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_70),
.B(n_55),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_75),
.B(n_76),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_65),
.Y(n_77)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_77),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_63),
.B(n_53),
.Y(n_78)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_71),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_80),
.A2(n_81),
.B1(n_71),
.B2(n_72),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_81),
.Y(n_90)
);

MAJx2_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_69),
.C(n_67),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_85),
.A2(n_76),
.B(n_62),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_79),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_88),
.B(n_89),
.C(n_91),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_90),
.A2(n_83),
.B1(n_62),
.B2(n_82),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_86),
.B(n_77),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_57),
.C(n_59),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_92),
.A2(n_2),
.B(n_21),
.Y(n_96)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_94),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_89),
.A2(n_85),
.B1(n_73),
.B2(n_57),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_95),
.A2(n_40),
.B1(n_60),
.B2(n_16),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_23),
.C(n_16),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_97),
.A2(n_98),
.B(n_51),
.Y(n_101)
);

O2A1O1Ixp33_ASAP7_75t_SL g100 ( 
.A1(n_99),
.A2(n_95),
.B(n_93),
.C(n_15),
.Y(n_100)
);

AOI322xp5_ASAP7_75t_L g102 ( 
.A1(n_100),
.A2(n_101),
.A3(n_40),
.B1(n_61),
.B2(n_15),
.C1(n_8),
.C2(n_10),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_102),
.B(n_8),
.Y(n_103)
);


endmodule