module fake_jpeg_31230_n_36 (n_3, n_2, n_1, n_0, n_4, n_5, n_36);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_36;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

OR2x2_ASAP7_75t_SL g6 ( 
.A(n_5),
.B(n_4),
.Y(n_6)
);

INVx8_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_SL g8 ( 
.A(n_4),
.B(n_2),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx1_ASAP7_75t_SL g10 ( 
.A(n_1),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_L g13 ( 
.A1(n_12),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_13)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_13),
.A2(n_11),
.B1(n_9),
.B2(n_6),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g14 ( 
.A(n_10),
.B(n_0),
.Y(n_14)
);

MAJx2_ASAP7_75t_L g25 ( 
.A(n_14),
.B(n_18),
.C(n_6),
.Y(n_25)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

NAND2xp33_ASAP7_75t_SL g21 ( 
.A(n_15),
.B(n_17),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_8),
.B(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx6p67_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_10),
.B(n_2),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_8),
.B(n_11),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

HB1xp67_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_14),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_26),
.A2(n_14),
.B1(n_18),
.B2(n_19),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_27),
.A2(n_28),
.B1(n_29),
.B2(n_23),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_22),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_30),
.A2(n_23),
.B(n_17),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_31),
.A2(n_13),
.B1(n_25),
.B2(n_17),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_32),
.B(n_33),
.Y(n_34)
);

AOI332xp33_ASAP7_75t_SL g35 ( 
.A1(n_34),
.A2(n_17),
.A3(n_6),
.B1(n_21),
.B2(n_20),
.B3(n_15),
.C1(n_7),
.C2(n_24),
.Y(n_35)
);

AOI221xp5_ASAP7_75t_L g36 ( 
.A1(n_35),
.A2(n_7),
.B1(n_9),
.B2(n_15),
.C(n_33),
.Y(n_36)
);


endmodule