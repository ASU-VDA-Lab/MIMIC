module fake_jpeg_10516_n_105 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_105);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_105;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_27),
.Y(n_30)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_30),
.B(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_32),
.Y(n_41)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_35),
.Y(n_43)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_0),
.C(n_1),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_39),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_14),
.B(n_16),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_14),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_19),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_46),
.Y(n_66)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_47),
.B(n_51),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_40),
.B(n_17),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_52),
.B(n_47),
.Y(n_57)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_36),
.A2(n_21),
.B1(n_19),
.B2(n_20),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_55),
.A2(n_21),
.B1(n_20),
.B2(n_18),
.Y(n_62)
);

AND2x6_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_1),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_SL g74 ( 
.A(n_56),
.B(n_69),
.C(n_73),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_59),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_35),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_50),
.B(n_35),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_55),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_65),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_62),
.A2(n_64),
.B1(n_68),
.B2(n_71),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_42),
.A2(n_39),
.B1(n_30),
.B2(n_31),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_27),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_72),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_42),
.A2(n_39),
.B1(n_28),
.B2(n_26),
.Y(n_68)
);

AND2x6_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_2),
.Y(n_69)
);

INVx6_ASAP7_75t_SL g70 ( 
.A(n_45),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_70),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_46),
.A2(n_28),
.B1(n_26),
.B2(n_24),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_49),
.A2(n_28),
.B1(n_26),
.B2(n_24),
.Y(n_72)
);

NOR2x1_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_29),
.Y(n_73)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_78),
.B(n_79),
.Y(n_82)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_83),
.B(n_85),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_74),
.A2(n_75),
.B(n_58),
.C(n_76),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_84),
.B(n_86),
.Y(n_90)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_78),
.B(n_60),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

AO21x1_ASAP7_75t_L g91 ( 
.A1(n_87),
.A2(n_48),
.B(n_63),
.Y(n_91)
);

OA21x2_ASAP7_75t_L g89 ( 
.A1(n_85),
.A2(n_81),
.B(n_72),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_89),
.A2(n_91),
.B1(n_82),
.B2(n_83),
.Y(n_95)
);

NAND2x1p5_ASAP7_75t_R g92 ( 
.A(n_87),
.B(n_48),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_93),
.B(n_94),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_92),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_96),
.Y(n_98)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_100),
.Y(n_101)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_98),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_13),
.B(n_5),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_4),
.C(n_6),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_4),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_4),
.Y(n_105)
);


endmodule