module fake_jpeg_2175_n_404 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_404);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_404;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_14),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_40),
.Y(n_44)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_44),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_24),
.B(n_0),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_45),
.B(n_60),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_46),
.Y(n_106)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_17),
.Y(n_47)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_47),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_24),
.B(n_15),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_48),
.B(n_71),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_49),
.Y(n_131)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_51),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_52),
.Y(n_107)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_54),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_56),
.Y(n_133)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_57),
.Y(n_123)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_59),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_15),
.B(n_0),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_62),
.B(n_70),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_63),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_64),
.Y(n_110)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_66),
.Y(n_134)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_67),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_68),
.Y(n_135)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_69),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_26),
.B(n_1),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_72),
.B(n_74),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_73),
.B(n_75),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_26),
.B(n_31),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_38),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_76),
.B(n_77),
.Y(n_130)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

AOI21xp33_ASAP7_75t_L g78 ( 
.A1(n_30),
.A2(n_1),
.B(n_2),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_78),
.B(n_84),
.Y(n_87)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_79),
.A2(n_43),
.B1(n_20),
.B2(n_22),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_81),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_85),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_86),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_33),
.B(n_2),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

CKINVDCx5p33_ASAP7_75t_R g86 ( 
.A(n_28),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_69),
.A2(n_37),
.B1(n_43),
.B2(n_28),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_89),
.A2(n_94),
.B1(n_128),
.B2(n_65),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_91),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_55),
.A2(n_39),
.B1(n_32),
.B2(n_31),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_58),
.A2(n_25),
.B1(n_20),
.B2(n_22),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_96),
.A2(n_97),
.B1(n_101),
.B2(n_109),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_50),
.A2(n_25),
.B1(n_20),
.B2(n_22),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_56),
.A2(n_16),
.B1(n_39),
.B2(n_32),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_98),
.A2(n_108),
.B1(n_114),
.B2(n_132),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_67),
.A2(n_42),
.B(n_35),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_99),
.A2(n_104),
.B(n_100),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_44),
.A2(n_25),
.B1(n_23),
.B2(n_42),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_79),
.A2(n_35),
.B1(n_27),
.B2(n_16),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_61),
.A2(n_37),
.B1(n_27),
.B2(n_23),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_51),
.A2(n_23),
.B1(n_17),
.B2(n_21),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_64),
.B(n_37),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_111),
.B(n_120),
.Y(n_176)
);

OAI22xp33_ASAP7_75t_L g114 ( 
.A1(n_66),
.A2(n_17),
.B1(n_21),
.B2(n_5),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_68),
.B(n_2),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_70),
.A2(n_21),
.B1(n_4),
.B2(n_6),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_122),
.A2(n_127),
.B1(n_46),
.B2(n_63),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_70),
.A2(n_2),
.B1(n_6),
.B2(n_8),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_71),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_73),
.A2(n_83),
.B1(n_81),
.B2(n_80),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_108),
.A2(n_99),
.B1(n_120),
.B2(n_111),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_137),
.A2(n_146),
.B1(n_161),
.B2(n_104),
.Y(n_192)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_136),
.Y(n_138)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_138),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_105),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_139),
.B(n_144),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_117),
.B(n_49),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_140),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_49),
.Y(n_141)
);

AND2x2_ASAP7_75t_SL g223 ( 
.A(n_141),
.B(n_156),
.Y(n_223)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_136),
.Y(n_142)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_142),
.Y(n_194)
);

INVx3_ASAP7_75t_SL g143 ( 
.A(n_126),
.Y(n_143)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_143),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_121),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_135),
.A2(n_75),
.B1(n_92),
.B2(n_100),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_135),
.Y(n_148)
);

BUFx2_ASAP7_75t_SL g188 ( 
.A(n_148),
.Y(n_188)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_149),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_93),
.Y(n_150)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_150),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_116),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_151),
.B(n_152),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_90),
.Y(n_152)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_119),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_153),
.B(n_158),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_L g155 ( 
.A1(n_88),
.A2(n_65),
.B1(n_46),
.B2(n_52),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_155),
.A2(n_165),
.B1(n_170),
.B2(n_106),
.Y(n_208)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_90),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_156),
.B(n_163),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_157),
.A2(n_128),
.B1(n_89),
.B2(n_114),
.Y(n_190)
);

NAND3xp33_ASAP7_75t_L g158 ( 
.A(n_87),
.B(n_102),
.C(n_130),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g159 ( 
.A(n_119),
.Y(n_159)
);

INVx13_ASAP7_75t_L g196 ( 
.A(n_159),
.Y(n_196)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_112),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_160),
.B(n_162),
.Y(n_202)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_112),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_90),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_164),
.B(n_166),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_87),
.A2(n_63),
.B1(n_54),
.B2(n_52),
.Y(n_165)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_113),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_103),
.B(n_54),
.C(n_10),
.Y(n_167)
);

MAJx2_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_133),
.C(n_93),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g168 ( 
.A(n_107),
.B(n_129),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_168),
.B(n_172),
.Y(n_184)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_110),
.Y(n_169)
);

INVx13_ASAP7_75t_L g222 ( 
.A(n_169),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_88),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_103),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_171),
.B(n_178),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_107),
.B(n_10),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_113),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_173),
.B(n_175),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_123),
.B(n_11),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_174),
.B(n_177),
.Y(n_203)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_115),
.Y(n_175)
);

AOI21xp33_ASAP7_75t_L g177 ( 
.A1(n_123),
.A2(n_12),
.B(n_13),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_124),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_129),
.B(n_124),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_179),
.B(n_12),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_115),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_180),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_125),
.B(n_12),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_181),
.B(n_182),
.Y(n_210)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_125),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_134),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_183),
.B(n_118),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_176),
.B(n_139),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_185),
.B(n_214),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_187),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_190),
.A2(n_217),
.B1(n_153),
.B2(n_169),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_192),
.A2(n_200),
.B1(n_205),
.B2(n_206),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_145),
.A2(n_95),
.B1(n_93),
.B2(n_133),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_197),
.A2(n_220),
.B1(n_205),
.B2(n_215),
.Y(n_251)
);

AOI21xp33_ASAP7_75t_L g198 ( 
.A1(n_164),
.A2(n_106),
.B(n_131),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_198),
.A2(n_212),
.B(n_204),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_199),
.B(n_175),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_176),
.A2(n_161),
.B1(n_147),
.B2(n_154),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_147),
.A2(n_126),
.B1(n_133),
.B2(n_110),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_144),
.A2(n_141),
.B1(n_155),
.B2(n_148),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_208),
.Y(n_230)
);

AND2x6_ASAP7_75t_L g211 ( 
.A(n_141),
.B(n_131),
.Y(n_211)
);

A2O1A1O1Ixp25_ASAP7_75t_L g228 ( 
.A1(n_211),
.A2(n_163),
.B(n_149),
.C(n_183),
.D(n_159),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_179),
.A2(n_95),
.B(n_13),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_138),
.B(n_110),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_223),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_143),
.A2(n_110),
.B1(n_12),
.B2(n_13),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_172),
.A2(n_173),
.B1(n_168),
.B2(n_166),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_218),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g220 ( 
.A1(n_142),
.A2(n_152),
.B1(n_178),
.B2(n_171),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_167),
.B(n_182),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_224),
.B(n_223),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_201),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_227),
.B(n_252),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_228),
.A2(n_241),
.B(n_256),
.Y(n_267)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_213),
.Y(n_229)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_229),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_185),
.B(n_180),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_231),
.B(n_234),
.C(n_243),
.Y(n_290)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_213),
.Y(n_232)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_232),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_204),
.A2(n_143),
.B1(n_150),
.B2(n_160),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_233),
.A2(n_245),
.B1(n_253),
.B2(n_259),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_162),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_235),
.B(n_201),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_236),
.A2(n_219),
.B1(n_196),
.B2(n_193),
.Y(n_277)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_188),
.Y(n_238)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_238),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_239),
.B(n_254),
.Y(n_283)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_188),
.Y(n_242)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_242),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_199),
.B(n_187),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_243),
.B(n_235),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_207),
.B(n_186),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_244),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_200),
.A2(n_190),
.B1(n_208),
.B2(n_211),
.Y(n_245)
);

OA21x2_ASAP7_75t_L g247 ( 
.A1(n_206),
.A2(n_211),
.B(n_212),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_247),
.A2(n_257),
.B(n_258),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_186),
.B(n_184),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_248),
.B(n_250),
.Y(n_260)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_194),
.Y(n_249)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_249),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_184),
.B(n_210),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_251),
.A2(n_233),
.B1(n_238),
.B2(n_242),
.Y(n_287)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_221),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_218),
.A2(n_203),
.B1(n_198),
.B2(n_199),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_221),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_221),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_255),
.B(n_254),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_203),
.A2(n_195),
.B1(n_210),
.B2(n_216),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_209),
.A2(n_191),
.B(n_195),
.Y(n_257)
);

O2A1O1Ixp33_ASAP7_75t_L g258 ( 
.A1(n_214),
.A2(n_223),
.B(n_209),
.C(n_194),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_223),
.A2(n_191),
.B1(n_202),
.B2(n_221),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_261),
.B(n_268),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_225),
.B(n_202),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_262),
.B(n_265),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_225),
.B(n_201),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_246),
.A2(n_217),
.B1(n_215),
.B2(n_201),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_266),
.A2(n_278),
.B1(n_287),
.B2(n_236),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_226),
.B(n_189),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_270),
.B(n_272),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_226),
.B(n_189),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_241),
.A2(n_196),
.B(n_222),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_273),
.A2(n_288),
.B(n_269),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_247),
.B(n_193),
.Y(n_275)
);

NAND2x1_ASAP7_75t_SL g294 ( 
.A(n_275),
.B(n_277),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_227),
.B(n_193),
.Y(n_276)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_276),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_230),
.A2(n_219),
.B1(n_222),
.B2(n_196),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_252),
.B(n_219),
.Y(n_280)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_280),
.Y(n_299)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_237),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_281),
.B(n_237),
.Y(n_296)
);

OA21x2_ASAP7_75t_L g282 ( 
.A1(n_245),
.A2(n_222),
.B(n_253),
.Y(n_282)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_282),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_285),
.B(n_240),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_246),
.A2(n_247),
.B(n_258),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_290),
.B(n_272),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_290),
.B(n_234),
.C(n_239),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_291),
.B(n_292),
.C(n_302),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_290),
.B(n_231),
.C(n_259),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_289),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_293),
.B(n_297),
.Y(n_319)
);

CKINVDCx14_ASAP7_75t_R g338 ( 
.A(n_296),
.Y(n_338)
);

NOR3xp33_ASAP7_75t_SL g297 ( 
.A(n_260),
.B(n_256),
.C(n_257),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_280),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_300),
.B(n_304),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_268),
.B(n_255),
.C(n_247),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_263),
.Y(n_303)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_303),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_260),
.B(n_229),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_305),
.A2(n_277),
.B1(n_281),
.B2(n_286),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_306),
.A2(n_275),
.B1(n_274),
.B2(n_266),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_268),
.B(n_240),
.C(n_232),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_307),
.B(n_308),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_261),
.B(n_228),
.C(n_249),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_263),
.Y(n_309)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_309),
.Y(n_328)
);

AOI32xp33_ASAP7_75t_L g310 ( 
.A1(n_269),
.A2(n_251),
.A3(n_288),
.B1(n_279),
.B2(n_267),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_313),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_283),
.B(n_285),
.C(n_286),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_311),
.B(n_265),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_262),
.B(n_283),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_270),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_315),
.A2(n_288),
.B(n_273),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_316),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_317),
.B(n_337),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_318),
.A2(n_320),
.B1(n_299),
.B2(n_295),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_301),
.A2(n_282),
.B1(n_274),
.B2(n_269),
.Y(n_320)
);

AOI21x1_ASAP7_75t_L g353 ( 
.A1(n_322),
.A2(n_315),
.B(n_294),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_325),
.B(n_336),
.Y(n_342)
);

OR2x2_ASAP7_75t_L g348 ( 
.A(n_326),
.B(n_298),
.Y(n_348)
);

INVxp33_ASAP7_75t_L g327 ( 
.A(n_306),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_327),
.B(n_329),
.Y(n_345)
);

OA21x2_ASAP7_75t_L g329 ( 
.A1(n_301),
.A2(n_275),
.B(n_273),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_314),
.B(n_267),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_330),
.B(n_331),
.Y(n_341)
);

XOR2x2_ASAP7_75t_L g331 ( 
.A(n_302),
.B(n_282),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_334),
.B(n_311),
.Y(n_346)
);

AOI321xp33_ASAP7_75t_L g335 ( 
.A1(n_297),
.A2(n_282),
.A3(n_264),
.B1(n_276),
.B2(n_266),
.C(n_271),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_335),
.A2(n_316),
.B(n_294),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_291),
.B(n_264),
.Y(n_336)
);

OA22x2_ASAP7_75t_L g337 ( 
.A1(n_298),
.A2(n_287),
.B1(n_278),
.B2(n_284),
.Y(n_337)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_321),
.Y(n_339)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_339),
.Y(n_364)
);

BUFx12_ASAP7_75t_L g340 ( 
.A(n_331),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_340),
.B(n_349),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_336),
.B(n_292),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_344),
.B(n_346),
.Y(n_361)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_323),
.Y(n_347)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_347),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_348),
.A2(n_351),
.B1(n_352),
.B2(n_355),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_333),
.B(n_307),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_328),
.Y(n_350)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_350),
.Y(n_369)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_327),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_319),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_353),
.A2(n_354),
.B(n_324),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_320),
.A2(n_299),
.B1(n_295),
.B2(n_308),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_356),
.A2(n_338),
.B1(n_335),
.B2(n_318),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_349),
.B(n_344),
.C(n_342),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_357),
.B(n_358),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_342),
.B(n_333),
.C(n_332),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_SL g359 ( 
.A(n_341),
.B(n_330),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_359),
.B(n_362),
.Y(n_381)
);

NOR2xp67_ASAP7_75t_L g363 ( 
.A(n_341),
.B(n_334),
.Y(n_363)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_363),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_365),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_355),
.B(n_332),
.C(n_325),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_367),
.B(n_370),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_353),
.B(n_322),
.C(n_312),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_362),
.A2(n_343),
.B(n_340),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_371),
.B(n_374),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_360),
.A2(n_340),
.B(n_345),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_366),
.A2(n_345),
.B(n_354),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_375),
.B(n_376),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_357),
.B(n_348),
.C(n_337),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_364),
.B(n_289),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_378),
.B(n_271),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_369),
.B(n_303),
.Y(n_380)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_380),
.Y(n_384)
);

AO21x1_ASAP7_75t_L g382 ( 
.A1(n_372),
.A2(n_373),
.B(n_376),
.Y(n_382)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_382),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_377),
.B(n_368),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_383),
.B(n_387),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_379),
.B(n_358),
.C(n_367),
.Y(n_387)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_388),
.Y(n_394)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_372),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_SL g392 ( 
.A(n_389),
.B(n_381),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_387),
.B(n_361),
.C(n_381),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_390),
.B(n_385),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_392),
.A2(n_393),
.B(n_384),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_386),
.A2(n_361),
.B(n_370),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_395),
.B(n_382),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_396),
.A2(n_398),
.B1(n_399),
.B2(n_390),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_397),
.Y(n_400)
);

AOI322xp5_ASAP7_75t_L g399 ( 
.A1(n_391),
.A2(n_293),
.A3(n_337),
.B1(n_329),
.B2(n_284),
.C1(n_359),
.C2(n_312),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_401),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_402),
.A2(n_400),
.B(n_394),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_403),
.B(n_337),
.C(n_329),
.Y(n_404)
);


endmodule