module real_jpeg_24317_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_364, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_364;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_1),
.A2(n_58),
.B1(n_59),
.B2(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_1),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_1),
.A2(n_77),
.B(n_82),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_1),
.B(n_91),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_1),
.A2(n_123),
.B1(n_147),
.B2(n_153),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_1),
.A2(n_36),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_1),
.B(n_48),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_2),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_44)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_2),
.A2(n_36),
.B1(n_37),
.B2(n_46),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_2),
.A2(n_46),
.B1(n_58),
.B2(n_59),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_2),
.A2(n_46),
.B1(n_81),
.B2(n_82),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_3),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_4),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_5),
.A2(n_58),
.B1(n_59),
.B2(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_5),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_5),
.A2(n_81),
.B1(n_82),
.B2(n_111),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_5),
.A2(n_36),
.B1(n_37),
.B2(n_111),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_5),
.A2(n_23),
.B1(n_26),
.B2(n_111),
.Y(n_237)
);

INVx8_ASAP7_75t_SL g35 ( 
.A(n_6),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_7),
.A2(n_24),
.B1(n_29),
.B2(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_7),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_7),
.A2(n_72),
.B1(n_81),
.B2(n_82),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_7),
.A2(n_58),
.B1(n_59),
.B2(n_72),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_7),
.A2(n_36),
.B1(n_37),
.B2(n_72),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_8),
.A2(n_23),
.B1(n_27),
.B2(n_28),
.Y(n_22)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_8),
.A2(n_27),
.B1(n_36),
.B2(n_37),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_8),
.A2(n_27),
.B1(n_81),
.B2(n_82),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_8),
.A2(n_27),
.B1(n_58),
.B2(n_59),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_9),
.A2(n_28),
.B1(n_45),
.B2(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_9),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_9),
.A2(n_70),
.B1(n_81),
.B2(n_82),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_9),
.A2(n_58),
.B1(n_59),
.B2(n_70),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g292 ( 
.A1(n_9),
.A2(n_36),
.B1(n_37),
.B2(n_70),
.Y(n_292)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_11),
.A2(n_58),
.B1(n_59),
.B2(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_11),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_11),
.A2(n_81),
.B1(n_82),
.B2(n_120),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_11),
.A2(n_36),
.B1(n_37),
.B2(n_120),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_11),
.A2(n_23),
.B1(n_41),
.B2(n_120),
.Y(n_249)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_13),
.A2(n_81),
.B1(n_82),
.B2(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_13),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_13),
.A2(n_58),
.B1(n_59),
.B2(n_128),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_13),
.A2(n_36),
.B1(n_37),
.B2(n_128),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_13),
.A2(n_23),
.B1(n_26),
.B2(n_128),
.Y(n_266)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_14),
.Y(n_60)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_15),
.Y(n_126)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_15),
.Y(n_132)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_15),
.Y(n_140)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_15),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_94),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_93),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_49),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_20),
.B(n_49),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_43),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_21),
.A2(n_32),
.B(n_69),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_30),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_22),
.B(n_48),
.Y(n_88)
);

OAI21xp33_ASAP7_75t_L g236 ( 
.A1(n_23),
.A2(n_107),
.B(n_217),
.Y(n_236)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI32xp33_ASAP7_75t_L g216 ( 
.A1(n_24),
.A2(n_33),
.A3(n_37),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_30),
.A2(n_48),
.B1(n_68),
.B2(n_71),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_30),
.A2(n_71),
.B(n_87),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_30),
.A2(n_48),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_30),
.A2(n_48),
.B1(n_237),
.B2(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_31),
.A2(n_32),
.B1(n_249),
.B2(n_266),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_31),
.A2(n_43),
.B(n_266),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_31),
.A2(n_88),
.B(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_40),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_32),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_34),
.B1(n_36),
.B2(n_37),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_34),
.B1(n_41),
.B2(n_42),
.Y(n_40)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_34),
.B(n_36),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_36),
.A2(n_37),
.B1(n_57),
.B2(n_61),
.Y(n_65)
);

OAI32xp33_ASAP7_75t_L g174 ( 
.A1(n_36),
.A2(n_57),
.A3(n_59),
.B1(n_166),
.B2(n_175),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_37),
.B(n_107),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_48),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_44),
.Y(n_315)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_45),
.B(n_107),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_86),
.C(n_89),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_50),
.A2(n_51),
.B1(n_357),
.B2(n_359),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_67),
.C(n_73),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_52),
.A2(n_53),
.B1(n_73),
.B2(n_74),
.Y(n_345)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_63),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_55),
.A2(n_64),
.B(n_231),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_62),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_56),
.A2(n_164),
.B1(n_167),
.B2(n_168),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_56),
.A2(n_63),
.B(n_292),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_59),
.B2(n_61),
.Y(n_56)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

OAI22xp33_ASAP7_75t_L g76 ( 
.A1(n_58),
.A2(n_59),
.B1(n_77),
.B2(n_79),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_58),
.B(n_61),
.Y(n_175)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_SL g112 ( 
.A1(n_59),
.A2(n_79),
.B(n_107),
.C(n_113),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_62),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_62),
.A2(n_167),
.B(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_66),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_64),
.A2(n_91),
.B(n_92),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_64),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_64),
.A2(n_91),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_64),
.A2(n_91),
.B1(n_192),
.B2(n_231),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_64),
.A2(n_91),
.B1(n_305),
.B2(n_306),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_64),
.A2(n_306),
.B(n_337),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_66),
.B(n_91),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g344 ( 
.A(n_67),
.B(n_345),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_73),
.A2(n_74),
.B1(n_336),
.B2(n_338),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_74),
.B(n_334),
.C(n_336),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_84),
.B(n_85),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_75),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_75),
.A2(n_84),
.B1(n_110),
.B2(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_75),
.A2(n_84),
.B1(n_119),
.B2(n_170),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_75),
.A2(n_85),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_75),
.B(n_257),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_80),
.Y(n_75)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_77),
.A2(n_79),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

BUFx24_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_80),
.A2(n_106),
.B1(n_108),
.B2(n_109),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_80),
.B(n_107),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_80),
.B(n_234),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_80),
.A2(n_255),
.B(n_256),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_80),
.A2(n_108),
.B1(n_255),
.B2(n_273),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_81),
.B(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_81),
.B(n_155),
.Y(n_154)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_84),
.B(n_85),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_86),
.A2(n_89),
.B1(n_90),
.B2(n_358),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_86),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_355),
.B(n_361),
.Y(n_94)
);

OAI321xp33_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_330),
.A3(n_348),
.B1(n_353),
.B2(n_354),
.C(n_364),
.Y(n_95)
);

AOI311xp33_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_283),
.A3(n_320),
.B(n_324),
.C(n_325),
.Y(n_96)
);

NOR3xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_239),
.C(n_278),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_211),
.B(n_238),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_185),
.B(n_210),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_159),
.B(n_184),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_133),
.B(n_158),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_114),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_103),
.B(n_114),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_112),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_104),
.A2(n_105),
.B1(n_112),
.B2(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_107),
.B(n_132),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_108),
.A2(n_206),
.B(n_207),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_108),
.A2(n_273),
.B(n_298),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_112),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_122),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_118),
.B2(n_121),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_116),
.B(n_121),
.C(n_122),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_118),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_127),
.B(n_129),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_123),
.A2(n_137),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_123),
.A2(n_177),
.B(n_178),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_123),
.A2(n_178),
.B(n_253),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_123),
.A2(n_148),
.B(n_177),
.Y(n_295)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_124),
.A2(n_136),
.B1(n_138),
.B2(n_139),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_124),
.B(n_181),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_124),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_219)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_127),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_129),
.B(n_201),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_130),
.Y(n_177)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_132),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_143),
.B(n_157),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_141),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_135),
.B(n_141),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_151),
.B(n_156),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_145),
.B(n_146),
.Y(n_156)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_148),
.Y(n_221)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_150),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_154),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_160),
.B(n_161),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_173),
.B1(n_182),
.B2(n_183),
.Y(n_161)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_162),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_169),
.B1(n_171),
.B2(n_172),
.Y(n_162)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_163),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_168),
.Y(n_191)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_169),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_172),
.C(n_182),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_170),
.Y(n_206)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_173),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_174),
.B(n_176),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_180),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_186),
.B(n_187),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_202),
.B2(n_203),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_188),
.B(n_205),
.C(n_208),
.Y(n_212)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_193),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_195),
.C(n_196),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_200),
.B(n_201),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_200),
.Y(n_220)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_208),
.B2(n_209),
.Y(n_203)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_204),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_205),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_207),
.B(n_256),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_212),
.B(n_213),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_228),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_225),
.B1(n_226),
.B2(n_227),
.Y(n_214)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_215),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_215),
.B(n_227),
.C(n_228),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_219),
.B1(n_223),
.B2(n_224),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_216),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_216),
.B(n_223),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_219),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_222),
.Y(n_253)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_225),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_235),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_232),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_232),
.C(n_235),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_233),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_234),
.Y(n_257)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

AOI21xp33_ASAP7_75t_L g326 ( 
.A1(n_240),
.A2(n_327),
.B(n_328),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_258),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_241),
.B(n_258),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_250),
.C(n_251),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_242),
.A2(n_243),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_244),
.B(n_246),
.C(n_247),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_250),
.B(n_251),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_254),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_254),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_259),
.A2(n_275),
.B1(n_276),
.B2(n_277),
.Y(n_258)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_259),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_270),
.B2(n_274),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_260),
.B(n_274),
.C(n_277),
.Y(n_322)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_264),
.B2(n_269),
.Y(n_261)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_262),
.Y(n_269)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_265),
.B(n_267),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_265),
.B(n_267),
.C(n_269),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_268),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_270),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_272),
.Y(n_288)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_275),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_279),
.B(n_280),
.Y(n_327)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

O2A1O1Ixp33_ASAP7_75t_SL g325 ( 
.A1(n_284),
.A2(n_321),
.B(n_326),
.C(n_329),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_301),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g324 ( 
.A(n_285),
.B(n_301),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_294),
.C(n_300),
.Y(n_285)
);

FAx1_ASAP7_75t_SL g323 ( 
.A(n_286),
.B(n_294),
.CI(n_300),
.CON(n_323),
.SN(n_323)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_289),
.B2(n_293),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_287),
.B(n_290),
.C(n_291),
.Y(n_319)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_289),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_292),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_297),
.B2(n_299),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_295),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_297),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_295),
.A2(n_299),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_299),
.A2(n_310),
.B(n_314),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_319),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_309),
.B1(n_317),
.B2(n_318),
.Y(n_302)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_303),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_307),
.B(n_308),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_304),
.B(n_307),
.Y(n_308)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_308),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_308),
.A2(n_332),
.B1(n_340),
.B2(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_309),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_309),
.B(n_317),
.C(n_319),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_311),
.B1(n_312),
.B2(n_316),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_312),
.Y(n_316)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_322),
.B(n_323),
.Y(n_329)
);

BUFx24_ASAP7_75t_SL g363 ( 
.A(n_323),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_342),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_331),
.B(n_342),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_340),
.C(n_341),
.Y(n_331)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_332),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_333),
.A2(n_334),
.B1(n_335),
.B2(n_339),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_333),
.A2(n_334),
.B1(n_344),
.B2(n_346),
.Y(n_343)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_334),
.B(n_346),
.C(n_347),
.Y(n_360)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_335),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_336),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_341),
.B(n_351),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_347),
.Y(n_342)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_344),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_349),
.B(n_350),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_360),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_356),
.B(n_360),
.Y(n_361)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_357),
.Y(n_359)
);


endmodule