module fake_jpeg_14972_n_396 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_396);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_396;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_11),
.B(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_39),
.Y(n_80)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_40),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_27),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_41),
.B(n_45),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

BUFx4f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_43),
.Y(n_113)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_23),
.B(n_38),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_52),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_14),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_49),
.B(n_54),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_0),
.Y(n_50)
);

AO22x1_ASAP7_75t_L g85 ( 
.A1(n_50),
.A2(n_33),
.B1(n_19),
.B2(n_15),
.Y(n_85)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_14),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_0),
.Y(n_56)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_21),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_60),
.Y(n_77)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_28),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_61),
.B(n_62),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_21),
.B(n_1),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_29),
.B(n_1),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_1),
.Y(n_96)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_16),
.Y(n_66)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_68),
.Y(n_119)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_18),
.Y(n_70)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_65),
.A2(n_26),
.B1(n_36),
.B2(n_32),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_71),
.A2(n_86),
.B(n_93),
.Y(n_148)
);

INVx13_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_74),
.B(n_79),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_43),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_75),
.A2(n_116),
.B1(n_112),
.B2(n_103),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_39),
.Y(n_79)
);

BUFx16f_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx13_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_48),
.Y(n_83)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_83),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_85),
.B(n_96),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_69),
.A2(n_32),
.B1(n_36),
.B2(n_53),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_41),
.B(n_22),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_87),
.B(n_100),
.Y(n_127)
);

BUFx4f_ASAP7_75t_SL g90 ( 
.A(n_48),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_90),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_55),
.A2(n_25),
.B1(n_24),
.B2(n_37),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_64),
.A2(n_37),
.B1(n_35),
.B2(n_20),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_94),
.A2(n_97),
.B1(n_118),
.B2(n_15),
.Y(n_146)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_70),
.A2(n_37),
.B1(n_35),
.B2(n_33),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_60),
.B(n_40),
.Y(n_100)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_52),
.Y(n_107)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_107),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_51),
.B(n_21),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_110),
.B(n_111),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_63),
.B(n_19),
.Y(n_111)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_42),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_112),
.B(n_116),
.Y(n_149)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_42),
.Y(n_114)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_47),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_47),
.Y(n_117)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_67),
.A2(n_35),
.B1(n_33),
.B2(n_19),
.Y(n_118)
);

CKINVDCx6p67_ASAP7_75t_R g120 ( 
.A(n_68),
.Y(n_120)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_120),
.Y(n_133)
);

AND2x4_ASAP7_75t_L g122 ( 
.A(n_50),
.B(n_33),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_1),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_124),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_125),
.B(n_155),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_100),
.B(n_50),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_128),
.B(n_132),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_73),
.Y(n_130)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_130),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_122),
.A2(n_66),
.B1(n_59),
.B2(n_68),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_131),
.A2(n_91),
.B1(n_89),
.B2(n_104),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_88),
.B(n_57),
.Y(n_132)
);

NAND2x1p5_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_18),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_135),
.B(n_144),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_103),
.A2(n_46),
.B1(n_70),
.B2(n_15),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_136),
.A2(n_93),
.B1(n_91),
.B2(n_95),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_18),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_142),
.B(n_151),
.Y(n_183)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_82),
.Y(n_143)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_146),
.A2(n_167),
.B1(n_6),
.B2(n_7),
.Y(n_215)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_74),
.Y(n_147)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_147),
.Y(n_198)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_99),
.Y(n_150)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_150),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_80),
.B(n_18),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_84),
.B(n_3),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_152),
.B(n_171),
.Y(n_213)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_78),
.Y(n_153)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_153),
.Y(n_187)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_92),
.Y(n_154)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_101),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_85),
.B(n_3),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_156),
.A2(n_102),
.B1(n_92),
.B2(n_83),
.Y(n_179)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_157),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_71),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_158),
.A2(n_12),
.B1(n_8),
.B2(n_9),
.Y(n_218)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_75),
.Y(n_159)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_159),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_81),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_161),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_113),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_76),
.Y(n_162)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_162),
.Y(n_209)
);

INVx11_ASAP7_75t_L g163 ( 
.A(n_76),
.Y(n_163)
);

INVx11_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_77),
.B(n_4),
.Y(n_164)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_164),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_109),
.B(n_4),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_6),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_119),
.Y(n_166)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_166),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_86),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_168),
.B(n_170),
.Y(n_211)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_98),
.Y(n_169)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_169),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_90),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_105),
.B(n_5),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_115),
.B(n_5),
.Y(n_172)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_172),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_97),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_173),
.B(n_119),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_124),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_175),
.B(n_192),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_135),
.B(n_90),
.C(n_107),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_177),
.B(n_195),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_178),
.A2(n_155),
.B(n_139),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_179),
.B(n_187),
.Y(n_254)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_181),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_191),
.A2(n_144),
.B1(n_123),
.B2(n_125),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_174),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_140),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_193),
.B(n_196),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_135),
.B(n_104),
.Y(n_195)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_157),
.Y(n_199)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_199),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g200 ( 
.A(n_134),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_200),
.Y(n_225)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_138),
.Y(n_202)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_202),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_149),
.Y(n_203)
);

INVxp33_ASAP7_75t_L g258 ( 
.A(n_203),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_204),
.A2(n_215),
.B1(n_219),
.B2(n_126),
.Y(n_248)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_138),
.Y(n_205)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_205),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_130),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_206),
.A2(n_207),
.B1(n_217),
.B2(n_163),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_173),
.A2(n_89),
.B1(n_120),
.B2(n_8),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_148),
.A2(n_120),
.B1(n_113),
.B2(n_8),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_212),
.A2(n_218),
.B1(n_126),
.B2(n_9),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_123),
.B(n_6),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_216),
.B(n_127),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_162),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_147),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_194),
.A2(n_148),
.B(n_159),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_221),
.A2(n_223),
.B(n_246),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_222),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_211),
.A2(n_156),
.B(n_144),
.Y(n_223)
);

OA21x2_ASAP7_75t_L g227 ( 
.A1(n_212),
.A2(n_156),
.B(n_151),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_227),
.B(n_229),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_180),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_228),
.B(n_231),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_176),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_230),
.A2(n_234),
.B1(n_251),
.B2(n_179),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_180),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_202),
.Y(n_232)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_232),
.Y(n_261)
);

AO21x1_ASAP7_75t_L g233 ( 
.A1(n_189),
.A2(n_142),
.B(n_165),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_233),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_197),
.A2(n_123),
.B1(n_169),
.B2(n_153),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_195),
.B(n_141),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_236),
.B(n_249),
.Y(n_273)
);

OA22x2_ASAP7_75t_L g237 ( 
.A1(n_204),
.A2(n_133),
.B1(n_154),
.B2(n_137),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_237),
.A2(n_254),
.B1(n_257),
.B2(n_214),
.Y(n_272)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_205),
.Y(n_238)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_238),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_240),
.B(n_242),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_182),
.A2(n_133),
.B1(n_134),
.B2(n_143),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_244),
.A2(n_198),
.B1(n_182),
.B2(n_217),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_197),
.A2(n_150),
.B(n_160),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_183),
.B(n_139),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_247),
.B(n_248),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_183),
.B(n_174),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_185),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_250),
.B(n_253),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_197),
.A2(n_166),
.B1(n_9),
.B2(n_10),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_177),
.A2(n_129),
.B(n_9),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_252),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_186),
.Y(n_253)
);

CKINVDCx6p67_ASAP7_75t_R g255 ( 
.A(n_190),
.Y(n_255)
);

INVx3_ASAP7_75t_SL g275 ( 
.A(n_255),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_203),
.B(n_129),
.Y(n_256)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_256),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_188),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_259),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_213),
.B(n_196),
.Y(n_260)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_260),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_262),
.A2(n_201),
.B1(n_209),
.B2(n_225),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_263),
.B(n_285),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_235),
.B(n_184),
.C(n_208),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_264),
.B(n_271),
.C(n_287),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_221),
.A2(n_218),
.B1(n_193),
.B2(n_210),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_265),
.A2(n_280),
.B1(n_288),
.B2(n_292),
.Y(n_304)
);

AOI22x1_ASAP7_75t_L g269 ( 
.A1(n_227),
.A2(n_219),
.B1(n_206),
.B2(n_198),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_269),
.A2(n_256),
.B1(n_237),
.B2(n_231),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_235),
.B(n_220),
.C(n_175),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_272),
.A2(n_278),
.B(n_242),
.Y(n_299)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_226),
.Y(n_277)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_277),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_234),
.B(n_7),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_254),
.A2(n_227),
.B1(n_247),
.B2(n_249),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_245),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_226),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_286),
.B(n_241),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_236),
.B(n_181),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_230),
.A2(n_246),
.B1(n_237),
.B2(n_254),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_233),
.B(n_199),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_251),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_237),
.A2(n_201),
.B1(n_209),
.B2(n_214),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_239),
.Y(n_293)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_293),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_294),
.A2(n_298),
.B1(n_306),
.B2(n_275),
.Y(n_324)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_266),
.Y(n_295)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_295),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_274),
.A2(n_257),
.B1(n_250),
.B2(n_252),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_296),
.A2(n_272),
.B1(n_270),
.B2(n_288),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_297),
.B(n_311),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_299),
.A2(n_313),
.B(n_319),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_260),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_300),
.B(n_303),
.Y(n_321)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_261),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_283),
.A2(n_224),
.B1(n_228),
.B2(n_238),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_267),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_307),
.B(n_308),
.Y(n_326)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_290),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_268),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_309),
.B(n_310),
.Y(n_329)
);

A2O1A1Ixp33_ASAP7_75t_L g310 ( 
.A1(n_276),
.A2(n_223),
.B(n_258),
.C(n_232),
.Y(n_310)
);

OAI32xp33_ASAP7_75t_L g311 ( 
.A1(n_291),
.A2(n_269),
.A3(n_280),
.B1(n_281),
.B2(n_284),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_292),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_312),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_284),
.A2(n_243),
.B(n_239),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_278),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_315),
.B(n_317),
.Y(n_336)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_286),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_316),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_282),
.B(n_241),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_318),
.B(n_285),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_274),
.A2(n_10),
.B(n_12),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_283),
.A2(n_255),
.B(n_190),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_320),
.A2(n_278),
.B(n_255),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_305),
.B(n_287),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_322),
.B(n_332),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_323),
.B(n_328),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_324),
.A2(n_336),
.B1(n_321),
.B2(n_333),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_312),
.A2(n_301),
.B1(n_298),
.B2(n_319),
.Y(n_327)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_327),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_296),
.A2(n_270),
.B1(n_265),
.B2(n_263),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_328),
.A2(n_331),
.B1(n_311),
.B2(n_314),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_304),
.A2(n_271),
.B1(n_264),
.B2(n_289),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_305),
.B(n_273),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_297),
.B(n_273),
.C(n_275),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_334),
.B(n_341),
.C(n_322),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_302),
.Y(n_338)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_338),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_339),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_340),
.A2(n_309),
.B(n_310),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_306),
.B(n_255),
.C(n_300),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_340),
.A2(n_313),
.B(n_320),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_342),
.B(n_353),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_343),
.B(n_347),
.C(n_349),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_332),
.B(n_295),
.C(n_304),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_348),
.A2(n_359),
.B1(n_350),
.B2(n_346),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_334),
.B(n_331),
.C(n_341),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_330),
.B(n_299),
.C(n_315),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_350),
.B(n_351),
.C(n_349),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_330),
.B(n_308),
.C(n_307),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_352),
.B(n_337),
.Y(n_371)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_326),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_326),
.B(n_303),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_354),
.B(n_356),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_355),
.B(n_358),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_329),
.B(n_316),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_329),
.B(n_325),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_362),
.B(n_369),
.C(n_357),
.Y(n_378)
);

A2O1A1Ixp33_ASAP7_75t_SL g364 ( 
.A1(n_359),
.A2(n_321),
.B(n_335),
.C(n_323),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_364),
.A2(n_370),
.B1(n_366),
.B2(n_361),
.Y(n_380)
);

INVxp33_ASAP7_75t_SL g366 ( 
.A(n_356),
.Y(n_366)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_366),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_343),
.B(n_347),
.C(n_351),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_367),
.B(n_371),
.Y(n_375)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_345),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_368),
.B(n_355),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_357),
.B(n_335),
.Y(n_369)
);

A2O1A1Ixp33_ASAP7_75t_SL g370 ( 
.A1(n_348),
.A2(n_337),
.B(n_344),
.C(n_358),
.Y(n_370)
);

CKINVDCx14_ASAP7_75t_R g377 ( 
.A(n_372),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_373),
.B(n_374),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_363),
.B(n_352),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_378),
.B(n_379),
.C(n_380),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_365),
.B(n_361),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_375),
.B(n_360),
.C(n_364),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_382),
.B(n_383),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_378),
.B(n_364),
.C(n_370),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_377),
.A2(n_364),
.B(n_370),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_385),
.B(n_370),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_381),
.B(n_380),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_386),
.A2(n_376),
.B(n_374),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_387),
.Y(n_389)
);

NOR2xp67_ASAP7_75t_SL g391 ( 
.A(n_390),
.B(n_386),
.Y(n_391)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_391),
.Y(n_392)
);

CKINVDCx14_ASAP7_75t_R g393 ( 
.A(n_392),
.Y(n_393)
);

OAI21x1_ASAP7_75t_L g394 ( 
.A1(n_393),
.A2(n_388),
.B(n_389),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_394),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_395),
.B(n_384),
.Y(n_396)
);


endmodule