module fake_jpeg_3868_n_309 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_309);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_309;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_SL g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_36),
.Y(n_51)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_42),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_17),
.B(n_12),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_38),
.B(n_45),
.Y(n_84)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_21),
.B(n_33),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_21),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_17),
.Y(n_68)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_23),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_28),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_47),
.B(n_30),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_49),
.A2(n_14),
.B1(n_19),
.B2(n_16),
.Y(n_70)
);

NAND2x1_ASAP7_75t_SL g50 ( 
.A(n_42),
.B(n_20),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_50),
.A2(n_76),
.B(n_98),
.C(n_34),
.Y(n_108)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_55),
.B(n_57),
.Y(n_101)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_58),
.Y(n_127)
);

CKINVDCx12_ASAP7_75t_R g59 ( 
.A(n_47),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_33),
.Y(n_60)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_23),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_62),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_24),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_63),
.B(n_69),
.Y(n_105)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_65),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

HB1xp67_ASAP7_75t_SL g117 ( 
.A(n_66),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_68),
.B(n_79),
.Y(n_116)
);

CKINVDCx9p33_ASAP7_75t_R g69 ( 
.A(n_47),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_70),
.A2(n_75),
.B1(n_91),
.B2(n_77),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_47),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_71),
.B(n_72),
.Y(n_112)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_74),
.B(n_78),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_41),
.A2(n_14),
.B1(n_19),
.B2(n_16),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_35),
.A2(n_32),
.B(n_30),
.Y(n_76)
);

AO22x2_ASAP7_75t_L g77 ( 
.A1(n_41),
.A2(n_22),
.B1(n_34),
.B2(n_26),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_77),
.A2(n_90),
.B1(n_95),
.B2(n_96),
.Y(n_118)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_31),
.Y(n_79)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_81),
.B(n_82),
.Y(n_120)
);

CKINVDCx12_ASAP7_75t_R g82 ( 
.A(n_44),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_43),
.B(n_18),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_83),
.B(n_92),
.Y(n_123)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_85),
.B(n_86),
.Y(n_121)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

CKINVDCx6p67_ASAP7_75t_R g87 ( 
.A(n_44),
.Y(n_87)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_87),
.Y(n_128)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_49),
.A2(n_24),
.B1(n_18),
.B2(n_25),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_35),
.B(n_31),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_36),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_99),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_36),
.B(n_25),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_97),
.Y(n_125)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_37),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_49),
.B(n_20),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_42),
.A2(n_20),
.B(n_22),
.C(n_30),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_67),
.B(n_22),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_109),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_108),
.A2(n_76),
.B1(n_70),
.B2(n_75),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_32),
.Y(n_109)
);

AND2x2_ASAP7_75t_SL g111 ( 
.A(n_50),
.B(n_0),
.Y(n_111)
);

OAI21xp33_ASAP7_75t_L g150 ( 
.A1(n_111),
.A2(n_1),
.B(n_2),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_115),
.B(n_77),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_51),
.B(n_1),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_91),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_54),
.Y(n_129)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_129),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_116),
.B(n_83),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_130),
.B(n_153),
.Y(n_168)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_131),
.B(n_137),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_108),
.A2(n_115),
.B1(n_109),
.B2(n_118),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_132),
.A2(n_134),
.B1(n_148),
.B2(n_160),
.Y(n_167)
);

NOR2x1_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_77),
.Y(n_133)
);

NAND3xp33_ASAP7_75t_L g174 ( 
.A(n_133),
.B(n_105),
.C(n_69),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_136),
.B(n_164),
.Y(n_176)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_122),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_139),
.Y(n_173)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_121),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_144),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_141),
.B(n_151),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_81),
.Y(n_142)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_142),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_111),
.A2(n_84),
.B(n_66),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_143),
.A2(n_136),
.B(n_154),
.Y(n_183)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_122),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_113),
.B(n_128),
.Y(n_145)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_145),
.Y(n_184)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_101),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_146),
.B(n_147),
.Y(n_179)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_101),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_104),
.A2(n_80),
.B1(n_56),
.B2(n_74),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_103),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_149),
.B(n_152),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_150),
.A2(n_3),
.B(n_4),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_87),
.Y(n_151)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_112),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_116),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_102),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_113),
.B(n_72),
.Y(n_155)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_155),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_123),
.B(n_87),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_162),
.Y(n_181)
);

OA22x2_ASAP7_75t_L g157 ( 
.A1(n_117),
.A2(n_111),
.B1(n_80),
.B2(n_73),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_157),
.A2(n_158),
.B1(n_105),
.B2(n_110),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_125),
.A2(n_56),
.B1(n_73),
.B2(n_90),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_65),
.Y(n_159)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_159),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_116),
.A2(n_53),
.B1(n_88),
.B2(n_96),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_125),
.A2(n_53),
.B1(n_95),
.B2(n_57),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_161),
.A2(n_102),
.B1(n_112),
.B2(n_106),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_100),
.Y(n_162)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_100),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_163),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_123),
.B(n_10),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_157),
.A2(n_106),
.B1(n_123),
.B2(n_125),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_165),
.B(n_9),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_148),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_166),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_169),
.B(n_185),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_171),
.A2(n_186),
.B1(n_194),
.B2(n_15),
.Y(n_220)
);

CKINVDCx12_ASAP7_75t_R g172 ( 
.A(n_157),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_172),
.B(n_192),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_174),
.B(n_168),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_157),
.A2(n_114),
.B1(n_124),
.B2(n_58),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_177),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_183),
.A2(n_193),
.B(n_199),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_135),
.B(n_124),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_133),
.A2(n_134),
.B1(n_132),
.B2(n_135),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_151),
.B(n_120),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_190),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_143),
.B(n_120),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_160),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_161),
.B(n_26),
.Y(n_193)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_158),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_195),
.B(n_198),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_150),
.B(n_1),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_3),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_162),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_196),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_218),
.Y(n_226)
);

A2O1A1O1Ixp25_ASAP7_75t_L g204 ( 
.A1(n_188),
.A2(n_134),
.B(n_15),
.C(n_34),
.D(n_26),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_204),
.B(n_194),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_149),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_206),
.B(n_208),
.C(n_210),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_114),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_198),
.B(n_152),
.Y(n_209)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_209),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_187),
.B(n_144),
.C(n_137),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_211),
.B(n_214),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_183),
.B(n_163),
.C(n_114),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_167),
.C(n_181),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_180),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_185),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_215),
.B(n_223),
.Y(n_240)
);

NAND2xp33_ASAP7_75t_SL g237 ( 
.A(n_216),
.B(n_221),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_175),
.B(n_15),
.Y(n_217)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_217),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_178),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_220),
.A2(n_224),
.B1(n_199),
.B2(n_168),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_9),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_176),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_175),
.B(n_191),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_192),
.A2(n_127),
.B1(n_4),
.B2(n_5),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_197),
.A2(n_3),
.B(n_4),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_225),
.A2(n_181),
.B(n_193),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_233),
.C(n_241),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_212),
.A2(n_166),
.B1(n_195),
.B2(n_193),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_229),
.A2(n_238),
.B1(n_245),
.B2(n_189),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_203),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_230),
.B(n_244),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_232),
.A2(n_179),
.B1(n_214),
.B2(n_180),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_247),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_200),
.B(n_169),
.Y(n_235)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_235),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_212),
.A2(n_171),
.B1(n_167),
.B2(n_172),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_206),
.B(n_176),
.C(n_182),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_246),
.C(n_208),
.Y(n_251)
);

AOI221xp5_ASAP7_75t_L g243 ( 
.A1(n_219),
.A2(n_207),
.B1(n_201),
.B2(n_204),
.C(n_220),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_173),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_210),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_219),
.A2(n_205),
.B1(n_213),
.B2(n_215),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_207),
.B(n_182),
.C(n_191),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_200),
.B(n_184),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_236),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_257),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_253),
.C(n_256),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_221),
.C(n_222),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_211),
.Y(n_255)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_255),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_227),
.B(n_184),
.C(n_224),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_226),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_247),
.B(n_225),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_258),
.A2(n_263),
.B(n_231),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_260),
.Y(n_273)
);

NAND3xp33_ASAP7_75t_SL g260 ( 
.A(n_238),
.B(n_205),
.C(n_189),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_261),
.A2(n_232),
.B1(n_228),
.B2(n_237),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_239),
.B(n_170),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_240),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_254),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_264),
.A2(n_265),
.B(n_267),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_263),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_248),
.A2(n_229),
.B1(n_245),
.B2(n_234),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_266),
.A2(n_271),
.B1(n_250),
.B2(n_255),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_248),
.A2(n_244),
.B(n_233),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_270),
.A2(n_4),
.B(n_5),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_258),
.A2(n_246),
.B1(n_252),
.B2(n_261),
.Y(n_271)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_274),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_242),
.C(n_241),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_253),
.C(n_127),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_276),
.A2(n_250),
.B(n_256),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_5),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_280),
.A2(n_267),
.B(n_276),
.Y(n_288)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_269),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_282),
.Y(n_294)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_270),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_272),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_283),
.A2(n_284),
.B(n_286),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_265),
.B(n_259),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_285),
.B(n_268),
.C(n_127),
.Y(n_290)
);

NOR3xp33_ASAP7_75t_L g287 ( 
.A(n_273),
.B(n_10),
.C(n_12),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_6),
.Y(n_296)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_288),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_280),
.A2(n_268),
.B(n_275),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_289),
.B(n_293),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_291),
.Y(n_299)
);

XNOR2x1_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_10),
.Y(n_292)
);

OAI21xp33_ASAP7_75t_L g302 ( 
.A1(n_292),
.A2(n_6),
.B(n_286),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_12),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_296),
.Y(n_301)
);

INVxp33_ASAP7_75t_SL g297 ( 
.A(n_292),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_297),
.B(n_302),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_298),
.B(n_290),
.C(n_285),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_303),
.A2(n_304),
.B(n_295),
.Y(n_306)
);

NOR2xp67_ASAP7_75t_L g304 ( 
.A(n_299),
.B(n_293),
.Y(n_304)
);

AO221x1_ASAP7_75t_L g308 ( 
.A1(n_306),
.A2(n_307),
.B1(n_291),
.B2(n_300),
.C(n_294),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_305),
.B(n_279),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_301),
.C(n_6),
.Y(n_309)
);


endmodule