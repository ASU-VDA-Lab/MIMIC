module real_jpeg_4722_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_323;
wire n_176;
wire n_215;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_155;
wire n_120;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_0),
.A2(n_134),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_0),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_0),
.A2(n_204),
.B1(n_211),
.B2(n_233),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g323 ( 
.A1(n_0),
.A2(n_164),
.B1(n_233),
.B2(n_324),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_0),
.A2(n_33),
.B1(n_145),
.B2(n_233),
.Y(n_451)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_1),
.A2(n_48),
.B1(n_52),
.B2(n_53),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_1),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_1),
.A2(n_53),
.B1(n_332),
.B2(n_335),
.Y(n_331)
);

OAI22xp33_ASAP7_75t_SL g409 ( 
.A1(n_1),
.A2(n_53),
.B1(n_191),
.B2(n_410),
.Y(n_409)
);

AOI22xp33_ASAP7_75t_SL g423 ( 
.A1(n_1),
.A2(n_53),
.B1(n_96),
.B2(n_424),
.Y(n_423)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_2),
.A2(n_95),
.B1(n_99),
.B2(n_101),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_2),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_2),
.A2(n_101),
.B1(n_131),
.B2(n_133),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_2),
.A2(n_101),
.B1(n_405),
.B2(n_406),
.Y(n_404)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_3),
.A2(n_88),
.B1(n_91),
.B2(n_92),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_3),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_3),
.A2(n_92),
.B1(n_143),
.B2(n_144),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_SL g401 ( 
.A1(n_3),
.A2(n_92),
.B1(n_402),
.B2(n_403),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_3),
.A2(n_92),
.B1(n_303),
.B2(n_434),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_4),
.A2(n_188),
.B1(n_190),
.B2(n_191),
.Y(n_187)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_4),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_4),
.A2(n_190),
.B1(n_224),
.B2(n_228),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_4),
.A2(n_90),
.B1(n_100),
.B2(n_190),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_4),
.A2(n_190),
.B1(n_357),
.B2(n_381),
.Y(n_380)
);

BUFx5_ASAP7_75t_L g216 ( 
.A(n_5),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_5),
.Y(n_222)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_5),
.Y(n_246)
);

INVx8_ASAP7_75t_L g261 ( 
.A(n_5),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_5),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_5),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g156 ( 
.A(n_6),
.Y(n_156)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_6),
.Y(n_358)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_6),
.Y(n_383)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_7),
.Y(n_354)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_8),
.Y(n_530)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_9),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_9),
.Y(n_121)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_10),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_11),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_11),
.Y(n_125)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_11),
.Y(n_209)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_12),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_13),
.A2(n_57),
.B1(n_59),
.B2(n_61),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_13),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_13),
.A2(n_61),
.B1(n_164),
.B2(n_166),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g364 ( 
.A1(n_13),
.A2(n_61),
.B1(n_365),
.B2(n_369),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_13),
.A2(n_61),
.B1(n_412),
.B2(n_414),
.Y(n_411)
);

OAI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_14),
.A2(n_204),
.B1(n_210),
.B2(n_211),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_14),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_14),
.A2(n_131),
.B1(n_210),
.B2(n_273),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g386 ( 
.A1(n_14),
.A2(n_210),
.B1(n_355),
.B2(n_387),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_14),
.A2(n_210),
.B1(n_427),
.B2(n_428),
.Y(n_426)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_16),
.A2(n_182),
.B1(n_184),
.B2(n_185),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_16),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_16),
.B(n_199),
.C(n_200),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_16),
.B(n_78),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_16),
.B(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_16),
.B(n_129),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_16),
.B(n_286),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_17),
.Y(n_533)
);

OAI22xp33_ASAP7_75t_L g154 ( 
.A1(n_18),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_18),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g293 ( 
.A1(n_18),
.A2(n_155),
.B1(n_294),
.B2(n_296),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g390 ( 
.A1(n_18),
.A2(n_155),
.B1(n_191),
.B2(n_391),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_18),
.A2(n_155),
.B1(n_301),
.B2(n_419),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_528),
.B(n_531),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_171),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_169),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_146),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_23),
.B(n_146),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_136),
.B2(n_137),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_62),
.C(n_102),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_26),
.B(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_47),
.B1(n_54),
.B2(n_56),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_27),
.A2(n_54),
.B1(n_56),
.B2(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_27),
.A2(n_47),
.B1(n_54),
.B2(n_153),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_27),
.A2(n_379),
.B(n_426),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_27),
.A2(n_37),
.B1(n_426),
.B2(n_451),
.Y(n_450)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_28),
.A2(n_377),
.B(n_378),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_28),
.B(n_380),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_37),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g427 ( 
.A(n_33),
.Y(n_427)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_34),
.Y(n_145)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_34),
.Y(n_157)
);

INVx3_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_37),
.B(n_185),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_42),
.B2(n_44),
.Y(n_37)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_40),
.Y(n_302)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_41),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_41),
.Y(n_388)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx6_ASAP7_75t_L g350 ( 
.A(n_43),
.Y(n_350)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI32xp33_ASAP7_75t_L g346 ( 
.A1(n_45),
.A2(n_347),
.A3(n_351),
.B1(n_352),
.B2(n_356),
.Y(n_346)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_52),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_54),
.A2(n_451),
.B(n_473),
.Y(n_483)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_55),
.B(n_380),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_55),
.B(n_154),
.Y(n_472)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_62),
.A2(n_102),
.B1(n_103),
.B2(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_62),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_87),
.B1(n_93),
.B2(n_94),
.Y(n_62)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_63),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_63),
.A2(n_87),
.B1(n_93),
.B2(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_63),
.A2(n_93),
.B1(n_323),
.B2(n_386),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_63),
.A2(n_93),
.B1(n_418),
.B2(n_423),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_78),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_68),
.B1(n_72),
.B2(n_77),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_66),
.Y(n_308)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_67),
.Y(n_312)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_71),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_71),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_71),
.Y(n_422)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_78),
.A2(n_139),
.B(n_140),
.Y(n_138)
);

AOI22x1_ASAP7_75t_L g452 ( 
.A1(n_78),
.A2(n_139),
.B1(n_327),
.B2(n_453),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_78),
.A2(n_139),
.B1(n_163),
.B2(n_461),
.Y(n_460)
);

AO22x2_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_81),
.B2(n_86),
.Y(n_78)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_SL g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g415 ( 
.A(n_82),
.Y(n_415)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_84),
.Y(n_86)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_84),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_84),
.Y(n_184)
);

INVx5_ASAP7_75t_L g305 ( 
.A(n_84),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_84),
.Y(n_410)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_85),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g193 ( 
.A(n_85),
.Y(n_193)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_85),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_85),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_86),
.Y(n_183)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_93),
.B(n_289),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_93),
.A2(n_323),
.B(n_326),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_94),
.Y(n_140)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx4_ASAP7_75t_SL g96 ( 
.A(n_97),
.Y(n_96)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_102),
.B(n_152),
.C(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_102),
.A2(n_103),
.B1(n_160),
.B2(n_161),
.Y(n_517)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_128),
.B(n_130),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_104),
.A2(n_181),
.B(n_186),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_104),
.A2(n_128),
.B1(n_232),
.B2(n_272),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_104),
.A2(n_186),
.B(n_272),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_104),
.A2(n_128),
.B1(n_390),
.B2(n_445),
.Y(n_444)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_105),
.B(n_187),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_105),
.A2(n_129),
.B1(n_409),
.B2(n_411),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_105),
.A2(n_129),
.B1(n_411),
.B2(n_433),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_105),
.A2(n_129),
.B1(n_433),
.B2(n_464),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_118),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_110),
.B1(n_113),
.B2(n_116),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_109),
.Y(n_197)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_109),
.Y(n_436)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_112),
.Y(n_115)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_117),
.Y(n_235)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_118),
.A2(n_232),
.B(n_236),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_122),
.B1(n_124),
.B2(n_126),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_120),
.Y(n_199)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g200 ( 
.A(n_123),
.Y(n_200)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_123),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_123),
.Y(n_296)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_123),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_123),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g335 ( 
.A(n_124),
.Y(n_335)
);

BUFx8_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g295 ( 
.A(n_125),
.Y(n_295)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_125),
.Y(n_368)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_128),
.A2(n_236),
.B(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_129),
.B(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_130),
.Y(n_464)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp33_ASAP7_75t_SL g309 ( 
.A(n_133),
.B(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_141),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_139),
.A2(n_280),
.B(n_288),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_139),
.B(n_327),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_139),
.A2(n_288),
.B(n_486),
.Y(n_485)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_151),
.C(n_158),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_147),
.A2(n_148),
.B1(n_151),
.B2(n_152),
.Y(n_523)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_151),
.A2(n_152),
.B1(n_517),
.B2(n_518),
.Y(n_516)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx3_ASAP7_75t_L g351 ( 
.A(n_156),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g521 ( 
.A1(n_158),
.A2(n_159),
.B1(n_522),
.B2(n_523),
.Y(n_521)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_168),
.Y(n_283)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_168),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_168),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_512),
.B(n_525),
.Y(n_172)
);

OAI311xp33_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_395),
.A3(n_488),
.B1(n_506),
.C1(n_511),
.Y(n_173)
);

AOI21x1_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_340),
.B(n_394),
.Y(n_174)
);

AO21x1_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_314),
.B(n_339),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_266),
.B(n_313),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_239),
.B(n_265),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_201),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_179),
.B(n_201),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_194),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_180),
.A2(n_194),
.B1(n_195),
.B2(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_180),
.Y(n_263)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx11_ASAP7_75t_L g189 ( 
.A(n_184),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_185),
.A2(n_214),
.B(n_220),
.Y(n_247)
);

OAI21xp33_ASAP7_75t_SL g280 ( 
.A1(n_185),
.A2(n_281),
.B(n_284),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_185),
.B(n_357),
.Y(n_356)
);

OAI21xp33_ASAP7_75t_SL g377 ( 
.A1(n_185),
.A2(n_356),
.B(n_357),
.Y(n_377)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_198),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_229),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_202),
.B(n_230),
.C(n_238),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_214),
.B(n_220),
.Y(n_202)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_203),
.Y(n_258)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_208),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_209),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g334 ( 
.A(n_209),
.Y(n_334)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_211),
.Y(n_243)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_213),
.Y(n_228)
);

INVx4_ASAP7_75t_L g407 ( 
.A(n_213),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_214),
.A2(n_361),
.B1(n_362),
.B2(n_363),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_214),
.A2(n_362),
.B1(n_401),
.B2(n_404),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_214),
.A2(n_404),
.B(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_215),
.B(n_223),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_215),
.A2(n_257),
.B1(n_258),
.B2(n_259),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_215),
.A2(n_293),
.B1(n_331),
.B2(n_336),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_215),
.A2(n_364),
.B1(n_447),
.B2(n_448),
.Y(n_446)
);

OR2x2_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_223),
.Y(n_220)
);

INVx4_ASAP7_75t_L g362 ( 
.A(n_221),
.Y(n_362)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_237),
.B2(n_238),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_255),
.B(n_264),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_248),
.B(n_254),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_247),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_246),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_253),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_249),
.B(n_253),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_251),
.B(n_252),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_250),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_252),
.A2(n_292),
.B(n_297),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_262),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_262),
.Y(n_264)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_267),
.B(n_268),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_290),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_278),
.B2(n_279),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_271),
.B(n_278),
.C(n_290),
.Y(n_315)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx5_ASAP7_75t_SL g274 ( 
.A(n_275),
.Y(n_274)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_281),
.Y(n_424)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVxp33_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

AOI32xp33_ASAP7_75t_L g300 ( 
.A1(n_285),
.A2(n_301),
.A3(n_303),
.B1(n_306),
.B2(n_309),
.Y(n_300)
);

INVx6_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_289),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_300),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_291),
.B(n_300),
.Y(n_320)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx3_ASAP7_75t_SL g297 ( 
.A(n_298),
.Y(n_297)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_299),
.Y(n_337)
);

INVx8_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx5_ASAP7_75t_L g392 ( 
.A(n_305),
.Y(n_392)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_315),
.B(n_316),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_318),
.B1(n_321),
.B2(n_338),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_319),
.B(n_320),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_319),
.B(n_320),
.C(n_338),
.Y(n_341)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_321),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_322),
.B(n_328),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_322),
.B(n_329),
.C(n_330),
.Y(n_371)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_331),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_333),
.Y(n_332)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_334),
.Y(n_370)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_334),
.Y(n_402)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_341),
.B(n_342),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_374),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_344),
.A2(n_371),
.B1(n_372),
.B2(n_373),
.Y(n_343)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_344),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_345),
.A2(n_346),
.B1(n_359),
.B2(n_360),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_346),
.B(n_359),
.Y(n_484)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_355),
.Y(n_352)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx6_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

BUFx2_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_371),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_371),
.B(n_372),
.C(n_374),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_375),
.A2(n_376),
.B1(n_384),
.B2(n_393),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_375),
.B(n_385),
.C(n_389),
.Y(n_497)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx4_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_383),
.Y(n_429)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_384),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_SL g384 ( 
.A(n_385),
.B(n_389),
.Y(n_384)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_386),
.Y(n_486)
);

INVx6_ASAP7_75t_SL g387 ( 
.A(n_388),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

NAND2xp33_ASAP7_75t_SL g395 ( 
.A(n_396),
.B(n_474),
.Y(n_395)
);

A2O1A1Ixp33_ASAP7_75t_SL g506 ( 
.A1(n_396),
.A2(n_474),
.B(n_507),
.C(n_510),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_454),
.Y(n_396)
);

OR2x2_ASAP7_75t_L g511 ( 
.A(n_397),
.B(n_454),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_430),
.C(n_442),
.Y(n_397)
);

FAx1_ASAP7_75t_SL g487 ( 
.A(n_398),
.B(n_430),
.CI(n_442),
.CON(n_487),
.SN(n_487)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_416),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_399),
.B(n_417),
.C(n_425),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_408),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_400),
.B(n_408),
.Y(n_480)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_401),
.Y(n_447)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_409),
.Y(n_445)
);

INVx5_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_425),
.Y(n_416)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_418),
.Y(n_453)
);

INVx1_ASAP7_75t_SL g419 ( 
.A(n_420),
.Y(n_419)
);

INVx5_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_423),
.Y(n_461)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_431),
.A2(n_432),
.B1(n_437),
.B2(n_441),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_432),
.B(n_437),
.Y(n_468)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_437),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_437),
.A2(n_441),
.B1(n_470),
.B2(n_471),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g515 ( 
.A1(n_437),
.A2(n_468),
.B(n_471),
.Y(n_515)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_440),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_449),
.C(n_452),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_443),
.B(n_478),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_444),
.B(n_446),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_444),
.B(n_446),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_449),
.A2(n_450),
.B1(n_452),
.B2(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_452),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_456),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_455),
.B(n_458),
.C(n_466),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_457),
.A2(n_458),
.B1(n_466),
.B2(n_467),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_459),
.A2(n_462),
.B(n_465),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_460),
.B(n_463),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

FAx1_ASAP7_75t_SL g514 ( 
.A(n_465),
.B(n_515),
.CI(n_516),
.CON(n_514),
.SN(n_514)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_465),
.B(n_515),
.C(n_516),
.Y(n_524)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_469),
.Y(n_467)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_473),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_487),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_475),
.B(n_487),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_480),
.C(n_481),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_476),
.A2(n_477),
.B1(n_480),
.B2(n_500),
.Y(n_499)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_480),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_481),
.B(n_499),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_484),
.C(n_485),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_482),
.A2(n_483),
.B1(n_485),
.B2(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_484),
.B(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_485),
.Y(n_494)
);

BUFx24_ASAP7_75t_SL g535 ( 
.A(n_487),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_489),
.B(n_501),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_490),
.A2(n_508),
.B(n_509),
.Y(n_507)
);

NOR2x1_ASAP7_75t_L g490 ( 
.A(n_491),
.B(n_498),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_491),
.B(n_498),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_495),
.C(n_497),
.Y(n_491)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_492),
.B(n_504),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_495),
.A2(n_496),
.B1(n_497),
.B2(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_497),
.Y(n_505)
);

OR2x2_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_503),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_502),
.B(n_503),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_513),
.B(n_520),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_514),
.B(n_519),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_514),
.B(n_519),
.Y(n_526)
);

BUFx24_ASAP7_75t_SL g536 ( 
.A(n_514),
.Y(n_536)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_517),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_520),
.A2(n_526),
.B(n_527),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_521),
.B(n_524),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_521),
.B(n_524),
.Y(n_527)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

INVx13_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

INVx5_ASAP7_75t_L g532 ( 
.A(n_530),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_532),
.B(n_533),
.Y(n_531)
);


endmodule