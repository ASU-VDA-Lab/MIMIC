module fake_netlist_1_5263_n_543 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_543);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_543;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g78 ( .A(n_53), .Y(n_78) );
CKINVDCx16_ASAP7_75t_R g79 ( .A(n_71), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_47), .Y(n_80) );
CKINVDCx16_ASAP7_75t_R g81 ( .A(n_66), .Y(n_81) );
BUFx3_ASAP7_75t_L g82 ( .A(n_32), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_20), .Y(n_83) );
BUFx2_ASAP7_75t_L g84 ( .A(n_12), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_63), .Y(n_85) );
BUFx6f_ASAP7_75t_L g86 ( .A(n_76), .Y(n_86) );
CKINVDCx20_ASAP7_75t_R g87 ( .A(n_73), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_69), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_40), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_16), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_36), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_28), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_9), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_77), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_60), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_3), .Y(n_96) );
NOR2xp67_ASAP7_75t_L g97 ( .A(n_56), .B(n_34), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_72), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_65), .Y(n_99) );
INVxp67_ASAP7_75t_L g100 ( .A(n_59), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_55), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_0), .Y(n_102) );
CKINVDCx14_ASAP7_75t_R g103 ( .A(n_75), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_70), .Y(n_104) );
BUFx2_ASAP7_75t_L g105 ( .A(n_23), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_6), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_10), .Y(n_107) );
BUFx6f_ASAP7_75t_L g108 ( .A(n_10), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_45), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_5), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_21), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_0), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_1), .Y(n_113) );
BUFx2_ASAP7_75t_L g114 ( .A(n_84), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_105), .Y(n_115) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_86), .Y(n_116) );
BUFx6f_ASAP7_75t_L g117 ( .A(n_86), .Y(n_117) );
AOI22xp5_ASAP7_75t_L g118 ( .A1(n_84), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_105), .B(n_2), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_112), .B(n_4), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_93), .Y(n_121) );
AND2x4_ASAP7_75t_L g122 ( .A(n_82), .B(n_4), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_112), .B(n_5), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_111), .Y(n_124) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_86), .Y(n_125) );
BUFx3_ASAP7_75t_L g126 ( .A(n_82), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_103), .B(n_6), .Y(n_127) );
BUFx2_ASAP7_75t_L g128 ( .A(n_113), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_86), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_96), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_86), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_111), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_88), .Y(n_133) );
BUFx2_ASAP7_75t_L g134 ( .A(n_113), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_88), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_80), .Y(n_136) );
AND2x2_ASAP7_75t_L g137 ( .A(n_114), .B(n_103), .Y(n_137) );
BUFx3_ASAP7_75t_L g138 ( .A(n_126), .Y(n_138) );
INVx3_ASAP7_75t_L g139 ( .A(n_122), .Y(n_139) );
BUFx10_ASAP7_75t_L g140 ( .A(n_115), .Y(n_140) );
AND2x2_ASAP7_75t_L g141 ( .A(n_114), .B(n_79), .Y(n_141) );
INVx2_ASAP7_75t_SL g142 ( .A(n_126), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_133), .B(n_83), .Y(n_143) );
NAND2xp33_ASAP7_75t_L g144 ( .A(n_127), .B(n_78), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_124), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_116), .Y(n_146) );
NOR2xp33_ASAP7_75t_L g147 ( .A(n_128), .B(n_100), .Y(n_147) );
AOI22xp33_ASAP7_75t_L g148 ( .A1(n_127), .A2(n_110), .B1(n_102), .B2(n_107), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_133), .B(n_109), .Y(n_149) );
NOR2xp33_ASAP7_75t_SL g150 ( .A(n_122), .B(n_81), .Y(n_150) );
AOI22xp33_ASAP7_75t_L g151 ( .A1(n_122), .A2(n_106), .B1(n_108), .B2(n_104), .Y(n_151) );
INVx6_ASAP7_75t_L g152 ( .A(n_117), .Y(n_152) );
AND2x2_ASAP7_75t_L g153 ( .A(n_128), .B(n_78), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_135), .B(n_94), .Y(n_154) );
INVx1_ASAP7_75t_SL g155 ( .A(n_134), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_135), .B(n_92), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_124), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_116), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_136), .B(n_95), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_134), .B(n_121), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_116), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_132), .Y(n_162) );
CKINVDCx5p33_ASAP7_75t_R g163 ( .A(n_155), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_160), .B(n_119), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_139), .A2(n_136), .B(n_132), .Y(n_165) );
INVx3_ASAP7_75t_L g166 ( .A(n_139), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_137), .B(n_130), .Y(n_167) );
AOI22xp33_ASAP7_75t_L g168 ( .A1(n_139), .A2(n_123), .B1(n_120), .B2(n_108), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_145), .Y(n_169) );
BUFx12f_ASAP7_75t_L g170 ( .A(n_140), .Y(n_170) );
INVx3_ASAP7_75t_L g171 ( .A(n_139), .Y(n_171) );
AND2x6_ASAP7_75t_SL g172 ( .A(n_141), .B(n_85), .Y(n_172) );
AOI22xp33_ASAP7_75t_L g173 ( .A1(n_153), .A2(n_108), .B1(n_118), .B2(n_87), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_137), .B(n_153), .Y(n_174) );
OR2x6_ASAP7_75t_L g175 ( .A(n_153), .B(n_108), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_140), .B(n_89), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_145), .Y(n_177) );
AO22x1_ASAP7_75t_L g178 ( .A1(n_137), .A2(n_89), .B1(n_99), .B2(n_90), .Y(n_178) );
OAI22xp5_ASAP7_75t_L g179 ( .A1(n_148), .A2(n_87), .B1(n_108), .B2(n_101), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_157), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_140), .B(n_91), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_157), .Y(n_182) );
INVxp67_ASAP7_75t_L g183 ( .A(n_155), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_140), .B(n_98), .Y(n_184) );
INVx2_ASAP7_75t_SL g185 ( .A(n_141), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_162), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_150), .B(n_97), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_147), .B(n_131), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_150), .B(n_131), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_162), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_144), .B(n_41), .Y(n_191) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_142), .B(n_39), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_143), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_146), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_151), .B(n_131), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_166), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_193), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_193), .B(n_159), .Y(n_198) );
AND2x4_ASAP7_75t_L g199 ( .A(n_183), .B(n_159), .Y(n_199) );
INVx3_ASAP7_75t_SL g200 ( .A(n_163), .Y(n_200) );
AND2x4_ASAP7_75t_L g201 ( .A(n_175), .B(n_143), .Y(n_201) );
INVx3_ASAP7_75t_L g202 ( .A(n_170), .Y(n_202) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_170), .B(n_138), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_170), .B(n_138), .Y(n_204) );
BUFx3_ASAP7_75t_L g205 ( .A(n_175), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_181), .A2(n_142), .B(n_138), .Y(n_206) );
A2O1A1Ixp33_ASAP7_75t_L g207 ( .A1(n_177), .A2(n_149), .B(n_156), .C(n_154), .Y(n_207) );
AOI221xp5_ASAP7_75t_L g208 ( .A1(n_174), .A2(n_156), .B1(n_154), .B2(n_149), .C(n_142), .Y(n_208) );
AOI22xp33_ASAP7_75t_L g209 ( .A1(n_175), .A2(n_131), .B1(n_117), .B2(n_129), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_169), .B(n_125), .Y(n_210) );
A2O1A1Ixp33_ASAP7_75t_L g211 ( .A1(n_177), .A2(n_125), .B(n_116), .C(n_129), .Y(n_211) );
BUFx12f_ASAP7_75t_L g212 ( .A(n_172), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_166), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_184), .A2(n_161), .B(n_158), .Y(n_214) );
NOR3xp33_ASAP7_75t_L g215 ( .A(n_178), .B(n_161), .C(n_158), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_166), .Y(n_216) );
NOR2x1_ASAP7_75t_R g217 ( .A(n_185), .B(n_7), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_166), .Y(n_218) );
OR2x2_ASAP7_75t_L g219 ( .A(n_185), .B(n_7), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_164), .B(n_8), .Y(n_220) );
OAI22xp5_ASAP7_75t_L g221 ( .A1(n_175), .A2(n_129), .B1(n_117), .B2(n_116), .Y(n_221) );
HB1xp67_ASAP7_75t_L g222 ( .A(n_175), .Y(n_222) );
BUFx2_ASAP7_75t_L g223 ( .A(n_172), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_165), .A2(n_161), .B(n_158), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_167), .A2(n_146), .B(n_125), .Y(n_225) );
NAND2x1_ASAP7_75t_L g226 ( .A(n_171), .B(n_152), .Y(n_226) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_169), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_178), .B(n_8), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_198), .A2(n_189), .B(n_176), .Y(n_229) );
NAND2x1_ASAP7_75t_L g230 ( .A(n_197), .B(n_169), .Y(n_230) );
OAI21x1_ASAP7_75t_SL g231 ( .A1(n_220), .A2(n_186), .B(n_180), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_227), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_199), .B(n_173), .Y(n_233) );
OAI22xp5_ASAP7_75t_L g234 ( .A1(n_201), .A2(n_179), .B1(n_180), .B2(n_186), .Y(n_234) );
BUFx3_ASAP7_75t_L g235 ( .A(n_202), .Y(n_235) );
BUFx12f_ASAP7_75t_L g236 ( .A(n_212), .Y(n_236) );
NOR2xp33_ASAP7_75t_SL g237 ( .A(n_200), .B(n_179), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_227), .Y(n_238) );
O2A1O1Ixp33_ASAP7_75t_SL g239 ( .A1(n_211), .A2(n_187), .B(n_192), .C(n_191), .Y(n_239) );
OR2x6_ASAP7_75t_L g240 ( .A(n_202), .B(n_186), .Y(n_240) );
AOI221xp5_ASAP7_75t_SL g241 ( .A1(n_207), .A2(n_168), .B1(n_188), .B2(n_182), .C(n_190), .Y(n_241) );
CKINVDCx20_ASAP7_75t_R g242 ( .A(n_200), .Y(n_242) );
OAI21x1_ASAP7_75t_L g243 ( .A1(n_206), .A2(n_182), .B(n_180), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_L g244 ( .A1(n_228), .A2(n_171), .B(n_190), .C(n_195), .Y(n_244) );
BUFx6f_ASAP7_75t_L g245 ( .A(n_227), .Y(n_245) );
AOI22xp5_ASAP7_75t_L g246 ( .A1(n_199), .A2(n_171), .B1(n_190), .B2(n_194), .Y(n_246) );
BUFx3_ASAP7_75t_L g247 ( .A(n_227), .Y(n_247) );
NOR2xp33_ASAP7_75t_SL g248 ( .A(n_217), .B(n_171), .Y(n_248) );
INVx1_ASAP7_75t_SL g249 ( .A(n_205), .Y(n_249) );
A2O1A1Ixp33_ASAP7_75t_L g250 ( .A1(n_228), .A2(n_194), .B(n_125), .C(n_129), .Y(n_250) );
AO21x2_ASAP7_75t_L g251 ( .A1(n_215), .A2(n_194), .B(n_146), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_223), .B(n_9), .Y(n_252) );
BUFx4f_ASAP7_75t_L g253 ( .A(n_201), .Y(n_253) );
A2O1A1Ixp33_ASAP7_75t_L g254 ( .A1(n_208), .A2(n_125), .B(n_117), .C(n_13), .Y(n_254) );
OAI22xp33_ASAP7_75t_L g255 ( .A1(n_219), .A2(n_11), .B1(n_12), .B2(n_13), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_253), .B(n_222), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_243), .Y(n_257) );
A2O1A1Ixp33_ASAP7_75t_L g258 ( .A1(n_254), .A2(n_215), .B(n_225), .C(n_222), .Y(n_258) );
BUFx3_ASAP7_75t_L g259 ( .A(n_253), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_239), .A2(n_214), .B(n_224), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_233), .B(n_216), .Y(n_261) );
OAI221xp5_ASAP7_75t_L g262 ( .A1(n_248), .A2(n_209), .B1(n_218), .B2(n_203), .C(n_204), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_230), .Y(n_263) );
AOI22xp33_ASAP7_75t_SL g264 ( .A1(n_237), .A2(n_221), .B1(n_213), .B2(n_196), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_239), .A2(n_210), .B(n_204), .Y(n_265) );
AOI221xp5_ASAP7_75t_L g266 ( .A1(n_255), .A2(n_203), .B1(n_209), .B2(n_210), .C(n_226), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g267 ( .A1(n_252), .A2(n_152), .B1(n_14), .B2(n_15), .Y(n_267) );
INVx3_ASAP7_75t_L g268 ( .A(n_247), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_241), .B(n_11), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_234), .B(n_246), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_229), .A2(n_152), .B(n_43), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_249), .B(n_14), .Y(n_272) );
OAI22xp5_ASAP7_75t_L g273 ( .A1(n_254), .A2(n_15), .B1(n_152), .B2(n_18), .Y(n_273) );
OAI21x1_ASAP7_75t_L g274 ( .A1(n_243), .A2(n_231), .B(n_232), .Y(n_274) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_242), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_244), .A2(n_152), .B(n_19), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_250), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_257), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_269), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_269), .Y(n_280) );
INVx3_ASAP7_75t_L g281 ( .A(n_274), .Y(n_281) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_257), .Y(n_282) );
AOI21xp5_ASAP7_75t_SL g283 ( .A1(n_273), .A2(n_250), .B(n_240), .Y(n_283) );
OR2x2_ASAP7_75t_L g284 ( .A(n_270), .B(n_240), .Y(n_284) );
INVx3_ASAP7_75t_L g285 ( .A(n_274), .Y(n_285) );
INVx3_ASAP7_75t_L g286 ( .A(n_268), .Y(n_286) );
OA21x2_ASAP7_75t_L g287 ( .A1(n_260), .A2(n_238), .B(n_232), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_261), .B(n_251), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_277), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_261), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_277), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_263), .Y(n_292) );
INVx3_ASAP7_75t_L g293 ( .A(n_268), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_263), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_270), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_268), .Y(n_296) );
OR2x2_ASAP7_75t_L g297 ( .A(n_256), .B(n_240), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g298 ( .A1(n_273), .A2(n_235), .B1(n_251), .B2(n_242), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_259), .Y(n_299) );
AOI22xp5_ASAP7_75t_L g300 ( .A1(n_295), .A2(n_267), .B1(n_256), .B2(n_259), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_278), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_288), .B(n_258), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_288), .B(n_247), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_292), .Y(n_304) );
HB1xp67_ASAP7_75t_L g305 ( .A(n_299), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_288), .B(n_238), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_290), .B(n_259), .Y(n_307) );
BUFx2_ASAP7_75t_L g308 ( .A(n_282), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_278), .Y(n_309) );
INVx5_ASAP7_75t_SL g310 ( .A(n_299), .Y(n_310) );
BUFx2_ASAP7_75t_L g311 ( .A(n_282), .Y(n_311) );
BUFx2_ASAP7_75t_L g312 ( .A(n_278), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_281), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_292), .Y(n_314) );
AND2x4_ASAP7_75t_L g315 ( .A(n_294), .B(n_265), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_290), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_295), .B(n_245), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_294), .Y(n_318) );
AO22x1_ASAP7_75t_L g319 ( .A1(n_279), .A2(n_275), .B1(n_235), .B2(n_272), .Y(n_319) );
AOI221xp5_ASAP7_75t_L g320 ( .A1(n_279), .A2(n_262), .B1(n_266), .B2(n_271), .C(n_276), .Y(n_320) );
INVx2_ASAP7_75t_SL g321 ( .A(n_299), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_289), .Y(n_322) );
NOR2x1_ASAP7_75t_L g323 ( .A(n_283), .B(n_245), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_289), .B(n_245), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_289), .B(n_245), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_291), .Y(n_326) );
INVx2_ASAP7_75t_L g327 ( .A(n_281), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_284), .Y(n_328) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_297), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_302), .B(n_291), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_304), .Y(n_331) );
AND2x4_ASAP7_75t_L g332 ( .A(n_315), .B(n_281), .Y(n_332) );
INVx2_ASAP7_75t_SL g333 ( .A(n_308), .Y(n_333) );
OAI211xp5_ASAP7_75t_L g334 ( .A1(n_300), .A2(n_298), .B(n_284), .C(n_280), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_302), .B(n_291), .Y(n_335) );
NAND2x1_ASAP7_75t_L g336 ( .A(n_323), .B(n_281), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_304), .Y(n_337) );
BUFx3_ASAP7_75t_L g338 ( .A(n_308), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_301), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_306), .B(n_280), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_301), .Y(n_341) );
NAND2xp5_ASAP7_75t_SL g342 ( .A(n_310), .B(n_298), .Y(n_342) );
BUFx2_ASAP7_75t_L g343 ( .A(n_311), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_306), .B(n_281), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_316), .B(n_236), .Y(n_345) );
INVx1_ASAP7_75t_SL g346 ( .A(n_311), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_309), .Y(n_347) );
BUFx2_ASAP7_75t_L g348 ( .A(n_312), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_314), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_328), .B(n_284), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_307), .B(n_296), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_314), .Y(n_352) );
AND2x4_ASAP7_75t_L g353 ( .A(n_315), .B(n_285), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_303), .B(n_285), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_318), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_303), .B(n_285), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_318), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_312), .B(n_285), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_322), .B(n_296), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_322), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_307), .B(n_296), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_326), .Y(n_362) );
OAI21xp33_ASAP7_75t_L g363 ( .A1(n_321), .A2(n_264), .B(n_297), .Y(n_363) );
NAND2xp5_ASAP7_75t_SL g364 ( .A(n_310), .B(n_293), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_326), .B(n_287), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_309), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_305), .B(n_287), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_313), .Y(n_368) );
AND2x4_ASAP7_75t_L g369 ( .A(n_315), .B(n_293), .Y(n_369) );
NAND2x1p5_ASAP7_75t_L g370 ( .A(n_321), .B(n_293), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_313), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_317), .B(n_287), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_327), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_317), .B(n_287), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_340), .B(n_329), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_339), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_331), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_331), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_344), .B(n_327), .Y(n_379) );
INVxp67_ASAP7_75t_L g380 ( .A(n_345), .Y(n_380) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_343), .Y(n_381) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_342), .A2(n_297), .B1(n_320), .B2(n_286), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_339), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_350), .B(n_236), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_346), .B(n_310), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_344), .B(n_325), .Y(n_386) );
NOR2x1_ASAP7_75t_L g387 ( .A(n_364), .B(n_293), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_354), .B(n_325), .Y(n_388) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_343), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_337), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_354), .B(n_324), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_337), .Y(n_392) );
AOI22xp5_ASAP7_75t_L g393 ( .A1(n_363), .A2(n_319), .B1(n_310), .B2(n_286), .Y(n_393) );
NOR2x1p5_ASAP7_75t_L g394 ( .A(n_338), .B(n_286), .Y(n_394) );
OR2x2_ASAP7_75t_L g395 ( .A(n_333), .B(n_319), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_349), .Y(n_396) );
NOR2xp33_ASAP7_75t_L g397 ( .A(n_351), .B(n_286), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_339), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_356), .B(n_324), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_363), .A2(n_287), .B1(n_22), .B2(n_24), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_341), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_340), .B(n_17), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_330), .B(n_25), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_356), .B(n_26), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_372), .B(n_27), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_349), .Y(n_406) );
AND2x4_ASAP7_75t_L g407 ( .A(n_332), .B(n_29), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_330), .B(n_30), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_341), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_352), .Y(n_410) );
OR2x2_ASAP7_75t_L g411 ( .A(n_333), .B(n_31), .Y(n_411) );
NOR2xp67_ASAP7_75t_L g412 ( .A(n_338), .B(n_33), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_352), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_372), .B(n_35), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_355), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_355), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_357), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_357), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_335), .B(n_37), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_360), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_374), .B(n_38), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_341), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_360), .Y(n_423) );
OR2x2_ASAP7_75t_L g424 ( .A(n_335), .B(n_42), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_362), .B(n_44), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_374), .B(n_46), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_390), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_390), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_392), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_392), .Y(n_430) );
NAND2xp33_ASAP7_75t_SL g431 ( .A(n_394), .B(n_348), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_406), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_375), .B(n_348), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_406), .Y(n_434) );
NAND4xp25_ASAP7_75t_SL g435 ( .A(n_382), .B(n_334), .C(n_361), .D(n_367), .Y(n_435) );
NAND2x1_ASAP7_75t_L g436 ( .A(n_393), .B(n_362), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_416), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_388), .B(n_338), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_388), .B(n_358), .Y(n_439) );
INVx1_ASAP7_75t_SL g440 ( .A(n_385), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_376), .Y(n_441) );
OAI21xp5_ASAP7_75t_L g442 ( .A1(n_412), .A2(n_370), .B(n_336), .Y(n_442) );
OR2x2_ASAP7_75t_L g443 ( .A(n_381), .B(n_367), .Y(n_443) );
BUFx3_ASAP7_75t_L g444 ( .A(n_385), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_391), .B(n_358), .Y(n_445) );
OR2x2_ASAP7_75t_L g446 ( .A(n_389), .B(n_366), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_416), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_420), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_391), .B(n_332), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_377), .B(n_365), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_376), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_386), .B(n_366), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_420), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_399), .B(n_369), .Y(n_454) );
INVx1_ASAP7_75t_SL g455 ( .A(n_405), .Y(n_455) );
INVx3_ASAP7_75t_L g456 ( .A(n_395), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_378), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_396), .Y(n_458) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_383), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_399), .B(n_332), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_410), .B(n_365), .Y(n_461) );
INVx2_ASAP7_75t_SL g462 ( .A(n_395), .Y(n_462) );
INVxp67_ASAP7_75t_L g463 ( .A(n_405), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_386), .B(n_347), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_379), .B(n_332), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_413), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_415), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_417), .Y(n_468) );
OAI22xp5_ASAP7_75t_L g469 ( .A1(n_380), .A2(n_370), .B1(n_369), .B2(n_336), .Y(n_469) );
INVx2_ASAP7_75t_SL g470 ( .A(n_387), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_418), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_431), .A2(n_426), .B(n_421), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_446), .Y(n_473) );
OAI21xp33_ASAP7_75t_L g474 ( .A1(n_435), .A2(n_384), .B(n_421), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_452), .Y(n_475) );
AOI22xp5_ASAP7_75t_L g476 ( .A1(n_463), .A2(n_397), .B1(n_379), .B2(n_426), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_450), .B(n_423), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_461), .B(n_383), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_427), .Y(n_479) );
INVx1_ASAP7_75t_SL g480 ( .A(n_438), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_462), .B(n_401), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_428), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_429), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_431), .B(n_407), .Y(n_484) );
OAI22xp5_ASAP7_75t_L g485 ( .A1(n_463), .A2(n_424), .B1(n_411), .B2(n_407), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_430), .Y(n_486) );
OAI22xp5_ASAP7_75t_L g487 ( .A1(n_455), .A2(n_424), .B1(n_411), .B2(n_407), .Y(n_487) );
INVxp67_ASAP7_75t_L g488 ( .A(n_462), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_439), .B(n_401), .Y(n_489) );
INVx1_ASAP7_75t_SL g490 ( .A(n_440), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_432), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g492 ( .A1(n_436), .A2(n_414), .B(n_404), .C(n_402), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_434), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_439), .B(n_398), .Y(n_494) );
OAI21xp33_ASAP7_75t_SL g495 ( .A1(n_470), .A2(n_414), .B(n_404), .Y(n_495) );
O2A1O1Ixp33_ASAP7_75t_SL g496 ( .A1(n_469), .A2(n_403), .B(n_419), .C(n_408), .Y(n_496) );
AOI221xp5_ASAP7_75t_L g497 ( .A1(n_456), .A2(n_400), .B1(n_425), .B2(n_409), .C(n_422), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_437), .Y(n_498) );
AOI21xp33_ASAP7_75t_L g499 ( .A1(n_470), .A2(n_353), .B(n_369), .Y(n_499) );
INVxp33_ASAP7_75t_L g500 ( .A(n_433), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_447), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_479), .Y(n_502) );
NAND3xp33_ASAP7_75t_SL g503 ( .A(n_474), .B(n_484), .C(n_472), .Y(n_503) );
AOI32xp33_ASAP7_75t_L g504 ( .A1(n_495), .A2(n_456), .A3(n_444), .B1(n_449), .B2(n_460), .Y(n_504) );
OAI221xp5_ASAP7_75t_L g505 ( .A1(n_484), .A2(n_456), .B1(n_444), .B2(n_443), .C(n_442), .Y(n_505) );
NOR2x1_ASAP7_75t_L g506 ( .A(n_492), .B(n_471), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_496), .A2(n_459), .B(n_449), .Y(n_507) );
OAI21xp33_ASAP7_75t_L g508 ( .A1(n_500), .A2(n_460), .B(n_465), .Y(n_508) );
NOR3xp33_ASAP7_75t_L g509 ( .A(n_497), .B(n_468), .C(n_467), .Y(n_509) );
AOI221xp5_ASAP7_75t_L g510 ( .A1(n_488), .A2(n_466), .B1(n_457), .B2(n_458), .C(n_445), .Y(n_510) );
NAND4xp25_ASAP7_75t_L g511 ( .A(n_499), .B(n_369), .C(n_353), .D(n_454), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_480), .B(n_465), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_473), .B(n_445), .Y(n_513) );
OAI22xp33_ASAP7_75t_L g514 ( .A1(n_485), .A2(n_464), .B1(n_459), .B2(n_370), .Y(n_514) );
NOR3x1_ASAP7_75t_L g515 ( .A(n_487), .B(n_453), .C(n_448), .Y(n_515) );
AO22x1_ASAP7_75t_L g516 ( .A1(n_488), .A2(n_451), .B1(n_441), .B2(n_353), .Y(n_516) );
AOI211xp5_ASAP7_75t_SL g517 ( .A1(n_476), .A2(n_353), .B(n_359), .C(n_451), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_482), .Y(n_518) );
AOI221xp5_ASAP7_75t_L g519 ( .A1(n_503), .A2(n_490), .B1(n_477), .B2(n_475), .C(n_493), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g520 ( .A1(n_511), .A2(n_501), .B1(n_498), .B2(n_483), .Y(n_520) );
OAI211xp5_ASAP7_75t_L g521 ( .A1(n_504), .A2(n_481), .B(n_489), .C(n_494), .Y(n_521) );
OAI211xp5_ASAP7_75t_SL g522 ( .A1(n_505), .A2(n_491), .B(n_486), .C(n_478), .Y(n_522) );
AOI221xp5_ASAP7_75t_L g523 ( .A1(n_510), .A2(n_441), .B1(n_422), .B2(n_409), .C(n_398), .Y(n_523) );
OR2x2_ASAP7_75t_L g524 ( .A(n_513), .B(n_373), .Y(n_524) );
AOI221xp5_ASAP7_75t_L g525 ( .A1(n_514), .A2(n_359), .B1(n_371), .B2(n_373), .C(n_368), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_509), .B(n_373), .Y(n_526) );
AOI22xp5_ASAP7_75t_L g527 ( .A1(n_506), .A2(n_508), .B1(n_507), .B2(n_518), .Y(n_527) );
NOR3xp33_ASAP7_75t_L g528 ( .A(n_519), .B(n_516), .C(n_502), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_520), .B(n_515), .Y(n_529) );
OR5x1_ASAP7_75t_L g530 ( .A(n_522), .B(n_517), .C(n_512), .D(n_50), .E(n_51), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g531 ( .A(n_527), .B(n_517), .Y(n_531) );
A2O1A1Ixp33_ASAP7_75t_L g532 ( .A1(n_521), .A2(n_371), .B(n_368), .C(n_347), .Y(n_532) );
NAND3xp33_ASAP7_75t_L g533 ( .A(n_531), .B(n_525), .C(n_523), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_529), .B(n_526), .Y(n_534) );
AND3x4_ASAP7_75t_L g535 ( .A(n_528), .B(n_524), .C(n_371), .Y(n_535) );
NOR3xp33_ASAP7_75t_SL g536 ( .A(n_533), .B(n_532), .C(n_530), .Y(n_536) );
NAND4xp25_ASAP7_75t_L g537 ( .A(n_534), .B(n_347), .C(n_49), .D(n_52), .Y(n_537) );
XNOR2xp5_ASAP7_75t_L g538 ( .A(n_536), .B(n_537), .Y(n_538) );
INVx1_ASAP7_75t_SL g539 ( .A(n_538), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_539), .B(n_535), .Y(n_540) );
AOI22x1_ASAP7_75t_L g541 ( .A1(n_540), .A2(n_48), .B1(n_54), .B2(n_57), .Y(n_541) );
OAI31xp33_ASAP7_75t_L g542 ( .A1(n_541), .A2(n_74), .A3(n_61), .B(n_62), .Y(n_542) );
OAI221xp5_ASAP7_75t_L g543 ( .A1(n_542), .A2(n_58), .B1(n_64), .B2(n_67), .C(n_68), .Y(n_543) );
endmodule