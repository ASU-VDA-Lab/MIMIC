module fake_netlist_6_1167_n_1945 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1945);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1945;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_268;
wire n_1760;
wire n_1927;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1848;
wire n_763;
wire n_1147;
wire n_1785;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_827;
wire n_531;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_81),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_66),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_115),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_124),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_162),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_141),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_174),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_18),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_86),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_189),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_28),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_87),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_56),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_127),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_16),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_4),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_56),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_16),
.Y(n_212)
);

BUFx10_ASAP7_75t_L g213 ( 
.A(n_143),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_31),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_106),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_163),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_180),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_35),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_120),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_102),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_76),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_107),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_11),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_129),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_1),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_42),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_175),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_32),
.Y(n_228)
);

BUFx10_ASAP7_75t_L g229 ( 
.A(n_73),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_193),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_6),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_68),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_50),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_74),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_172),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_80),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_85),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_118),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_105),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_146),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_156),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_99),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_12),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_89),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_170),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_190),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_157),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_114),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_55),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_48),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_3),
.Y(n_251)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_21),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_131),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_109),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_154),
.Y(n_255)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_84),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_44),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_184),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_179),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_128),
.Y(n_260)
);

BUFx5_ASAP7_75t_L g261 ( 
.A(n_50),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_33),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_192),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_45),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_165),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_19),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_8),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_123),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_31),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_37),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_69),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_71),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_98),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_149),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_14),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_60),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_13),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_104),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_153),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_49),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_138),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_52),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_72),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_11),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_158),
.Y(n_285)
);

BUFx10_ASAP7_75t_L g286 ( 
.A(n_125),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_91),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_20),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_187),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_92),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_95),
.Y(n_291)
);

BUFx10_ASAP7_75t_L g292 ( 
.A(n_37),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_67),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_22),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_150),
.Y(n_295)
);

BUFx2_ASAP7_75t_L g296 ( 
.A(n_24),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_151),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_185),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_10),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_164),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_194),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_155),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_34),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_5),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_15),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_168),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_88),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_161),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_7),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_182),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_43),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_113),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_70),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_110),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_160),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_173),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_41),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_100),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_101),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_94),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_22),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_7),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_167),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_142),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_108),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_58),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_32),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_169),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_1),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_54),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_116),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_36),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_178),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_61),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_83),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_111),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_35),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_134),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_96),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_119),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_97),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_171),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_77),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_21),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_47),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_52),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_188),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_36),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_45),
.Y(n_349)
);

INVx2_ASAP7_75t_SL g350 ( 
.A(n_57),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_40),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_112),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_117),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_18),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_26),
.Y(n_355)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_177),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_191),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_135),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g359 ( 
.A(n_6),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_2),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_20),
.Y(n_361)
);

INVx2_ASAP7_75t_SL g362 ( 
.A(n_24),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_30),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_103),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_183),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_126),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_57),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_75),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_39),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_44),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_63),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_51),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_121),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_147),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_90),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_9),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_8),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_54),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_65),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_34),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_4),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_148),
.Y(n_382)
);

INVx1_ASAP7_75t_SL g383 ( 
.A(n_49),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_139),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_30),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_181),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_51),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_93),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_122),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_39),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_195),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_284),
.B(n_0),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_296),
.Y(n_393)
);

INVxp33_ASAP7_75t_L g394 ( 
.A(n_296),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_261),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_199),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_261),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_227),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_204),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_261),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_261),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_200),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_261),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_204),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_245),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_261),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_206),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_261),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_205),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_290),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_261),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_208),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_310),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_261),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_326),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_338),
.Y(n_416)
);

CKINVDCx16_ASAP7_75t_R g417 ( 
.A(n_240),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_216),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_382),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_220),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_326),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_326),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_222),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_224),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_326),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_326),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_278),
.B(n_246),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_232),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_202),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_250),
.Y(n_430)
);

INVxp67_ASAP7_75t_SL g431 ( 
.A(n_313),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_237),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_238),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_241),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_250),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_262),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_262),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_242),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_244),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_278),
.B(n_0),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_247),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_248),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_351),
.Y(n_443)
);

INVxp67_ASAP7_75t_SL g444 ( 
.A(n_253),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_255),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_351),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_258),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_259),
.Y(n_448)
);

INVxp67_ASAP7_75t_SL g449 ( 
.A(n_253),
.Y(n_449)
);

INVxp67_ASAP7_75t_SL g450 ( 
.A(n_256),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_263),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_265),
.Y(n_452)
);

INVxp67_ASAP7_75t_SL g453 ( 
.A(n_256),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_390),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_196),
.B(n_2),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_274),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_205),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_390),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_385),
.Y(n_459)
);

NOR2xp67_ASAP7_75t_L g460 ( 
.A(n_350),
.B(n_3),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_279),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_281),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_292),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_283),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_385),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_385),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_212),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_246),
.B(n_306),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_287),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g470 ( 
.A(n_212),
.Y(n_470)
);

INVxp67_ASAP7_75t_SL g471 ( 
.A(n_324),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_293),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_214),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_295),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_297),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_298),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_302),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_307),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_196),
.B(n_5),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_308),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_214),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_218),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_218),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_315),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_197),
.B(n_9),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_319),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_325),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_225),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_460),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_401),
.Y(n_490)
);

AND2x6_ASAP7_75t_L g491 ( 
.A(n_395),
.B(n_254),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_401),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_415),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_415),
.Y(n_494)
);

INVx2_ASAP7_75t_SL g495 ( 
.A(n_399),
.Y(n_495)
);

INVx5_ASAP7_75t_L g496 ( 
.A(n_399),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_421),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_427),
.B(n_350),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_421),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_422),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_395),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_397),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_397),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_400),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_391),
.B(n_215),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_400),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_422),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_403),
.Y(n_508)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_444),
.B(n_252),
.Y(n_509)
);

OAI21x1_ASAP7_75t_L g510 ( 
.A1(n_403),
.A2(n_203),
.B(n_201),
.Y(n_510)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_425),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_449),
.B(n_389),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_396),
.B(n_402),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_406),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_406),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_450),
.B(n_252),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_425),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_408),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_408),
.Y(n_519)
);

INVx1_ASAP7_75t_SL g520 ( 
.A(n_398),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_426),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_411),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_411),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_453),
.B(n_328),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_414),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_414),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_426),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_467),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_417),
.B(n_213),
.Y(n_529)
);

BUFx8_ASAP7_75t_L g530 ( 
.A(n_404),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_430),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_430),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_435),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_435),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_436),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_467),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_471),
.B(n_331),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_436),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_405),
.Y(n_539)
);

INVxp67_ASAP7_75t_L g540 ( 
.A(n_429),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_437),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_482),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_482),
.Y(n_543)
);

OA21x2_ASAP7_75t_L g544 ( 
.A1(n_437),
.A2(n_198),
.B(n_197),
.Y(n_544)
);

AND2x4_ASAP7_75t_L g545 ( 
.A(n_459),
.B(n_246),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_459),
.B(n_333),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_483),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_483),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_465),
.B(n_306),
.Y(n_549)
);

BUFx3_ASAP7_75t_L g550 ( 
.A(n_404),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_465),
.B(n_306),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_488),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_417),
.B(n_463),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_488),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_466),
.B(n_339),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_443),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_410),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_443),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_446),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_446),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_454),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_454),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_458),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_458),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_466),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_SL g566 ( 
.A(n_440),
.B(n_292),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_468),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_501),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_567),
.B(n_407),
.Y(n_569)
);

BUFx4f_ASAP7_75t_L g570 ( 
.A(n_544),
.Y(n_570)
);

INVx4_ASAP7_75t_L g571 ( 
.A(n_496),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_490),
.Y(n_572)
);

INVx2_ASAP7_75t_SL g573 ( 
.A(n_489),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_567),
.B(n_431),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_505),
.B(n_412),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_565),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_550),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_L g578 ( 
.A1(n_567),
.A2(n_392),
.B1(n_479),
.B2(n_455),
.Y(n_578)
);

BUFx4f_ASAP7_75t_L g579 ( 
.A(n_544),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_490),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_501),
.Y(n_581)
);

AND2x4_ASAP7_75t_L g582 ( 
.A(n_545),
.B(n_549),
.Y(n_582)
);

INVxp33_ASAP7_75t_L g583 ( 
.A(n_509),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_489),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_490),
.Y(n_585)
);

BUFx10_ASAP7_75t_L g586 ( 
.A(n_513),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_501),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_509),
.B(n_516),
.Y(n_588)
);

INVx2_ASAP7_75t_SL g589 ( 
.A(n_550),
.Y(n_589)
);

BUFx4f_ASAP7_75t_L g590 ( 
.A(n_544),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_566),
.B(n_418),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_516),
.B(n_394),
.Y(n_592)
);

INVx2_ASAP7_75t_SL g593 ( 
.A(n_550),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_504),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_565),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_502),
.Y(n_596)
);

BUFx10_ASAP7_75t_L g597 ( 
.A(n_545),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_504),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_504),
.Y(n_599)
);

NAND3xp33_ASAP7_75t_L g600 ( 
.A(n_566),
.B(n_393),
.C(n_420),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_490),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_512),
.B(n_423),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_540),
.B(n_424),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_508),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_545),
.B(n_409),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_490),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_524),
.B(n_428),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_490),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_508),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_498),
.A2(n_485),
.B1(n_460),
.B2(n_362),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_490),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_540),
.B(n_432),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_508),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_498),
.Y(n_614)
);

INVx8_ASAP7_75t_L g615 ( 
.A(n_545),
.Y(n_615)
);

INVx2_ASAP7_75t_SL g616 ( 
.A(n_495),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_502),
.Y(n_617)
);

BUFx2_ASAP7_75t_L g618 ( 
.A(n_495),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_502),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_502),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_492),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_506),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_514),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_514),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_524),
.B(n_433),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_537),
.B(n_434),
.Y(n_626)
);

INVx2_ASAP7_75t_SL g627 ( 
.A(n_495),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_530),
.B(n_439),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_514),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_539),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_530),
.B(n_441),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_537),
.B(n_445),
.Y(n_632)
);

INVxp67_ASAP7_75t_L g633 ( 
.A(n_529),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_530),
.B(n_447),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_530),
.B(n_448),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_515),
.Y(n_636)
);

INVx4_ASAP7_75t_L g637 ( 
.A(n_496),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_515),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_546),
.B(n_451),
.Y(n_639)
);

OAI21xp33_ASAP7_75t_SL g640 ( 
.A1(n_510),
.A2(n_362),
.B(n_359),
.Y(n_640)
);

NAND2x1p5_ASAP7_75t_L g641 ( 
.A(n_544),
.B(n_324),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_492),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_492),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_492),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_515),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_523),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_546),
.B(n_456),
.Y(n_647)
);

BUFx2_ASAP7_75t_L g648 ( 
.A(n_555),
.Y(n_648)
);

BUFx4f_ASAP7_75t_L g649 ( 
.A(n_544),
.Y(n_649)
);

BUFx4f_ASAP7_75t_L g650 ( 
.A(n_503),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_523),
.Y(n_651)
);

AND2x6_ASAP7_75t_L g652 ( 
.A(n_506),
.B(n_201),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_492),
.Y(n_653)
);

BUFx8_ASAP7_75t_SL g654 ( 
.A(n_557),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_523),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_526),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_526),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_526),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_559),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_520),
.Y(n_660)
);

INVx4_ASAP7_75t_L g661 ( 
.A(n_496),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_555),
.B(n_464),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_559),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_506),
.B(n_469),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_492),
.Y(n_665)
);

OAI22xp33_ASAP7_75t_L g666 ( 
.A1(n_553),
.A2(n_463),
.B1(n_383),
.B2(n_228),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_549),
.B(n_551),
.Y(n_667)
);

BUFx6f_ASAP7_75t_SL g668 ( 
.A(n_549),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_549),
.B(n_474),
.Y(n_669)
);

NAND2xp33_ASAP7_75t_SL g670 ( 
.A(n_551),
.B(n_359),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_506),
.Y(n_671)
);

INVx5_ASAP7_75t_L g672 ( 
.A(n_491),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_492),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_559),
.Y(n_674)
);

INVx4_ASAP7_75t_L g675 ( 
.A(n_496),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_519),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_559),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_559),
.Y(n_678)
);

AND2x4_ASAP7_75t_L g679 ( 
.A(n_551),
.B(n_341),
.Y(n_679)
);

NAND2xp33_ASAP7_75t_L g680 ( 
.A(n_491),
.B(n_254),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_519),
.B(n_475),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_551),
.B(n_477),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_559),
.Y(n_683)
);

OAI21xp33_ASAP7_75t_SL g684 ( 
.A1(n_510),
.A2(n_219),
.B(n_198),
.Y(n_684)
);

AND3x1_ASAP7_75t_L g685 ( 
.A(n_528),
.B(n_231),
.C(n_225),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_503),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_519),
.B(n_478),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_519),
.B(n_480),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_522),
.B(n_484),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_522),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_522),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_522),
.B(n_486),
.Y(n_692)
);

INVx4_ASAP7_75t_L g693 ( 
.A(n_496),
.Y(n_693)
);

INVxp33_ASAP7_75t_SL g694 ( 
.A(n_520),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_496),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_493),
.Y(n_696)
);

INVx3_ASAP7_75t_L g697 ( 
.A(n_503),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_494),
.Y(n_698)
);

INVx5_ASAP7_75t_L g699 ( 
.A(n_491),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_496),
.B(n_487),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_494),
.Y(n_701)
);

NOR2x1p5_ASAP7_75t_L g702 ( 
.A(n_528),
.B(n_376),
.Y(n_702)
);

INVx1_ASAP7_75t_SL g703 ( 
.A(n_536),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_497),
.Y(n_704)
);

INVx1_ASAP7_75t_SL g705 ( 
.A(n_536),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_497),
.Y(n_706)
);

BUFx6f_ASAP7_75t_SL g707 ( 
.A(n_542),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_542),
.B(n_438),
.Y(n_708)
);

BUFx10_ASAP7_75t_L g709 ( 
.A(n_543),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_499),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_543),
.B(n_442),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_503),
.B(n_341),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_547),
.B(n_452),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_547),
.B(n_461),
.Y(n_714)
);

OAI22x1_ASAP7_75t_L g715 ( 
.A1(n_548),
.A2(n_327),
.B1(n_251),
.B2(n_282),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_510),
.Y(n_716)
);

NOR3xp33_ASAP7_75t_L g717 ( 
.A(n_548),
.B(n_470),
.C(n_457),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_667),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_583),
.B(n_462),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_667),
.Y(n_720)
);

NOR3xp33_ASAP7_75t_L g721 ( 
.A(n_666),
.B(n_481),
.C(n_473),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_582),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_602),
.B(n_503),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_607),
.B(n_503),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_648),
.B(n_639),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_701),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_582),
.B(n_503),
.Y(n_727)
);

INVx3_ASAP7_75t_L g728 ( 
.A(n_582),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_701),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_576),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_704),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_576),
.Y(n_732)
);

BUFx8_ASAP7_75t_L g733 ( 
.A(n_707),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_595),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_595),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_615),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_592),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_706),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_706),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_710),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_648),
.B(n_575),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_696),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_588),
.B(n_518),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_588),
.B(n_518),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_696),
.Y(n_745)
);

NOR2xp67_ASAP7_75t_L g746 ( 
.A(n_633),
.B(n_552),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_570),
.B(n_518),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_592),
.B(n_413),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_710),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_573),
.B(n_416),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_698),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_569),
.B(n_573),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_625),
.B(n_518),
.Y(n_753)
);

INVx4_ASAP7_75t_L g754 ( 
.A(n_615),
.Y(n_754)
);

NAND3xp33_ASAP7_75t_L g755 ( 
.A(n_578),
.B(n_476),
.C(n_472),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_626),
.B(n_518),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_698),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_568),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_632),
.B(n_525),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_L g760 ( 
.A1(n_570),
.A2(n_231),
.B1(n_344),
.B2(n_251),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_584),
.B(n_207),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_616),
.B(n_525),
.Y(n_762)
);

INVx2_ASAP7_75t_SL g763 ( 
.A(n_702),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_584),
.B(n_209),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_616),
.B(n_525),
.Y(n_765)
);

NOR3xp33_ASAP7_75t_L g766 ( 
.A(n_600),
.B(n_211),
.C(n_210),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_703),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_568),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_581),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_614),
.B(n_226),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_627),
.B(n_525),
.Y(n_771)
);

OAI22xp5_ASAP7_75t_L g772 ( 
.A1(n_614),
.A2(n_419),
.B1(n_300),
.B2(n_285),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_627),
.B(n_525),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_705),
.B(n_618),
.Y(n_774)
);

OR2x2_ASAP7_75t_L g775 ( 
.A(n_711),
.B(n_552),
.Y(n_775)
);

BUFx6f_ASAP7_75t_SL g776 ( 
.A(n_586),
.Y(n_776)
);

O2A1O1Ixp33_ASAP7_75t_L g777 ( 
.A1(n_640),
.A2(n_554),
.B(n_355),
.C(n_311),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_581),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_570),
.B(n_525),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_587),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_618),
.B(n_525),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_SL g782 ( 
.A(n_694),
.B(n_660),
.Y(n_782)
);

OAI221xp5_ASAP7_75t_L g783 ( 
.A1(n_610),
.A2(n_299),
.B1(n_329),
.B2(n_321),
.C(n_311),
.Y(n_783)
);

BUFx12f_ASAP7_75t_SL g784 ( 
.A(n_574),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_574),
.B(n_554),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_647),
.B(n_233),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_664),
.B(n_499),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_587),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_671),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_671),
.Y(n_790)
);

INVx1_ASAP7_75t_SL g791 ( 
.A(n_660),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_662),
.B(n_243),
.Y(n_792)
);

INVx2_ASAP7_75t_SL g793 ( 
.A(n_709),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_579),
.B(n_254),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_681),
.B(n_500),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_594),
.Y(n_796)
);

HB1xp67_ASAP7_75t_L g797 ( 
.A(n_715),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_690),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_687),
.B(n_500),
.Y(n_799)
);

AND2x2_ASAP7_75t_L g800 ( 
.A(n_605),
.B(n_556),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_594),
.Y(n_801)
);

OR2x6_ASAP7_75t_L g802 ( 
.A(n_628),
.B(n_376),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_688),
.B(n_507),
.Y(n_803)
);

OR2x2_ASAP7_75t_L g804 ( 
.A(n_714),
.B(n_708),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_689),
.B(n_507),
.Y(n_805)
);

AND2x6_ASAP7_75t_L g806 ( 
.A(n_690),
.B(n_219),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_692),
.B(n_517),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_598),
.Y(n_808)
);

NAND2xp33_ASAP7_75t_L g809 ( 
.A(n_641),
.B(n_254),
.Y(n_809)
);

OR2x6_ASAP7_75t_L g810 ( 
.A(n_631),
.B(n_634),
.Y(n_810)
);

NAND3xp33_ASAP7_75t_L g811 ( 
.A(n_713),
.B(n_257),
.C(n_249),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_589),
.B(n_593),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_589),
.B(n_517),
.Y(n_813)
);

AND2x4_ASAP7_75t_L g814 ( 
.A(n_593),
.B(n_356),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_579),
.B(n_254),
.Y(n_815)
);

OR2x2_ASAP7_75t_L g816 ( 
.A(n_603),
.B(n_264),
.Y(n_816)
);

INVx1_ASAP7_75t_SL g817 ( 
.A(n_694),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_579),
.A2(n_299),
.B1(n_329),
.B2(n_321),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_691),
.B(n_682),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_591),
.B(n_267),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_590),
.B(n_272),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_654),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_691),
.Y(n_823)
);

INVx3_ASAP7_75t_L g824 ( 
.A(n_597),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_590),
.B(n_272),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_709),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_598),
.Y(n_827)
);

INVx3_ASAP7_75t_L g828 ( 
.A(n_597),
.Y(n_828)
);

O2A1O1Ixp33_ASAP7_75t_L g829 ( 
.A1(n_684),
.A2(n_344),
.B(n_282),
.C(n_378),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_709),
.Y(n_830)
);

INVx2_ASAP7_75t_SL g831 ( 
.A(n_679),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_590),
.B(n_272),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_679),
.Y(n_833)
);

AND2x6_ASAP7_75t_L g834 ( 
.A(n_605),
.B(n_221),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_679),
.Y(n_835)
);

INVx2_ASAP7_75t_SL g836 ( 
.A(n_577),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_596),
.B(n_521),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_615),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_649),
.B(n_272),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_617),
.B(n_619),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_620),
.B(n_521),
.Y(n_841)
);

INVx8_ASAP7_75t_L g842 ( 
.A(n_707),
.Y(n_842)
);

INVx2_ASAP7_75t_SL g843 ( 
.A(n_577),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_649),
.B(n_272),
.Y(n_844)
);

BUFx6f_ASAP7_75t_SL g845 ( 
.A(n_586),
.Y(n_845)
);

INVx2_ASAP7_75t_SL g846 ( 
.A(n_669),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_599),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_615),
.Y(n_848)
);

BUFx3_ASAP7_75t_L g849 ( 
.A(n_597),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_599),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_L g851 ( 
.A1(n_649),
.A2(n_354),
.B1(n_355),
.B2(n_360),
.Y(n_851)
);

OAI221xp5_ASAP7_75t_L g852 ( 
.A1(n_670),
.A2(n_360),
.B1(n_354),
.B2(n_372),
.C(n_378),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_612),
.B(n_269),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_622),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_676),
.B(n_707),
.Y(n_855)
);

INVx1_ASAP7_75t_SL g856 ( 
.A(n_630),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_670),
.B(n_586),
.Y(n_857)
);

INVx2_ASAP7_75t_SL g858 ( 
.A(n_715),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_641),
.B(n_527),
.Y(n_859)
);

AOI22xp5_ASAP7_75t_L g860 ( 
.A1(n_668),
.A2(n_352),
.B1(n_353),
.B2(n_357),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_641),
.A2(n_372),
.B1(n_318),
.B2(n_236),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_604),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_604),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_654),
.Y(n_864)
);

NOR2xp67_ASAP7_75t_L g865 ( 
.A(n_635),
.B(n_560),
.Y(n_865)
);

OAI21xp5_ASAP7_75t_L g866 ( 
.A1(n_716),
.A2(n_650),
.B(n_624),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_609),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_609),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_672),
.B(n_203),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_712),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_716),
.B(n_527),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_613),
.Y(n_872)
);

INVxp67_ASAP7_75t_SL g873 ( 
.A(n_572),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_580),
.B(n_601),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_580),
.B(n_560),
.Y(n_875)
);

OR2x2_ASAP7_75t_L g876 ( 
.A(n_630),
.B(n_270),
.Y(n_876)
);

OAI22xp5_ASAP7_75t_L g877 ( 
.A1(n_668),
.A2(n_300),
.B1(n_285),
.B2(n_268),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_613),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_717),
.B(n_556),
.Y(n_879)
);

NOR2xp67_ASAP7_75t_L g880 ( 
.A(n_700),
.B(n_560),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_638),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_623),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_623),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_624),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_638),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_725),
.B(n_629),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_752),
.B(n_672),
.Y(n_887)
);

AOI21x1_ASAP7_75t_L g888 ( 
.A1(n_747),
.A2(n_636),
.B(n_629),
.Y(n_888)
);

INVx4_ASAP7_75t_L g889 ( 
.A(n_736),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_809),
.A2(n_650),
.B(n_601),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_809),
.A2(n_650),
.B(n_601),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_751),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_744),
.A2(n_606),
.B(n_580),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_751),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_794),
.A2(n_611),
.B(n_606),
.Y(n_895)
);

BUFx2_ASAP7_75t_SL g896 ( 
.A(n_817),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_748),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_752),
.B(n_636),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_785),
.B(n_655),
.Y(n_899)
);

O2A1O1Ixp33_ASAP7_75t_L g900 ( 
.A1(n_858),
.A2(n_797),
.B(n_741),
.C(n_743),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_794),
.A2(n_611),
.B(n_606),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_815),
.A2(n_643),
.B(n_611),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_815),
.A2(n_653),
.B(n_643),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_821),
.A2(n_653),
.B(n_643),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_774),
.B(n_672),
.Y(n_905)
);

A2O1A1Ixp33_ASAP7_75t_L g906 ( 
.A1(n_820),
.A2(n_235),
.B(n_230),
.C(n_312),
.Y(n_906)
);

AOI22xp5_ASAP7_75t_L g907 ( 
.A1(n_718),
.A2(n_668),
.B1(n_652),
.B2(n_697),
.Y(n_907)
);

O2A1O1Ixp33_ASAP7_75t_L g908 ( 
.A1(n_743),
.A2(n_680),
.B(n_655),
.C(n_651),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_804),
.B(n_223),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_819),
.B(n_653),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_720),
.Y(n_911)
);

OAI21xp5_ASAP7_75t_L g912 ( 
.A1(n_821),
.A2(n_646),
.B(n_645),
.Y(n_912)
);

OAI22x1_ASAP7_75t_L g913 ( 
.A1(n_791),
.A2(n_330),
.B1(n_294),
.B2(n_288),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_825),
.A2(n_665),
.B(n_646),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_825),
.A2(n_839),
.B(n_832),
.Y(n_915)
);

INVx3_ASAP7_75t_L g916 ( 
.A(n_728),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_789),
.Y(n_917)
);

O2A1O1Ixp33_ASAP7_75t_SL g918 ( 
.A1(n_832),
.A2(n_316),
.B(n_358),
.C(n_364),
.Y(n_918)
);

BUFx4f_ASAP7_75t_L g919 ( 
.A(n_842),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_839),
.A2(n_665),
.B(n_651),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_849),
.Y(n_921)
);

AND2x2_ASAP7_75t_L g922 ( 
.A(n_774),
.B(n_767),
.Y(n_922)
);

O2A1O1Ixp33_ASAP7_75t_L g923 ( 
.A1(n_783),
.A2(n_680),
.B(n_645),
.C(n_657),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_787),
.B(n_665),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_793),
.B(n_672),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_737),
.B(n_672),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_790),
.Y(n_927)
);

AND2x4_ASAP7_75t_L g928 ( 
.A(n_836),
.B(n_685),
.Y(n_928)
);

O2A1O1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_829),
.A2(n_656),
.B(n_657),
.C(n_658),
.Y(n_929)
);

OAI21xp5_ASAP7_75t_L g930 ( 
.A1(n_844),
.A2(n_658),
.B(n_656),
.Y(n_930)
);

OAI21xp5_ASAP7_75t_L g931 ( 
.A1(n_844),
.A2(n_697),
.B(n_686),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_746),
.B(n_699),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_795),
.B(n_686),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_859),
.A2(n_697),
.B(n_686),
.Y(n_934)
);

O2A1O1Ixp33_ASAP7_75t_SL g935 ( 
.A1(n_779),
.A2(n_316),
.B(n_291),
.C(n_301),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_779),
.A2(n_663),
.B(n_659),
.Y(n_936)
);

O2A1O1Ixp33_ASAP7_75t_L g937 ( 
.A1(n_777),
.A2(n_314),
.B(n_343),
.C(n_342),
.Y(n_937)
);

OAI21xp33_ASAP7_75t_L g938 ( 
.A1(n_761),
.A2(n_276),
.B(n_275),
.Y(n_938)
);

AND2x4_ASAP7_75t_L g939 ( 
.A(n_843),
.B(n_558),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_798),
.Y(n_940)
);

OAI21xp5_ASAP7_75t_L g941 ( 
.A1(n_866),
.A2(n_677),
.B(n_674),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_723),
.A2(n_677),
.B(n_674),
.Y(n_942)
);

INVxp67_ASAP7_75t_L g943 ( 
.A(n_782),
.Y(n_943)
);

AOI21x1_ASAP7_75t_L g944 ( 
.A1(n_727),
.A2(n_683),
.B(n_678),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_799),
.B(n_572),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_803),
.B(n_572),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_823),
.Y(n_947)
);

BUFx2_ASAP7_75t_L g948 ( 
.A(n_784),
.Y(n_948)
);

AOI22xp5_ASAP7_75t_L g949 ( 
.A1(n_722),
.A2(n_652),
.B1(n_678),
.B2(n_683),
.Y(n_949)
);

AOI22xp5_ASAP7_75t_L g950 ( 
.A1(n_834),
.A2(n_652),
.B1(n_572),
.B2(n_673),
.Y(n_950)
);

INVx2_ASAP7_75t_SL g951 ( 
.A(n_775),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_849),
.Y(n_952)
);

AO21x1_ASAP7_75t_L g953 ( 
.A1(n_724),
.A2(n_230),
.B(n_221),
.Y(n_953)
);

OAI21xp33_ASAP7_75t_L g954 ( 
.A1(n_761),
.A2(n_280),
.B(n_277),
.Y(n_954)
);

AOI21x1_ASAP7_75t_L g955 ( 
.A1(n_727),
.A2(n_535),
.B(n_534),
.Y(n_955)
);

BUFx12f_ASAP7_75t_L g956 ( 
.A(n_733),
.Y(n_956)
);

OAI21xp33_ASAP7_75t_L g957 ( 
.A1(n_764),
.A2(n_770),
.B(n_853),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_726),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_753),
.A2(n_608),
.B(n_585),
.Y(n_959)
);

BUFx8_ASAP7_75t_L g960 ( 
.A(n_776),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_756),
.A2(n_608),
.B(n_585),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_846),
.B(n_699),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_759),
.A2(n_608),
.B(n_585),
.Y(n_963)
);

OAI21xp33_ASAP7_75t_L g964 ( 
.A1(n_764),
.A2(n_304),
.B(n_303),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_L g965 ( 
.A(n_784),
.B(n_266),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_728),
.Y(n_966)
);

AOI21x1_ASAP7_75t_L g967 ( 
.A1(n_871),
.A2(n_535),
.B(n_534),
.Y(n_967)
);

BUFx3_ASAP7_75t_L g968 ( 
.A(n_733),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_729),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_781),
.A2(n_621),
.B(n_608),
.Y(n_970)
);

INVx4_ASAP7_75t_L g971 ( 
.A(n_736),
.Y(n_971)
);

INVx3_ASAP7_75t_L g972 ( 
.A(n_833),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_805),
.A2(n_642),
.B(n_621),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_719),
.B(n_332),
.Y(n_974)
);

INVx3_ASAP7_75t_L g975 ( 
.A(n_835),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_731),
.Y(n_976)
);

O2A1O1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_760),
.A2(n_314),
.B(n_320),
.C(n_312),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_807),
.B(n_621),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_822),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_800),
.B(n_292),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_826),
.B(n_699),
.Y(n_981)
);

AO21x2_ASAP7_75t_L g982 ( 
.A1(n_870),
.A2(n_236),
.B(n_235),
.Y(n_982)
);

NOR2x1_ASAP7_75t_L g983 ( 
.A(n_755),
.B(n_356),
.Y(n_983)
);

AOI21xp5_ASAP7_75t_L g984 ( 
.A1(n_861),
.A2(n_642),
.B(n_621),
.Y(n_984)
);

CKINVDCx5p33_ASAP7_75t_R g985 ( 
.A(n_864),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_830),
.B(n_699),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_861),
.A2(n_642),
.B(n_621),
.Y(n_987)
);

AOI22xp5_ASAP7_75t_L g988 ( 
.A1(n_834),
.A2(n_652),
.B1(n_644),
.B2(n_673),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_SL g989 ( 
.A(n_719),
.B(n_699),
.Y(n_989)
);

INVxp67_ASAP7_75t_L g990 ( 
.A(n_770),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_750),
.B(n_292),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_762),
.A2(n_642),
.B(n_644),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_730),
.B(n_642),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_732),
.B(n_644),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_734),
.B(n_644),
.Y(n_995)
);

XOR2xp5_ASAP7_75t_L g996 ( 
.A(n_856),
.B(n_340),
.Y(n_996)
);

AO21x1_ASAP7_75t_L g997 ( 
.A1(n_820),
.A2(n_335),
.B(n_239),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_735),
.B(n_644),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_SL g999 ( 
.A(n_776),
.B(n_213),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_876),
.B(n_673),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_742),
.B(n_673),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_786),
.B(n_673),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_786),
.B(n_792),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_765),
.A2(n_693),
.B(n_675),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_745),
.B(n_652),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_757),
.B(n_652),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_879),
.B(n_558),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_738),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_771),
.A2(n_693),
.B(n_675),
.Y(n_1009)
);

NAND2x1p5_ASAP7_75t_L g1010 ( 
.A(n_754),
.B(n_560),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_760),
.B(n_562),
.Y(n_1011)
);

OAI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_875),
.A2(n_695),
.B(n_491),
.Y(n_1012)
);

INVx3_ASAP7_75t_L g1013 ( 
.A(n_738),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_773),
.A2(n_693),
.B(n_675),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_818),
.B(n_562),
.Y(n_1015)
);

INVxp67_ASAP7_75t_L g1016 ( 
.A(n_853),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_739),
.Y(n_1017)
);

AOI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_834),
.A2(n_368),
.B1(n_371),
.B2(n_373),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_812),
.A2(n_661),
.B(n_637),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_818),
.B(n_851),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_874),
.A2(n_661),
.B(n_637),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_873),
.A2(n_661),
.B(n_637),
.Y(n_1022)
);

AO21x1_ASAP7_75t_L g1023 ( 
.A1(n_792),
.A2(n_273),
.B(n_239),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_739),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_857),
.B(n_305),
.Y(n_1025)
);

AOI22xp33_ASAP7_75t_L g1026 ( 
.A1(n_851),
.A2(n_323),
.B1(n_217),
.B2(n_234),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_721),
.B(n_561),
.Y(n_1027)
);

OR2x2_ASAP7_75t_L g1028 ( 
.A(n_816),
.B(n_561),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_840),
.A2(n_571),
.B(n_695),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_857),
.B(n_374),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_772),
.B(n_763),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_831),
.B(n_562),
.Y(n_1032)
);

BUFx2_ASAP7_75t_L g1033 ( 
.A(n_814),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_813),
.A2(n_571),
.B(n_388),
.Y(n_1034)
);

NAND3xp33_ASAP7_75t_SL g1035 ( 
.A(n_766),
.B(n_309),
.C(n_317),
.Y(n_1035)
);

OAI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_740),
.A2(n_491),
.B(n_260),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_740),
.Y(n_1037)
);

INVx3_ASAP7_75t_L g1038 ( 
.A(n_749),
.Y(n_1038)
);

AND2x2_ASAP7_75t_SL g1039 ( 
.A(n_855),
.B(n_260),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_837),
.A2(n_571),
.B(n_268),
.Y(n_1040)
);

BUFx3_ASAP7_75t_L g1041 ( 
.A(n_733),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_SL g1042 ( 
.A(n_845),
.B(n_213),
.Y(n_1042)
);

A2O1A1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_855),
.A2(n_271),
.B(n_273),
.C(n_289),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_758),
.Y(n_1044)
);

OR2x6_ASAP7_75t_L g1045 ( 
.A(n_842),
.B(n_365),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_814),
.B(n_322),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_854),
.B(n_562),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_841),
.A2(n_217),
.B(n_234),
.Y(n_1048)
);

OAI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_880),
.A2(n_491),
.B(n_289),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_824),
.Y(n_1050)
);

O2A1O1Ixp5_ASAP7_75t_L g1051 ( 
.A1(n_882),
.A2(n_323),
.B(n_366),
.C(n_379),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_814),
.B(n_802),
.Y(n_1052)
);

BUFx2_ASAP7_75t_L g1053 ( 
.A(n_842),
.Y(n_1053)
);

NOR3xp33_ASAP7_75t_L g1054 ( 
.A(n_811),
.B(n_364),
.C(n_301),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_834),
.B(n_271),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_834),
.B(n_291),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_824),
.B(n_318),
.Y(n_1057)
);

OAI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_828),
.A2(n_388),
.B1(n_379),
.B2(n_366),
.Y(n_1058)
);

BUFx8_ASAP7_75t_L g1059 ( 
.A(n_845),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_828),
.B(n_320),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_883),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_736),
.B(n_375),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_884),
.B(n_335),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_885),
.B(n_336),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_886),
.B(n_957),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_1007),
.B(n_865),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_1020),
.A2(n_810),
.B1(n_802),
.B2(n_852),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_892),
.Y(n_1068)
);

AOI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_1003),
.A2(n_810),
.B1(n_802),
.B2(n_860),
.Y(n_1069)
);

HB1xp67_ASAP7_75t_L g1070 ( 
.A(n_948),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_897),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_894),
.Y(n_1072)
);

NOR2x1_ASAP7_75t_R g1073 ( 
.A(n_956),
.B(n_334),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_990),
.B(n_1016),
.Y(n_1074)
);

BUFx12f_ASAP7_75t_L g1075 ( 
.A(n_960),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_1039),
.B(n_736),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_R g1077 ( 
.A(n_979),
.B(n_806),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_915),
.A2(n_754),
.B(n_838),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_L g1079 ( 
.A(n_909),
.B(n_810),
.Y(n_1079)
);

OR2x2_ASAP7_75t_L g1080 ( 
.A(n_951),
.B(n_768),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_1026),
.A2(n_898),
.B1(n_915),
.B2(n_899),
.Y(n_1081)
);

OAI21xp33_ASAP7_75t_SL g1082 ( 
.A1(n_1002),
.A2(n_754),
.B(n_869),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_945),
.A2(n_838),
.B(n_848),
.Y(n_1083)
);

AND2x2_ASAP7_75t_L g1084 ( 
.A(n_922),
.B(n_769),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_980),
.B(n_769),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_1025),
.A2(n_885),
.B(n_881),
.C(n_878),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_1027),
.B(n_881),
.Y(n_1087)
);

BUFx2_ASAP7_75t_R g1088 ( 
.A(n_896),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_911),
.B(n_778),
.Y(n_1089)
);

AOI22xp33_ASAP7_75t_L g1090 ( 
.A1(n_1054),
.A2(n_806),
.B1(n_877),
.B2(n_365),
.Y(n_1090)
);

A2O1A1Ixp33_ASAP7_75t_L g1091 ( 
.A1(n_900),
.A2(n_878),
.B(n_872),
.C(n_868),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1061),
.B(n_917),
.Y(n_1092)
);

BUFx2_ASAP7_75t_L g1093 ( 
.A(n_943),
.Y(n_1093)
);

OAI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_1011),
.A2(n_872),
.B1(n_778),
.B2(n_868),
.Y(n_1094)
);

OAI22x1_ASAP7_75t_L g1095 ( 
.A1(n_974),
.A2(n_380),
.B1(n_337),
.B2(n_345),
.Y(n_1095)
);

OAI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_936),
.A2(n_808),
.B(n_867),
.Y(n_1096)
);

INVx3_ASAP7_75t_L g1097 ( 
.A(n_889),
.Y(n_1097)
);

O2A1O1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_906),
.A2(n_358),
.B(n_347),
.C(n_343),
.Y(n_1098)
);

A2O1A1Ixp33_ASAP7_75t_SL g1099 ( 
.A1(n_1000),
.A2(n_796),
.B(n_867),
.C(n_863),
.Y(n_1099)
);

INVx3_ASAP7_75t_SL g1100 ( 
.A(n_985),
.Y(n_1100)
);

INVxp67_ASAP7_75t_L g1101 ( 
.A(n_991),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_958),
.Y(n_1102)
);

BUFx2_ASAP7_75t_L g1103 ( 
.A(n_1052),
.Y(n_1103)
);

OR2x2_ASAP7_75t_L g1104 ( 
.A(n_1028),
.B(n_780),
.Y(n_1104)
);

OAI22x1_ASAP7_75t_L g1105 ( 
.A1(n_965),
.A2(n_363),
.B1(n_377),
.B2(n_346),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_946),
.A2(n_838),
.B(n_848),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_927),
.B(n_780),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_969),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_978),
.A2(n_848),
.B(n_869),
.Y(n_1109)
);

OR2x6_ASAP7_75t_L g1110 ( 
.A(n_1053),
.B(n_848),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_890),
.A2(n_863),
.B(n_862),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_1031),
.B(n_788),
.Y(n_1112)
);

BUFx2_ASAP7_75t_L g1113 ( 
.A(n_928),
.Y(n_1113)
);

NOR2xp67_ASAP7_75t_L g1114 ( 
.A(n_1035),
.B(n_788),
.Y(n_1114)
);

INVx4_ASAP7_75t_L g1115 ( 
.A(n_921),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_960),
.Y(n_1116)
);

INVx2_ASAP7_75t_SL g1117 ( 
.A(n_928),
.Y(n_1117)
);

INVx2_ASAP7_75t_SL g1118 ( 
.A(n_1046),
.Y(n_1118)
);

A2O1A1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_938),
.A2(n_862),
.B(n_850),
.C(n_847),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_940),
.B(n_796),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1013),
.Y(n_1121)
);

OR2x2_ASAP7_75t_L g1122 ( 
.A(n_1033),
.B(n_801),
.Y(n_1122)
);

BUFx2_ASAP7_75t_L g1123 ( 
.A(n_921),
.Y(n_1123)
);

NAND3xp33_ASAP7_75t_SL g1124 ( 
.A(n_999),
.B(n_381),
.C(n_370),
.Y(n_1124)
);

O2A1O1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_1043),
.A2(n_347),
.B(n_342),
.C(n_336),
.Y(n_1125)
);

NOR3xp33_ASAP7_75t_SL g1126 ( 
.A(n_954),
.B(n_964),
.C(n_1030),
.Y(n_1126)
);

AOI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_983),
.A2(n_806),
.B1(n_384),
.B2(n_386),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_890),
.A2(n_847),
.B(n_827),
.Y(n_1128)
);

O2A1O1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_977),
.A2(n_827),
.B(n_808),
.C(n_541),
.Y(n_1129)
);

CKINVDCx14_ASAP7_75t_R g1130 ( 
.A(n_996),
.Y(n_1130)
);

O2A1O1Ixp33_ASAP7_75t_L g1131 ( 
.A1(n_977),
.A2(n_541),
.B(n_538),
.C(n_535),
.Y(n_1131)
);

BUFx12f_ASAP7_75t_L g1132 ( 
.A(n_1059),
.Y(n_1132)
);

AOI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_972),
.A2(n_806),
.B1(n_213),
.B2(n_229),
.Y(n_1133)
);

A2O1A1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_972),
.A2(n_349),
.B(n_361),
.C(n_367),
.Y(n_1134)
);

OAI21xp33_ASAP7_75t_L g1135 ( 
.A1(n_1042),
.A2(n_387),
.B(n_369),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_891),
.A2(n_511),
.B(n_538),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_891),
.A2(n_511),
.B(n_538),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_947),
.B(n_806),
.Y(n_1138)
);

OR2x2_ASAP7_75t_L g1139 ( 
.A(n_939),
.B(n_348),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_939),
.B(n_286),
.Y(n_1140)
);

AOI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_975),
.A2(n_229),
.B1(n_286),
.B2(n_491),
.Y(n_1141)
);

AOI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_1023),
.A2(n_229),
.B1(n_286),
.B2(n_491),
.Y(n_1142)
);

CKINVDCx14_ASAP7_75t_R g1143 ( 
.A(n_968),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_921),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_952),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_1059),
.Y(n_1146)
);

AOI21xp33_ASAP7_75t_L g1147 ( 
.A1(n_1055),
.A2(n_10),
.B(n_12),
.Y(n_1147)
);

BUFx4f_ASAP7_75t_SL g1148 ( 
.A(n_1041),
.Y(n_1148)
);

HB1xp67_ASAP7_75t_L g1149 ( 
.A(n_952),
.Y(n_1149)
);

BUFx3_ASAP7_75t_L g1150 ( 
.A(n_952),
.Y(n_1150)
);

O2A1O1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_1057),
.A2(n_229),
.B(n_286),
.C(n_15),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_975),
.B(n_13),
.Y(n_1152)
);

AOI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_1062),
.A2(n_491),
.B1(n_563),
.B2(n_533),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_L g1154 ( 
.A(n_919),
.Y(n_1154)
);

BUFx6f_ASAP7_75t_L g1155 ( 
.A(n_919),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_933),
.B(n_564),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_959),
.A2(n_564),
.B(n_563),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_913),
.B(n_1045),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_924),
.B(n_564),
.Y(n_1159)
);

A2O1A1Ixp33_ASAP7_75t_SL g1160 ( 
.A1(n_937),
.A2(n_564),
.B(n_563),
.C(n_533),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1015),
.A2(n_564),
.B1(n_563),
.B2(n_533),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_910),
.B(n_916),
.Y(n_1162)
);

OAI22x1_ASAP7_75t_L g1163 ( 
.A1(n_907),
.A2(n_14),
.B1(n_17),
.B2(n_19),
.Y(n_1163)
);

AND2x6_ASAP7_75t_L g1164 ( 
.A(n_1050),
.B(n_966),
.Y(n_1164)
);

AO21x1_ASAP7_75t_L g1165 ( 
.A1(n_1058),
.A2(n_17),
.B(n_23),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_L g1166 ( 
.A(n_916),
.B(n_23),
.Y(n_1166)
);

INVx2_ASAP7_75t_SL g1167 ( 
.A(n_1045),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_984),
.A2(n_564),
.B1(n_563),
.B2(n_533),
.Y(n_1168)
);

BUFx3_ASAP7_75t_L g1169 ( 
.A(n_1045),
.Y(n_1169)
);

INVxp67_ASAP7_75t_SL g1170 ( 
.A(n_1038),
.Y(n_1170)
);

INVxp67_ASAP7_75t_L g1171 ( 
.A(n_1063),
.Y(n_1171)
);

O2A1O1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_1060),
.A2(n_25),
.B(n_26),
.C(n_27),
.Y(n_1172)
);

AOI221xp5_ASAP7_75t_L g1173 ( 
.A1(n_997),
.A2(n_533),
.B1(n_532),
.B2(n_531),
.C(n_564),
.Y(n_1173)
);

HB1xp67_ASAP7_75t_L g1174 ( 
.A(n_976),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1044),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_959),
.A2(n_533),
.B(n_532),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1050),
.B(n_533),
.Y(n_1177)
);

AOI222xp33_ASAP7_75t_L g1178 ( 
.A1(n_1056),
.A2(n_1064),
.B1(n_905),
.B2(n_1008),
.C1(n_1037),
.C2(n_1024),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_971),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_961),
.A2(n_532),
.B(n_531),
.Y(n_1180)
);

AND2x4_ASAP7_75t_L g1181 ( 
.A(n_971),
.B(n_64),
.Y(n_1181)
);

OAI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_984),
.A2(n_532),
.B1(n_531),
.B2(n_28),
.Y(n_1182)
);

OA22x2_ASAP7_75t_L g1183 ( 
.A1(n_949),
.A2(n_986),
.B1(n_981),
.B2(n_1018),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_SL g1184 ( 
.A(n_1005),
.B(n_532),
.Y(n_1184)
);

AND2x2_ASAP7_75t_L g1185 ( 
.A(n_982),
.B(n_532),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_961),
.A2(n_532),
.B(n_531),
.Y(n_1186)
);

O2A1O1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_935),
.A2(n_25),
.B(n_27),
.C(n_29),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_963),
.A2(n_531),
.B(n_78),
.Y(n_1188)
);

OAI22x1_ASAP7_75t_L g1189 ( 
.A1(n_962),
.A2(n_29),
.B1(n_33),
.B2(n_38),
.Y(n_1189)
);

O2A1O1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_918),
.A2(n_38),
.B(n_40),
.C(n_41),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_963),
.A2(n_531),
.B(n_130),
.Y(n_1191)
);

NAND3xp33_ASAP7_75t_L g1192 ( 
.A(n_1048),
.B(n_531),
.C(n_43),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_1032),
.B(n_42),
.Y(n_1193)
);

O2A1O1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_1047),
.A2(n_46),
.B(n_47),
.C(n_48),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_987),
.A2(n_133),
.B(n_176),
.Y(n_1195)
);

BUFx2_ASAP7_75t_SL g1196 ( 
.A(n_1017),
.Y(n_1196)
);

OAI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_987),
.A2(n_46),
.B1(n_53),
.B2(n_55),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_1006),
.B(n_136),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_993),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_950),
.A2(n_53),
.B1(n_58),
.B2(n_59),
.Y(n_1200)
);

O2A1O1Ixp33_ASAP7_75t_L g1201 ( 
.A1(n_989),
.A2(n_59),
.B(n_60),
.C(n_61),
.Y(n_1201)
);

OAI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_988),
.A2(n_62),
.B1(n_79),
.B2(n_82),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_955),
.Y(n_1203)
);

BUFx12f_ASAP7_75t_L g1204 ( 
.A(n_1010),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_994),
.B(n_995),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_970),
.A2(n_145),
.B(n_132),
.Y(n_1206)
);

A2O1A1Ixp33_ASAP7_75t_L g1207 ( 
.A1(n_1079),
.A2(n_973),
.B(n_923),
.C(n_1049),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1102),
.Y(n_1208)
);

OAI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1081),
.A2(n_942),
.B(n_893),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1092),
.Y(n_1210)
);

AO31x2_ASAP7_75t_L g1211 ( 
.A1(n_1182),
.A2(n_953),
.A3(n_942),
.B(n_973),
.Y(n_1211)
);

INVx3_ASAP7_75t_L g1212 ( 
.A(n_1179),
.Y(n_1212)
);

INVx4_ASAP7_75t_L g1213 ( 
.A(n_1179),
.Y(n_1213)
);

OAI21x1_ASAP7_75t_L g1214 ( 
.A1(n_1111),
.A2(n_936),
.B(n_944),
.Y(n_1214)
);

OR2x2_ASAP7_75t_L g1215 ( 
.A(n_1104),
.B(n_1093),
.Y(n_1215)
);

INVx1_ASAP7_75t_SL g1216 ( 
.A(n_1088),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1108),
.Y(n_1217)
);

BUFx2_ASAP7_75t_L g1218 ( 
.A(n_1070),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1128),
.A2(n_1096),
.B(n_1078),
.Y(n_1219)
);

AO21x1_ASAP7_75t_L g1220 ( 
.A1(n_1182),
.A2(n_1048),
.B(n_887),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1082),
.A2(n_970),
.B(n_1010),
.Y(n_1221)
);

AO31x2_ASAP7_75t_L g1222 ( 
.A1(n_1081),
.A2(n_920),
.A3(n_914),
.B(n_895),
.Y(n_1222)
);

OAI22x1_ASAP7_75t_L g1223 ( 
.A1(n_1069),
.A2(n_925),
.B1(n_888),
.B2(n_926),
.Y(n_1223)
);

AO31x2_ASAP7_75t_L g1224 ( 
.A1(n_1161),
.A2(n_920),
.A3(n_914),
.B(n_902),
.Y(n_1224)
);

OAI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1086),
.A2(n_893),
.B(n_1051),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1084),
.B(n_1001),
.Y(n_1226)
);

AO31x2_ASAP7_75t_L g1227 ( 
.A1(n_1161),
.A2(n_901),
.A3(n_904),
.B(n_903),
.Y(n_1227)
);

O2A1O1Ixp5_ASAP7_75t_SL g1228 ( 
.A1(n_1197),
.A2(n_941),
.B(n_912),
.C(n_930),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1065),
.B(n_998),
.Y(n_1229)
);

A2O1A1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1126),
.A2(n_1034),
.B(n_908),
.C(n_1040),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1083),
.A2(n_931),
.B(n_992),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1096),
.A2(n_967),
.B(n_992),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_L g1233 ( 
.A(n_1074),
.B(n_1034),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1106),
.A2(n_1029),
.B(n_934),
.Y(n_1234)
);

AOI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1205),
.A2(n_1029),
.B(n_934),
.Y(n_1235)
);

BUFx10_ASAP7_75t_L g1236 ( 
.A(n_1154),
.Y(n_1236)
);

BUFx2_ASAP7_75t_R g1237 ( 
.A(n_1100),
.Y(n_1237)
);

NAND3xp33_ASAP7_75t_L g1238 ( 
.A(n_1067),
.B(n_1040),
.C(n_929),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1136),
.A2(n_904),
.B(n_903),
.Y(n_1239)
);

AO21x1_ASAP7_75t_L g1240 ( 
.A1(n_1197),
.A2(n_902),
.B(n_901),
.Y(n_1240)
);

AO31x2_ASAP7_75t_L g1241 ( 
.A1(n_1168),
.A2(n_895),
.A3(n_1019),
.B(n_1014),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1109),
.A2(n_1019),
.B(n_1022),
.Y(n_1242)
);

NAND2x1_ASAP7_75t_L g1243 ( 
.A(n_1164),
.B(n_1021),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1065),
.B(n_908),
.Y(n_1244)
);

A2O1A1Ixp33_ASAP7_75t_L g1245 ( 
.A1(n_1067),
.A2(n_929),
.B(n_1012),
.C(n_1036),
.Y(n_1245)
);

NAND2x1p5_ASAP7_75t_L g1246 ( 
.A(n_1115),
.B(n_932),
.Y(n_1246)
);

OAI21xp5_ASAP7_75t_SL g1247 ( 
.A1(n_1200),
.A2(n_1021),
.B(n_1014),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1174),
.Y(n_1248)
);

BUFx12f_ASAP7_75t_L g1249 ( 
.A(n_1075),
.Y(n_1249)
);

OAI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1119),
.A2(n_1009),
.B(n_1004),
.Y(n_1250)
);

A2O1A1Ixp33_ASAP7_75t_L g1251 ( 
.A1(n_1066),
.A2(n_1009),
.B(n_1004),
.C(n_1022),
.Y(n_1251)
);

OR2x2_ASAP7_75t_L g1252 ( 
.A(n_1103),
.B(n_62),
.Y(n_1252)
);

OAI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1137),
.A2(n_186),
.B(n_140),
.Y(n_1253)
);

NOR2xp33_ASAP7_75t_L g1254 ( 
.A(n_1171),
.B(n_166),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1156),
.A2(n_137),
.B(n_144),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1085),
.B(n_152),
.Y(n_1256)
);

CKINVDCx11_ASAP7_75t_R g1257 ( 
.A(n_1132),
.Y(n_1257)
);

CKINVDCx8_ASAP7_75t_R g1258 ( 
.A(n_1154),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1089),
.Y(n_1259)
);

NAND2xp5_ASAP7_75t_L g1260 ( 
.A(n_1112),
.B(n_159),
.Y(n_1260)
);

A2O1A1Ixp33_ASAP7_75t_L g1261 ( 
.A1(n_1193),
.A2(n_1114),
.B(n_1101),
.C(n_1140),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1159),
.A2(n_1162),
.B(n_1076),
.Y(n_1262)
);

O2A1O1Ixp33_ASAP7_75t_L g1263 ( 
.A1(n_1200),
.A2(n_1134),
.B(n_1151),
.C(n_1172),
.Y(n_1263)
);

AOI31xp67_ASAP7_75t_L g1264 ( 
.A1(n_1183),
.A2(n_1203),
.A3(n_1184),
.B(n_1198),
.Y(n_1264)
);

NAND2x1p5_ASAP7_75t_L g1265 ( 
.A(n_1115),
.B(n_1179),
.Y(n_1265)
);

O2A1O1Ixp33_ASAP7_75t_L g1266 ( 
.A1(n_1124),
.A2(n_1147),
.B(n_1194),
.C(n_1202),
.Y(n_1266)
);

AND2x4_ASAP7_75t_L g1267 ( 
.A(n_1117),
.B(n_1150),
.Y(n_1267)
);

INVx2_ASAP7_75t_SL g1268 ( 
.A(n_1144),
.Y(n_1268)
);

BUFx2_ASAP7_75t_L g1269 ( 
.A(n_1113),
.Y(n_1269)
);

O2A1O1Ixp5_ASAP7_75t_L g1270 ( 
.A1(n_1165),
.A2(n_1195),
.B(n_1188),
.C(n_1191),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1178),
.A2(n_1099),
.B(n_1183),
.Y(n_1271)
);

OR2x6_ASAP7_75t_L g1272 ( 
.A(n_1154),
.B(n_1155),
.Y(n_1272)
);

AO31x2_ASAP7_75t_L g1273 ( 
.A1(n_1168),
.A2(n_1091),
.A3(n_1094),
.B(n_1157),
.Y(n_1273)
);

AO31x2_ASAP7_75t_L g1274 ( 
.A1(n_1094),
.A2(n_1176),
.A3(n_1180),
.B(n_1186),
.Y(n_1274)
);

INVx4_ASAP7_75t_L g1275 ( 
.A(n_1144),
.Y(n_1275)
);

INVx3_ASAP7_75t_L g1276 ( 
.A(n_1164),
.Y(n_1276)
);

AOI221xp5_ASAP7_75t_L g1277 ( 
.A1(n_1095),
.A2(n_1105),
.B1(n_1147),
.B2(n_1135),
.C(n_1163),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_L g1278 ( 
.A(n_1118),
.B(n_1071),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1087),
.B(n_1199),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_L g1280 ( 
.A(n_1080),
.B(n_1139),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1122),
.B(n_1120),
.Y(n_1281)
);

INVxp67_ASAP7_75t_L g1282 ( 
.A(n_1149),
.Y(n_1282)
);

INVx1_ASAP7_75t_SL g1283 ( 
.A(n_1123),
.Y(n_1283)
);

OAI21x1_ASAP7_75t_L g1284 ( 
.A1(n_1177),
.A2(n_1129),
.B(n_1206),
.Y(n_1284)
);

A2O1A1Ixp33_ASAP7_75t_L g1285 ( 
.A1(n_1152),
.A2(n_1201),
.B(n_1138),
.C(n_1166),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1107),
.B(n_1068),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1185),
.A2(n_1131),
.B(n_1072),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_1145),
.Y(n_1288)
);

INVxp67_ASAP7_75t_L g1289 ( 
.A(n_1145),
.Y(n_1289)
);

NOR2xp33_ASAP7_75t_L g1290 ( 
.A(n_1130),
.B(n_1155),
.Y(n_1290)
);

CKINVDCx9p33_ASAP7_75t_R g1291 ( 
.A(n_1148),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_SL g1292 ( 
.A1(n_1202),
.A2(n_1187),
.B(n_1190),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1178),
.A2(n_1170),
.B(n_1097),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1097),
.A2(n_1181),
.B(n_1160),
.Y(n_1294)
);

BUFx12f_ASAP7_75t_L g1295 ( 
.A(n_1116),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1158),
.B(n_1167),
.Y(n_1296)
);

NAND3xp33_ASAP7_75t_L g1297 ( 
.A(n_1192),
.B(n_1098),
.C(n_1142),
.Y(n_1297)
);

BUFx12f_ASAP7_75t_L g1298 ( 
.A(n_1146),
.Y(n_1298)
);

A2O1A1Ixp33_ASAP7_75t_L g1299 ( 
.A1(n_1133),
.A2(n_1125),
.B(n_1127),
.C(n_1192),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1121),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1196),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1189),
.A2(n_1090),
.B1(n_1181),
.B2(n_1169),
.Y(n_1302)
);

AO31x2_ASAP7_75t_L g1303 ( 
.A1(n_1173),
.A2(n_1141),
.A3(n_1153),
.B(n_1164),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1110),
.A2(n_1155),
.B(n_1164),
.Y(n_1304)
);

OAI22xp5_ASAP7_75t_L g1305 ( 
.A1(n_1110),
.A2(n_1204),
.B1(n_1143),
.B2(n_1077),
.Y(n_1305)
);

AO21x1_ASAP7_75t_L g1306 ( 
.A1(n_1110),
.A2(n_1003),
.B(n_1182),
.Y(n_1306)
);

OAI22xp5_ASAP7_75t_L g1307 ( 
.A1(n_1073),
.A2(n_1020),
.B1(n_760),
.B2(n_851),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1078),
.A2(n_809),
.B(n_915),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1111),
.A2(n_1128),
.B(n_1096),
.Y(n_1309)
);

A2O1A1Ixp33_ASAP7_75t_L g1310 ( 
.A1(n_1079),
.A2(n_957),
.B(n_1003),
.C(n_1016),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1111),
.A2(n_1128),
.B(n_1096),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1078),
.A2(n_809),
.B(n_915),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1078),
.A2(n_809),
.B(n_915),
.Y(n_1313)
);

OR2x2_ASAP7_75t_L g1314 ( 
.A(n_1104),
.B(n_520),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1111),
.A2(n_1128),
.B(n_1096),
.Y(n_1315)
);

OAI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1069),
.A2(n_782),
.B1(n_566),
.B2(n_804),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1065),
.A2(n_1020),
.B1(n_760),
.B2(n_851),
.Y(n_1317)
);

INVx1_ASAP7_75t_SL g1318 ( 
.A(n_1088),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1078),
.A2(n_809),
.B(n_915),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1078),
.A2(n_809),
.B(n_915),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1078),
.A2(n_809),
.B(n_915),
.Y(n_1321)
);

O2A1O1Ixp33_ASAP7_75t_SL g1322 ( 
.A1(n_1076),
.A2(n_1003),
.B(n_1020),
.C(n_906),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1111),
.A2(n_1128),
.B(n_1096),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1111),
.A2(n_1128),
.B(n_1096),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1078),
.A2(n_809),
.B(n_915),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1065),
.B(n_1112),
.Y(n_1326)
);

OR2x2_ASAP7_75t_L g1327 ( 
.A(n_1104),
.B(n_520),
.Y(n_1327)
);

NOR2xp33_ASAP7_75t_L g1328 ( 
.A(n_1074),
.B(n_741),
.Y(n_1328)
);

BUFx3_ASAP7_75t_L g1329 ( 
.A(n_1100),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1111),
.A2(n_1128),
.B(n_1096),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1111),
.A2(n_1128),
.B(n_1096),
.Y(n_1331)
);

AO31x2_ASAP7_75t_L g1332 ( 
.A1(n_1182),
.A2(n_953),
.A3(n_1023),
.B(n_997),
.Y(n_1332)
);

HB1xp67_ASAP7_75t_L g1333 ( 
.A(n_1113),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1084),
.B(n_725),
.Y(n_1334)
);

A2O1A1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1079),
.A2(n_957),
.B(n_1003),
.C(n_1016),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_SL g1336 ( 
.A1(n_1165),
.A2(n_900),
.B(n_1195),
.Y(n_1336)
);

A2O1A1Ixp33_ASAP7_75t_L g1337 ( 
.A1(n_1079),
.A2(n_957),
.B(n_1003),
.C(n_1016),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1103),
.B(n_922),
.Y(n_1338)
);

INVxp67_ASAP7_75t_SL g1339 ( 
.A(n_1122),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1092),
.Y(n_1340)
);

BUFx2_ASAP7_75t_L g1341 ( 
.A(n_1093),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1111),
.A2(n_1128),
.B(n_1096),
.Y(n_1342)
);

OAI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1081),
.A2(n_915),
.B(n_1003),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1175),
.Y(n_1344)
);

AO31x2_ASAP7_75t_L g1345 ( 
.A1(n_1182),
.A2(n_953),
.A3(n_1023),
.B(n_997),
.Y(n_1345)
);

AO31x2_ASAP7_75t_L g1346 ( 
.A1(n_1182),
.A2(n_953),
.A3(n_1023),
.B(n_997),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_L g1347 ( 
.A(n_1074),
.B(n_741),
.Y(n_1347)
);

AO31x2_ASAP7_75t_L g1348 ( 
.A1(n_1182),
.A2(n_953),
.A3(n_1023),
.B(n_997),
.Y(n_1348)
);

INVx3_ASAP7_75t_SL g1349 ( 
.A(n_1100),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1078),
.A2(n_809),
.B(n_915),
.Y(n_1350)
);

NOR2xp67_ASAP7_75t_SL g1351 ( 
.A(n_1075),
.B(n_896),
.Y(n_1351)
);

AND2x4_ASAP7_75t_L g1352 ( 
.A(n_1117),
.B(n_1150),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1084),
.B(n_725),
.Y(n_1353)
);

AOI21xp5_ASAP7_75t_L g1354 ( 
.A1(n_1078),
.A2(n_809),
.B(n_915),
.Y(n_1354)
);

INVx1_ASAP7_75t_SL g1355 ( 
.A(n_1088),
.Y(n_1355)
);

OR2x2_ASAP7_75t_L g1356 ( 
.A(n_1104),
.B(n_520),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1103),
.B(n_922),
.Y(n_1357)
);

AOI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1078),
.A2(n_809),
.B(n_915),
.Y(n_1358)
);

NOR2xp33_ASAP7_75t_SL g1359 ( 
.A(n_1088),
.B(n_957),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_SL g1360 ( 
.A1(n_1285),
.A2(n_1335),
.B(n_1310),
.Y(n_1360)
);

INVxp67_ASAP7_75t_SL g1361 ( 
.A(n_1293),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1277),
.A2(n_1316),
.B1(n_1307),
.B2(n_1328),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1210),
.A2(n_1340),
.B1(n_1353),
.B2(n_1334),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1347),
.A2(n_1317),
.B1(n_1326),
.B2(n_1302),
.Y(n_1364)
);

CKINVDCx11_ASAP7_75t_R g1365 ( 
.A(n_1257),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1217),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_SL g1367 ( 
.A1(n_1337),
.A2(n_1299),
.B(n_1207),
.Y(n_1367)
);

BUFx12f_ASAP7_75t_L g1368 ( 
.A(n_1249),
.Y(n_1368)
);

AOI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1359),
.A2(n_1280),
.B1(n_1254),
.B2(n_1307),
.Y(n_1369)
);

NAND2x1p5_ASAP7_75t_L g1370 ( 
.A(n_1213),
.B(n_1276),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1306),
.A2(n_1292),
.B1(n_1233),
.B2(n_1297),
.Y(n_1371)
);

BUFx3_ASAP7_75t_L g1372 ( 
.A(n_1341),
.Y(n_1372)
);

OAI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1359),
.A2(n_1215),
.B1(n_1327),
.B2(n_1314),
.Y(n_1373)
);

CKINVDCx11_ASAP7_75t_R g1374 ( 
.A(n_1295),
.Y(n_1374)
);

INVx1_ASAP7_75t_SL g1375 ( 
.A(n_1338),
.Y(n_1375)
);

OAI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1356),
.A2(n_1279),
.B1(n_1318),
.B2(n_1355),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1297),
.A2(n_1317),
.B1(n_1357),
.B2(n_1296),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1269),
.A2(n_1333),
.B1(n_1253),
.B2(n_1260),
.Y(n_1378)
);

CKINVDCx11_ASAP7_75t_R g1379 ( 
.A(n_1298),
.Y(n_1379)
);

CKINVDCx11_ASAP7_75t_R g1380 ( 
.A(n_1258),
.Y(n_1380)
);

BUFx2_ASAP7_75t_SL g1381 ( 
.A(n_1329),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1344),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1339),
.B(n_1248),
.Y(n_1383)
);

INVx1_ASAP7_75t_SL g1384 ( 
.A(n_1283),
.Y(n_1384)
);

INVx3_ASAP7_75t_SL g1385 ( 
.A(n_1272),
.Y(n_1385)
);

AOI22xp33_ASAP7_75t_L g1386 ( 
.A1(n_1253),
.A2(n_1260),
.B1(n_1256),
.B2(n_1343),
.Y(n_1386)
);

OAI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1326),
.A2(n_1281),
.B1(n_1244),
.B2(n_1259),
.Y(n_1387)
);

INVx6_ASAP7_75t_L g1388 ( 
.A(n_1236),
.Y(n_1388)
);

INVxp67_ASAP7_75t_SL g1389 ( 
.A(n_1240),
.Y(n_1389)
);

OAI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1216),
.A2(n_1355),
.B1(n_1318),
.B2(n_1301),
.Y(n_1390)
);

BUFx6f_ASAP7_75t_L g1391 ( 
.A(n_1272),
.Y(n_1391)
);

BUFx10_ASAP7_75t_L g1392 ( 
.A(n_1290),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1300),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1343),
.A2(n_1218),
.B1(n_1336),
.B2(n_1252),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1238),
.A2(n_1271),
.B1(n_1223),
.B2(n_1278),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1286),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1238),
.A2(n_1283),
.B1(n_1226),
.B2(n_1220),
.Y(n_1397)
);

CKINVDCx11_ASAP7_75t_R g1398 ( 
.A(n_1216),
.Y(n_1398)
);

INVx6_ASAP7_75t_L g1399 ( 
.A(n_1213),
.Y(n_1399)
);

BUFx6f_ASAP7_75t_L g1400 ( 
.A(n_1272),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1286),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_L g1402 ( 
.A1(n_1282),
.A2(n_1267),
.B1(n_1352),
.B2(n_1351),
.Y(n_1402)
);

OAI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1229),
.A2(n_1245),
.B1(n_1261),
.B2(n_1266),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1267),
.A2(n_1352),
.B1(n_1262),
.B2(n_1305),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1212),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1212),
.Y(n_1406)
);

BUFx12f_ASAP7_75t_L g1407 ( 
.A(n_1288),
.Y(n_1407)
);

BUFx2_ASAP7_75t_L g1408 ( 
.A(n_1289),
.Y(n_1408)
);

OAI21xp5_ASAP7_75t_SL g1409 ( 
.A1(n_1263),
.A2(n_1247),
.B(n_1305),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1308),
.A2(n_1313),
.B(n_1354),
.Y(n_1410)
);

BUFx10_ASAP7_75t_L g1411 ( 
.A(n_1268),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1255),
.A2(n_1209),
.B1(n_1294),
.B2(n_1287),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_L g1413 ( 
.A1(n_1209),
.A2(n_1304),
.B1(n_1235),
.B2(n_1250),
.Y(n_1413)
);

BUFx3_ASAP7_75t_L g1414 ( 
.A(n_1265),
.Y(n_1414)
);

BUFx3_ASAP7_75t_L g1415 ( 
.A(n_1275),
.Y(n_1415)
);

BUFx6f_ASAP7_75t_L g1416 ( 
.A(n_1275),
.Y(n_1416)
);

OAI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1247),
.A2(n_1276),
.B1(n_1243),
.B2(n_1246),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1322),
.B(n_1230),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1250),
.A2(n_1231),
.B1(n_1325),
.B2(n_1319),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1222),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1222),
.Y(n_1421)
);

INVx6_ASAP7_75t_L g1422 ( 
.A(n_1237),
.Y(n_1422)
);

BUFx12f_ASAP7_75t_L g1423 ( 
.A(n_1270),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1312),
.A2(n_1358),
.B1(n_1320),
.B2(n_1321),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_SL g1425 ( 
.A1(n_1350),
.A2(n_1225),
.B1(n_1219),
.B2(n_1221),
.Y(n_1425)
);

AOI22xp5_ASAP7_75t_SL g1426 ( 
.A1(n_1234),
.A2(n_1225),
.B1(n_1242),
.B2(n_1264),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_SL g1427 ( 
.A1(n_1309),
.A2(n_1324),
.B1(n_1342),
.B2(n_1331),
.Y(n_1427)
);

INVx3_ASAP7_75t_L g1428 ( 
.A(n_1222),
.Y(n_1428)
);

CKINVDCx11_ASAP7_75t_R g1429 ( 
.A(n_1228),
.Y(n_1429)
);

CKINVDCx11_ASAP7_75t_R g1430 ( 
.A(n_1332),
.Y(n_1430)
);

CKINVDCx16_ASAP7_75t_R g1431 ( 
.A(n_1332),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_SL g1432 ( 
.A1(n_1311),
.A2(n_1315),
.B1(n_1323),
.B2(n_1330),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1284),
.A2(n_1239),
.B1(n_1232),
.B2(n_1214),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1332),
.A2(n_1348),
.B1(n_1346),
.B2(n_1345),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_SL g1435 ( 
.A1(n_1345),
.A2(n_1348),
.B1(n_1346),
.B2(n_1303),
.Y(n_1435)
);

BUFx12f_ASAP7_75t_L g1436 ( 
.A(n_1251),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1345),
.A2(n_1348),
.B1(n_1346),
.B2(n_1303),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1227),
.Y(n_1438)
);

NAND2x1p5_ASAP7_75t_L g1439 ( 
.A(n_1241),
.B(n_1274),
.Y(n_1439)
);

BUFx2_ASAP7_75t_SL g1440 ( 
.A(n_1224),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1303),
.A2(n_1211),
.B1(n_1241),
.B2(n_1273),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_SL g1442 ( 
.A1(n_1273),
.A2(n_1211),
.B1(n_1241),
.B2(n_1274),
.Y(n_1442)
);

AOI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1211),
.A2(n_1273),
.B1(n_1274),
.B2(n_1224),
.Y(n_1443)
);

INVx6_ASAP7_75t_L g1444 ( 
.A(n_1236),
.Y(n_1444)
);

NAND2x1p5_ASAP7_75t_L g1445 ( 
.A(n_1213),
.B(n_889),
.Y(n_1445)
);

CKINVDCx20_ASAP7_75t_R g1446 ( 
.A(n_1291),
.Y(n_1446)
);

CKINVDCx20_ASAP7_75t_R g1447 ( 
.A(n_1291),
.Y(n_1447)
);

BUFx6f_ASAP7_75t_L g1448 ( 
.A(n_1258),
.Y(n_1448)
);

INVx4_ASAP7_75t_L g1449 ( 
.A(n_1272),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1277),
.A2(n_957),
.B1(n_974),
.B2(n_1003),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_SL g1451 ( 
.A1(n_1307),
.A2(n_566),
.B1(n_909),
.B2(n_974),
.Y(n_1451)
);

BUFx6f_ASAP7_75t_L g1452 ( 
.A(n_1258),
.Y(n_1452)
);

AOI22xp5_ASAP7_75t_SL g1453 ( 
.A1(n_1328),
.A2(n_974),
.B1(n_1016),
.B2(n_1079),
.Y(n_1453)
);

INVx4_ASAP7_75t_L g1454 ( 
.A(n_1272),
.Y(n_1454)
);

CKINVDCx16_ASAP7_75t_R g1455 ( 
.A(n_1249),
.Y(n_1455)
);

OAI21xp5_ASAP7_75t_SL g1456 ( 
.A1(n_1316),
.A2(n_974),
.B(n_909),
.Y(n_1456)
);

OAI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1359),
.A2(n_566),
.B1(n_1020),
.B2(n_725),
.Y(n_1457)
);

OAI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1271),
.A2(n_1003),
.B(n_957),
.Y(n_1458)
);

BUFx10_ASAP7_75t_L g1459 ( 
.A(n_1290),
.Y(n_1459)
);

BUFx10_ASAP7_75t_L g1460 ( 
.A(n_1290),
.Y(n_1460)
);

BUFx8_ASAP7_75t_L g1461 ( 
.A(n_1249),
.Y(n_1461)
);

BUFx10_ASAP7_75t_L g1462 ( 
.A(n_1290),
.Y(n_1462)
);

INVx1_ASAP7_75t_SL g1463 ( 
.A(n_1215),
.Y(n_1463)
);

CKINVDCx6p67_ASAP7_75t_R g1464 ( 
.A(n_1291),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1326),
.B(n_1279),
.Y(n_1465)
);

AOI22xp5_ASAP7_75t_SL g1466 ( 
.A1(n_1328),
.A2(n_974),
.B1(n_1016),
.B2(n_1079),
.Y(n_1466)
);

BUFx6f_ASAP7_75t_L g1467 ( 
.A(n_1258),
.Y(n_1467)
);

OAI21xp5_ASAP7_75t_SL g1468 ( 
.A1(n_1316),
.A2(n_974),
.B(n_909),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1208),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1326),
.B(n_1279),
.Y(n_1470)
);

CKINVDCx14_ASAP7_75t_R g1471 ( 
.A(n_1257),
.Y(n_1471)
);

BUFx3_ASAP7_75t_L g1472 ( 
.A(n_1341),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1277),
.A2(n_957),
.B1(n_974),
.B2(n_1003),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_SL g1474 ( 
.A1(n_1307),
.A2(n_566),
.B1(n_909),
.B2(n_974),
.Y(n_1474)
);

INVx6_ASAP7_75t_L g1475 ( 
.A(n_1236),
.Y(n_1475)
);

CKINVDCx20_ASAP7_75t_R g1476 ( 
.A(n_1291),
.Y(n_1476)
);

INVx1_ASAP7_75t_SL g1477 ( 
.A(n_1215),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1277),
.A2(n_957),
.B1(n_974),
.B2(n_1003),
.Y(n_1478)
);

OAI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1210),
.A2(n_1020),
.B1(n_760),
.B2(n_851),
.Y(n_1479)
);

CKINVDCx20_ASAP7_75t_R g1480 ( 
.A(n_1291),
.Y(n_1480)
);

INVx3_ASAP7_75t_SL g1481 ( 
.A(n_1349),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1208),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_SL g1483 ( 
.A1(n_1307),
.A2(n_566),
.B1(n_909),
.B2(n_974),
.Y(n_1483)
);

OAI21xp5_ASAP7_75t_SL g1484 ( 
.A1(n_1316),
.A2(n_974),
.B(n_909),
.Y(n_1484)
);

CKINVDCx20_ASAP7_75t_R g1485 ( 
.A(n_1291),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1208),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1277),
.A2(n_957),
.B1(n_974),
.B2(n_1003),
.Y(n_1487)
);

OAI22x1_ASAP7_75t_SL g1488 ( 
.A1(n_1216),
.A2(n_822),
.B1(n_864),
.B2(n_1116),
.Y(n_1488)
);

OAI22xp33_ASAP7_75t_L g1489 ( 
.A1(n_1359),
.A2(n_566),
.B1(n_804),
.B2(n_782),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_SL g1490 ( 
.A1(n_1307),
.A2(n_566),
.B1(n_909),
.B2(n_974),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1277),
.A2(n_957),
.B1(n_974),
.B2(n_1003),
.Y(n_1491)
);

INVx4_ASAP7_75t_L g1492 ( 
.A(n_1272),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1421),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1410),
.A2(n_1433),
.B(n_1424),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1465),
.B(n_1470),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1465),
.B(n_1470),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1420),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1363),
.B(n_1463),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1366),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1431),
.B(n_1361),
.Y(n_1500)
);

INVx2_ASAP7_75t_SL g1501 ( 
.A(n_1399),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1361),
.B(n_1437),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1438),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1363),
.B(n_1463),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1371),
.B(n_1377),
.Y(n_1505)
);

HB1xp67_ASAP7_75t_L g1506 ( 
.A(n_1383),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1435),
.B(n_1430),
.Y(n_1507)
);

INVx2_ASAP7_75t_SL g1508 ( 
.A(n_1399),
.Y(n_1508)
);

OA21x2_ASAP7_75t_L g1509 ( 
.A1(n_1410),
.A2(n_1389),
.B(n_1434),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1428),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1428),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1389),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1384),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1443),
.Y(n_1514)
);

INVx2_ASAP7_75t_SL g1515 ( 
.A(n_1399),
.Y(n_1515)
);

OAI21x1_ASAP7_75t_L g1516 ( 
.A1(n_1419),
.A2(n_1439),
.B(n_1412),
.Y(n_1516)
);

BUFx12f_ASAP7_75t_L g1517 ( 
.A(n_1365),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1440),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1418),
.Y(n_1519)
);

AO31x2_ASAP7_75t_L g1520 ( 
.A1(n_1403),
.A2(n_1418),
.A3(n_1364),
.B(n_1387),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1442),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1442),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1441),
.B(n_1387),
.Y(n_1523)
);

BUFx3_ASAP7_75t_L g1524 ( 
.A(n_1407),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_1384),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1469),
.Y(n_1526)
);

CKINVDCx20_ASAP7_75t_R g1527 ( 
.A(n_1446),
.Y(n_1527)
);

INVx3_ASAP7_75t_L g1528 ( 
.A(n_1436),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1458),
.B(n_1395),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1482),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1403),
.Y(n_1531)
);

OR2x6_ASAP7_75t_L g1532 ( 
.A(n_1367),
.B(n_1360),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1486),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1393),
.Y(n_1534)
);

CKINVDCx16_ASAP7_75t_R g1535 ( 
.A(n_1455),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1458),
.B(n_1397),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1362),
.B(n_1375),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1451),
.A2(n_1474),
.B1(n_1483),
.B2(n_1490),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1375),
.B(n_1396),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1477),
.B(n_1401),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1426),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1477),
.B(n_1453),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1466),
.B(n_1364),
.Y(n_1543)
);

OA21x2_ASAP7_75t_L g1544 ( 
.A1(n_1413),
.A2(n_1386),
.B(n_1409),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1450),
.B(n_1473),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1394),
.B(n_1429),
.Y(n_1546)
);

BUFx2_ASAP7_75t_L g1547 ( 
.A(n_1423),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1382),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1378),
.B(n_1369),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1373),
.B(n_1376),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1427),
.Y(n_1551)
);

INVx2_ASAP7_75t_SL g1552 ( 
.A(n_1391),
.Y(n_1552)
);

AO21x2_ASAP7_75t_L g1553 ( 
.A1(n_1417),
.A2(n_1456),
.B(n_1468),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1427),
.Y(n_1554)
);

OAI21x1_ASAP7_75t_L g1555 ( 
.A1(n_1404),
.A2(n_1370),
.B(n_1479),
.Y(n_1555)
);

OAI21xp5_ASAP7_75t_L g1556 ( 
.A1(n_1484),
.A2(n_1474),
.B(n_1451),
.Y(n_1556)
);

OAI21x1_ASAP7_75t_L g1557 ( 
.A1(n_1370),
.A2(n_1479),
.B(n_1432),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1432),
.Y(n_1558)
);

BUFx2_ASAP7_75t_L g1559 ( 
.A(n_1449),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1425),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1425),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1483),
.B(n_1490),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1405),
.B(n_1406),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1400),
.Y(n_1564)
);

BUFx3_ASAP7_75t_L g1565 ( 
.A(n_1448),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1478),
.B(n_1491),
.Y(n_1566)
);

INVx2_ASAP7_75t_SL g1567 ( 
.A(n_1388),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1390),
.B(n_1457),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1454),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1492),
.Y(n_1570)
);

OAI21x1_ASAP7_75t_L g1571 ( 
.A1(n_1487),
.A2(n_1445),
.B(n_1402),
.Y(n_1571)
);

INVx1_ASAP7_75t_SL g1572 ( 
.A(n_1372),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1457),
.Y(n_1573)
);

BUFx3_ASAP7_75t_L g1574 ( 
.A(n_1448),
.Y(n_1574)
);

INVx1_ASAP7_75t_SL g1575 ( 
.A(n_1472),
.Y(n_1575)
);

AOI21x1_ASAP7_75t_L g1576 ( 
.A1(n_1408),
.A2(n_1385),
.B(n_1489),
.Y(n_1576)
);

INVx1_ASAP7_75t_SL g1577 ( 
.A(n_1380),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1385),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1414),
.Y(n_1579)
);

AO31x2_ASAP7_75t_L g1580 ( 
.A1(n_1411),
.A2(n_1416),
.A3(n_1459),
.B(n_1392),
.Y(n_1580)
);

NAND2x1_ASAP7_75t_L g1581 ( 
.A(n_1388),
.B(n_1444),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1392),
.B(n_1460),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1411),
.Y(n_1583)
);

AOI22xp33_ASAP7_75t_L g1584 ( 
.A1(n_1422),
.A2(n_1481),
.B1(n_1462),
.B2(n_1459),
.Y(n_1584)
);

AO21x2_ASAP7_75t_L g1585 ( 
.A1(n_1460),
.A2(n_1462),
.B(n_1475),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1398),
.B(n_1488),
.Y(n_1586)
);

BUFx6f_ASAP7_75t_L g1587 ( 
.A(n_1448),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1415),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1452),
.B(n_1467),
.Y(n_1589)
);

OAI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1422),
.A2(n_1481),
.B1(n_1452),
.B2(n_1467),
.Y(n_1590)
);

NAND2x1_ASAP7_75t_L g1591 ( 
.A(n_1444),
.B(n_1475),
.Y(n_1591)
);

CKINVDCx20_ASAP7_75t_R g1592 ( 
.A(n_1447),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1500),
.B(n_1381),
.Y(n_1593)
);

CKINVDCx10_ASAP7_75t_R g1594 ( 
.A(n_1535),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1500),
.B(n_1464),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1495),
.B(n_1452),
.Y(n_1596)
);

INVxp67_ASAP7_75t_L g1597 ( 
.A(n_1513),
.Y(n_1597)
);

AOI211xp5_ASAP7_75t_L g1598 ( 
.A1(n_1556),
.A2(n_1467),
.B(n_1422),
.C(n_1471),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1521),
.B(n_1522),
.Y(n_1599)
);

AOI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1532),
.A2(n_1485),
.B1(n_1480),
.B2(n_1476),
.Y(n_1600)
);

INVx4_ASAP7_75t_L g1601 ( 
.A(n_1585),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1521),
.B(n_1374),
.Y(n_1602)
);

AND2x2_ASAP7_75t_L g1603 ( 
.A(n_1522),
.B(n_1379),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1560),
.B(n_1368),
.Y(n_1604)
);

O2A1O1Ixp33_ASAP7_75t_L g1605 ( 
.A1(n_1545),
.A2(n_1461),
.B(n_1566),
.C(n_1543),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1560),
.B(n_1561),
.Y(n_1606)
);

AO21x2_ASAP7_75t_L g1607 ( 
.A1(n_1494),
.A2(n_1518),
.B(n_1516),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1561),
.B(n_1514),
.Y(n_1608)
);

AO21x2_ASAP7_75t_L g1609 ( 
.A1(n_1518),
.A2(n_1516),
.B(n_1541),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1502),
.B(n_1551),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1498),
.B(n_1504),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1502),
.B(n_1551),
.Y(n_1612)
);

OAI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1538),
.A2(n_1532),
.B1(n_1550),
.B2(n_1568),
.Y(n_1613)
);

BUFx2_ASAP7_75t_L g1614 ( 
.A(n_1585),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1499),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1554),
.B(n_1558),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1506),
.B(n_1542),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1554),
.B(n_1558),
.Y(n_1618)
);

HB1xp67_ASAP7_75t_L g1619 ( 
.A(n_1525),
.Y(n_1619)
);

BUFx3_ASAP7_75t_L g1620 ( 
.A(n_1580),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1496),
.B(n_1539),
.Y(n_1621)
);

NOR3xp33_ASAP7_75t_SL g1622 ( 
.A(n_1590),
.B(n_1586),
.C(n_1578),
.Y(n_1622)
);

AOI21xp5_ASAP7_75t_L g1623 ( 
.A1(n_1544),
.A2(n_1509),
.B(n_1512),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1539),
.B(n_1540),
.Y(n_1624)
);

AOI21xp5_ASAP7_75t_L g1625 ( 
.A1(n_1544),
.A2(n_1509),
.B(n_1553),
.Y(n_1625)
);

NOR2x1_ASAP7_75t_L g1626 ( 
.A(n_1585),
.B(n_1528),
.Y(n_1626)
);

INVxp67_ASAP7_75t_L g1627 ( 
.A(n_1563),
.Y(n_1627)
);

OA21x2_ASAP7_75t_L g1628 ( 
.A1(n_1557),
.A2(n_1541),
.B(n_1555),
.Y(n_1628)
);

OR2x2_ASAP7_75t_L g1629 ( 
.A(n_1523),
.B(n_1534),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1507),
.B(n_1529),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1507),
.B(n_1529),
.Y(n_1631)
);

AOI22xp5_ASAP7_75t_SL g1632 ( 
.A1(n_1562),
.A2(n_1528),
.B1(n_1547),
.B2(n_1546),
.Y(n_1632)
);

AO21x1_ASAP7_75t_L g1633 ( 
.A1(n_1568),
.A2(n_1531),
.B(n_1549),
.Y(n_1633)
);

CKINVDCx5p33_ASAP7_75t_R g1634 ( 
.A(n_1527),
.Y(n_1634)
);

OAI21xp5_ASAP7_75t_L g1635 ( 
.A1(n_1549),
.A2(n_1571),
.B(n_1550),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1493),
.Y(n_1636)
);

AO32x2_ASAP7_75t_L g1637 ( 
.A1(n_1552),
.A2(n_1567),
.A3(n_1508),
.B1(n_1501),
.B2(n_1515),
.Y(n_1637)
);

BUFx4f_ASAP7_75t_SL g1638 ( 
.A(n_1517),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1536),
.B(n_1544),
.Y(n_1639)
);

AND2x4_ASAP7_75t_L g1640 ( 
.A(n_1569),
.B(n_1570),
.Y(n_1640)
);

AOI21xp5_ASAP7_75t_L g1641 ( 
.A1(n_1544),
.A2(n_1509),
.B(n_1553),
.Y(n_1641)
);

OAI21xp5_ASAP7_75t_L g1642 ( 
.A1(n_1571),
.A2(n_1536),
.B(n_1576),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1573),
.B(n_1509),
.Y(n_1643)
);

OA21x2_ASAP7_75t_L g1644 ( 
.A1(n_1493),
.A2(n_1511),
.B(n_1510),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1531),
.B(n_1573),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1526),
.B(n_1530),
.Y(n_1646)
);

HB1xp67_ASAP7_75t_L g1647 ( 
.A(n_1526),
.Y(n_1647)
);

BUFx3_ASAP7_75t_L g1648 ( 
.A(n_1580),
.Y(n_1648)
);

HB1xp67_ASAP7_75t_L g1649 ( 
.A(n_1619),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_SL g1650 ( 
.A(n_1605),
.B(n_1528),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1610),
.B(n_1497),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1611),
.B(n_1520),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1636),
.Y(n_1653)
);

HB1xp67_ASAP7_75t_L g1654 ( 
.A(n_1647),
.Y(n_1654)
);

HB1xp67_ASAP7_75t_L g1655 ( 
.A(n_1629),
.Y(n_1655)
);

NAND2xp67_ASAP7_75t_L g1656 ( 
.A(n_1604),
.B(n_1582),
.Y(n_1656)
);

INVx1_ASAP7_75t_SL g1657 ( 
.A(n_1594),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1644),
.Y(n_1658)
);

AOI22xp33_ASAP7_75t_L g1659 ( 
.A1(n_1635),
.A2(n_1553),
.B1(n_1505),
.B2(n_1546),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1643),
.B(n_1503),
.Y(n_1660)
);

NAND4xp25_ASAP7_75t_L g1661 ( 
.A(n_1598),
.B(n_1584),
.C(n_1537),
.D(n_1505),
.Y(n_1661)
);

INVx1_ASAP7_75t_SL g1662 ( 
.A(n_1595),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1644),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1621),
.B(n_1520),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1624),
.B(n_1520),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1643),
.B(n_1520),
.Y(n_1666)
);

AND2x4_ASAP7_75t_L g1667 ( 
.A(n_1620),
.B(n_1564),
.Y(n_1667)
);

OR2x6_ASAP7_75t_L g1668 ( 
.A(n_1625),
.B(n_1581),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1612),
.B(n_1520),
.Y(n_1669)
);

INVxp67_ASAP7_75t_L g1670 ( 
.A(n_1617),
.Y(n_1670)
);

BUFx2_ASAP7_75t_L g1671 ( 
.A(n_1637),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1615),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1615),
.Y(n_1673)
);

BUFx2_ASAP7_75t_L g1674 ( 
.A(n_1637),
.Y(n_1674)
);

NOR2xp33_ASAP7_75t_L g1675 ( 
.A(n_1596),
.B(n_1547),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1597),
.B(n_1533),
.Y(n_1676)
);

AOI22xp5_ASAP7_75t_L g1677 ( 
.A1(n_1613),
.A2(n_1537),
.B1(n_1582),
.B2(n_1575),
.Y(n_1677)
);

AOI22xp5_ASAP7_75t_L g1678 ( 
.A1(n_1622),
.A2(n_1572),
.B1(n_1589),
.B2(n_1517),
.Y(n_1678)
);

OAI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1632),
.A2(n_1600),
.B1(n_1604),
.B2(n_1602),
.Y(n_1679)
);

INVx4_ASAP7_75t_L g1680 ( 
.A(n_1638),
.Y(n_1680)
);

AND2x2_ASAP7_75t_SL g1681 ( 
.A(n_1639),
.B(n_1559),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1612),
.B(n_1639),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1646),
.Y(n_1683)
);

BUFx6f_ASAP7_75t_L g1684 ( 
.A(n_1648),
.Y(n_1684)
);

INVx2_ASAP7_75t_SL g1685 ( 
.A(n_1640),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1666),
.B(n_1609),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1682),
.B(n_1628),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1672),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1658),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1682),
.B(n_1628),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1671),
.B(n_1628),
.Y(n_1691)
);

OAI33xp33_ASAP7_75t_L g1692 ( 
.A1(n_1679),
.A2(n_1645),
.A3(n_1519),
.B1(n_1548),
.B2(n_1579),
.B3(n_1627),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1672),
.Y(n_1693)
);

BUFx6f_ASAP7_75t_L g1694 ( 
.A(n_1684),
.Y(n_1694)
);

INVxp67_ASAP7_75t_L g1695 ( 
.A(n_1654),
.Y(n_1695)
);

AOI221xp5_ASAP7_75t_L g1696 ( 
.A1(n_1659),
.A2(n_1642),
.B1(n_1633),
.B2(n_1641),
.C(n_1631),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1671),
.B(n_1616),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1674),
.B(n_1616),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1674),
.B(n_1618),
.Y(n_1699)
);

NAND4xp25_ASAP7_75t_L g1700 ( 
.A(n_1661),
.B(n_1603),
.C(n_1602),
.D(n_1623),
.Y(n_1700)
);

NOR2xp33_ASAP7_75t_L g1701 ( 
.A(n_1680),
.B(n_1638),
.Y(n_1701)
);

HB1xp67_ASAP7_75t_L g1702 ( 
.A(n_1663),
.Y(n_1702)
);

OAI33xp33_ASAP7_75t_L g1703 ( 
.A1(n_1652),
.A2(n_1650),
.A3(n_1664),
.B1(n_1665),
.B2(n_1676),
.B3(n_1670),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1681),
.B(n_1614),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1681),
.B(n_1630),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1655),
.B(n_1631),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1673),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1673),
.Y(n_1708)
);

BUFx2_ASAP7_75t_L g1709 ( 
.A(n_1684),
.Y(n_1709)
);

OAI22xp5_ASAP7_75t_L g1710 ( 
.A1(n_1677),
.A2(n_1599),
.B1(n_1603),
.B2(n_1606),
.Y(n_1710)
);

OAI22xp33_ASAP7_75t_L g1711 ( 
.A1(n_1678),
.A2(n_1591),
.B1(n_1581),
.B2(n_1626),
.Y(n_1711)
);

AOI221xp5_ASAP7_75t_L g1712 ( 
.A1(n_1669),
.A2(n_1633),
.B1(n_1606),
.B2(n_1608),
.C(n_1599),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1683),
.B(n_1607),
.Y(n_1713)
);

BUFx3_ASAP7_75t_L g1714 ( 
.A(n_1680),
.Y(n_1714)
);

INVx5_ASAP7_75t_L g1715 ( 
.A(n_1668),
.Y(n_1715)
);

NOR2x1_ASAP7_75t_L g1716 ( 
.A(n_1668),
.B(n_1601),
.Y(n_1716)
);

INVx4_ASAP7_75t_L g1717 ( 
.A(n_1680),
.Y(n_1717)
);

NAND3xp33_ASAP7_75t_L g1718 ( 
.A(n_1649),
.B(n_1675),
.C(n_1601),
.Y(n_1718)
);

INVx4_ASAP7_75t_L g1719 ( 
.A(n_1684),
.Y(n_1719)
);

NOR3xp33_ASAP7_75t_L g1720 ( 
.A(n_1657),
.B(n_1579),
.C(n_1588),
.Y(n_1720)
);

BUFx3_ASAP7_75t_L g1721 ( 
.A(n_1714),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1695),
.B(n_1669),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1695),
.B(n_1651),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1688),
.Y(n_1724)
);

NAND3xp33_ASAP7_75t_SL g1725 ( 
.A(n_1696),
.B(n_1662),
.C(n_1634),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1705),
.B(n_1697),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1705),
.B(n_1685),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1697),
.B(n_1684),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1688),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1687),
.B(n_1668),
.Y(n_1730)
);

OR2x2_ASAP7_75t_L g1731 ( 
.A(n_1686),
.B(n_1698),
.Y(n_1731)
);

BUFx2_ASAP7_75t_L g1732 ( 
.A(n_1719),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1693),
.Y(n_1733)
);

INVx3_ASAP7_75t_L g1734 ( 
.A(n_1694),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1687),
.B(n_1668),
.Y(n_1735)
);

HB1xp67_ASAP7_75t_L g1736 ( 
.A(n_1702),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1693),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1707),
.Y(n_1738)
);

NOR2xp33_ASAP7_75t_L g1739 ( 
.A(n_1701),
.B(n_1634),
.Y(n_1739)
);

INVxp67_ASAP7_75t_L g1740 ( 
.A(n_1703),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1707),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1689),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1708),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1689),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1689),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1699),
.B(n_1667),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1704),
.B(n_1687),
.Y(n_1747)
);

INVx2_ASAP7_75t_SL g1748 ( 
.A(n_1694),
.Y(n_1748)
);

INVx1_ASAP7_75t_SL g1749 ( 
.A(n_1709),
.Y(n_1749)
);

AND2x4_ASAP7_75t_L g1750 ( 
.A(n_1715),
.B(n_1667),
.Y(n_1750)
);

NOR2xp33_ASAP7_75t_L g1751 ( 
.A(n_1717),
.B(n_1577),
.Y(n_1751)
);

OR2x2_ASAP7_75t_L g1752 ( 
.A(n_1718),
.B(n_1660),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1712),
.B(n_1653),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1724),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1726),
.B(n_1690),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1742),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1730),
.B(n_1691),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1724),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1729),
.Y(n_1759)
);

INVx1_ASAP7_75t_SL g1760 ( 
.A(n_1732),
.Y(n_1760)
);

OR2x2_ASAP7_75t_L g1761 ( 
.A(n_1753),
.B(n_1752),
.Y(n_1761)
);

HB1xp67_ASAP7_75t_L g1762 ( 
.A(n_1736),
.Y(n_1762)
);

INVx3_ASAP7_75t_L g1763 ( 
.A(n_1750),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1729),
.Y(n_1764)
);

AND2x2_ASAP7_75t_L g1765 ( 
.A(n_1730),
.B(n_1691),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1742),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1730),
.B(n_1691),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1742),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1733),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1733),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1737),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1737),
.Y(n_1772)
);

OR2x2_ASAP7_75t_L g1773 ( 
.A(n_1753),
.B(n_1718),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1744),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1735),
.B(n_1715),
.Y(n_1775)
);

OR2x2_ASAP7_75t_L g1776 ( 
.A(n_1752),
.B(n_1713),
.Y(n_1776)
);

HB1xp67_ASAP7_75t_L g1777 ( 
.A(n_1736),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1744),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1740),
.B(n_1712),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1744),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1738),
.Y(n_1781)
);

INVx1_ASAP7_75t_SL g1782 ( 
.A(n_1732),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1738),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1741),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1745),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1735),
.B(n_1715),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_L g1787 ( 
.A(n_1740),
.B(n_1706),
.Y(n_1787)
);

OR2x2_ASAP7_75t_L g1788 ( 
.A(n_1722),
.B(n_1713),
.Y(n_1788)
);

INVx3_ASAP7_75t_L g1789 ( 
.A(n_1750),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1741),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1743),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1722),
.B(n_1706),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1743),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1745),
.Y(n_1794)
);

INVxp67_ASAP7_75t_L g1795 ( 
.A(n_1721),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1745),
.Y(n_1796)
);

AND2x4_ASAP7_75t_L g1797 ( 
.A(n_1750),
.B(n_1715),
.Y(n_1797)
);

INVx1_ASAP7_75t_SL g1798 ( 
.A(n_1749),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1775),
.B(n_1726),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1762),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1779),
.B(n_1721),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1775),
.B(n_1721),
.Y(n_1802)
);

HB1xp67_ASAP7_75t_L g1803 ( 
.A(n_1762),
.Y(n_1803)
);

OR2x2_ASAP7_75t_L g1804 ( 
.A(n_1787),
.B(n_1725),
.Y(n_1804)
);

OR2x2_ASAP7_75t_L g1805 ( 
.A(n_1787),
.B(n_1761),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1775),
.B(n_1747),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1779),
.B(n_1720),
.Y(n_1807)
);

OAI32xp33_ASAP7_75t_L g1808 ( 
.A1(n_1773),
.A2(n_1700),
.A3(n_1749),
.B1(n_1731),
.B2(n_1725),
.Y(n_1808)
);

INVx3_ASAP7_75t_L g1809 ( 
.A(n_1763),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1777),
.Y(n_1810)
);

A2O1A1Ixp33_ASAP7_75t_L g1811 ( 
.A1(n_1773),
.A2(n_1696),
.B(n_1700),
.C(n_1751),
.Y(n_1811)
);

OR2x2_ASAP7_75t_L g1812 ( 
.A(n_1761),
.B(n_1723),
.Y(n_1812)
);

NOR3xp33_ASAP7_75t_L g1813 ( 
.A(n_1795),
.B(n_1711),
.C(n_1703),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1795),
.B(n_1720),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1777),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1754),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1798),
.B(n_1760),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1786),
.B(n_1747),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1754),
.Y(n_1819)
);

OAI21xp33_ASAP7_75t_L g1820 ( 
.A1(n_1798),
.A2(n_1735),
.B(n_1656),
.Y(n_1820)
);

OR2x2_ASAP7_75t_L g1821 ( 
.A(n_1792),
.B(n_1723),
.Y(n_1821)
);

NOR2x1_ASAP7_75t_L g1822 ( 
.A(n_1760),
.B(n_1714),
.Y(n_1822)
);

INVxp67_ASAP7_75t_SL g1823 ( 
.A(n_1756),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1758),
.Y(n_1824)
);

INVx1_ASAP7_75t_SL g1825 ( 
.A(n_1782),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1782),
.B(n_1746),
.Y(n_1826)
);

AND2x4_ASAP7_75t_L g1827 ( 
.A(n_1786),
.B(n_1750),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1792),
.B(n_1746),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1786),
.B(n_1728),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1758),
.Y(n_1830)
);

NAND2x1p5_ASAP7_75t_L g1831 ( 
.A(n_1797),
.B(n_1715),
.Y(n_1831)
);

NAND2xp33_ASAP7_75t_SL g1832 ( 
.A(n_1797),
.B(n_1717),
.Y(n_1832)
);

INVx2_ASAP7_75t_SL g1833 ( 
.A(n_1763),
.Y(n_1833)
);

NAND2x1p5_ASAP7_75t_L g1834 ( 
.A(n_1797),
.B(n_1715),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1757),
.B(n_1727),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1809),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1803),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1803),
.Y(n_1838)
);

AOI222xp33_ASAP7_75t_L g1839 ( 
.A1(n_1807),
.A2(n_1692),
.B1(n_1710),
.B2(n_1739),
.C1(n_1714),
.C2(n_1717),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1800),
.B(n_1759),
.Y(n_1840)
);

OAI22xp5_ASAP7_75t_L g1841 ( 
.A1(n_1811),
.A2(n_1710),
.B1(n_1715),
.B2(n_1704),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1829),
.B(n_1797),
.Y(n_1842)
);

OR2x2_ASAP7_75t_L g1843 ( 
.A(n_1805),
.B(n_1776),
.Y(n_1843)
);

NAND2xp5_ASAP7_75t_L g1844 ( 
.A(n_1825),
.B(n_1757),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1816),
.Y(n_1845)
);

INVx1_ASAP7_75t_SL g1846 ( 
.A(n_1822),
.Y(n_1846)
);

AOI22xp5_ASAP7_75t_L g1847 ( 
.A1(n_1811),
.A2(n_1692),
.B1(n_1716),
.B2(n_1717),
.Y(n_1847)
);

OR2x2_ASAP7_75t_L g1848 ( 
.A(n_1801),
.B(n_1776),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1819),
.Y(n_1849)
);

AOI22xp5_ASAP7_75t_L g1850 ( 
.A1(n_1813),
.A2(n_1716),
.B1(n_1763),
.B2(n_1789),
.Y(n_1850)
);

AND2x4_ASAP7_75t_L g1851 ( 
.A(n_1802),
.B(n_1763),
.Y(n_1851)
);

OR2x2_ASAP7_75t_L g1852 ( 
.A(n_1817),
.B(n_1788),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1799),
.B(n_1789),
.Y(n_1853)
);

INVxp67_ASAP7_75t_L g1854 ( 
.A(n_1814),
.Y(n_1854)
);

OAI222xp33_ASAP7_75t_L g1855 ( 
.A1(n_1804),
.A2(n_1789),
.B1(n_1767),
.B2(n_1765),
.C1(n_1757),
.C2(n_1788),
.Y(n_1855)
);

OAI221xp5_ASAP7_75t_L g1856 ( 
.A1(n_1820),
.A2(n_1789),
.B1(n_1759),
.B2(n_1769),
.C(n_1793),
.Y(n_1856)
);

INVx2_ASAP7_75t_L g1857 ( 
.A(n_1809),
.Y(n_1857)
);

OAI21xp5_ASAP7_75t_L g1858 ( 
.A1(n_1808),
.A2(n_1748),
.B(n_1734),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1813),
.B(n_1765),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1827),
.B(n_1765),
.Y(n_1860)
);

AOI22xp5_ASAP7_75t_L g1861 ( 
.A1(n_1827),
.A2(n_1767),
.B1(n_1748),
.B2(n_1728),
.Y(n_1861)
);

O2A1O1Ixp33_ASAP7_75t_L g1862 ( 
.A1(n_1810),
.A2(n_1815),
.B(n_1834),
.C(n_1831),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1837),
.Y(n_1863)
);

INVx1_ASAP7_75t_SL g1864 ( 
.A(n_1846),
.Y(n_1864)
);

INVxp67_ASAP7_75t_SL g1865 ( 
.A(n_1862),
.Y(n_1865)
);

XNOR2xp5_ASAP7_75t_L g1866 ( 
.A(n_1841),
.B(n_1656),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1838),
.Y(n_1867)
);

A2O1A1Ixp33_ASAP7_75t_L g1868 ( 
.A1(n_1841),
.A2(n_1832),
.B(n_1812),
.C(n_1827),
.Y(n_1868)
);

NOR2xp33_ASAP7_75t_L g1869 ( 
.A(n_1854),
.B(n_1826),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1845),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1849),
.Y(n_1871)
);

OAI21xp5_ASAP7_75t_SL g1872 ( 
.A1(n_1839),
.A2(n_1834),
.B(n_1831),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1840),
.Y(n_1873)
);

AOI22xp5_ASAP7_75t_L g1874 ( 
.A1(n_1839),
.A2(n_1832),
.B1(n_1818),
.B2(n_1806),
.Y(n_1874)
);

INVx1_ASAP7_75t_SL g1875 ( 
.A(n_1846),
.Y(n_1875)
);

INVxp67_ASAP7_75t_SL g1876 ( 
.A(n_1844),
.Y(n_1876)
);

NOR2xp33_ASAP7_75t_L g1877 ( 
.A(n_1859),
.B(n_1806),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1860),
.B(n_1851),
.Y(n_1878)
);

NOR2xp67_ASAP7_75t_SL g1879 ( 
.A(n_1858),
.B(n_1524),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1851),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1842),
.B(n_1818),
.Y(n_1881)
);

NAND3xp33_ASAP7_75t_SL g1882 ( 
.A(n_1850),
.B(n_1835),
.C(n_1821),
.Y(n_1882)
);

NAND3xp33_ASAP7_75t_SL g1883 ( 
.A(n_1847),
.B(n_1830),
.C(n_1824),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1848),
.B(n_1828),
.Y(n_1884)
);

OAI221xp5_ASAP7_75t_L g1885 ( 
.A1(n_1872),
.A2(n_1858),
.B1(n_1856),
.B2(n_1861),
.C(n_1852),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1864),
.B(n_1853),
.Y(n_1886)
);

AOI21xp33_ASAP7_75t_L g1887 ( 
.A1(n_1865),
.A2(n_1843),
.B(n_1836),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1863),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1881),
.B(n_1857),
.Y(n_1889)
);

INVxp67_ASAP7_75t_L g1890 ( 
.A(n_1877),
.Y(n_1890)
);

AOI221xp5_ASAP7_75t_L g1891 ( 
.A1(n_1883),
.A2(n_1855),
.B1(n_1840),
.B2(n_1833),
.C(n_1823),
.Y(n_1891)
);

OR2x2_ASAP7_75t_L g1892 ( 
.A(n_1875),
.B(n_1833),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1877),
.B(n_1767),
.Y(n_1893)
);

AOI21xp33_ASAP7_75t_L g1894 ( 
.A1(n_1874),
.A2(n_1823),
.B(n_1809),
.Y(n_1894)
);

INVxp67_ASAP7_75t_SL g1895 ( 
.A(n_1879),
.Y(n_1895)
);

INVx3_ASAP7_75t_L g1896 ( 
.A(n_1880),
.Y(n_1896)
);

OAI221xp5_ASAP7_75t_SL g1897 ( 
.A1(n_1868),
.A2(n_1866),
.B1(n_1878),
.B2(n_1876),
.C(n_1869),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1867),
.Y(n_1898)
);

NAND3xp33_ASAP7_75t_L g1899 ( 
.A(n_1891),
.B(n_1897),
.C(n_1894),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1896),
.B(n_1880),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1896),
.B(n_1869),
.Y(n_1901)
);

AOI21xp33_ASAP7_75t_L g1902 ( 
.A1(n_1895),
.A2(n_1868),
.B(n_1873),
.Y(n_1902)
);

OR3x1_ASAP7_75t_L g1903 ( 
.A(n_1887),
.B(n_1882),
.C(n_1871),
.Y(n_1903)
);

INVx2_ASAP7_75t_L g1904 ( 
.A(n_1892),
.Y(n_1904)
);

NAND3xp33_ASAP7_75t_SL g1905 ( 
.A(n_1885),
.B(n_1884),
.C(n_1870),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_SL g1906 ( 
.A(n_1886),
.B(n_1748),
.Y(n_1906)
);

NOR2xp33_ASAP7_75t_L g1907 ( 
.A(n_1890),
.B(n_1592),
.Y(n_1907)
);

NAND2xp33_ASAP7_75t_L g1908 ( 
.A(n_1893),
.B(n_1734),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1889),
.B(n_1755),
.Y(n_1909)
);

NOR2x1_ASAP7_75t_L g1910 ( 
.A(n_1903),
.B(n_1888),
.Y(n_1910)
);

NOR2x1_ASAP7_75t_L g1911 ( 
.A(n_1899),
.B(n_1898),
.Y(n_1911)
);

OAI321xp33_ASAP7_75t_L g1912 ( 
.A1(n_1905),
.A2(n_1894),
.A3(n_1694),
.B1(n_1587),
.B2(n_1794),
.C(n_1796),
.Y(n_1912)
);

AOI211xp5_ASAP7_75t_SL g1913 ( 
.A1(n_1902),
.A2(n_1734),
.B(n_1583),
.C(n_1771),
.Y(n_1913)
);

OAI21xp5_ASAP7_75t_L g1914 ( 
.A1(n_1901),
.A2(n_1734),
.B(n_1764),
.Y(n_1914)
);

OAI21xp33_ASAP7_75t_L g1915 ( 
.A1(n_1909),
.A2(n_1766),
.B(n_1756),
.Y(n_1915)
);

O2A1O1Ixp33_ASAP7_75t_L g1916 ( 
.A1(n_1900),
.A2(n_1524),
.B(n_1756),
.C(n_1794),
.Y(n_1916)
);

OAI221xp5_ASAP7_75t_SL g1917 ( 
.A1(n_1916),
.A2(n_1904),
.B1(n_1907),
.B2(n_1908),
.C(n_1906),
.Y(n_1917)
);

AOI221xp5_ASAP7_75t_SL g1918 ( 
.A1(n_1914),
.A2(n_1796),
.B1(n_1766),
.B2(n_1794),
.C(n_1768),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1910),
.Y(n_1919)
);

AOI211xp5_ASAP7_75t_L g1920 ( 
.A1(n_1912),
.A2(n_1565),
.B(n_1574),
.C(n_1589),
.Y(n_1920)
);

AOI211xp5_ASAP7_75t_SL g1921 ( 
.A1(n_1915),
.A2(n_1764),
.B(n_1769),
.C(n_1793),
.Y(n_1921)
);

OAI211xp5_ASAP7_75t_SL g1922 ( 
.A1(n_1911),
.A2(n_1796),
.B(n_1766),
.C(n_1768),
.Y(n_1922)
);

BUFx4f_ASAP7_75t_L g1923 ( 
.A(n_1913),
.Y(n_1923)
);

OAI221xp5_ASAP7_75t_L g1924 ( 
.A1(n_1919),
.A2(n_1774),
.B1(n_1768),
.B2(n_1778),
.C(n_1785),
.Y(n_1924)
);

NOR2x1_ASAP7_75t_L g1925 ( 
.A(n_1922),
.B(n_1923),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1917),
.Y(n_1926)
);

NOR2x1_ASAP7_75t_L g1927 ( 
.A(n_1921),
.B(n_1565),
.Y(n_1927)
);

OAI221xp5_ASAP7_75t_L g1928 ( 
.A1(n_1920),
.A2(n_1778),
.B1(n_1774),
.B2(n_1780),
.C(n_1785),
.Y(n_1928)
);

NOR2x1_ASAP7_75t_L g1929 ( 
.A(n_1918),
.B(n_1574),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1925),
.Y(n_1930)
);

AOI221x1_ASAP7_75t_L g1931 ( 
.A1(n_1926),
.A2(n_1927),
.B1(n_1929),
.B2(n_1924),
.C(n_1784),
.Y(n_1931)
);

NOR3xp33_ASAP7_75t_L g1932 ( 
.A(n_1928),
.B(n_1719),
.C(n_1774),
.Y(n_1932)
);

INVxp67_ASAP7_75t_SL g1933 ( 
.A(n_1930),
.Y(n_1933)
);

AOI22xp5_ASAP7_75t_L g1934 ( 
.A1(n_1933),
.A2(n_1932),
.B1(n_1931),
.B2(n_1778),
.Y(n_1934)
);

AOI21xp33_ASAP7_75t_SL g1935 ( 
.A1(n_1934),
.A2(n_1785),
.B(n_1780),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1934),
.Y(n_1936)
);

OAI31xp33_ASAP7_75t_L g1937 ( 
.A1(n_1936),
.A2(n_1770),
.A3(n_1791),
.B(n_1790),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1935),
.B(n_1770),
.Y(n_1938)
);

OAI22xp5_ASAP7_75t_SL g1939 ( 
.A1(n_1938),
.A2(n_1587),
.B1(n_1591),
.B2(n_1780),
.Y(n_1939)
);

XNOR2xp5_ASAP7_75t_L g1940 ( 
.A(n_1937),
.B(n_1593),
.Y(n_1940)
);

AND2x4_ASAP7_75t_L g1941 ( 
.A(n_1940),
.B(n_1771),
.Y(n_1941)
);

OAI21xp5_ASAP7_75t_L g1942 ( 
.A1(n_1941),
.A2(n_1939),
.B(n_1781),
.Y(n_1942)
);

AOI21xp33_ASAP7_75t_L g1943 ( 
.A1(n_1942),
.A2(n_1781),
.B(n_1772),
.Y(n_1943)
);

AOI22xp5_ASAP7_75t_L g1944 ( 
.A1(n_1943),
.A2(n_1791),
.B1(n_1790),
.B2(n_1784),
.Y(n_1944)
);

AOI211xp5_ASAP7_75t_L g1945 ( 
.A1(n_1944),
.A2(n_1587),
.B(n_1783),
.C(n_1772),
.Y(n_1945)
);


endmodule