module fake_jpeg_23391_n_267 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_267);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_267;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_37),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_38),
.B(n_33),
.Y(n_44)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_26),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_42),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_24),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_33),
.B1(n_26),
.B2(n_20),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_43),
.A2(n_46),
.B1(n_53),
.B2(n_55),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_62),
.Y(n_75)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_48),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_35),
.A2(n_33),
.B1(n_29),
.B2(n_18),
.Y(n_46)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_30),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_22),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_35),
.A2(n_32),
.B1(n_18),
.B2(n_28),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_52),
.A2(n_54),
.B1(n_56),
.B2(n_60),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_35),
.A2(n_21),
.B1(n_27),
.B2(n_32),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_39),
.A2(n_32),
.B1(n_18),
.B2(n_28),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_27),
.B1(n_21),
.B2(n_29),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_38),
.B1(n_27),
.B2(n_21),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_28),
.Y(n_58)
);

OR2x2_ASAP7_75t_SL g89 ( 
.A(n_58),
.B(n_31),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_39),
.A2(n_30),
.B1(n_17),
.B2(n_29),
.Y(n_60)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_39),
.A2(n_30),
.B1(n_17),
.B2(n_31),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_63),
.A2(n_34),
.B1(n_42),
.B2(n_37),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_19),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_64),
.B(n_42),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_22),
.C(n_19),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_24),
.C(n_25),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_59),
.B(n_42),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_66),
.B(n_70),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_68),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_60),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_69),
.B(n_74),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_51),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_72),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_73),
.A2(n_92),
.B1(n_0),
.B2(n_1),
.Y(n_128)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_77),
.B(n_83),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_57),
.A2(n_34),
.B1(n_25),
.B2(n_31),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_37),
.Y(n_79)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_47),
.B(n_36),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_37),
.Y(n_84)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_84),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_85),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_36),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_91),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_40),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_88),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_44),
.B(n_10),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_89),
.B(n_97),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_60),
.B(n_10),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_95),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_53),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_58),
.A2(n_31),
.B1(n_23),
.B2(n_34),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_93),
.A2(n_94),
.B1(n_82),
.B2(n_48),
.Y(n_114)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_55),
.B(n_0),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_58),
.B(n_8),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_97),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_58),
.B(n_23),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_57),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_63),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_99),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_100),
.Y(n_106)
);

O2A1O1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_55),
.A2(n_46),
.B(n_56),
.C(n_43),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_101),
.A2(n_62),
.B(n_61),
.C(n_49),
.Y(n_112)
);

NOR2xp67_ASAP7_75t_R g110 ( 
.A(n_89),
.B(n_43),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_110),
.A2(n_112),
.B(n_124),
.Y(n_156)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_120),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_114),
.A2(n_121),
.B1(n_103),
.B2(n_127),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_93),
.A2(n_48),
.B1(n_61),
.B2(n_49),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

INVx2_ASAP7_75t_SL g120 ( 
.A(n_85),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_68),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_125),
.A2(n_95),
.B(n_69),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_128),
.A2(n_122),
.B1(n_117),
.B2(n_118),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_87),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_150),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_131),
.A2(n_149),
.B1(n_4),
.B2(n_5),
.Y(n_182)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_109),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_132),
.B(n_137),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_112),
.A2(n_80),
.B(n_86),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_133),
.A2(n_136),
.B(n_138),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_134),
.A2(n_140),
.B1(n_147),
.B2(n_135),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_124),
.B(n_97),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_109),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_L g138 ( 
.A1(n_108),
.A2(n_70),
.B(n_79),
.C(n_71),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_127),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_139),
.B(n_152),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_112),
.A2(n_71),
.B1(n_101),
.B2(n_80),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_108),
.A2(n_66),
.B(n_96),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_141),
.A2(n_144),
.B(n_145),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_127),
.A2(n_99),
.B1(n_75),
.B2(n_90),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_142),
.A2(n_158),
.B1(n_159),
.B2(n_5),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_104),
.B(n_74),
.C(n_75),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_115),
.C(n_106),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_116),
.A2(n_83),
.B(n_88),
.Y(n_144)
);

OAI21xp33_ASAP7_75t_L g145 ( 
.A1(n_102),
.A2(n_116),
.B(n_105),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_107),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_146),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_117),
.A2(n_104),
.B1(n_110),
.B2(n_107),
.Y(n_147)
);

AO21x1_ASAP7_75t_L g148 ( 
.A1(n_123),
.A2(n_73),
.B(n_67),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_148),
.A2(n_122),
.B(n_113),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_120),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_84),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_77),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_76),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_157),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_105),
.B(n_10),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_154),
.B(n_11),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_118),
.B(n_100),
.Y(n_155)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_155),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_113),
.B(n_85),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_128),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_151),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_161),
.B(n_171),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_162),
.A2(n_166),
.B1(n_182),
.B2(n_142),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_156),
.A2(n_113),
.B(n_126),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_163),
.A2(n_165),
.B(n_136),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_132),
.A2(n_122),
.B1(n_126),
.B2(n_120),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_168),
.C(n_181),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_106),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_130),
.B(n_11),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_173),
.B(n_175),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_149),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_174),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_133),
.B(n_12),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_137),
.B(n_111),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_178),
.B(n_180),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_158),
.A2(n_115),
.B1(n_111),
.B2(n_3),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_179),
.A2(n_183),
.B1(n_154),
.B2(n_134),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_150),
.B(n_4),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_157),
.B(n_4),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_146),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_185),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_155),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_186),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_191),
.A2(n_161),
.B1(n_172),
.B2(n_186),
.Y(n_218)
);

A2O1A1O1Ixp25_ASAP7_75t_L g192 ( 
.A1(n_160),
.A2(n_136),
.B(n_144),
.C(n_141),
.D(n_147),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_192),
.B(n_162),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_168),
.B(n_140),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_193),
.A2(n_207),
.B(n_163),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_169),
.B(n_143),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_195),
.B(n_199),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_143),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_200),
.C(n_204),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_205),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_167),
.B(n_136),
.C(n_145),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_166),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_179),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_149),
.Y(n_202)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_202),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_176),
.B(n_153),
.C(n_131),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_184),
.Y(n_205)
);

AOI21xp33_ASAP7_75t_L g206 ( 
.A1(n_176),
.A2(n_138),
.B(n_148),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_206),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_165),
.A2(n_139),
.B(n_148),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_160),
.B(n_152),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_181),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_211),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_212),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_164),
.Y(n_214)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_203),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_217),
.B(n_194),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_218),
.A2(n_219),
.B1(n_222),
.B2(n_224),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_201),
.A2(n_185),
.B1(n_164),
.B2(n_170),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_187),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_204),
.A2(n_170),
.B1(n_178),
.B2(n_138),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_223),
.B(n_226),
.C(n_197),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_207),
.A2(n_177),
.B(n_151),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_199),
.A2(n_175),
.B(n_159),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_225),
.A2(n_220),
.B1(n_218),
.B2(n_198),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_173),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_216),
.B(n_188),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_227),
.B(n_235),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_228),
.B(n_229),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_195),
.Y(n_229)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_231),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_205),
.Y(n_232)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_232),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_197),
.C(n_226),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_236),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_234),
.A2(n_224),
.B1(n_193),
.B2(n_222),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_208),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_213),
.B(n_193),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_200),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_223),
.Y(n_242)
);

NOR3xp33_ASAP7_75t_L g241 ( 
.A(n_239),
.B(n_225),
.C(n_210),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_230),
.Y(n_250)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_242),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_243),
.A2(n_248),
.B1(n_238),
.B2(n_6),
.Y(n_255)
);

OAI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_230),
.A2(n_192),
.B1(n_209),
.B2(n_3),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_250),
.A2(n_229),
.B1(n_240),
.B2(n_13),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_246),
.B(n_245),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_251),
.B(n_253),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_244),
.B(n_234),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_247),
.B(n_190),
.Y(n_253)
);

AO21x1_ASAP7_75t_L g254 ( 
.A1(n_248),
.A2(n_238),
.B(n_209),
.Y(n_254)
);

FAx1_ASAP7_75t_SL g258 ( 
.A(n_254),
.B(n_255),
.CI(n_252),
.CON(n_258),
.SN(n_258)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_257),
.A2(n_259),
.B1(n_5),
.B2(n_7),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_258),
.B(n_249),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_254),
.A2(n_240),
.B1(n_7),
.B2(n_13),
.Y(n_259)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_260),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_261),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_256),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_264),
.Y(n_265)
);

BUFx24_ASAP7_75t_SL g266 ( 
.A(n_265),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_266),
.B(n_263),
.Y(n_267)
);


endmodule