module fake_jpeg_31491_n_515 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_515);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_515;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_15),
.B(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_14),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_6),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_54),
.Y(n_104)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_55),
.Y(n_136)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_56),
.Y(n_141)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_58),
.B(n_68),
.Y(n_103)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_59),
.Y(n_138)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_61),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_21),
.B(n_1),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_62),
.B(n_99),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_21),
.B(n_17),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_63),
.B(n_79),
.Y(n_134)
);

INVx4_ASAP7_75t_SL g64 ( 
.A(n_19),
.Y(n_64)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_64),
.Y(n_156)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_65),
.Y(n_122)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_66),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_67),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_48),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_48),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_70),
.B(n_71),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_48),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_72),
.Y(n_140)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_73),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_19),
.Y(n_74)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_74),
.Y(n_121)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_76),
.Y(n_150)
);

BUFx12_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

BUFx4f_ASAP7_75t_SL g106 ( 
.A(n_77),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_78),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_24),
.B(n_1),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_31),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_80),
.B(n_82),
.Y(n_123)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_81),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_48),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_85),
.Y(n_125)
);

INVx13_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_86),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_34),
.Y(n_87)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_87),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_48),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_88),
.B(n_95),
.Y(n_135)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

NAND2xp33_ASAP7_75t_SL g90 ( 
.A(n_24),
.B(n_1),
.Y(n_90)
);

INVx4_ASAP7_75t_SL g146 ( 
.A(n_90),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_91),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_92),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_24),
.B(n_1),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_93),
.B(n_100),
.Y(n_115)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

INVx11_ASAP7_75t_L g151 ( 
.A(n_94),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_20),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_33),
.Y(n_96)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

INVx11_ASAP7_75t_L g158 ( 
.A(n_97),
.Y(n_158)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_23),
.Y(n_98)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_27),
.B(n_3),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_42),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_32),
.Y(n_101)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_101),
.Y(n_160)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_32),
.Y(n_102)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_99),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_112),
.B(n_113),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_74),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_87),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_119),
.B(n_155),
.Y(n_179)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_53),
.Y(n_137)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_137),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_62),
.B(n_26),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_139),
.B(n_145),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_75),
.Y(n_143)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_79),
.B(n_26),
.Y(n_145)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_57),
.Y(n_147)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_64),
.A2(n_42),
.B1(n_29),
.B2(n_50),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_148),
.A2(n_94),
.B1(n_102),
.B2(n_97),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_79),
.B(n_39),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_157),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g152 ( 
.A(n_86),
.Y(n_152)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_152),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_93),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_93),
.B(n_39),
.Y(n_157)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_61),
.Y(n_159)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_159),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_136),
.Y(n_164)
);

INVx4_ASAP7_75t_SL g219 ( 
.A(n_164),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_103),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_166),
.B(n_171),
.Y(n_228)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_151),
.Y(n_167)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_167),
.Y(n_261)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_111),
.Y(n_170)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_170),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_124),
.B(n_52),
.Y(n_171)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_116),
.Y(n_173)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_173),
.Y(n_224)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_107),
.Y(n_174)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_174),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_134),
.B(n_89),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_175),
.B(n_180),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_176),
.A2(n_199),
.B1(n_203),
.B2(n_109),
.Y(n_229)
);

OA22x2_ASAP7_75t_L g177 ( 
.A1(n_146),
.A2(n_90),
.B1(n_96),
.B2(n_66),
.Y(n_177)
);

AO22x1_ASAP7_75t_L g220 ( 
.A1(n_177),
.A2(n_152),
.B1(n_131),
.B2(n_143),
.Y(n_220)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_110),
.Y(n_178)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_178),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_123),
.B(n_77),
.Y(n_180)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_181),
.Y(n_233)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_114),
.Y(n_182)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_182),
.Y(n_258)
);

A2O1A1Ixp33_ASAP7_75t_L g183 ( 
.A1(n_146),
.A2(n_134),
.B(n_115),
.C(n_117),
.Y(n_183)
);

A2O1A1Ixp33_ASAP7_75t_L g216 ( 
.A1(n_183),
.A2(n_30),
.B(n_28),
.C(n_106),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_138),
.A2(n_101),
.B1(n_92),
.B2(n_65),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_184),
.A2(n_186),
.B1(n_213),
.B2(n_185),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_118),
.A2(n_67),
.B1(n_91),
.B2(n_85),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_185),
.A2(n_120),
.B1(n_125),
.B2(n_127),
.Y(n_234)
);

OAI22xp33_ASAP7_75t_L g186 ( 
.A1(n_158),
.A2(n_54),
.B1(n_84),
.B2(n_69),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_150),
.Y(n_187)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_187),
.Y(n_259)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_140),
.Y(n_188)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_188),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_121),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_189),
.Y(n_225)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_105),
.Y(n_190)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_190),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_153),
.B(n_37),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_194),
.Y(n_227)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_111),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_192),
.Y(n_253)
);

AND2x4_ASAP7_75t_L g193 ( 
.A(n_148),
.B(n_83),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_193),
.B(n_197),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_108),
.B(n_27),
.Y(n_194)
);

INVx13_ASAP7_75t_L g195 ( 
.A(n_156),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_195),
.B(n_196),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_135),
.B(n_77),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_128),
.A2(n_130),
.B1(n_43),
.B2(n_51),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_104),
.Y(n_198)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_198),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_144),
.A2(n_60),
.B1(n_56),
.B2(n_78),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_154),
.B(n_41),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_200),
.B(n_205),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_126),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_201),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_141),
.B(n_41),
.Y(n_203)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_105),
.Y(n_204)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_204),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_131),
.B(n_37),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_150),
.Y(n_206)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_206),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_133),
.A2(n_43),
.B1(n_33),
.B2(n_51),
.Y(n_207)
);

AOI32xp33_ASAP7_75t_L g218 ( 
.A1(n_207),
.A2(n_45),
.A3(n_35),
.B1(n_168),
.B2(n_179),
.Y(n_218)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_132),
.Y(n_208)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_208),
.Y(n_252)
);

INVx11_ASAP7_75t_L g209 ( 
.A(n_132),
.Y(n_209)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_209),
.Y(n_254)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_160),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_210),
.Y(n_222)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_160),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_211),
.Y(n_236)
);

CKINVDCx12_ASAP7_75t_R g212 ( 
.A(n_106),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_212),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_122),
.A2(n_76),
.B1(n_55),
.B2(n_36),
.Y(n_213)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_104),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_214),
.A2(n_118),
.B1(n_120),
.B2(n_125),
.Y(n_231)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_156),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_215),
.Y(n_240)
);

OR2x2_ASAP7_75t_SL g265 ( 
.A(n_216),
.B(n_202),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_SL g279 ( 
.A(n_218),
.B(n_250),
.C(n_131),
.Y(n_279)
);

AND2x4_ASAP7_75t_SL g280 ( 
.A(n_220),
.B(n_238),
.Y(n_280)
);

AOI22x1_ASAP7_75t_L g226 ( 
.A1(n_193),
.A2(n_177),
.B1(n_176),
.B2(n_183),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_226),
.A2(n_231),
.B1(n_243),
.B2(n_199),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_229),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_175),
.B(n_109),
.C(n_122),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_230),
.B(n_241),
.C(n_244),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g267 ( 
.A1(n_234),
.A2(n_247),
.B1(n_255),
.B2(n_257),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_193),
.A2(n_29),
.B1(n_127),
.B2(n_45),
.Y(n_238)
);

MAJx2_ASAP7_75t_L g241 ( 
.A(n_172),
.B(n_28),
.C(n_30),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_193),
.A2(n_129),
.B1(n_142),
.B2(n_158),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_177),
.B(n_129),
.C(n_142),
.Y(n_244)
);

NOR2x1_ASAP7_75t_L g250 ( 
.A(n_163),
.B(n_152),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_162),
.B(n_36),
.C(n_143),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_208),
.C(n_201),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_207),
.A2(n_36),
.B1(n_35),
.B2(n_28),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_197),
.A2(n_36),
.B1(n_30),
.B2(n_34),
.Y(n_257)
);

INVx13_ASAP7_75t_L g262 ( 
.A(n_232),
.Y(n_262)
);

INVx3_ASAP7_75t_SL g339 ( 
.A(n_262),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_263),
.A2(n_272),
.B1(n_290),
.B2(n_292),
.Y(n_308)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_219),
.Y(n_264)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_264),
.Y(n_310)
);

CKINVDCx14_ASAP7_75t_R g323 ( 
.A(n_265),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_220),
.A2(n_181),
.B1(n_167),
.B2(n_189),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_266),
.Y(n_316)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_219),
.Y(n_268)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_268),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_225),
.Y(n_269)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_269),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_228),
.B(n_215),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g333 ( 
.A(n_270),
.Y(n_333)
);

OAI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_220),
.A2(n_216),
.B1(n_249),
.B2(n_250),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_225),
.Y(n_273)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_273),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_274),
.B(n_49),
.Y(n_335)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_246),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_275),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_217),
.A2(n_190),
.B1(n_204),
.B2(n_170),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_276),
.A2(n_301),
.B1(n_223),
.B2(n_221),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_227),
.B(n_195),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_277),
.B(n_281),
.Y(n_311)
);

INVx6_ASAP7_75t_L g278 ( 
.A(n_261),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_278),
.B(n_283),
.Y(n_313)
);

NOR2xp67_ASAP7_75t_L g325 ( 
.A(n_279),
.B(n_17),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_260),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_246),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_282),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_233),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_235),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_284),
.B(n_294),
.Y(n_312)
);

INVxp33_ASAP7_75t_L g286 ( 
.A(n_240),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_286),
.B(n_288),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_235),
.B(n_165),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_287),
.B(n_291),
.Y(n_307)
);

OAI32xp33_ASAP7_75t_L g288 ( 
.A1(n_226),
.A2(n_213),
.A3(n_169),
.B1(n_78),
.B2(n_50),
.Y(n_288)
);

INVx6_ASAP7_75t_L g289 ( 
.A(n_261),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_289),
.B(n_295),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_244),
.A2(n_186),
.B1(n_214),
.B2(n_198),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_249),
.B(n_192),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_226),
.A2(n_164),
.B1(n_98),
.B2(n_209),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_247),
.A2(n_50),
.B1(n_25),
.B2(n_18),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_293),
.A2(n_237),
.B1(n_252),
.B2(n_254),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_227),
.B(n_202),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_224),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_242),
.B(n_161),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_296),
.B(n_297),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_222),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_254),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_303),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_256),
.B(n_161),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_299),
.B(n_300),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_239),
.B(n_50),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_217),
.A2(n_49),
.B1(n_50),
.B2(n_25),
.Y(n_301)
);

MAJx2_ASAP7_75t_L g302 ( 
.A(n_230),
.B(n_17),
.C(n_16),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_302),
.B(n_303),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_249),
.B(n_3),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_271),
.B(n_251),
.C(n_241),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_305),
.B(n_335),
.C(n_336),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_285),
.A2(n_238),
.B1(n_243),
.B2(n_231),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_306),
.A2(n_309),
.B1(n_327),
.B2(n_337),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_285),
.A2(n_234),
.B1(n_237),
.B2(n_223),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_318),
.A2(n_325),
.B(n_273),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_320),
.A2(n_322),
.B1(n_328),
.B2(n_329),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_291),
.B(n_252),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_321),
.B(n_268),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_263),
.A2(n_236),
.B1(n_233),
.B2(n_224),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_284),
.A2(n_258),
.B1(n_248),
.B2(n_245),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_292),
.A2(n_258),
.B1(n_248),
.B2(n_245),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_290),
.A2(n_253),
.B1(n_232),
.B2(n_259),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_287),
.B(n_259),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_330),
.B(n_264),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_265),
.A2(n_25),
.B(n_18),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_334),
.A2(n_280),
.B(n_279),
.Y(n_356)
);

MAJx2_ASAP7_75t_L g336 ( 
.A(n_271),
.B(n_49),
.C(n_18),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_267),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_337)
);

OAI32xp33_ASAP7_75t_L g340 ( 
.A1(n_280),
.A2(n_5),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_340)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_340),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_341),
.B(n_283),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_304),
.B(n_297),
.Y(n_343)
);

CKINVDCx14_ASAP7_75t_R g392 ( 
.A(n_343),
.Y(n_392)
);

INVx8_ASAP7_75t_L g344 ( 
.A(n_339),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g389 ( 
.A(n_344),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_345),
.B(n_350),
.Y(n_377)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_326),
.Y(n_346)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_346),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_347),
.B(n_351),
.Y(n_388)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_317),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_348),
.B(n_349),
.Y(n_395)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_310),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_334),
.B(n_280),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_312),
.B(n_274),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_304),
.B(n_295),
.Y(n_352)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_352),
.Y(n_378)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_310),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_353),
.B(n_355),
.Y(n_375)
);

CKINVDCx14_ASAP7_75t_R g355 ( 
.A(n_311),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_356),
.B(n_360),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_305),
.B(n_302),
.C(n_275),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_357),
.B(n_367),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_323),
.A2(n_280),
.B(n_288),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_359),
.A2(n_322),
.B(n_308),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_321),
.B(n_293),
.Y(n_360)
);

FAx1_ASAP7_75t_SL g362 ( 
.A(n_307),
.B(n_341),
.CI(n_314),
.CON(n_362),
.SN(n_362)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_362),
.B(n_364),
.Y(n_384)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_319),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_363),
.B(n_365),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_339),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_330),
.B(n_282),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_366),
.B(n_368),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_335),
.B(n_289),
.C(n_278),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_333),
.B(n_314),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_331),
.A2(n_283),
.B1(n_273),
.B2(n_269),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_369),
.A2(n_372),
.B1(n_309),
.B2(n_364),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_370),
.B(n_367),
.Y(n_396)
);

INVx4_ASAP7_75t_L g371 ( 
.A(n_339),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_371),
.B(n_374),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_308),
.A2(n_269),
.B1(n_262),
.B2(n_8),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_307),
.B(n_5),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_373),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_327),
.B(n_7),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_379),
.A2(n_381),
.B1(n_358),
.B2(n_369),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_360),
.A2(n_372),
.B1(n_361),
.B2(n_354),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_382),
.A2(n_359),
.B(n_365),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_350),
.A2(n_316),
.B(n_321),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g411 ( 
.A1(n_383),
.A2(n_393),
.B(n_400),
.Y(n_411)
);

NOR3xp33_ASAP7_75t_L g385 ( 
.A(n_361),
.B(n_340),
.C(n_316),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_385),
.B(n_404),
.Y(n_407)
);

BUFx24_ASAP7_75t_SL g390 ( 
.A(n_351),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_390),
.B(n_324),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_345),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_391),
.B(n_344),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_350),
.A2(n_306),
.B(n_328),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_396),
.B(n_398),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_342),
.B(n_357),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_356),
.A2(n_329),
.B(n_319),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_SL g401 ( 
.A(n_342),
.B(n_336),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_401),
.B(n_403),
.Y(n_412)
);

OR2x2_ASAP7_75t_L g402 ( 
.A(n_360),
.B(n_345),
.Y(n_402)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_402),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_362),
.B(n_320),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_347),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_405),
.A2(n_427),
.B1(n_408),
.B2(n_400),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_406),
.B(n_428),
.Y(n_448)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_379),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_408),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_402),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_409),
.B(n_410),
.Y(n_431)
);

CKINVDCx16_ASAP7_75t_R g410 ( 
.A(n_395),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_392),
.B(n_373),
.Y(n_414)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_414),
.Y(n_432)
);

OAI22xp33_ASAP7_75t_SL g415 ( 
.A1(n_378),
.A2(n_366),
.B1(n_363),
.B2(n_337),
.Y(n_415)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_415),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_393),
.A2(n_354),
.B1(n_358),
.B2(n_346),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_416),
.B(n_421),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_380),
.B(n_362),
.C(n_315),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_417),
.B(n_424),
.C(n_401),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_380),
.B(n_338),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_418),
.B(n_396),
.Y(n_430)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_394),
.Y(n_419)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_419),
.Y(n_440)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_394),
.Y(n_422)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_422),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_377),
.B(n_371),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_423),
.B(n_429),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_398),
.B(n_313),
.C(n_332),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_375),
.Y(n_425)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_425),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_426),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_381),
.A2(n_332),
.B1(n_326),
.B2(n_9),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_388),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_388),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_430),
.B(n_436),
.Y(n_461)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_433),
.Y(n_450)
);

FAx1_ASAP7_75t_SL g434 ( 
.A(n_412),
.B(n_403),
.CI(n_377),
.CON(n_434),
.SN(n_434)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_434),
.B(n_411),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_405),
.A2(n_399),
.B1(n_409),
.B2(n_413),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_420),
.B(n_384),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_437),
.B(n_439),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_420),
.B(n_391),
.C(n_399),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_444),
.B(n_447),
.C(n_417),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_SL g445 ( 
.A(n_412),
.B(n_377),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_445),
.B(n_447),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_424),
.B(n_399),
.C(n_383),
.Y(n_447)
);

XNOR2x1_ASAP7_75t_L g472 ( 
.A(n_451),
.B(n_455),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_452),
.B(n_456),
.Y(n_467)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_431),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_453),
.B(n_457),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_439),
.B(n_418),
.C(n_411),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_454),
.B(n_464),
.C(n_434),
.Y(n_470)
);

XNOR2x1_ASAP7_75t_L g456 ( 
.A(n_444),
.B(n_445),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_438),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_438),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_458),
.B(n_460),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_446),
.B(n_448),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_459),
.B(n_462),
.Y(n_480)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_438),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_437),
.B(n_430),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_436),
.B(n_423),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_432),
.Y(n_465)
);

INVx11_ASAP7_75t_L g475 ( 
.A(n_465),
.Y(n_475)
);

INVxp33_ASAP7_75t_L g468 ( 
.A(n_464),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_468),
.B(n_376),
.Y(n_486)
);

INVx6_ASAP7_75t_L g469 ( 
.A(n_450),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_469),
.B(n_397),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_470),
.B(n_427),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_454),
.B(n_433),
.C(n_435),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_471),
.B(n_473),
.C(n_474),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_463),
.B(n_434),
.C(n_449),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_463),
.B(n_416),
.C(n_426),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_SL g476 ( 
.A1(n_451),
.A2(n_407),
.B(n_386),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_476),
.A2(n_7),
.B(n_9),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_SL g477 ( 
.A1(n_461),
.A2(n_406),
.B(n_441),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_477),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_461),
.B(n_423),
.C(n_443),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_478),
.B(n_456),
.C(n_382),
.Y(n_487)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_481),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_467),
.B(n_478),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_482),
.B(n_486),
.Y(n_498)
);

AOI22xp33_ASAP7_75t_SL g483 ( 
.A1(n_469),
.A2(n_442),
.B1(n_440),
.B2(n_389),
.Y(n_483)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_483),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_480),
.B(n_376),
.Y(n_485)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_485),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_487),
.B(n_490),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_488),
.B(n_489),
.Y(n_494)
);

MAJx2_ASAP7_75t_L g489 ( 
.A(n_473),
.B(n_387),
.C(n_389),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_466),
.A2(n_387),
.B1(n_8),
.B2(n_9),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_492),
.A2(n_477),
.B(n_475),
.Y(n_493)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_493),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_491),
.B(n_475),
.Y(n_497)
);

AO21x1_ASAP7_75t_L g502 ( 
.A1(n_497),
.A2(n_483),
.B(n_468),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_498),
.B(n_479),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_501),
.B(n_502),
.Y(n_506)
);

AOI322xp5_ASAP7_75t_L g503 ( 
.A1(n_496),
.A2(n_489),
.A3(n_488),
.B1(n_471),
.B2(n_474),
.C1(n_472),
.C2(n_487),
.Y(n_503)
);

NAND2x1_ASAP7_75t_SL g507 ( 
.A(n_503),
.B(n_484),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_500),
.B(n_484),
.C(n_472),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_505),
.B(n_494),
.Y(n_508)
);

AOI322xp5_ASAP7_75t_L g509 ( 
.A1(n_507),
.A2(n_508),
.A3(n_504),
.B1(n_503),
.B2(n_497),
.C1(n_499),
.C2(n_495),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_509),
.B(n_510),
.Y(n_511)
);

AOI322xp5_ASAP7_75t_L g510 ( 
.A1(n_506),
.A2(n_7),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C1(n_470),
.C2(n_508),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_511),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_512),
.B(n_10),
.C(n_11),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_513),
.B(n_10),
.Y(n_514)
);

BUFx24_ASAP7_75t_SL g515 ( 
.A(n_514),
.Y(n_515)
);


endmodule