module fake_jpeg_31139_n_188 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_188);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_188;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_31),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_22),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_9),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_47),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_2),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_13),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_9),
.Y(n_72)
);

BUFx10_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

BUFx4f_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_61),
.B(n_0),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_84),
.Y(n_90)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

INVx6_ASAP7_75t_SL g84 ( 
.A(n_75),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_76),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_50),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_68),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_96),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_85),
.Y(n_92)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_79),
.A2(n_58),
.B1(n_72),
.B2(n_60),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_95),
.A2(n_98),
.B1(n_65),
.B2(n_82),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_80),
.B(n_67),
.Y(n_96)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_81),
.A2(n_72),
.B1(n_60),
.B2(n_65),
.Y(n_98)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_102),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_104),
.B(n_107),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_98),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_105),
.B(n_113),
.Y(n_123)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_90),
.B(n_59),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_67),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_111),
.Y(n_125)
);

OR2x2_ASAP7_75t_SL g109 ( 
.A(n_97),
.B(n_52),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_116),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

INVxp33_ASAP7_75t_L g142 ( 
.A(n_110),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_59),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_101),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_54),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_119),
.Y(n_138)
);

A2O1A1Ixp33_ASAP7_75t_L g116 ( 
.A1(n_87),
.A2(n_62),
.B(n_56),
.C(n_73),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_116),
.B(n_1),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_117),
.A2(n_118),
.B1(n_28),
.B2(n_45),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_88),
.A2(n_83),
.B1(n_71),
.B2(n_70),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_73),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_112),
.A2(n_63),
.B1(n_64),
.B2(n_66),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_124),
.A2(n_127),
.B1(n_134),
.B2(n_139),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_102),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_126),
.A2(n_135),
.B1(n_140),
.B2(n_21),
.Y(n_158)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_121),
.Y(n_130)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_12),
.Y(n_150)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_141),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_110),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_133),
.B(n_137),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_103),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_134)
);

NOR2x1_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_4),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_114),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_105),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_106),
.Y(n_141)
);

AO21x2_ASAP7_75t_L g145 ( 
.A1(n_137),
.A2(n_32),
.B(n_44),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_145),
.A2(n_157),
.B(n_162),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_138),
.A2(n_8),
.B(n_11),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_146),
.A2(n_126),
.B(n_140),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_125),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_150),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_33),
.C(n_16),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_163),
.C(n_36),
.Y(n_172)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_128),
.Y(n_152)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_152),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_122),
.B(n_12),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_155),
.B(n_158),
.Y(n_170)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_136),
.Y(n_156)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_156),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_123),
.A2(n_18),
.B(n_19),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_143),
.Y(n_160)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_160),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_142),
.B(n_25),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_161),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_26),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_144),
.B(n_29),
.C(n_34),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_171),
.Y(n_174)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_161),
.Y(n_171)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_172),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_165),
.A2(n_153),
.B(n_148),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_175),
.B(n_176),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_170),
.A2(n_147),
.B1(n_145),
.B2(n_154),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g178 ( 
.A(n_173),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_173),
.C(n_162),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_179),
.B(n_174),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_181),
.A2(n_180),
.B(n_177),
.Y(n_182)
);

AOI322xp5_ASAP7_75t_L g183 ( 
.A1(n_182),
.A2(n_169),
.A3(n_178),
.B1(n_168),
.B2(n_145),
.C1(n_171),
.C2(n_147),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_183),
.B(n_164),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_184),
.A2(n_145),
.B1(n_159),
.B2(n_167),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_185),
.B(n_172),
.C(n_39),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_37),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_41),
.Y(n_188)
);


endmodule