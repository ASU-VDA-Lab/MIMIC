module fake_jpeg_2538_n_182 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_182);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_182;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_25),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_16),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

BUFx12_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_14),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_1),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_1),
.B(n_9),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

AND2x2_ASAP7_75t_SL g63 ( 
.A(n_45),
.B(n_22),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_65),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_0),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_0),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_50),
.Y(n_74)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_67),
.Y(n_77)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_68),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_47),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_SL g95 ( 
.A(n_69),
.B(n_61),
.Y(n_95)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_75),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_46),
.Y(n_75)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_62),
.A2(n_54),
.B1(n_59),
.B2(n_52),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_80),
.A2(n_64),
.B1(n_59),
.B2(n_58),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_78),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_86),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_69),
.B(n_65),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_72),
.Y(n_108)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_70),
.B(n_63),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_2),
.Y(n_115)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_47),
.Y(n_86)
);

NOR3xp33_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_63),
.C(n_55),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_91),
.Y(n_103)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_73),
.A2(n_52),
.B(n_48),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_95),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_71),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_55),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_57),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_93),
.A2(n_72),
.B1(n_79),
.B2(n_71),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_76),
.B(n_48),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_53),
.Y(n_106)
);

INVxp33_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_94),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_106),
.Y(n_130)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_90),
.Y(n_105)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_84),
.A2(n_67),
.B1(n_56),
.B2(n_58),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_107),
.A2(n_113),
.B1(n_96),
.B2(n_82),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_116),
.Y(n_119)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_109),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_114),
.Y(n_131)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

OAI21xp33_ASAP7_75t_SL g112 ( 
.A1(n_89),
.A2(n_50),
.B(n_67),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_115),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_84),
.A2(n_60),
.B1(n_51),
.B2(n_4),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_26),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_117),
.B(n_128),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_88),
.C(n_85),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_123),
.C(n_98),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_100),
.A2(n_60),
.B1(n_51),
.B2(n_24),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_121),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_115),
.B(n_60),
.C(n_51),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_108),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_126),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_3),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_116),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_135),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_113),
.A2(n_27),
.B1(n_42),
.B2(n_41),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_132),
.A2(n_133),
.B(n_31),
.Y(n_144)
);

A2O1A1O1Ixp25_ASAP7_75t_L g133 ( 
.A1(n_115),
.A2(n_44),
.B(n_40),
.C(n_38),
.D(n_36),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_103),
.A2(n_5),
.B(n_7),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_134),
.A2(n_7),
.B(n_8),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_5),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_127),
.Y(n_137)
);

NAND3xp33_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_140),
.C(n_143),
.Y(n_161)
);

AOI21x1_ASAP7_75t_L g138 ( 
.A1(n_120),
.A2(n_114),
.B(n_102),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_138),
.A2(n_150),
.B(n_152),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_118),
.B(n_107),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_28),
.C(n_29),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_144),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_122),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_145),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_124),
.A2(n_109),
.B1(n_9),
.B2(n_10),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_146),
.A2(n_17),
.B1(n_19),
.B2(n_147),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_124),
.A2(n_35),
.B(n_34),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_147),
.A2(n_148),
.B(n_123),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_120),
.A2(n_8),
.B(n_10),
.Y(n_148)
);

OAI321xp33_ASAP7_75t_L g154 ( 
.A1(n_149),
.A2(n_126),
.A3(n_132),
.B1(n_133),
.B2(n_20),
.C(n_18),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_151),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_15),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_142),
.A2(n_117),
.B1(n_130),
.B2(n_121),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_153),
.A2(n_154),
.B1(n_149),
.B2(n_150),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_156),
.A2(n_159),
.B(n_148),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_158),
.B(n_156),
.C(n_145),
.Y(n_166)
);

A2O1A1O1Ixp25_ASAP7_75t_L g159 ( 
.A1(n_136),
.A2(n_30),
.B(n_32),
.C(n_20),
.D(n_17),
.Y(n_159)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_160),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_161),
.Y(n_164)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_164),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_157),
.B(n_139),
.Y(n_165)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_165),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_166),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_168),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_163),
.A2(n_151),
.B(n_141),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_153),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_175),
.B(n_176),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_159),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_172),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_155),
.Y(n_179)
);

AOI322xp5_ASAP7_75t_L g180 ( 
.A1(n_179),
.A2(n_162),
.A3(n_174),
.B1(n_169),
.B2(n_170),
.C1(n_158),
.C2(n_140),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_174),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_181),
.A2(n_170),
.B(n_19),
.Y(n_182)
);


endmodule