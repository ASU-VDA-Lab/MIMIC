module fake_jpeg_28788_n_467 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_467);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_467;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_393;
wire n_288;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_14),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_6),
.B(n_15),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_49),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_7),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_50),
.B(n_75),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_51),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx5_ASAP7_75t_SL g142 ( 
.A(n_52),
.Y(n_142)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_56),
.Y(n_134)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_57),
.Y(n_120)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_58),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_59),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_60),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_61),
.Y(n_140)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_63),
.Y(n_132)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_64),
.Y(n_143)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_65),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_66),
.Y(n_127)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_39),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_67),
.B(n_80),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_16),
.Y(n_71)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_73),
.Y(n_108)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_16),
.Y(n_74)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_7),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_78),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_79),
.Y(n_148)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_39),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_81),
.Y(n_129)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_82),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

INVx6_ASAP7_75t_SL g133 ( 
.A(n_83),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_18),
.B(n_7),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_84),
.B(n_85),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_8),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_86),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_87),
.B(n_88),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx11_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_93),
.Y(n_114)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

NAND2xp33_ASAP7_75t_SL g111 ( 
.A(n_90),
.B(n_91),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_92),
.Y(n_115)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_38),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_18),
.B(n_8),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_94),
.B(n_95),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_20),
.B(n_8),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_28),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_96),
.A2(n_21),
.B1(n_28),
.B2(n_30),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_105),
.A2(n_151),
.B1(n_40),
.B2(n_29),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_51),
.A2(n_44),
.B1(n_20),
.B2(n_24),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_116),
.A2(n_122),
.B1(n_128),
.B2(n_131),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_84),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_35),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_91),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_119),
.B(n_124),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_59),
.A2(n_44),
.B1(n_24),
.B2(n_34),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_95),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_67),
.A2(n_21),
.B1(n_47),
.B2(n_41),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_80),
.A2(n_47),
.B1(n_41),
.B2(n_28),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_61),
.A2(n_34),
.B1(n_35),
.B2(n_40),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_135),
.A2(n_136),
.B1(n_138),
.B2(n_141),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_L g136 ( 
.A1(n_68),
.A2(n_23),
.B1(n_33),
.B2(n_29),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_69),
.A2(n_77),
.B1(n_70),
.B2(n_72),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_76),
.A2(n_47),
.B1(n_41),
.B2(n_28),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_78),
.A2(n_47),
.B1(n_41),
.B2(n_30),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_144),
.A2(n_63),
.B1(n_53),
.B2(n_30),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_92),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_150),
.B(n_56),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_79),
.A2(n_43),
.B1(n_19),
.B2(n_23),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_152),
.B(n_153),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_102),
.B(n_49),
.Y(n_153)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_97),
.Y(n_154)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_154),
.Y(n_205)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_106),
.Y(n_155)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_155),
.Y(n_226)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_106),
.Y(n_157)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_157),
.Y(n_232)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_125),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_158),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_125),
.Y(n_159)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_159),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_160),
.A2(n_186),
.B1(n_194),
.B2(n_200),
.Y(n_234)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_123),
.Y(n_161)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_161),
.Y(n_203)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_109),
.Y(n_162)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_162),
.Y(n_210)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_109),
.Y(n_163)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_163),
.Y(n_236)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_98),
.Y(n_164)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_164),
.Y(n_242)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_97),
.Y(n_165)
);

INVx4_ASAP7_75t_SL g224 ( 
.A(n_165),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_110),
.B(n_113),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_166),
.B(n_183),
.Y(n_216)
);

OAI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_136),
.A2(n_83),
.B1(n_55),
.B2(n_73),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_167),
.A2(n_168),
.B1(n_104),
.B2(n_99),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_133),
.A2(n_88),
.B1(n_87),
.B2(n_86),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_130),
.Y(n_169)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_169),
.Y(n_241)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_100),
.Y(n_170)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_170),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_121),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_171),
.B(n_181),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_132),
.Y(n_172)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_172),
.Y(n_238)
);

AND2x2_ASAP7_75t_SL g173 ( 
.A(n_118),
.B(n_96),
.Y(n_173)
);

FAx1_ASAP7_75t_SL g233 ( 
.A(n_173),
.B(n_117),
.CI(n_98),
.CON(n_233),
.SN(n_233)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_100),
.Y(n_174)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_174),
.Y(n_213)
);

OA22x2_ASAP7_75t_L g235 ( 
.A1(n_175),
.A2(n_201),
.B1(n_99),
.B2(n_104),
.Y(n_235)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_101),
.Y(n_176)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_176),
.Y(n_214)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_101),
.Y(n_177)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_177),
.Y(n_218)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_142),
.Y(n_179)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_179),
.Y(n_222)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_146),
.Y(n_180)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_180),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_121),
.Y(n_181)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_142),
.Y(n_182)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_182),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_114),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_139),
.B(n_33),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_184),
.B(n_197),
.Y(n_229)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_146),
.Y(n_185)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_185),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_133),
.A2(n_43),
.B1(n_19),
.B2(n_52),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_139),
.B(n_60),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_189),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_134),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_190),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_145),
.B(n_60),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_129),
.Y(n_190)
);

MAJx2_ASAP7_75t_L g191 ( 
.A(n_111),
.B(n_56),
.C(n_52),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_191),
.B(n_173),
.C(n_178),
.Y(n_225)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_148),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_192),
.Y(n_227)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_148),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_195),
.Y(n_208)
);

INVx4_ASAP7_75t_SL g194 ( 
.A(n_134),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_103),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_115),
.B(n_49),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_120),
.Y(n_202)
);

O2A1O1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_111),
.A2(n_30),
.B(n_8),
.C(n_9),
.Y(n_199)
);

OA22x2_ASAP7_75t_L g240 ( 
.A1(n_199),
.A2(n_127),
.B1(n_112),
.B2(n_130),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_132),
.A2(n_6),
.B1(n_12),
.B2(n_11),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_103),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_202),
.B(n_233),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_108),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_204),
.B(n_225),
.C(n_230),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_211),
.A2(n_217),
.B1(n_220),
.B2(n_196),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_161),
.A2(n_138),
.B1(n_107),
.B2(n_126),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_191),
.A2(n_147),
.B(n_143),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_219),
.A2(n_137),
.B(n_165),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_175),
.A2(n_126),
.B1(n_117),
.B2(n_107),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_152),
.B(n_147),
.C(n_143),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_235),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_184),
.B(n_112),
.C(n_149),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_239),
.B(n_137),
.Y(n_275)
);

OAI21xp33_ASAP7_75t_SL g279 ( 
.A1(n_240),
.A2(n_127),
.B(n_194),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_215),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_243),
.B(n_249),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_225),
.A2(n_203),
.B1(n_235),
.B2(n_234),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_244),
.A2(n_253),
.B1(n_269),
.B2(n_279),
.Y(n_282)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_210),
.Y(n_246)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_246),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_247),
.A2(n_227),
.B1(n_209),
.B2(n_221),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_220),
.A2(n_183),
.B1(n_199),
.B2(n_164),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_248),
.B(n_229),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_206),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_241),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_250),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_235),
.A2(n_190),
.B1(n_162),
.B2(n_170),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_251),
.A2(n_254),
.B1(n_255),
.B2(n_256),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_219),
.A2(n_189),
.B(n_156),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_252),
.A2(n_276),
.B(n_188),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_235),
.A2(n_140),
.B1(n_177),
.B2(n_176),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_217),
.A2(n_174),
.B1(n_155),
.B2(n_157),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_202),
.A2(n_163),
.B1(n_193),
.B2(n_140),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_204),
.A2(n_201),
.B1(n_195),
.B2(n_192),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_206),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_257),
.B(n_259),
.Y(n_302)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_212),
.Y(n_258)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_258),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_206),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_208),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_260),
.B(n_261),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_208),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_233),
.B(n_185),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_266),
.Y(n_283)
);

INVxp33_ASAP7_75t_L g263 ( 
.A(n_224),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_263),
.B(n_264),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_208),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_213),
.Y(n_265)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_265),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_233),
.B(n_180),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_230),
.B(n_182),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_267),
.B(n_277),
.Y(n_308)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_214),
.Y(n_268)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_268),
.Y(n_295)
);

OAI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_240),
.A2(n_158),
.B1(n_172),
.B2(n_169),
.Y(n_269)
);

AO21x2_ASAP7_75t_L g270 ( 
.A1(n_240),
.A2(n_159),
.B(n_179),
.Y(n_270)
);

AO22x1_ASAP7_75t_SL g285 ( 
.A1(n_270),
.A2(n_279),
.B1(n_253),
.B2(n_240),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_238),
.Y(n_273)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_273),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_238),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_274),
.Y(n_284)
);

XNOR2x1_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_231),
.Y(n_296)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_223),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_226),
.Y(n_278)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_278),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_245),
.A2(n_276),
.B(n_266),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_280),
.A2(n_301),
.B(n_245),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_239),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_281),
.B(n_296),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_285),
.B(n_299),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_272),
.A2(n_216),
.B1(n_242),
.B2(n_218),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_287),
.A2(n_251),
.B1(n_247),
.B2(n_255),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_272),
.A2(n_229),
.B1(n_207),
.B2(n_242),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_290),
.A2(n_303),
.B1(n_311),
.B2(n_304),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_291),
.B(n_298),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_246),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_292),
.B(n_307),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_248),
.B(n_262),
.Y(n_298)
);

OA21x2_ASAP7_75t_L g299 ( 
.A1(n_270),
.A2(n_222),
.B(n_237),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_272),
.A2(n_209),
.B1(n_241),
.B2(n_221),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_271),
.B(n_228),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_305),
.B(n_252),
.C(n_256),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_258),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_265),
.Y(n_309)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_309),
.Y(n_317)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_268),
.Y(n_312)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_312),
.Y(n_335)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_274),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_313),
.A2(n_286),
.B1(n_297),
.B2(n_306),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_314),
.A2(n_334),
.B1(n_287),
.B2(n_298),
.Y(n_346)
);

OAI32xp33_ASAP7_75t_L g315 ( 
.A1(n_283),
.A2(n_267),
.A3(n_245),
.B1(n_275),
.B2(n_277),
.Y(n_315)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_315),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_316),
.B(n_341),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_318),
.A2(n_319),
.B1(n_327),
.B2(n_329),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_282),
.A2(n_244),
.B1(n_270),
.B2(n_264),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_310),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_321),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_280),
.A2(n_260),
.B(n_261),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_322),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_323),
.B(n_330),
.C(n_332),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_304),
.A2(n_270),
.B1(n_254),
.B2(n_250),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_325),
.A2(n_326),
.B1(n_336),
.B2(n_295),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_290),
.A2(n_270),
.B1(n_250),
.B2(n_224),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_282),
.A2(n_270),
.B1(n_278),
.B2(n_273),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_300),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_328),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_285),
.A2(n_273),
.B1(n_205),
.B2(n_232),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_305),
.B(n_205),
.C(n_232),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_331),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_281),
.B(n_236),
.C(n_226),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_285),
.A2(n_236),
.B1(n_1),
.B2(n_2),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_333),
.B(n_338),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_SL g334 ( 
.A1(n_286),
.A2(n_9),
.B1(n_12),
.B2(n_3),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_298),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_299),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_337),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_308),
.A2(n_0),
.B1(n_4),
.B2(n_9),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_283),
.A2(n_0),
.B(n_4),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_291),
.A2(n_0),
.B1(n_10),
.B2(n_11),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_342),
.B(n_343),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_291),
.A2(n_14),
.B1(n_10),
.B2(n_12),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_340),
.B(n_308),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_344),
.B(n_351),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_346),
.A2(n_368),
.B1(n_327),
.B2(n_329),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_321),
.B(n_289),
.Y(n_348)
);

CKINVDCx14_ASAP7_75t_R g393 ( 
.A(n_348),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_340),
.B(n_296),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_349),
.B(n_352),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_323),
.B(n_301),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_315),
.B(n_302),
.Y(n_352)
);

INVx4_ASAP7_75t_L g354 ( 
.A(n_328),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_354),
.Y(n_376)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_324),
.Y(n_359)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_359),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_324),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_360),
.B(n_309),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_316),
.B(n_294),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_362),
.B(n_363),
.C(n_367),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_332),
.B(n_284),
.C(n_313),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_337),
.B(n_299),
.Y(n_365)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_365),
.Y(n_382)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_317),
.Y(n_366)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_366),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_330),
.B(n_284),
.C(n_312),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_339),
.B(n_295),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_370),
.B(n_342),
.C(n_336),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_365),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_371),
.B(n_373),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_347),
.B(n_333),
.Y(n_372)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_372),
.Y(n_400)
);

NOR2xp67_ASAP7_75t_L g373 ( 
.A(n_352),
.B(n_339),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_353),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_374),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g375 ( 
.A1(n_361),
.A2(n_339),
.B(n_322),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_375),
.A2(n_361),
.B(n_355),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_378),
.A2(n_364),
.B1(n_369),
.B2(n_350),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_364),
.A2(n_320),
.B1(n_326),
.B2(n_314),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_379),
.A2(n_370),
.B1(n_355),
.B2(n_362),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_357),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_380),
.B(n_388),
.Y(n_397)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_383),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_384),
.B(n_344),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_358),
.B(n_319),
.C(n_318),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_386),
.B(n_391),
.C(n_367),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_354),
.B(n_320),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_368),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_389),
.B(n_338),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_345),
.B(n_317),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_390),
.B(n_341),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_358),
.B(n_335),
.C(n_325),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_394),
.A2(n_375),
.B(n_380),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_395),
.A2(n_401),
.B1(n_409),
.B2(n_379),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_396),
.B(n_403),
.C(n_404),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_392),
.B(n_351),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_398),
.B(n_411),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_378),
.A2(n_369),
.B1(n_345),
.B2(n_356),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_381),
.B(n_363),
.C(n_391),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_406),
.A2(n_408),
.B1(n_384),
.B2(n_372),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_385),
.B(n_349),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_407),
.B(n_385),
.C(n_381),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_389),
.A2(n_355),
.B1(n_303),
.B2(n_343),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_382),
.A2(n_356),
.B1(n_335),
.B2(n_341),
.Y(n_409)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_410),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_SL g427 ( 
.A(n_413),
.B(n_418),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_399),
.A2(n_388),
.B(n_382),
.Y(n_414)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_414),
.A2(n_394),
.B(n_377),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_405),
.B(n_374),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_415),
.B(n_420),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_417),
.A2(n_395),
.B1(n_410),
.B2(n_407),
.Y(n_436)
);

AOI22xp33_ASAP7_75t_SL g419 ( 
.A1(n_400),
.A2(n_377),
.B1(n_393),
.B2(n_387),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_419),
.A2(n_297),
.B1(n_288),
.B2(n_293),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_402),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_396),
.B(n_386),
.C(n_392),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_421),
.B(n_424),
.C(n_404),
.Y(n_431)
);

OR2x2_ASAP7_75t_L g422 ( 
.A(n_397),
.B(n_371),
.Y(n_422)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_422),
.Y(n_439)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_409),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_423),
.B(n_411),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_403),
.B(n_376),
.C(n_390),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_425),
.A2(n_408),
.B1(n_401),
.B2(n_373),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_412),
.Y(n_429)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_429),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_430),
.B(n_434),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_431),
.B(n_433),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_416),
.B(n_398),
.C(n_406),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_432),
.B(n_438),
.C(n_421),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_422),
.A2(n_410),
.B1(n_376),
.B2(n_387),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_435),
.B(n_437),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_436),
.A2(n_288),
.B1(n_293),
.B2(n_294),
.Y(n_448)
);

INVxp33_ASAP7_75t_L g437 ( 
.A(n_413),
.Y(n_437)
);

AOI21x1_ASAP7_75t_L g440 ( 
.A1(n_437),
.A2(n_414),
.B(n_426),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_L g450 ( 
.A1(n_440),
.A2(n_436),
.B(n_433),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_439),
.A2(n_425),
.B1(n_424),
.B2(n_416),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_441),
.B(n_442),
.C(n_445),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_431),
.B(n_418),
.C(n_306),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_448),
.A2(n_10),
.B(n_14),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g449 ( 
.A(n_428),
.B(n_432),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_449),
.B(n_427),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_450),
.A2(n_453),
.B(n_454),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_451),
.B(n_452),
.Y(n_457)
);

INVx6_ASAP7_75t_L g452 ( 
.A(n_443),
.Y(n_452)
);

NOR2x1_ASAP7_75t_L g453 ( 
.A(n_448),
.B(n_427),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_440),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_455),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_SL g459 ( 
.A(n_456),
.B(n_446),
.Y(n_459)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_459),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_457),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_462),
.B(n_447),
.Y(n_463)
);

OAI311xp33_ASAP7_75t_L g464 ( 
.A1(n_463),
.A2(n_460),
.A3(n_461),
.B1(n_458),
.C1(n_454),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_464),
.A2(n_442),
.B(n_444),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_465),
.B(n_445),
.C(n_453),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_466),
.B(n_14),
.Y(n_467)
);


endmodule