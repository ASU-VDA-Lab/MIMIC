module fake_jpeg_29316_n_514 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_514);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_514;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_11),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_11),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_7),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_52),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_53),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_54),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_55),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_58),
.Y(n_141)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_59),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_17),
.B(n_9),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_60),
.B(n_97),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_61),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_62),
.Y(n_150)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

INVx3_ASAP7_75t_SL g64 ( 
.A(n_51),
.Y(n_64)
);

INVx1_ASAP7_75t_SL g108 ( 
.A(n_64),
.Y(n_108)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_65),
.Y(n_125)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_66),
.Y(n_112)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_67),
.Y(n_118)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_68),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_70),
.Y(n_133)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_72),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_73),
.Y(n_139)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_77),
.Y(n_130)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_78),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_17),
.B(n_9),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_79),
.B(n_95),
.Y(n_123)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_80),
.Y(n_142)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_38),
.Y(n_81)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_82),
.Y(n_107)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_83),
.Y(n_103)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_25),
.Y(n_84)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_85),
.Y(n_149)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_86),
.Y(n_152)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_87),
.Y(n_154)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_88),
.Y(n_155)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_90),
.Y(n_124)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_49),
.Y(n_92)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_92),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_93),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_23),
.Y(n_94)
);

BUFx10_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_20),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_96),
.B(n_98),
.Y(n_102)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_39),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_39),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_20),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_23),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_28),
.B(n_10),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_100),
.B(n_30),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_60),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_104),
.B(n_109),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_100),
.B(n_44),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_95),
.A2(n_50),
.B1(n_47),
.B2(n_28),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_113),
.A2(n_120),
.B1(n_126),
.B2(n_140),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_66),
.B(n_50),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_115),
.B(n_24),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_93),
.A2(n_47),
.B1(n_33),
.B2(n_44),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_53),
.A2(n_33),
.B1(n_19),
.B2(n_24),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_70),
.B(n_25),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_127),
.B(n_147),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_138),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_64),
.A2(n_46),
.B1(n_20),
.B2(n_23),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_74),
.A2(n_46),
.B1(n_20),
.B2(n_23),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_144),
.A2(n_157),
.B1(n_32),
.B2(n_75),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_72),
.B(n_19),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_52),
.A2(n_46),
.B1(n_23),
.B2(n_40),
.Y(n_157)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_158),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_137),
.A2(n_32),
.B(n_22),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_159),
.A2(n_195),
.B(n_32),
.Y(n_223)
);

BUFx10_ASAP7_75t_L g160 ( 
.A(n_111),
.Y(n_160)
);

INVx11_ASAP7_75t_L g234 ( 
.A(n_160),
.Y(n_234)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_110),
.Y(n_161)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_161),
.Y(n_212)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_163),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_137),
.A2(n_40),
.B1(n_42),
.B2(n_34),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_164),
.B(n_165),
.Y(n_249)
);

OA22x2_ASAP7_75t_L g165 ( 
.A1(n_115),
.A2(n_80),
.B1(n_91),
.B2(n_88),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_101),
.Y(n_166)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_166),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_141),
.Y(n_167)
);

NAND2xp33_ASAP7_75t_SL g242 ( 
.A(n_167),
.B(n_203),
.Y(n_242)
);

AO22x2_ASAP7_75t_L g168 ( 
.A1(n_144),
.A2(n_92),
.B1(n_85),
.B2(n_77),
.Y(n_168)
);

NOR2x1_ASAP7_75t_L g213 ( 
.A(n_168),
.B(n_140),
.Y(n_213)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_142),
.Y(n_169)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_169),
.Y(n_250)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_124),
.Y(n_171)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_171),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_172),
.A2(n_187),
.B1(n_188),
.B2(n_197),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_119),
.Y(n_173)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_173),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_157),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_174),
.Y(n_246)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_154),
.Y(n_175)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_175),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_122),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_176),
.B(n_183),
.Y(n_248)
);

INVx11_ASAP7_75t_L g178 ( 
.A(n_131),
.Y(n_178)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_178),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_152),
.Y(n_179)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_179),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_143),
.Y(n_180)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_180),
.Y(n_252)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_131),
.Y(n_181)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_181),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

BUFx4f_ASAP7_75t_L g245 ( 
.A(n_182),
.Y(n_245)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_106),
.Y(n_183)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_184),
.B(n_185),
.Y(n_254)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_118),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_150),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_186),
.B(n_190),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_151),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_153),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_129),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_189),
.B(n_191),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_138),
.B(n_123),
.Y(n_190)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_132),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_146),
.A2(n_76),
.B1(n_73),
.B2(n_69),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_192),
.A2(n_105),
.B1(n_117),
.B2(n_130),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_102),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_193),
.B(n_194),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_103),
.A2(n_45),
.B1(n_30),
.B2(n_34),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_134),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_196),
.Y(n_247)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_148),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_112),
.B(n_125),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_198),
.B(n_207),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_108),
.B(n_107),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_199),
.B(n_32),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_153),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_200),
.A2(n_201),
.B1(n_202),
.B2(n_204),
.Y(n_221)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_136),
.Y(n_201)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_156),
.Y(n_202)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_143),
.Y(n_203)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_114),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_114),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_205),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_150),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_145),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_208),
.A2(n_209),
.B1(n_103),
.B2(n_107),
.Y(n_222)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_133),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_206),
.A2(n_146),
.B1(n_135),
.B2(n_156),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_210),
.A2(n_225),
.B1(n_227),
.B2(n_239),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_213),
.A2(n_214),
.B1(n_243),
.B2(n_181),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_159),
.A2(n_108),
.B(n_22),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_216),
.A2(n_195),
.B(n_184),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_177),
.B(n_162),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_217),
.B(n_224),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_222),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_223),
.A2(n_178),
.B(n_191),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_162),
.B(n_149),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_174),
.A2(n_105),
.B1(n_117),
.B2(n_130),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_168),
.A2(n_55),
.B1(n_62),
.B2(n_61),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_164),
.B(n_54),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_228),
.B(n_231),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_165),
.B(n_45),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_165),
.B(n_42),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_232),
.B(n_236),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_235),
.B(n_241),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_170),
.B(n_139),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_168),
.A2(n_139),
.B1(n_116),
.B2(n_141),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_199),
.B(n_111),
.C(n_112),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_240),
.B(n_183),
.C(n_204),
.Y(n_272)
);

AND2x2_ASAP7_75t_SL g241 ( 
.A(n_161),
.B(n_0),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_172),
.A2(n_111),
.B1(n_46),
.B2(n_2),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_251),
.A2(n_167),
.B1(n_180),
.B2(n_203),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_256),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_257),
.A2(n_243),
.B(n_221),
.Y(n_300)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_238),
.Y(n_258)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_258),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_259),
.A2(n_260),
.B1(n_274),
.B2(n_275),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_249),
.A2(n_168),
.B1(n_192),
.B2(n_202),
.Y(n_260)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_252),
.Y(n_261)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_261),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_263),
.B(n_293),
.Y(n_312)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_238),
.Y(n_264)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_264),
.Y(n_308)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_229),
.Y(n_269)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_269),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_231),
.A2(n_158),
.B1(n_169),
.B2(n_200),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_270),
.A2(n_278),
.B1(n_281),
.B2(n_291),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_211),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_271),
.B(n_273),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_272),
.B(n_280),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g273 ( 
.A(n_211),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g274 ( 
.A1(n_246),
.A2(n_205),
.B1(n_188),
.B2(n_187),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_249),
.A2(n_182),
.B1(n_173),
.B2(n_11),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_249),
.A2(n_160),
.B(n_10),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_276),
.A2(n_283),
.B(n_225),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_226),
.B(n_6),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_277),
.B(n_287),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_232),
.A2(n_160),
.B1(n_1),
.B2(n_2),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_224),
.B(n_6),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_279),
.B(n_284),
.C(n_296),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_217),
.B(n_12),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_213),
.A2(n_5),
.B1(n_15),
.B2(n_3),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_223),
.A2(n_213),
.B(n_216),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_282),
.A2(n_295),
.B(n_234),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_239),
.A2(n_5),
.B(n_14),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_218),
.B(n_3),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_236),
.B(n_3),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_285),
.B(n_289),
.Y(n_301)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_220),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_286),
.Y(n_316)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_229),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_212),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_288),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_248),
.B(n_4),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_254),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_290),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_227),
.A2(n_210),
.B1(n_228),
.B2(n_215),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_230),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_230),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_297),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_240),
.A2(n_4),
.B(n_13),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_235),
.B(n_0),
.C(n_1),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_233),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_266),
.B(n_265),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_299),
.B(n_303),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_300),
.A2(n_314),
.B(n_245),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_266),
.B(n_241),
.C(n_253),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_265),
.B(n_233),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_305),
.B(n_332),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_292),
.B(n_267),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_311),
.B(n_319),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_291),
.A2(n_214),
.B1(n_241),
.B2(n_247),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_315),
.A2(n_318),
.B1(n_321),
.B2(n_326),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_262),
.A2(n_247),
.B1(n_253),
.B2(n_242),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_292),
.B(n_255),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_262),
.A2(n_242),
.B1(n_220),
.B2(n_244),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_290),
.B(n_237),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_323),
.B(n_325),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_280),
.B(n_237),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_270),
.A2(n_220),
.B1(n_244),
.B2(n_212),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_288),
.Y(n_327)
);

OR2x2_ASAP7_75t_L g357 ( 
.A(n_327),
.B(n_333),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_267),
.B(n_278),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_328),
.B(n_329),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_279),
.B(n_250),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_257),
.A2(n_245),
.B1(n_250),
.B2(n_219),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_330),
.A2(n_275),
.B1(n_260),
.B2(n_268),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_331),
.A2(n_276),
.B(n_263),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_282),
.B(n_245),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_269),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_287),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_334),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_304),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_338),
.Y(n_389)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_304),
.Y(n_339)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_339),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_317),
.A2(n_283),
.B1(n_268),
.B2(n_259),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_340),
.A2(n_351),
.B1(n_367),
.B2(n_321),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_341),
.B(n_331),
.Y(n_378)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_306),
.Y(n_342)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_342),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_344),
.A2(n_349),
.B1(n_320),
.B2(n_305),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_323),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_345),
.B(n_364),
.Y(n_399)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_306),
.Y(n_347)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_347),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_302),
.A2(n_281),
.B1(n_272),
.B2(n_295),
.Y(n_349)
);

NOR2xp67_ASAP7_75t_L g350 ( 
.A(n_322),
.B(n_284),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_350),
.B(n_369),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_317),
.A2(n_297),
.B1(n_294),
.B2(n_293),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_299),
.B(n_296),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_353),
.B(n_298),
.C(n_320),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_311),
.B(n_264),
.Y(n_354)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_354),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_319),
.B(n_258),
.Y(n_355)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_355),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_SL g376 ( 
.A(n_356),
.B(n_360),
.Y(n_376)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_308),
.Y(n_358)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_358),
.Y(n_390)
);

OAI32xp33_ASAP7_75t_L g359 ( 
.A1(n_328),
.A2(n_313),
.A3(n_315),
.B1(n_322),
.B2(n_318),
.Y(n_359)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_359),
.Y(n_394)
);

XNOR2x1_ASAP7_75t_L g360 ( 
.A(n_303),
.B(n_261),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_307),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_361),
.B(n_363),
.Y(n_370)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_308),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_313),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g365 ( 
.A1(n_312),
.A2(n_286),
.B(n_252),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_365),
.B(n_332),
.Y(n_375)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_324),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_366),
.B(n_309),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_310),
.A2(n_219),
.B1(n_234),
.B2(n_13),
.Y(n_367)
);

OA21x2_ASAP7_75t_L g368 ( 
.A1(n_314),
.A2(n_4),
.B(n_13),
.Y(n_368)
);

AO22x1_ASAP7_75t_SL g374 ( 
.A1(n_368),
.A2(n_300),
.B1(n_324),
.B2(n_330),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_335),
.B(n_14),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_372),
.A2(n_344),
.B1(n_349),
.B2(n_364),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_373),
.B(n_379),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_374),
.B(n_338),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_375),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_377),
.A2(n_382),
.B1(n_392),
.B2(n_351),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_SL g419 ( 
.A(n_378),
.B(n_398),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_348),
.B(n_337),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_343),
.A2(n_312),
.B1(n_302),
.B2(n_333),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_348),
.B(n_298),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_385),
.B(n_387),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_340),
.A2(n_335),
.B1(n_301),
.B2(n_334),
.Y(n_386)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_386),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_337),
.B(n_329),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_345),
.A2(n_301),
.B1(n_326),
.B2(n_312),
.Y(n_388)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_388),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_353),
.B(n_325),
.C(n_307),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_391),
.B(n_397),
.C(n_354),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_343),
.A2(n_309),
.B1(n_327),
.B2(n_316),
.Y(n_392)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_393),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_360),
.B(n_16),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_395),
.B(n_346),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_352),
.B(n_0),
.C(n_16),
.Y(n_397)
);

XNOR2x2_ASAP7_75t_SL g398 ( 
.A(n_355),
.B(n_0),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_400),
.B(n_382),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_405),
.B(n_411),
.C(n_418),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_394),
.Y(n_407)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_407),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_399),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_408),
.B(n_422),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_396),
.B(n_362),
.Y(n_409)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_409),
.Y(n_429)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_393),
.Y(n_410)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_410),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_385),
.B(n_352),
.C(n_339),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_412),
.B(n_415),
.Y(n_426)
);

AOI22xp33_ASAP7_75t_SL g413 ( 
.A1(n_389),
.A2(n_356),
.B1(n_336),
.B2(n_371),
.Y(n_413)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_413),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_414),
.A2(n_383),
.B1(n_380),
.B2(n_374),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_380),
.A2(n_359),
.B1(n_362),
.B2(n_336),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_SL g436 ( 
.A(n_416),
.B(n_418),
.Y(n_436)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_370),
.Y(n_417)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_417),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_387),
.B(n_346),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_379),
.B(n_341),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_420),
.B(n_378),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_377),
.B(n_365),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_421),
.B(n_376),
.C(n_395),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_391),
.B(n_357),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_381),
.Y(n_423)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_423),
.Y(n_443)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_370),
.Y(n_424)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_424),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_430),
.B(n_432),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_431),
.B(n_433),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_402),
.B(n_373),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_402),
.B(n_376),
.C(n_375),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_434),
.B(n_441),
.C(n_442),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_436),
.B(n_425),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_438),
.A2(n_400),
.B1(n_392),
.B2(n_403),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_406),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_439),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_404),
.B(n_383),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_404),
.B(n_374),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_412),
.B(n_357),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_444),
.B(n_415),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_447),
.B(n_452),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_448),
.B(n_458),
.Y(n_466)
);

INVxp67_ASAP7_75t_SL g449 ( 
.A(n_444),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_449),
.B(n_439),
.Y(n_467)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_450),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_438),
.A2(n_401),
.B1(n_437),
.B2(n_426),
.Y(n_451)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_451),
.Y(n_471)
);

XOR2x2_ASAP7_75t_L g452 ( 
.A(n_442),
.B(n_420),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_431),
.A2(n_421),
.B1(n_425),
.B2(n_416),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_457),
.B(n_433),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_446),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_428),
.B(n_411),
.C(n_405),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_459),
.B(n_462),
.C(n_463),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_427),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_460),
.B(n_461),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_429),
.B(n_423),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_428),
.B(n_419),
.C(n_361),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_432),
.B(n_419),
.C(n_390),
.Y(n_463)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_467),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_459),
.B(n_441),
.C(n_430),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_468),
.B(n_476),
.C(n_453),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_455),
.A2(n_431),
.B(n_435),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_469),
.A2(n_472),
.B(n_358),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_470),
.B(n_457),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_455),
.A2(n_426),
.B(n_440),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_451),
.B(n_445),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_474),
.B(n_477),
.Y(n_487)
);

OR2x2_ASAP7_75t_L g475 ( 
.A(n_456),
.B(n_443),
.Y(n_475)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_475),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_453),
.B(n_434),
.C(n_436),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_456),
.B(n_397),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_475),
.B(n_462),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_479),
.B(n_482),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_464),
.A2(n_398),
.B1(n_452),
.B2(n_384),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_480),
.A2(n_486),
.B1(n_367),
.B2(n_368),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_481),
.B(n_485),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_466),
.B(n_463),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_465),
.B(n_454),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_483),
.B(n_491),
.Y(n_500)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_471),
.A2(n_363),
.B1(n_342),
.B2(n_347),
.Y(n_486)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_488),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_478),
.B(n_469),
.Y(n_489)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_489),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_465),
.B(n_454),
.C(n_366),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_488),
.A2(n_470),
.B(n_472),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_493),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_484),
.A2(n_491),
.B(n_481),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_494),
.B(n_495),
.Y(n_502)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_487),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_497),
.B(n_490),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_501),
.B(n_505),
.Y(n_506)
);

O2A1O1Ixp33_ASAP7_75t_SL g503 ( 
.A1(n_499),
.A2(n_486),
.B(n_480),
.C(n_473),
.Y(n_503)
);

CKINVDCx16_ASAP7_75t_R g507 ( 
.A(n_503),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_498),
.B(n_485),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_SL g508 ( 
.A1(n_502),
.A2(n_500),
.B(n_496),
.Y(n_508)
);

AO21x2_ASAP7_75t_L g510 ( 
.A1(n_508),
.A2(n_504),
.B(n_493),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_506),
.B(n_498),
.Y(n_509)
);

OAI21xp33_ASAP7_75t_L g511 ( 
.A1(n_509),
.A2(n_510),
.B(n_507),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_511),
.A2(n_492),
.B(n_468),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_512),
.B(n_476),
.C(n_473),
.Y(n_513)
);

AOI21xp5_ASAP7_75t_L g514 ( 
.A1(n_513),
.A2(n_368),
.B(n_0),
.Y(n_514)
);


endmodule