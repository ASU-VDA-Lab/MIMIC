module real_jpeg_6241_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_0),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_0),
.Y(n_232)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_0),
.Y(n_244)
);

BUFx5_ASAP7_75t_L g287 ( 
.A(n_0),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_0),
.Y(n_324)
);

INVx8_ASAP7_75t_L g431 ( 
.A(n_0),
.Y(n_431)
);

OAI22xp33_ASAP7_75t_L g141 ( 
.A1(n_1),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_1),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_1),
.A2(n_142),
.B1(n_285),
.B2(n_286),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_SL g377 ( 
.A1(n_1),
.A2(n_142),
.B1(n_169),
.B2(n_217),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_1),
.A2(n_68),
.B1(n_142),
.B2(n_403),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_2),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_2),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_2),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g348 ( 
.A(n_2),
.Y(n_348)
);

INVx6_ASAP7_75t_L g363 ( 
.A(n_2),
.Y(n_363)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_2),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_3),
.A2(n_82),
.B1(n_84),
.B2(n_87),
.Y(n_81)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_3),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_3),
.A2(n_87),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g386 ( 
.A1(n_3),
.A2(n_87),
.B1(n_115),
.B2(n_197),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_3),
.A2(n_87),
.B1(n_417),
.B2(n_418),
.Y(n_416)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_4),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_5),
.A2(n_48),
.B1(n_50),
.B2(n_52),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_5),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_5),
.A2(n_52),
.B1(n_318),
.B2(n_321),
.Y(n_317)
);

OAI22xp33_ASAP7_75t_SL g391 ( 
.A1(n_5),
.A2(n_52),
.B1(n_392),
.B2(n_393),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_SL g404 ( 
.A1(n_5),
.A2(n_52),
.B1(n_289),
.B2(n_405),
.Y(n_404)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_6),
.A2(n_169),
.B1(n_171),
.B2(n_173),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_6),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_6),
.B(n_112),
.C(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_6),
.B(n_73),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_6),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_6),
.B(n_178),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_6),
.B(n_92),
.Y(n_274)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_7),
.Y(n_513)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_8),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_8),
.Y(n_107)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_9),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_10),
.A2(n_90),
.B1(n_94),
.B2(n_95),
.Y(n_89)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_10),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_10),
.A2(n_95),
.B1(n_101),
.B2(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_10),
.A2(n_95),
.B1(n_388),
.B2(n_389),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_11),
.A2(n_216),
.B1(n_218),
.B2(n_219),
.Y(n_215)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_11),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_11),
.A2(n_218),
.B1(n_237),
.B2(n_240),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_11),
.A2(n_92),
.B1(n_218),
.B2(n_309),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_11),
.A2(n_48),
.B1(n_218),
.B2(n_367),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_12),
.Y(n_116)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_12),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_12),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_13),
.A2(n_101),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_13),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_13),
.A2(n_177),
.B1(n_207),
.B2(n_211),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_13),
.A2(n_177),
.B1(n_277),
.B2(n_279),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_13),
.A2(n_177),
.B1(n_367),
.B2(n_368),
.Y(n_366)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_14),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_15),
.A2(n_192),
.B1(n_196),
.B2(n_197),
.Y(n_191)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_15),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_15),
.A2(n_196),
.B1(n_266),
.B2(n_267),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g372 ( 
.A1(n_15),
.A2(n_196),
.B1(n_309),
.B2(n_373),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_15),
.A2(n_51),
.B1(n_196),
.B2(n_411),
.Y(n_410)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_16),
.A2(n_56),
.B1(n_57),
.B2(n_60),
.Y(n_55)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_16),
.A2(n_60),
.B1(n_152),
.B2(n_154),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g353 ( 
.A1(n_16),
.A2(n_60),
.B1(n_184),
.B2(n_354),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_16),
.A2(n_60),
.B1(n_123),
.B2(n_397),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_17),
.Y(n_516)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_511),
.B(n_514),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_158),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_156),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_133),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_23),
.B(n_133),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_124),
.B2(n_125),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_61),
.C(n_96),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_26),
.B(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_47),
.B1(n_53),
.B2(n_55),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_27),
.A2(n_53),
.B1(n_55),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_27),
.A2(n_47),
.B1(n_53),
.B2(n_140),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_27),
.A2(n_365),
.B(n_410),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_27),
.A2(n_37),
.B1(n_410),
.B2(n_434),
.Y(n_433)
);

INVx3_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_28),
.A2(n_361),
.B(n_364),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_28),
.B(n_366),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_37),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_SL g46 ( 
.A(n_32),
.Y(n_46)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_35),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_35),
.Y(n_369)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_37),
.B(n_173),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_39),
.B1(n_43),
.B2(n_46),
.Y(n_37)
);

OAI32xp33_ASAP7_75t_L g333 ( 
.A1(n_38),
.A2(n_334),
.A3(n_337),
.B1(n_340),
.B2(n_345),
.Y(n_333)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_41),
.Y(n_155)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_42),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_42),
.Y(n_280)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g403 ( 
.A(n_45),
.Y(n_403)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_53),
.A2(n_434),
.B(n_456),
.Y(n_466)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_54),
.B(n_366),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_54),
.B(n_141),
.Y(n_455)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_61),
.A2(n_96),
.B1(n_97),
.B2(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_61),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_81),
.B1(n_88),
.B2(n_89),
.Y(n_61)
);

INVx3_ASAP7_75t_SL g127 ( 
.A(n_62),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_62),
.A2(n_81),
.B1(n_88),
.B2(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_62),
.A2(n_88),
.B1(n_308),
.B2(n_372),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_62),
.A2(n_88),
.B1(n_402),
.B2(n_404),
.Y(n_401)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_73),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_68),
.B1(n_69),
.B2(n_71),
.Y(n_63)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_64),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_67),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_70),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_72),
.Y(n_153)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_72),
.Y(n_272)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_72),
.Y(n_336)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_72),
.Y(n_344)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_72),
.Y(n_408)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_73),
.A2(n_127),
.B(n_128),
.Y(n_126)
);

AOI22x1_ASAP7_75t_L g435 ( 
.A1(n_73),
.A2(n_127),
.B1(n_313),
.B2(n_436),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_73),
.A2(n_127),
.B1(n_151),
.B2(n_444),
.Y(n_443)
);

AO22x2_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_78),
.B2(n_80),
.Y(n_73)
);

INVx8_ASAP7_75t_L g291 ( 
.A(n_75),
.Y(n_291)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_76),
.Y(n_217)
);

INVx6_ASAP7_75t_L g399 ( 
.A(n_76),
.Y(n_399)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g172 ( 
.A(n_77),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_77),
.Y(n_220)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_77),
.Y(n_395)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_88),
.B(n_276),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_88),
.A2(n_308),
.B(n_312),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx5_ASAP7_75t_L g311 ( 
.A(n_93),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_96),
.B(n_139),
.C(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_96),
.A2(n_97),
.B1(n_148),
.B2(n_149),
.Y(n_500)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_111),
.B(n_122),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_98),
.A2(n_168),
.B(n_174),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_98),
.A2(n_215),
.B1(n_264),
.B2(n_265),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_98),
.A2(n_174),
.B(n_265),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_98),
.A2(n_264),
.B1(n_377),
.B2(n_425),
.Y(n_424)
);

INVx2_ASAP7_75t_SL g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_99),
.B(n_175),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_99),
.A2(n_178),
.B1(n_391),
.B2(n_396),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_99),
.A2(n_178),
.B1(n_396),
.B2(n_416),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_99),
.A2(n_178),
.B1(n_416),
.B2(n_447),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_111),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_103),
.B1(n_106),
.B2(n_108),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_102),
.Y(n_176)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_105),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_108),
.Y(n_181)
);

INVx5_ASAP7_75t_SL g268 ( 
.A(n_108),
.Y(n_268)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_109),
.Y(n_170)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_111),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_111),
.A2(n_215),
.B(n_221),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_111),
.A2(n_221),
.B(n_377),
.Y(n_376)
);

AOI22x1_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_114),
.B1(n_117),
.B2(n_119),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_SL g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_116),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_116),
.Y(n_211)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_122),
.Y(n_447)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_123),
.Y(n_266)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_127),
.A2(n_271),
.B(n_275),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_127),
.B(n_313),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_127),
.A2(n_275),
.B(n_469),
.Y(n_468)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_131),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_138),
.C(n_146),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_134),
.A2(n_135),
.B1(n_138),
.B2(n_139),
.Y(n_506)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_138),
.A2(n_139),
.B1(n_500),
.B2(n_501),
.Y(n_499)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx8_ASAP7_75t_L g339 ( 
.A(n_143),
.Y(n_339)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_146),
.A2(n_147),
.B1(n_505),
.B2(n_506),
.Y(n_504)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_154),
.Y(n_289)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx5_ASAP7_75t_L g375 ( 
.A(n_155),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_495),
.B(n_508),
.Y(n_159)
);

OAI311xp33_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_380),
.A3(n_471),
.B1(n_489),
.C1(n_494),
.Y(n_160)
);

AOI21x1_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_327),
.B(n_379),
.Y(n_161)
);

AO21x1_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_299),
.B(n_326),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_258),
.B(n_298),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_224),
.B(n_257),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_189),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_166),
.B(n_189),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_179),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_167),
.A2(n_179),
.B1(n_180),
.B2(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_167),
.Y(n_255)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NAND2xp33_ASAP7_75t_SL g296 ( 
.A(n_171),
.B(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_171),
.Y(n_418)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx3_ASAP7_75t_SL g417 ( 
.A(n_172),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_173),
.A2(n_199),
.B(n_204),
.Y(n_233)
);

OAI21xp33_ASAP7_75t_SL g271 ( 
.A1(n_173),
.A2(n_272),
.B(n_273),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_173),
.B(n_346),
.Y(n_345)
);

OAI21xp33_ASAP7_75t_SL g361 ( 
.A1(n_173),
.A2(n_345),
.B(n_362),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_178),
.Y(n_174)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_178),
.Y(n_264)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_188),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_212),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_190),
.B(n_213),
.C(n_223),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_199),
.B(n_204),
.Y(n_190)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_191),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_193),
.Y(n_192)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_194),
.Y(n_322)
);

BUFx5_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_195),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_195),
.Y(n_203)
);

BUFx8_ASAP7_75t_L g242 ( 
.A(n_195),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_198),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_199),
.A2(n_230),
.B1(n_351),
.B2(n_352),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_199),
.A2(n_253),
.B1(n_386),
.B2(n_387),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g419 ( 
.A1(n_199),
.A2(n_387),
.B(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_200),
.B(n_206),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_200),
.A2(n_250),
.B1(n_251),
.B2(n_252),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_200),
.A2(n_284),
.B1(n_317),
.B2(n_323),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_200),
.A2(n_353),
.B1(n_427),
.B2(n_428),
.Y(n_426)
);

OR2x2_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_201),
.Y(n_205)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_202),
.Y(n_286)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_205),
.Y(n_253)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_207),
.Y(n_228)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx4_ASAP7_75t_L g388 ( 
.A(n_209),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_210),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_222),
.B2(n_223),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx11_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_248),
.B(n_256),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_234),
.B(n_247),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_233),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_246),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_235),
.B(n_246),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_243),
.B(n_245),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_236),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g389 ( 
.A(n_237),
.Y(n_389)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx8_ASAP7_75t_L g285 ( 
.A(n_242),
.Y(n_285)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_245),
.A2(n_283),
.B(n_287),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_254),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_254),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_253),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_259),
.B(n_260),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_281),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_262),
.A2(n_263),
.B1(n_269),
.B2(n_270),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_263),
.B(n_269),
.C(n_281),
.Y(n_300)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVxp33_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

AOI32xp33_ASAP7_75t_L g288 ( 
.A1(n_274),
.A2(n_289),
.A3(n_290),
.B1(n_292),
.B2(n_296),
.Y(n_288)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_276),
.Y(n_313)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx6_ASAP7_75t_SL g279 ( 
.A(n_280),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_288),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_282),
.B(n_288),
.Y(n_305)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_285),
.Y(n_354)
);

INVx3_ASAP7_75t_SL g290 ( 
.A(n_291),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_291),
.Y(n_392)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx8_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_300),
.B(n_301),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_303),
.B1(n_306),
.B2(n_325),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_304),
.B(n_305),
.C(n_325),
.Y(n_328)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_306),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_314),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_307),
.B(n_315),
.C(n_316),
.Y(n_355)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_317),
.Y(n_351)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

CKINVDCx14_ASAP7_75t_R g321 ( 
.A(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_323),
.Y(n_420)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_328),
.B(n_329),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_358),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_331),
.A2(n_355),
.B1(n_356),
.B2(n_357),
.Y(n_330)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_331),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_332),
.A2(n_333),
.B1(n_349),
.B2(n_350),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_333),
.B(n_349),
.Y(n_467)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx4_ASAP7_75t_L g367 ( 
.A(n_339),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_343),
.Y(n_340)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx4_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_355),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_355),
.B(n_356),
.C(n_358),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_360),
.B1(n_370),
.B2(n_378),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_359),
.B(n_371),
.C(n_376),
.Y(n_480)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx8_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_370),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_371),
.B(n_376),
.Y(n_370)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_372),
.Y(n_469)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx4_ASAP7_75t_SL g374 ( 
.A(n_375),
.Y(n_374)
);

NAND2xp33_ASAP7_75t_SL g380 ( 
.A(n_381),
.B(n_457),
.Y(n_380)
);

A2O1A1Ixp33_ASAP7_75t_SL g489 ( 
.A1(n_381),
.A2(n_457),
.B(n_490),
.C(n_493),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_437),
.Y(n_381)
);

OR2x2_ASAP7_75t_L g494 ( 
.A(n_382),
.B(n_437),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_413),
.C(n_422),
.Y(n_382)
);

FAx1_ASAP7_75t_SL g470 ( 
.A(n_383),
.B(n_413),
.CI(n_422),
.CON(n_470),
.SN(n_470)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_400),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_384),
.B(n_401),
.C(n_409),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_390),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_385),
.B(n_390),
.Y(n_463)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_386),
.Y(n_427)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_391),
.Y(n_425)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

BUFx3_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx6_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_409),
.Y(n_400)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_402),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_404),
.Y(n_444)
);

INVx1_ASAP7_75t_SL g405 ( 
.A(n_406),
.Y(n_405)
);

INVx5_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx4_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_414),
.A2(n_415),
.B1(n_419),
.B2(n_421),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_415),
.B(n_419),
.Y(n_451)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_419),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_419),
.A2(n_421),
.B1(n_453),
.B2(n_454),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g498 ( 
.A1(n_419),
.A2(n_451),
.B(n_454),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_432),
.C(n_435),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_423),
.B(n_461),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_424),
.B(n_426),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_424),
.B(n_426),
.Y(n_479)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx8_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_432),
.A2(n_433),
.B1(n_435),
.B2(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_SL g462 ( 
.A(n_435),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_439),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_438),
.B(n_441),
.C(n_449),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_440),
.A2(n_441),
.B1(n_449),
.B2(n_450),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_442),
.A2(n_445),
.B(n_448),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_443),
.B(n_446),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

FAx1_ASAP7_75t_SL g497 ( 
.A(n_448),
.B(n_498),
.CI(n_499),
.CON(n_497),
.SN(n_497)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_448),
.B(n_498),
.C(n_499),
.Y(n_507)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_452),
.Y(n_450)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_456),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_470),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_458),
.B(n_470),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_463),
.C(n_464),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_459),
.A2(n_460),
.B1(n_463),
.B2(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_463),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_464),
.B(n_482),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_467),
.C(n_468),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_465),
.A2(n_466),
.B1(n_468),
.B2(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_467),
.B(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_468),
.Y(n_477)
);

BUFx24_ASAP7_75t_SL g517 ( 
.A(n_470),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_472),
.B(n_484),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_473),
.A2(n_491),
.B(n_492),
.Y(n_490)
);

NOR2x1_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_481),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_474),
.B(n_481),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_475),
.B(n_478),
.C(n_480),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_475),
.B(n_487),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_478),
.A2(n_479),
.B1(n_480),
.B2(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_480),
.Y(n_488)
);

OR2x2_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_486),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_485),
.B(n_486),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_496),
.B(n_503),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_SL g496 ( 
.A(n_497),
.B(n_502),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_497),
.B(n_502),
.Y(n_509)
);

BUFx24_ASAP7_75t_SL g518 ( 
.A(n_497),
.Y(n_518)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_500),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_503),
.A2(n_509),
.B(n_510),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_504),
.B(n_507),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_504),
.B(n_507),
.Y(n_510)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

BUFx4f_ASAP7_75t_SL g511 ( 
.A(n_512),
.Y(n_511)
);

INVx13_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVx5_ASAP7_75t_L g515 ( 
.A(n_513),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_515),
.B(n_516),
.Y(n_514)
);


endmodule