module fake_jpeg_31570_n_500 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_500);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_500;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_13),
.B(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

BUFx8_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_51),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_53),
.Y(n_123)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_54),
.Y(n_119)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_56),
.Y(n_132)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_58),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_29),
.B(n_7),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_59),
.B(n_61),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_60),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_29),
.B(n_7),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_62),
.Y(n_134)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_63),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_64),
.Y(n_126)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_28),
.Y(n_65)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_65),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_7),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_66),
.B(n_72),
.Y(n_107)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_67),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_68),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_18),
.B(n_38),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_69),
.B(n_25),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

CKINVDCx6p67_ASAP7_75t_R g145 ( 
.A(n_70),
.Y(n_145)
);

NAND2x1_ASAP7_75t_L g71 ( 
.A(n_37),
.B(n_48),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_71),
.A2(n_48),
.B(n_14),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_25),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_73),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx8_ASAP7_75t_L g137 ( 
.A(n_74),
.Y(n_137)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_75),
.Y(n_130)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_76),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g77 ( 
.A(n_19),
.Y(n_77)
);

INVx4_ASAP7_75t_SL g116 ( 
.A(n_77),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_18),
.B(n_9),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_80),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_79),
.Y(n_160)
);

INVx6_ASAP7_75t_SL g80 ( 
.A(n_45),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_81),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_17),
.Y(n_83)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_83),
.Y(n_143)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_84),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_85),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_24),
.B(n_9),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_100),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_87),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_88),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_89),
.Y(n_150)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_19),
.Y(n_90)
);

INVx2_ASAP7_75t_SL g140 ( 
.A(n_90),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_91),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_92),
.Y(n_161)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_93),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

BUFx10_ASAP7_75t_L g153 ( 
.A(n_94),
.Y(n_153)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_95),
.Y(n_155)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_96),
.Y(n_156)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_27),
.Y(n_97)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_40),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_99),
.A2(n_44),
.B1(n_25),
.B2(n_47),
.Y(n_147)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_41),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_31),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_101),
.B(n_102),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_24),
.B(n_9),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_63),
.A2(n_31),
.B1(n_35),
.B2(n_34),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_103),
.A2(n_108),
.B1(n_113),
.B2(n_118),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_78),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_106),
.B(n_79),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_66),
.A2(n_38),
.B1(n_36),
.B2(n_39),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_52),
.A2(n_35),
.B1(n_34),
.B2(n_39),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_SL g114 ( 
.A(n_87),
.Y(n_114)
);

INVx11_ASAP7_75t_L g208 ( 
.A(n_114),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_86),
.A2(n_33),
.B1(n_32),
.B2(n_36),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_58),
.A2(n_35),
.B1(n_33),
.B2(n_43),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_121),
.A2(n_157),
.B1(n_64),
.B2(n_91),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_127),
.B(n_88),
.Y(n_175)
);

AOI21xp33_ASAP7_75t_SL g133 ( 
.A1(n_71),
.A2(n_44),
.B(n_25),
.Y(n_133)
);

XNOR2x1_ASAP7_75t_SL g197 ( 
.A(n_133),
.B(n_151),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_136),
.B(n_152),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_147),
.A2(n_94),
.B1(n_79),
.B2(n_47),
.Y(n_185)
);

AOI21xp33_ASAP7_75t_L g151 ( 
.A1(n_102),
.A2(n_55),
.B(n_44),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_77),
.B(n_44),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_60),
.A2(n_43),
.B1(n_20),
.B2(n_12),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_89),
.A2(n_10),
.B1(n_16),
.B2(n_15),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_158),
.A2(n_12),
.B1(n_16),
.B2(n_15),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_162),
.Y(n_244)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_163),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_153),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_164),
.B(n_169),
.Y(n_237)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_105),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_165),
.Y(n_225)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_149),
.Y(n_166)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_166),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_62),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_167),
.B(n_168),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_117),
.B(n_82),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_145),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_122),
.B(n_74),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_170),
.B(n_177),
.Y(n_226)
);

INVx4_ASAP7_75t_SL g171 ( 
.A(n_104),
.Y(n_171)
);

BUFx2_ASAP7_75t_SL g246 ( 
.A(n_171),
.Y(n_246)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_150),
.Y(n_172)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_172),
.Y(n_250)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_154),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_173),
.Y(n_229)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_156),
.Y(n_174)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_174),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_175),
.A2(n_207),
.B1(n_140),
.B2(n_126),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_107),
.B(n_99),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_176),
.B(n_192),
.C(n_198),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_111),
.B(n_68),
.Y(n_177)
);

BUFx12f_ASAP7_75t_L g178 ( 
.A(n_145),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_178),
.Y(n_222)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_131),
.Y(n_179)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_179),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_145),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_180),
.B(n_194),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_112),
.Y(n_181)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_181),
.Y(n_227)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_116),
.Y(n_182)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_182),
.Y(n_241)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_148),
.Y(n_183)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_183),
.Y(n_251)
);

FAx1_ASAP7_75t_SL g184 ( 
.A(n_110),
.B(n_70),
.CI(n_94),
.CON(n_184),
.SN(n_184)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_184),
.B(n_202),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_185),
.A2(n_187),
.B1(n_205),
.B2(n_158),
.Y(n_240)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_116),
.Y(n_186)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_186),
.Y(n_252)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_137),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_188),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_132),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_189),
.Y(n_216)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_146),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_190),
.Y(n_224)
);

AND2x2_ASAP7_75t_SL g192 ( 
.A(n_115),
.B(n_0),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_114),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_193),
.Y(n_236)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_125),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_124),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_195),
.B(n_196),
.Y(n_233)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_143),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_123),
.B(n_92),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_109),
.B(n_70),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_199),
.B(n_140),
.C(n_144),
.Y(n_235)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_120),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_200),
.B(n_201),
.Y(n_234)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_120),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_153),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_147),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_203),
.B(n_204),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_159),
.A2(n_20),
.B1(n_47),
.B2(n_12),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_153),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_209),
.B(n_210),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_160),
.B(n_47),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_155),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_211),
.B(n_212),
.Y(n_253)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_135),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_126),
.B(n_5),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_113),
.Y(n_219)
);

INVx4_ASAP7_75t_SL g214 ( 
.A(n_130),
.Y(n_214)
);

AND2x2_ASAP7_75t_SL g232 ( 
.A(n_214),
.B(n_141),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_215),
.A2(n_247),
.B1(n_248),
.B2(n_170),
.Y(n_264)
);

XNOR2x1_ASAP7_75t_L g272 ( 
.A(n_219),
.B(n_235),
.Y(n_272)
);

AOI32xp33_ASAP7_75t_L g223 ( 
.A1(n_197),
.A2(n_142),
.A3(n_138),
.B1(n_119),
.B2(n_161),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_223),
.B(n_245),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_184),
.A2(n_135),
.B1(n_159),
.B2(n_161),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_230),
.A2(n_240),
.B1(n_249),
.B2(n_254),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_232),
.Y(n_279)
);

AOI32xp33_ASAP7_75t_L g245 ( 
.A1(n_197),
.A2(n_144),
.A3(n_103),
.B1(n_121),
.B2(n_141),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_206),
.A2(n_134),
.B1(n_129),
.B2(n_128),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_206),
.A2(n_134),
.B1(n_129),
.B2(n_128),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_187),
.A2(n_112),
.B1(n_1),
.B2(n_2),
.Y(n_249)
);

OAI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_184),
.A2(n_16),
.B1(n_5),
.B2(n_4),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_191),
.B(n_0),
.C(n_1),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_255),
.B(n_192),
.C(n_175),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_257),
.B(n_258),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_220),
.B(n_175),
.C(n_176),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_245),
.A2(n_163),
.B1(n_214),
.B2(n_188),
.Y(n_260)
);

OAI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_260),
.A2(n_232),
.B1(n_246),
.B2(n_256),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_226),
.B(n_218),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_261),
.B(n_269),
.Y(n_294)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_253),
.Y(n_262)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_262),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_220),
.B(n_176),
.C(n_199),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_263),
.B(n_266),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g307 ( 
.A1(n_264),
.A2(n_271),
.B1(n_261),
.B2(n_268),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_253),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_265),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_228),
.A2(n_177),
.B(n_167),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_240),
.A2(n_198),
.B1(n_192),
.B2(n_199),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_267),
.A2(n_274),
.B1(n_284),
.B2(n_286),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_218),
.B(n_168),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_228),
.A2(n_185),
.B(n_183),
.Y(n_270)
);

OA21x2_ASAP7_75t_L g295 ( 
.A1(n_270),
.A2(n_276),
.B(n_232),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_233),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_271),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_226),
.B(n_213),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_273),
.B(n_277),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_219),
.A2(n_198),
.B1(n_190),
.B2(n_179),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_234),
.Y(n_275)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_275),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_238),
.A2(n_172),
.B(n_178),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_247),
.A2(n_181),
.B1(n_201),
.B2(n_212),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_233),
.B(n_166),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_278),
.B(n_281),
.Y(n_317)
);

OAI32xp33_ASAP7_75t_L g280 ( 
.A1(n_238),
.A2(n_178),
.A3(n_200),
.B1(n_162),
.B2(n_196),
.Y(n_280)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_280),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_242),
.B(n_189),
.Y(n_281)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_231),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g318 ( 
.A(n_282),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_248),
.A2(n_208),
.B1(n_193),
.B2(n_171),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_283),
.B(n_285),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_249),
.A2(n_208),
.B1(n_1),
.B2(n_2),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_241),
.B(n_4),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_223),
.A2(n_4),
.B1(n_6),
.B2(n_14),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_234),
.Y(n_287)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_287),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_215),
.A2(n_4),
.B1(n_6),
.B2(n_14),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_288),
.A2(n_227),
.B1(n_216),
.B2(n_225),
.Y(n_309)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_217),
.Y(n_289)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_289),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_242),
.A2(n_15),
.B(n_0),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_237),
.Y(n_299)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_217),
.Y(n_291)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_291),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_255),
.B(n_235),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_292),
.B(n_252),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_295),
.A2(n_304),
.B(n_276),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_298),
.B(n_260),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_299),
.B(n_272),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_272),
.B(n_243),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_301),
.B(n_305),
.Y(n_332)
);

NAND2xp33_ASAP7_75t_SL g304 ( 
.A(n_278),
.B(n_241),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_270),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_306),
.B(n_308),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_307),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_L g308 ( 
.A1(n_268),
.A2(n_231),
.B1(n_225),
.B2(n_252),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_309),
.B(n_316),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_265),
.B(n_224),
.Y(n_316)
);

CKINVDCx14_ASAP7_75t_R g320 ( 
.A(n_281),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_323),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_259),
.A2(n_275),
.B1(n_287),
.B2(n_286),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_321),
.A2(n_259),
.B1(n_267),
.B2(n_315),
.Y(n_337)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_289),
.Y(n_322)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_322),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_269),
.B(n_224),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_285),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_324),
.B(n_290),
.Y(n_336)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_291),
.Y(n_325)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_325),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_316),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_326),
.B(n_347),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_309),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_327),
.B(n_345),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_317),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_329),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_314),
.B(n_272),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_333),
.B(n_340),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_295),
.A2(n_302),
.B(n_319),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g382 ( 
.A1(n_335),
.A2(n_355),
.B(n_303),
.Y(n_382)
);

CKINVDCx14_ASAP7_75t_R g366 ( 
.A(n_336),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_337),
.A2(n_341),
.B1(n_354),
.B2(n_303),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_339),
.B(n_305),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_314),
.B(n_258),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_342),
.B(n_295),
.Y(n_357)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_311),
.Y(n_344)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_344),
.Y(n_360)
);

CKINVDCx14_ASAP7_75t_R g345 ( 
.A(n_319),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_311),
.Y(n_346)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_346),
.Y(n_361)
);

INVxp33_ASAP7_75t_L g347 ( 
.A(n_317),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_324),
.B(n_266),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_348),
.B(n_320),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_297),
.B(n_273),
.Y(n_349)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_349),
.Y(n_374)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_312),
.Y(n_350)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_350),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_297),
.B(n_262),
.Y(n_351)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_351),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_313),
.B(n_274),
.Y(n_352)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_352),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_313),
.B(n_276),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_353),
.B(n_356),
.Y(n_367)
);

OAI22x1_ASAP7_75t_L g354 ( 
.A1(n_295),
.A2(n_280),
.B1(n_279),
.B2(n_283),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_302),
.A2(n_258),
.B(n_222),
.Y(n_355)
);

OR2x2_ASAP7_75t_L g356 ( 
.A(n_321),
.B(n_264),
.Y(n_356)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_357),
.A2(n_382),
.B(n_341),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_359),
.A2(n_356),
.B1(n_345),
.B2(n_327),
.Y(n_388)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_362),
.Y(n_391)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_338),
.Y(n_365)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_365),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_333),
.B(n_340),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_368),
.B(n_372),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_339),
.B(n_296),
.C(n_301),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_369),
.B(n_383),
.C(n_385),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_332),
.B(n_296),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_335),
.Y(n_373)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_373),
.Y(n_409)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_338),
.Y(n_376)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_376),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_SL g405 ( 
.A(n_377),
.B(n_331),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_332),
.B(n_299),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_378),
.B(n_351),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_349),
.B(n_323),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_379),
.B(n_326),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_348),
.B(n_315),
.Y(n_381)
);

CKINVDCx16_ASAP7_75t_R g404 ( 
.A(n_381),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_355),
.B(n_292),
.C(n_257),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_336),
.B(n_294),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g397 ( 
.A(n_384),
.B(n_329),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_337),
.B(n_257),
.C(n_263),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_330),
.B(n_263),
.C(n_294),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_386),
.B(n_352),
.C(n_310),
.Y(n_408)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_387),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_388),
.A2(n_393),
.B1(n_402),
.B2(n_375),
.Y(n_422)
);

XOR2x1_ASAP7_75t_L g389 ( 
.A(n_357),
.B(n_342),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_SL g412 ( 
.A(n_389),
.B(n_403),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_366),
.A2(n_354),
.B1(n_357),
.B2(n_380),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_390),
.A2(n_383),
.B1(n_310),
.B2(n_300),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_359),
.A2(n_356),
.B1(n_328),
.B2(n_354),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_394),
.B(n_399),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_371),
.B(n_331),
.Y(n_396)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_396),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_397),
.B(n_410),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_363),
.B(n_353),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_401),
.A2(n_407),
.B(n_411),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_358),
.A2(n_380),
.B1(n_367),
.B2(n_328),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_363),
.B(n_368),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_SL g431 ( 
.A(n_405),
.B(n_406),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_369),
.B(n_334),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_SL g407 ( 
.A(n_382),
.B(n_334),
.C(n_304),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_408),
.B(n_372),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_379),
.B(n_293),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_358),
.A2(n_350),
.B(n_346),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_391),
.B(n_386),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_413),
.B(n_418),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g418 ( 
.A(n_404),
.B(n_374),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_419),
.B(n_322),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_403),
.B(n_400),
.C(n_392),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_420),
.B(n_428),
.C(n_429),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_408),
.B(n_370),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_421),
.B(n_426),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_422),
.B(n_424),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_390),
.A2(n_374),
.B1(n_375),
.B2(n_367),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_423),
.A2(n_407),
.B1(n_393),
.B2(n_388),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_401),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_396),
.B(n_293),
.Y(n_427)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_427),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_400),
.B(n_385),
.C(n_377),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_392),
.B(n_378),
.C(n_300),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_409),
.B(n_364),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_430),
.B(n_395),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_415),
.B(n_399),
.Y(n_432)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_432),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_436),
.A2(n_437),
.B1(n_417),
.B2(n_416),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_417),
.A2(n_402),
.B1(n_411),
.B2(n_398),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_420),
.B(n_394),
.C(n_406),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_438),
.B(n_443),
.C(n_444),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_426),
.A2(n_387),
.B(n_389),
.Y(n_440)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_440),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_441),
.B(n_424),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_428),
.B(n_405),
.C(n_410),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_419),
.B(n_360),
.C(n_361),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_425),
.B(n_398),
.C(n_344),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_445),
.B(n_446),
.C(n_416),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_425),
.B(n_343),
.C(n_325),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_412),
.B(n_343),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_447),
.B(n_448),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_446),
.B(n_429),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_451),
.B(n_452),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_445),
.B(n_443),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_442),
.A2(n_415),
.B(n_414),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_453),
.B(n_457),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_455),
.B(n_288),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_433),
.B(n_412),
.C(n_422),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_456),
.B(n_435),
.C(n_447),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_439),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_458),
.B(n_459),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_433),
.B(n_431),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_460),
.B(n_463),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_444),
.B(n_431),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_461),
.B(n_438),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_434),
.B(n_435),
.Y(n_463)
);

OR2x2_ASAP7_75t_L g482 ( 
.A(n_465),
.B(n_469),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_466),
.B(n_475),
.Y(n_479)
);

AOI22xp33_ASAP7_75t_SL g467 ( 
.A1(n_462),
.A2(n_282),
.B1(n_318),
.B2(n_231),
.Y(n_467)
);

AOI21x1_ASAP7_75t_SL g484 ( 
.A1(n_467),
.A2(n_284),
.B(n_236),
.Y(n_484)
);

OAI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_454),
.A2(n_318),
.B(n_312),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_468),
.A2(n_449),
.B(n_222),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_452),
.B(n_454),
.C(n_455),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_470),
.B(n_473),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_450),
.A2(n_282),
.B1(n_277),
.B2(n_216),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_472),
.B(n_284),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_461),
.A2(n_227),
.B1(n_256),
.B2(n_251),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_451),
.B(n_251),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_477),
.B(n_480),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_469),
.B(n_456),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_481),
.B(n_483),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_476),
.B(n_474),
.Y(n_483)
);

AOI31xp33_ASAP7_75t_L g490 ( 
.A1(n_484),
.A2(n_236),
.A3(n_244),
.B(n_229),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_466),
.B(n_221),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_485),
.B(n_250),
.C(n_221),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_482),
.A2(n_471),
.B(n_464),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_SL g493 ( 
.A1(n_488),
.A2(n_489),
.B(n_486),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_479),
.A2(n_472),
.B(n_467),
.Y(n_489)
);

AO21x1_ASAP7_75t_L g494 ( 
.A1(n_490),
.A2(n_491),
.B(n_477),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g492 ( 
.A(n_487),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_492),
.A2(n_493),
.B(n_494),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_SL g496 ( 
.A1(n_492),
.A2(n_478),
.B(n_250),
.Y(n_496)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_496),
.A2(n_478),
.B(n_244),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_497),
.A2(n_495),
.B(n_239),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_498),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_499),
.B(n_239),
.Y(n_500)
);


endmodule