module fake_ariane_1033_n_1138 (n_83, n_8, n_233, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_240, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_269, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_237, n_172, n_69, n_259, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_242, n_260, n_274, n_115, n_272, n_133, n_66, n_205, n_236, n_265, n_71, n_267, n_24, n_7, n_109, n_208, n_245, n_96, n_156, n_209, n_49, n_262, n_20, n_174, n_275, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_235, n_200, n_51, n_166, n_253, n_76, n_218, n_103, n_79, n_26, n_244, n_226, n_3, n_246, n_271, n_46, n_220, n_0, n_84, n_247, n_261, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_263, n_201, n_229, n_70, n_250, n_222, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_256, n_6, n_214, n_227, n_48, n_94, n_101, n_243, n_4, n_134, n_188, n_185, n_2, n_32, n_249, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_264, n_129, n_126, n_137, n_255, n_278, n_122, n_268, n_257, n_266, n_198, n_148, n_232, n_164, n_52, n_277, n_157, n_248, n_184, n_177, n_135, n_258, n_73, n_77, n_171, n_228, n_15, n_118, n_93, n_121, n_276, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_241, n_29, n_254, n_238, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_231, n_192, n_28, n_80, n_146, n_234, n_230, n_211, n_270, n_194, n_97, n_154, n_215, n_252, n_142, n_251, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_239, n_223, n_35, n_273, n_54, n_25, n_1138);

input n_83;
input n_8;
input n_233;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_240;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_269;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_237;
input n_172;
input n_69;
input n_259;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_242;
input n_260;
input n_274;
input n_115;
input n_272;
input n_133;
input n_66;
input n_205;
input n_236;
input n_265;
input n_71;
input n_267;
input n_24;
input n_7;
input n_109;
input n_208;
input n_245;
input n_96;
input n_156;
input n_209;
input n_49;
input n_262;
input n_20;
input n_174;
input n_275;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_235;
input n_200;
input n_51;
input n_166;
input n_253;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_244;
input n_226;
input n_3;
input n_246;
input n_271;
input n_46;
input n_220;
input n_0;
input n_84;
input n_247;
input n_261;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_263;
input n_201;
input n_229;
input n_70;
input n_250;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_256;
input n_6;
input n_214;
input n_227;
input n_48;
input n_94;
input n_101;
input n_243;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_264;
input n_129;
input n_126;
input n_137;
input n_255;
input n_278;
input n_122;
input n_268;
input n_257;
input n_266;
input n_198;
input n_148;
input n_232;
input n_164;
input n_52;
input n_277;
input n_157;
input n_248;
input n_184;
input n_177;
input n_135;
input n_258;
input n_73;
input n_77;
input n_171;
input n_228;
input n_15;
input n_118;
input n_93;
input n_121;
input n_276;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_241;
input n_29;
input n_254;
input n_238;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_231;
input n_192;
input n_28;
input n_80;
input n_146;
input n_234;
input n_230;
input n_211;
input n_270;
input n_194;
input n_97;
input n_154;
input n_215;
input n_252;
input n_142;
input n_251;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_239;
input n_223;
input n_35;
input n_273;
input n_54;
input n_25;

output n_1138;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_1127;
wire n_1072;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_1137;
wire n_646;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_1118;
wire n_678;
wire n_1058;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_1042;
wire n_961;
wire n_469;
wire n_1046;
wire n_479;
wire n_726;
wire n_603;
wire n_1123;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_752;
wire n_341;
wire n_1029;
wire n_985;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_1109;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_643;
wire n_679;
wire n_924;
wire n_927;
wire n_781;
wire n_1095;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_1096;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_1130;
wire n_524;
wire n_634;
wire n_391;
wire n_349;
wire n_756;
wire n_466;
wire n_1016;
wire n_346;
wire n_940;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_1077;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_956;
wire n_949;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_1131;
wire n_891;
wire n_737;
wire n_885;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_1088;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_958;
wire n_945;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_1067;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_1064;
wire n_633;
wire n_900;
wire n_1133;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_1093;
wire n_473;
wire n_801;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_903;
wire n_315;
wire n_871;
wire n_1073;
wire n_594;
wire n_311;
wire n_402;
wire n_1052;
wire n_1068;
wire n_829;
wire n_1062;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_1117;
wire n_422;
wire n_1106;
wire n_648;
wire n_784;
wire n_597;
wire n_816;
wire n_1018;
wire n_855;
wire n_1047;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_1076;
wire n_753;
wire n_1050;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_1125;
wire n_625;
wire n_405;
wire n_557;
wire n_1107;
wire n_858;
wire n_645;
wire n_989;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_1134;
wire n_485;
wire n_401;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_1053;
wire n_1084;
wire n_398;
wire n_1090;
wire n_529;
wire n_502;
wire n_561;
wire n_770;
wire n_821;
wire n_839;
wire n_1099;
wire n_928;
wire n_465;
wire n_507;
wire n_486;
wire n_901;
wire n_759;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_1103;
wire n_971;
wire n_369;
wire n_787;
wire n_894;
wire n_1105;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_1061;
wire n_1045;
wire n_831;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_874;
wire n_323;
wire n_550;
wire n_1023;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_1116;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1113;
wire n_1034;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_467;
wire n_1085;
wire n_432;
wire n_545;
wire n_1015;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_325;
wire n_688;
wire n_1074;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_1098;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_352;
wire n_538;
wire n_899;
wire n_1080;
wire n_576;
wire n_843;
wire n_920;
wire n_511;
wire n_1086;
wire n_611;
wire n_1092;
wire n_365;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_1104;
wire n_638;
wire n_334;
wire n_1128;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_1048;
wire n_775;
wire n_667;
wire n_1122;
wire n_1049;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_1132;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_1059;
wire n_314;
wire n_684;
wire n_1120;
wire n_440;
wire n_627;
wire n_1039;
wire n_305;
wire n_539;
wire n_312;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_321;
wire n_911;
wire n_1136;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_1065;
wire n_453;
wire n_1119;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_1055;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_601;
wire n_683;
wire n_565;
wire n_1089;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_1121;
wire n_490;
wire n_743;
wire n_907;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_1112;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_747;
wire n_741;
wire n_772;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1114;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_1038;
wire n_572;
wire n_343;
wire n_865;
wire n_1041;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_1097;
wire n_710;
wire n_860;
wire n_534;
wire n_1108;
wire n_355;
wire n_444;
wire n_609;
wire n_851;
wire n_1043;
wire n_560;
wire n_450;
wire n_890;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_468;
wire n_1056;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_1040;
wire n_674;
wire n_1081;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_832;
wire n_535;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_629;
wire n_664;
wire n_1075;
wire n_454;
wire n_992;
wire n_966;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_1091;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_1063;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_1126;
wire n_395;
wire n_621;
wire n_606;
wire n_951;
wire n_1026;
wire n_938;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_509;
wire n_583;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_1100;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_622;
wire n_697;
wire n_967;
wire n_998;
wire n_1083;
wire n_999;
wire n_472;
wire n_937;
wire n_296;
wire n_746;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_1079;
wire n_704;
wire n_1060;
wire n_1044;
wire n_751;
wire n_615;
wire n_1027;
wire n_1070;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_1082;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_517;
wire n_925;
wire n_530;
wire n_1094;
wire n_792;
wire n_1001;
wire n_1115;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_1051;
wire n_719;
wire n_434;
wire n_360;
wire n_1101;
wire n_975;
wire n_1102;
wire n_1129;
wire n_563;
wire n_394;
wire n_923;
wire n_1124;
wire n_932;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_1110;
wire n_317;
wire n_867;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_1078;
wire n_972;
wire n_470;
wire n_457;
wire n_1087;
wire n_632;
wire n_477;
wire n_364;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_1054;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1071;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_736;
wire n_767;
wire n_1025;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_1057;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_1069;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_191),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_50),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_25),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_153),
.Y(n_282)
);

BUFx10_ASAP7_75t_L g283 ( 
.A(n_135),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_24),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_261),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_59),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_242),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_115),
.Y(n_288)
);

BUFx2_ASAP7_75t_SL g289 ( 
.A(n_174),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_73),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_23),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_92),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_187),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_83),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_183),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_235),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_124),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_139),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_194),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_111),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_155),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_166),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_217),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_21),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_199),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_247),
.Y(n_306)
);

BUFx10_ASAP7_75t_L g307 ( 
.A(n_42),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_227),
.Y(n_308)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_210),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_136),
.Y(n_310)
);

BUFx10_ASAP7_75t_L g311 ( 
.A(n_176),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_46),
.Y(n_312)
);

INVx2_ASAP7_75t_SL g313 ( 
.A(n_254),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_35),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_169),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_249),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_215),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_145),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_25),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_165),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_119),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_154),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_221),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_88),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_232),
.Y(n_325)
);

BUFx10_ASAP7_75t_L g326 ( 
.A(n_56),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_17),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_43),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_102),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_184),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_59),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_189),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_157),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_70),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_126),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_140),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_26),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_150),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_182),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_222),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_277),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_89),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_55),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_57),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_266),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_156),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_281),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_309),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_285),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_337),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_291),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_344),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_283),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_283),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_285),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_283),
.Y(n_356)
);

OR2x2_ASAP7_75t_L g357 ( 
.A(n_284),
.B(n_0),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_332),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_280),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_286),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_282),
.Y(n_361)
);

INVxp33_ASAP7_75t_L g362 ( 
.A(n_288),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_332),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_340),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_311),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_311),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_311),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_307),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_307),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_304),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_340),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_307),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_291),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_326),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_326),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_326),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_279),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_279),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_292),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_312),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_300),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_314),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_306),
.B(n_0),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_317),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_319),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_327),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_320),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_328),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_331),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_343),
.Y(n_390)
);

INVxp67_ASAP7_75t_SL g391 ( 
.A(n_313),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_361),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g393 ( 
.A(n_351),
.Y(n_393)
);

OAI21x1_ASAP7_75t_L g394 ( 
.A1(n_361),
.A2(n_324),
.B(n_322),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_355),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_355),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_359),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_358),
.Y(n_398)
);

AND2x2_ASAP7_75t_SL g399 ( 
.A(n_357),
.B(n_329),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_379),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_353),
.B(n_313),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_358),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_360),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_R g404 ( 
.A(n_377),
.B(n_378),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_364),
.Y(n_405)
);

NOR2xp67_ASAP7_75t_L g406 ( 
.A(n_377),
.B(n_287),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_347),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_350),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_391),
.B(n_330),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_352),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_R g411 ( 
.A(n_378),
.B(n_290),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_381),
.Y(n_412)
);

OA21x2_ASAP7_75t_L g413 ( 
.A1(n_384),
.A2(n_334),
.B(n_333),
.Y(n_413)
);

AND3x1_ASAP7_75t_L g414 ( 
.A(n_383),
.B(n_369),
.C(n_368),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_387),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_364),
.Y(n_416)
);

AND2x4_ASAP7_75t_L g417 ( 
.A(n_354),
.B(n_342),
.Y(n_417)
);

BUFx8_ASAP7_75t_L g418 ( 
.A(n_372),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_356),
.B(n_293),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_375),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_365),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_366),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_367),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_376),
.Y(n_424)
);

OAI21x1_ASAP7_75t_L g425 ( 
.A1(n_362),
.A2(n_289),
.B(n_321),
.Y(n_425)
);

OAI21x1_ASAP7_75t_L g426 ( 
.A1(n_370),
.A2(n_321),
.B(n_295),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_348),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_348),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_380),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_380),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_382),
.B(n_294),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_382),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_385),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_349),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_385),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_386),
.B(n_321),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_363),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_386),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_371),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_R g440 ( 
.A(n_388),
.B(n_296),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_388),
.B(n_297),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_389),
.B(n_321),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_390),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_436),
.B(n_389),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_422),
.B(n_298),
.Y(n_445)
);

BUFx10_ASAP7_75t_L g446 ( 
.A(n_431),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_422),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_422),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_SL g449 ( 
.A(n_399),
.B(n_374),
.Y(n_449)
);

NOR2x1p5_ASAP7_75t_L g450 ( 
.A(n_430),
.B(n_299),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_436),
.B(n_301),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_430),
.B(n_302),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_392),
.Y(n_453)
);

INVx2_ASAP7_75t_SL g454 ( 
.A(n_430),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_393),
.B(n_373),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_407),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_443),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_442),
.B(n_303),
.Y(n_458)
);

OR2x2_ASAP7_75t_L g459 ( 
.A(n_428),
.B(n_427),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_443),
.Y(n_460)
);

OR2x6_ASAP7_75t_L g461 ( 
.A(n_403),
.B(n_1),
.Y(n_461)
);

INVx2_ASAP7_75t_SL g462 ( 
.A(n_430),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_392),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_408),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_394),
.Y(n_465)
);

AND2x6_ASAP7_75t_L g466 ( 
.A(n_442),
.B(n_61),
.Y(n_466)
);

INVx5_ASAP7_75t_L g467 ( 
.A(n_422),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_394),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_427),
.B(n_428),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_422),
.B(n_346),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_413),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_423),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_410),
.Y(n_473)
);

O2A1O1Ixp33_ASAP7_75t_L g474 ( 
.A1(n_424),
.A2(n_3),
.B(n_1),
.C(n_2),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_413),
.Y(n_475)
);

AND2x6_ASAP7_75t_L g476 ( 
.A(n_430),
.B(n_62),
.Y(n_476)
);

INVx5_ASAP7_75t_L g477 ( 
.A(n_423),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_400),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_423),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_397),
.B(n_305),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_423),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_404),
.Y(n_482)
);

AND2x4_ASAP7_75t_L g483 ( 
.A(n_432),
.B(n_417),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_421),
.B(n_308),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_438),
.B(n_399),
.Y(n_485)
);

BUFx10_ASAP7_75t_L g486 ( 
.A(n_441),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_413),
.Y(n_487)
);

AO22x2_ASAP7_75t_L g488 ( 
.A1(n_417),
.A2(n_4),
.B1(n_2),
.B2(n_3),
.Y(n_488)
);

AND2x6_ASAP7_75t_L g489 ( 
.A(n_438),
.B(n_63),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_413),
.Y(n_490)
);

BUFx2_ASAP7_75t_L g491 ( 
.A(n_395),
.Y(n_491)
);

AND2x6_ASAP7_75t_L g492 ( 
.A(n_438),
.B(n_64),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_400),
.Y(n_493)
);

AND2x4_ASAP7_75t_L g494 ( 
.A(n_417),
.B(n_4),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_412),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_SL g496 ( 
.A(n_429),
.B(n_310),
.Y(n_496)
);

INVx5_ASAP7_75t_L g497 ( 
.A(n_423),
.Y(n_497)
);

INVx2_ASAP7_75t_SL g498 ( 
.A(n_438),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_415),
.Y(n_499)
);

INVx1_ASAP7_75t_SL g500 ( 
.A(n_434),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_421),
.B(n_315),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_419),
.B(n_345),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_424),
.Y(n_503)
);

AND2x6_ASAP7_75t_L g504 ( 
.A(n_438),
.B(n_65),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_432),
.B(n_316),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_425),
.Y(n_506)
);

OR2x2_ASAP7_75t_L g507 ( 
.A(n_433),
.B(n_5),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_395),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_425),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_420),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_418),
.B(n_318),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_496),
.B(n_433),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_483),
.B(n_435),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_502),
.B(n_469),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_502),
.B(n_409),
.Y(n_515)
);

BUFx6f_ASAP7_75t_SL g516 ( 
.A(n_461),
.Y(n_516)
);

INVx2_ASAP7_75t_SL g517 ( 
.A(n_455),
.Y(n_517)
);

O2A1O1Ixp5_ASAP7_75t_L g518 ( 
.A1(n_485),
.A2(n_505),
.B(n_465),
.C(n_468),
.Y(n_518)
);

NAND3xp33_ASAP7_75t_SL g519 ( 
.A(n_508),
.B(n_398),
.C(n_396),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_456),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_483),
.B(n_503),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_451),
.A2(n_426),
.B(n_401),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_485),
.B(n_406),
.Y(n_523)
);

BUFx3_ASAP7_75t_L g524 ( 
.A(n_482),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_453),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_L g526 ( 
.A1(n_488),
.A2(n_418),
.B1(n_426),
.B2(n_398),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_444),
.B(n_418),
.Y(n_527)
);

AOI21xp5_ASAP7_75t_L g528 ( 
.A1(n_458),
.A2(n_414),
.B(n_325),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_510),
.B(n_459),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_505),
.A2(n_335),
.B(n_323),
.Y(n_530)
);

NAND2xp33_ASAP7_75t_L g531 ( 
.A(n_482),
.B(n_411),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_464),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_446),
.B(n_396),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_510),
.B(n_440),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_454),
.B(n_336),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_L g536 ( 
.A1(n_488),
.A2(n_405),
.B1(n_416),
.B2(n_402),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_473),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_452),
.A2(n_405),
.B1(n_416),
.B2(n_402),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_462),
.B(n_338),
.Y(n_539)
);

NAND2x1_ASAP7_75t_L g540 ( 
.A(n_466),
.B(n_66),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_498),
.B(n_339),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_495),
.B(n_341),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_499),
.B(n_5),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_446),
.B(n_6),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_478),
.Y(n_545)
);

AND2x2_ASAP7_75t_SL g546 ( 
.A(n_494),
.B(n_449),
.Y(n_546)
);

OAI221xp5_ASAP7_75t_L g547 ( 
.A1(n_507),
.A2(n_439),
.B1(n_437),
.B2(n_434),
.C(n_9),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_493),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_494),
.B(n_437),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_486),
.B(n_6),
.Y(n_550)
);

A2O1A1Ixp33_ASAP7_75t_L g551 ( 
.A1(n_494),
.A2(n_439),
.B(n_9),
.C(n_7),
.Y(n_551)
);

BUFx2_ASAP7_75t_L g552 ( 
.A(n_460),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_453),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_480),
.B(n_7),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_506),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_486),
.B(n_8),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_491),
.B(n_8),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_488),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_463),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_463),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_508),
.B(n_10),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_484),
.B(n_11),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_506),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_501),
.B(n_12),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_452),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_447),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_448),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_445),
.B(n_13),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_448),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_466),
.A2(n_16),
.B1(n_14),
.B2(n_15),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_445),
.B(n_16),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_447),
.B(n_17),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_466),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_573)
);

OAI221xp5_ASAP7_75t_L g574 ( 
.A1(n_461),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.C(n_21),
.Y(n_574)
);

AOI22xp33_ASAP7_75t_L g575 ( 
.A1(n_466),
.A2(n_475),
.B1(n_487),
.B2(n_471),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_470),
.B(n_22),
.Y(n_576)
);

INVxp67_ASAP7_75t_L g577 ( 
.A(n_500),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_511),
.B(n_22),
.Y(n_578)
);

AOI21xp5_ASAP7_75t_L g579 ( 
.A1(n_465),
.A2(n_68),
.B(n_67),
.Y(n_579)
);

INVx1_ASAP7_75t_SL g580 ( 
.A(n_457),
.Y(n_580)
);

A2O1A1Ixp33_ASAP7_75t_SL g581 ( 
.A1(n_470),
.A2(n_26),
.B(n_23),
.C(n_24),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_472),
.B(n_27),
.Y(n_582)
);

AND3x1_ASAP7_75t_L g583 ( 
.A(n_474),
.B(n_27),
.C(n_28),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_472),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_466),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_585)
);

OAI22x1_ASAP7_75t_L g586 ( 
.A1(n_460),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_586)
);

AND2x4_ASAP7_75t_L g587 ( 
.A(n_524),
.B(n_450),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_520),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_514),
.B(n_506),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_515),
.B(n_461),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_R g591 ( 
.A(n_519),
.B(n_506),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_527),
.B(n_479),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_532),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_525),
.Y(n_594)
);

AND2x4_ASAP7_75t_L g595 ( 
.A(n_513),
.B(n_467),
.Y(n_595)
);

INVx4_ASAP7_75t_L g596 ( 
.A(n_555),
.Y(n_596)
);

INVx6_ASAP7_75t_L g597 ( 
.A(n_546),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_527),
.B(n_479),
.Y(n_598)
);

NAND3xp33_ASAP7_75t_L g599 ( 
.A(n_536),
.B(n_481),
.C(n_479),
.Y(n_599)
);

AOI22xp33_ASAP7_75t_L g600 ( 
.A1(n_558),
.A2(n_471),
.B1(n_487),
.B2(n_475),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_546),
.A2(n_481),
.B1(n_479),
.B2(n_509),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_529),
.B(n_490),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_521),
.B(n_537),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_534),
.B(n_490),
.Y(n_604)
);

INVx5_ASAP7_75t_L g605 ( 
.A(n_555),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_512),
.B(n_481),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_533),
.B(n_481),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_533),
.B(n_509),
.Y(n_608)
);

CKINVDCx20_ASAP7_75t_R g609 ( 
.A(n_552),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_544),
.B(n_467),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_580),
.B(n_468),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_545),
.Y(n_612)
);

AND2x4_ASAP7_75t_SL g613 ( 
.A(n_517),
.B(n_476),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_548),
.Y(n_614)
);

INVx4_ASAP7_75t_L g615 ( 
.A(n_555),
.Y(n_615)
);

NOR3xp33_ASAP7_75t_SL g616 ( 
.A(n_574),
.B(n_31),
.C(n_32),
.Y(n_616)
);

OR2x2_ASAP7_75t_SL g617 ( 
.A(n_536),
.B(n_476),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_553),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_544),
.B(n_467),
.Y(n_619)
);

AND3x1_ASAP7_75t_SL g620 ( 
.A(n_547),
.B(n_32),
.C(n_33),
.Y(n_620)
);

AND2x4_ASAP7_75t_L g621 ( 
.A(n_549),
.B(n_467),
.Y(n_621)
);

BUFx2_ASAP7_75t_L g622 ( 
.A(n_577),
.Y(n_622)
);

INVx1_ASAP7_75t_SL g623 ( 
.A(n_561),
.Y(n_623)
);

NAND3xp33_ASAP7_75t_SL g624 ( 
.A(n_538),
.B(n_489),
.C(n_476),
.Y(n_624)
);

BUFx2_ASAP7_75t_L g625 ( 
.A(n_557),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_516),
.Y(n_626)
);

HB1xp67_ASAP7_75t_L g627 ( 
.A(n_572),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_559),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_555),
.Y(n_629)
);

NOR3xp33_ASAP7_75t_SL g630 ( 
.A(n_550),
.B(n_556),
.C(n_551),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_563),
.B(n_575),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_566),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_560),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_550),
.B(n_556),
.Y(n_634)
);

BUFx2_ASAP7_75t_L g635 ( 
.A(n_554),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_531),
.B(n_477),
.Y(n_636)
);

NAND3xp33_ASAP7_75t_SL g637 ( 
.A(n_573),
.B(n_489),
.C(n_476),
.Y(n_637)
);

AO22x1_ASAP7_75t_L g638 ( 
.A1(n_558),
.A2(n_489),
.B1(n_492),
.B2(n_476),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_543),
.Y(n_639)
);

AOI22xp5_ASAP7_75t_L g640 ( 
.A1(n_526),
.A2(n_492),
.B1(n_489),
.B2(n_504),
.Y(n_640)
);

OR2x2_ASAP7_75t_L g641 ( 
.A(n_542),
.B(n_33),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_516),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_567),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g644 ( 
.A(n_566),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_523),
.B(n_477),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_563),
.Y(n_646)
);

NAND2xp33_ASAP7_75t_R g647 ( 
.A(n_523),
.B(n_489),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_528),
.B(n_477),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_564),
.B(n_477),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_584),
.Y(n_650)
);

OR2x4_ASAP7_75t_L g651 ( 
.A(n_572),
.B(n_34),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_578),
.Y(n_652)
);

AOI21xp5_ASAP7_75t_L g653 ( 
.A1(n_589),
.A2(n_563),
.B(n_522),
.Y(n_653)
);

OAI21x1_ASAP7_75t_L g654 ( 
.A1(n_589),
.A2(n_518),
.B(n_540),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_590),
.B(n_634),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_590),
.B(n_526),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_SL g657 ( 
.A1(n_637),
.A2(n_631),
.B(n_563),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_SL g658 ( 
.A1(n_631),
.A2(n_571),
.B(n_568),
.Y(n_658)
);

AOI21xp5_ASAP7_75t_L g659 ( 
.A1(n_608),
.A2(n_575),
.B(n_576),
.Y(n_659)
);

AO31x2_ASAP7_75t_L g660 ( 
.A1(n_604),
.A2(n_608),
.A3(n_645),
.B(n_602),
.Y(n_660)
);

BUFx2_ASAP7_75t_SL g661 ( 
.A(n_609),
.Y(n_661)
);

INVx8_ASAP7_75t_L g662 ( 
.A(n_626),
.Y(n_662)
);

OAI21x1_ASAP7_75t_L g663 ( 
.A1(n_646),
.A2(n_579),
.B(n_582),
.Y(n_663)
);

HB1xp67_ASAP7_75t_L g664 ( 
.A(n_622),
.Y(n_664)
);

OAI21x1_ASAP7_75t_L g665 ( 
.A1(n_648),
.A2(n_562),
.B(n_569),
.Y(n_665)
);

OAI21x1_ASAP7_75t_L g666 ( 
.A1(n_640),
.A2(n_570),
.B(n_573),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_627),
.B(n_535),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_603),
.B(n_585),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_644),
.Y(n_669)
);

OAI21x1_ASAP7_75t_L g670 ( 
.A1(n_649),
.A2(n_585),
.B(n_541),
.Y(n_670)
);

AOI21x1_ASAP7_75t_L g671 ( 
.A1(n_610),
.A2(n_539),
.B(n_530),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_627),
.B(n_586),
.Y(n_672)
);

OAI21xp33_ASAP7_75t_L g673 ( 
.A1(n_630),
.A2(n_565),
.B(n_583),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_623),
.B(n_34),
.Y(n_674)
);

AOI21x1_ASAP7_75t_L g675 ( 
.A1(n_619),
.A2(n_581),
.B(n_497),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_594),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_628),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_605),
.B(n_497),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_625),
.B(n_35),
.Y(n_679)
);

OAI21x1_ASAP7_75t_L g680 ( 
.A1(n_646),
.A2(n_504),
.B(n_492),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_611),
.B(n_497),
.Y(n_681)
);

BUFx3_ASAP7_75t_L g682 ( 
.A(n_587),
.Y(n_682)
);

BUFx2_ASAP7_75t_L g683 ( 
.A(n_642),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_639),
.B(n_497),
.Y(n_684)
);

INVx3_ASAP7_75t_L g685 ( 
.A(n_644),
.Y(n_685)
);

NOR2x1_ASAP7_75t_SL g686 ( 
.A(n_605),
.B(n_492),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_588),
.Y(n_687)
);

INVx5_ASAP7_75t_L g688 ( 
.A(n_597),
.Y(n_688)
);

OAI21x1_ASAP7_75t_L g689 ( 
.A1(n_624),
.A2(n_504),
.B(n_492),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_L g690 ( 
.A1(n_607),
.A2(n_605),
.B(n_598),
.Y(n_690)
);

OAI21x1_ASAP7_75t_L g691 ( 
.A1(n_606),
.A2(n_504),
.B(n_71),
.Y(n_691)
);

NOR2x1_ASAP7_75t_SL g692 ( 
.A(n_605),
.B(n_504),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_635),
.B(n_36),
.Y(n_693)
);

AOI21xp5_ASAP7_75t_L g694 ( 
.A1(n_592),
.A2(n_598),
.B(n_629),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_633),
.Y(n_695)
);

AOI21xp5_ASAP7_75t_L g696 ( 
.A1(n_592),
.A2(n_72),
.B(n_69),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_593),
.Y(n_697)
);

AOI21xp5_ASAP7_75t_L g698 ( 
.A1(n_629),
.A2(n_75),
.B(n_74),
.Y(n_698)
);

AOI21x1_ASAP7_75t_SL g699 ( 
.A1(n_636),
.A2(n_621),
.B(n_587),
.Y(n_699)
);

AOI21x1_ASAP7_75t_L g700 ( 
.A1(n_638),
.A2(n_77),
.B(n_76),
.Y(n_700)
);

OR2x2_ASAP7_75t_L g701 ( 
.A(n_612),
.B(n_36),
.Y(n_701)
);

OAI21x1_ASAP7_75t_L g702 ( 
.A1(n_601),
.A2(n_79),
.B(n_78),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_629),
.B(n_591),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_618),
.Y(n_704)
);

AOI21xp5_ASAP7_75t_L g705 ( 
.A1(n_629),
.A2(n_81),
.B(n_80),
.Y(n_705)
);

AOI21xp5_ASAP7_75t_L g706 ( 
.A1(n_596),
.A2(n_84),
.B(n_82),
.Y(n_706)
);

INVx3_ASAP7_75t_SL g707 ( 
.A(n_652),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_614),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_597),
.B(n_37),
.Y(n_709)
);

NOR2x1_ASAP7_75t_SL g710 ( 
.A(n_596),
.B(n_278),
.Y(n_710)
);

AOI211x1_ASAP7_75t_L g711 ( 
.A1(n_643),
.A2(n_37),
.B(n_38),
.C(n_39),
.Y(n_711)
);

AOI21xp33_ASAP7_75t_L g712 ( 
.A1(n_599),
.A2(n_38),
.B(n_39),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_R g713 ( 
.A(n_647),
.B(n_276),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_597),
.B(n_40),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_650),
.Y(n_715)
);

BUFx6f_ASAP7_75t_L g716 ( 
.A(n_615),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_641),
.Y(n_717)
);

NOR2xp67_ASAP7_75t_L g718 ( 
.A(n_664),
.B(n_688),
.Y(n_718)
);

NOR2xp67_ASAP7_75t_L g719 ( 
.A(n_664),
.B(n_632),
.Y(n_719)
);

OAI21x1_ASAP7_75t_L g720 ( 
.A1(n_653),
.A2(n_632),
.B(n_600),
.Y(n_720)
);

OAI21x1_ASAP7_75t_L g721 ( 
.A1(n_663),
.A2(n_600),
.B(n_647),
.Y(n_721)
);

HB1xp67_ASAP7_75t_L g722 ( 
.A(n_714),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_661),
.Y(n_723)
);

OAI21xp5_ASAP7_75t_L g724 ( 
.A1(n_655),
.A2(n_630),
.B(n_616),
.Y(n_724)
);

OAI22xp5_ASAP7_75t_L g725 ( 
.A1(n_655),
.A2(n_617),
.B1(n_651),
.B2(n_616),
.Y(n_725)
);

OAI21x1_ASAP7_75t_L g726 ( 
.A1(n_654),
.A2(n_615),
.B(n_613),
.Y(n_726)
);

AOI22xp33_ASAP7_75t_L g727 ( 
.A1(n_673),
.A2(n_621),
.B1(n_595),
.B2(n_591),
.Y(n_727)
);

OR2x2_ASAP7_75t_L g728 ( 
.A(n_682),
.B(n_595),
.Y(n_728)
);

A2O1A1Ixp33_ASAP7_75t_L g729 ( 
.A1(n_666),
.A2(n_620),
.B(n_651),
.C(n_42),
.Y(n_729)
);

AND2x4_ASAP7_75t_L g730 ( 
.A(n_688),
.B(n_85),
.Y(n_730)
);

HB1xp67_ASAP7_75t_L g731 ( 
.A(n_709),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_676),
.Y(n_732)
);

OAI21x1_ASAP7_75t_L g733 ( 
.A1(n_702),
.A2(n_620),
.B(n_87),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_688),
.Y(n_734)
);

OAI22xp5_ASAP7_75t_L g735 ( 
.A1(n_667),
.A2(n_40),
.B1(n_41),
.B2(n_43),
.Y(n_735)
);

BUFx3_ASAP7_75t_L g736 ( 
.A(n_682),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_679),
.B(n_41),
.Y(n_737)
);

INVx2_ASAP7_75t_L g738 ( 
.A(n_676),
.Y(n_738)
);

AND2x4_ASAP7_75t_L g739 ( 
.A(n_688),
.B(n_86),
.Y(n_739)
);

INVx3_ASAP7_75t_L g740 ( 
.A(n_716),
.Y(n_740)
);

INVx2_ASAP7_75t_SL g741 ( 
.A(n_662),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_687),
.Y(n_742)
);

AO21x2_ASAP7_75t_L g743 ( 
.A1(n_658),
.A2(n_91),
.B(n_90),
.Y(n_743)
);

AOI22x1_ASAP7_75t_L g744 ( 
.A1(n_659),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_744)
);

AOI222xp33_ASAP7_75t_L g745 ( 
.A1(n_672),
.A2(n_668),
.B1(n_656),
.B2(n_717),
.C1(n_674),
.C2(n_697),
.Y(n_745)
);

AOI221xp5_ASAP7_75t_L g746 ( 
.A1(n_693),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.C(n_48),
.Y(n_746)
);

AOI22xp5_ASAP7_75t_L g747 ( 
.A1(n_667),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_708),
.Y(n_748)
);

OAI21x1_ASAP7_75t_SL g749 ( 
.A1(n_686),
.A2(n_49),
.B(n_50),
.Y(n_749)
);

OR2x2_ASAP7_75t_L g750 ( 
.A(n_701),
.B(n_51),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_707),
.B(n_51),
.Y(n_751)
);

OAI21x1_ASAP7_75t_SL g752 ( 
.A1(n_692),
.A2(n_52),
.B(n_53),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_677),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_677),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_704),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_704),
.Y(n_756)
);

AO21x2_ASAP7_75t_L g757 ( 
.A1(n_671),
.A2(n_675),
.B(n_657),
.Y(n_757)
);

INVx3_ASAP7_75t_L g758 ( 
.A(n_716),
.Y(n_758)
);

OAI21x1_ASAP7_75t_L g759 ( 
.A1(n_702),
.A2(n_94),
.B(n_93),
.Y(n_759)
);

BUFx12f_ASAP7_75t_L g760 ( 
.A(n_683),
.Y(n_760)
);

OAI21x1_ASAP7_75t_L g761 ( 
.A1(n_691),
.A2(n_96),
.B(n_95),
.Y(n_761)
);

INVx3_ASAP7_75t_L g762 ( 
.A(n_716),
.Y(n_762)
);

O2A1O1Ixp33_ASAP7_75t_SL g763 ( 
.A1(n_703),
.A2(n_52),
.B(n_53),
.C(n_54),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_707),
.B(n_54),
.Y(n_764)
);

OAI21x1_ASAP7_75t_L g765 ( 
.A1(n_691),
.A2(n_98),
.B(n_97),
.Y(n_765)
);

OAI22xp5_ASAP7_75t_L g766 ( 
.A1(n_684),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_766)
);

OAI21x1_ASAP7_75t_L g767 ( 
.A1(n_689),
.A2(n_100),
.B(n_99),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_715),
.B(n_669),
.Y(n_768)
);

OAI22xp5_ASAP7_75t_L g769 ( 
.A1(n_684),
.A2(n_58),
.B1(n_60),
.B2(n_101),
.Y(n_769)
);

NAND2x1p5_ASAP7_75t_L g770 ( 
.A(n_703),
.B(n_103),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_L g771 ( 
.A1(n_666),
.A2(n_58),
.B1(n_60),
.B2(n_104),
.Y(n_771)
);

OAI21x1_ASAP7_75t_L g772 ( 
.A1(n_689),
.A2(n_105),
.B(n_106),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_662),
.A2(n_107),
.B1(n_108),
.B2(n_109),
.Y(n_773)
);

OAI21x1_ASAP7_75t_L g774 ( 
.A1(n_665),
.A2(n_110),
.B(n_112),
.Y(n_774)
);

OR2x6_ASAP7_75t_L g775 ( 
.A(n_694),
.B(n_113),
.Y(n_775)
);

BUFx6f_ASAP7_75t_SL g776 ( 
.A(n_716),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_695),
.Y(n_777)
);

OAI22xp33_ASAP7_75t_L g778 ( 
.A1(n_725),
.A2(n_712),
.B1(n_681),
.B2(n_662),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_745),
.A2(n_695),
.B1(n_713),
.B2(n_696),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_737),
.B(n_669),
.Y(n_780)
);

INVx4_ASAP7_75t_L g781 ( 
.A(n_734),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_SL g782 ( 
.A1(n_724),
.A2(n_713),
.B1(n_710),
.B2(n_680),
.Y(n_782)
);

OAI21x1_ASAP7_75t_L g783 ( 
.A1(n_774),
.A2(n_700),
.B(n_665),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_729),
.B(n_685),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_722),
.B(n_685),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_727),
.A2(n_690),
.B1(n_678),
.B2(n_680),
.Y(n_786)
);

OAI22xp5_ASAP7_75t_L g787 ( 
.A1(n_729),
.A2(n_711),
.B1(n_678),
.B2(n_706),
.Y(n_787)
);

BUFx6f_ASAP7_75t_L g788 ( 
.A(n_734),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_742),
.B(n_660),
.Y(n_789)
);

AOI222xp33_ASAP7_75t_L g790 ( 
.A1(n_746),
.A2(n_670),
.B1(n_699),
.B2(n_660),
.C1(n_705),
.C2(n_698),
.Y(n_790)
);

OAI22xp5_ASAP7_75t_L g791 ( 
.A1(n_747),
.A2(n_670),
.B1(n_660),
.B2(n_117),
.Y(n_791)
);

AOI22xp5_ASAP7_75t_L g792 ( 
.A1(n_727),
.A2(n_660),
.B1(n_116),
.B2(n_118),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_732),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_764),
.B(n_114),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_748),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_755),
.Y(n_796)
);

NOR2xp67_ASAP7_75t_L g797 ( 
.A(n_741),
.B(n_120),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_756),
.B(n_275),
.Y(n_798)
);

OAI21x1_ASAP7_75t_L g799 ( 
.A1(n_774),
.A2(n_121),
.B(n_122),
.Y(n_799)
);

HB1xp67_ASAP7_75t_L g800 ( 
.A(n_768),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_735),
.A2(n_123),
.B1(n_125),
.B2(n_127),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_777),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_731),
.B(n_274),
.Y(n_803)
);

INVxp67_ASAP7_75t_L g804 ( 
.A(n_750),
.Y(n_804)
);

AND2x4_ASAP7_75t_L g805 ( 
.A(n_730),
.B(n_739),
.Y(n_805)
);

BUFx3_ASAP7_75t_L g806 ( 
.A(n_736),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_751),
.B(n_128),
.Y(n_807)
);

INVx1_ASAP7_75t_SL g808 ( 
.A(n_723),
.Y(n_808)
);

INVx4_ASAP7_75t_L g809 ( 
.A(n_734),
.Y(n_809)
);

INVx2_ASAP7_75t_SL g810 ( 
.A(n_736),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_730),
.B(n_129),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_732),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_738),
.Y(n_813)
);

NAND2xp33_ASAP7_75t_R g814 ( 
.A(n_775),
.B(n_130),
.Y(n_814)
);

INVx6_ASAP7_75t_L g815 ( 
.A(n_734),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_753),
.Y(n_816)
);

INVx3_ASAP7_75t_L g817 ( 
.A(n_775),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_753),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_719),
.B(n_273),
.Y(n_819)
);

OAI22xp5_ASAP7_75t_L g820 ( 
.A1(n_771),
.A2(n_751),
.B1(n_744),
.B2(n_723),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_754),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_718),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_728),
.B(n_741),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_754),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_757),
.Y(n_825)
);

INVx2_ASAP7_75t_SL g826 ( 
.A(n_760),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_760),
.B(n_740),
.Y(n_827)
);

CKINVDCx6p67_ASAP7_75t_R g828 ( 
.A(n_776),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_740),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_775),
.A2(n_131),
.B(n_132),
.Y(n_830)
);

A2O1A1Ixp33_ASAP7_75t_L g831 ( 
.A1(n_771),
.A2(n_133),
.B(n_134),
.C(n_137),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_740),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_758),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_776),
.Y(n_834)
);

BUFx2_ASAP7_75t_L g835 ( 
.A(n_758),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_757),
.Y(n_836)
);

OAI221xp5_ASAP7_75t_L g837 ( 
.A1(n_766),
.A2(n_272),
.B1(n_141),
.B2(n_142),
.C(n_143),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_720),
.Y(n_838)
);

BUFx2_ASAP7_75t_L g839 ( 
.A(n_758),
.Y(n_839)
);

CKINVDCx20_ASAP7_75t_R g840 ( 
.A(n_762),
.Y(n_840)
);

OAI211xp5_ASAP7_75t_SL g841 ( 
.A1(n_769),
.A2(n_763),
.B(n_773),
.C(n_762),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_762),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_730),
.B(n_138),
.Y(n_843)
);

AND2x4_ASAP7_75t_L g844 ( 
.A(n_739),
.B(n_144),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_800),
.B(n_775),
.Y(n_845)
);

AO31x2_ASAP7_75t_L g846 ( 
.A1(n_791),
.A2(n_743),
.A3(n_721),
.B(n_759),
.Y(n_846)
);

INVxp67_ASAP7_75t_L g847 ( 
.A(n_789),
.Y(n_847)
);

INVx5_ASAP7_75t_SL g848 ( 
.A(n_828),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_795),
.Y(n_849)
);

OAI221xp5_ASAP7_75t_L g850 ( 
.A1(n_820),
.A2(n_763),
.B1(n_770),
.B2(n_733),
.C(n_749),
.Y(n_850)
);

AOI221xp5_ASAP7_75t_L g851 ( 
.A1(n_804),
.A2(n_778),
.B1(n_831),
.B2(n_807),
.C(n_784),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_831),
.A2(n_743),
.B(n_733),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_SL g853 ( 
.A1(n_814),
.A2(n_770),
.B1(n_739),
.B2(n_759),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_780),
.B(n_720),
.Y(n_854)
);

OAI211xp5_ASAP7_75t_L g855 ( 
.A1(n_801),
.A2(n_765),
.B(n_761),
.C(n_752),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_796),
.Y(n_856)
);

AOI222xp33_ASAP7_75t_L g857 ( 
.A1(n_779),
.A2(n_721),
.B1(n_765),
.B2(n_761),
.C1(n_767),
.C2(n_772),
.Y(n_857)
);

AOI21x1_ASAP7_75t_L g858 ( 
.A1(n_830),
.A2(n_772),
.B(n_767),
.Y(n_858)
);

BUFx2_ASAP7_75t_L g859 ( 
.A(n_806),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_L g860 ( 
.A1(n_779),
.A2(n_726),
.B1(n_147),
.B2(n_148),
.Y(n_860)
);

AO22x1_ASAP7_75t_L g861 ( 
.A1(n_811),
.A2(n_726),
.B1(n_149),
.B2(n_151),
.Y(n_861)
);

OAI22xp5_ASAP7_75t_L g862 ( 
.A1(n_801),
.A2(n_146),
.B1(n_152),
.B2(n_158),
.Y(n_862)
);

OAI22xp5_ASAP7_75t_L g863 ( 
.A1(n_784),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_SL g864 ( 
.A1(n_808),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_864)
);

INVx1_ASAP7_75t_SL g865 ( 
.A(n_827),
.Y(n_865)
);

OAI21xp33_ASAP7_75t_L g866 ( 
.A1(n_841),
.A2(n_167),
.B(n_168),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_802),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_812),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_813),
.Y(n_869)
);

HB1xp67_ASAP7_75t_L g870 ( 
.A(n_838),
.Y(n_870)
);

A2O1A1Ixp33_ASAP7_75t_L g871 ( 
.A1(n_792),
.A2(n_170),
.B(n_171),
.C(n_172),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_793),
.Y(n_872)
);

BUFx2_ASAP7_75t_L g873 ( 
.A(n_806),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_810),
.B(n_785),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_793),
.Y(n_875)
);

OAI22xp33_ASAP7_75t_L g876 ( 
.A1(n_814),
.A2(n_173),
.B1(n_175),
.B2(n_177),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_810),
.B(n_178),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_L g878 ( 
.A1(n_805),
.A2(n_179),
.B1(n_180),
.B2(n_181),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_L g879 ( 
.A1(n_805),
.A2(n_185),
.B1(n_186),
.B2(n_188),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_L g880 ( 
.A1(n_805),
.A2(n_190),
.B1(n_192),
.B2(n_193),
.Y(n_880)
);

OAI22xp5_ASAP7_75t_L g881 ( 
.A1(n_837),
.A2(n_782),
.B1(n_811),
.B2(n_844),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_823),
.B(n_195),
.Y(n_882)
);

OAI22xp5_ASAP7_75t_L g883 ( 
.A1(n_811),
.A2(n_196),
.B1(n_197),
.B2(n_198),
.Y(n_883)
);

AOI221xp5_ASAP7_75t_L g884 ( 
.A1(n_787),
.A2(n_794),
.B1(n_803),
.B2(n_844),
.C(n_817),
.Y(n_884)
);

OR2x2_ASAP7_75t_L g885 ( 
.A(n_835),
.B(n_200),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_816),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_817),
.A2(n_844),
.B(n_783),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_817),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_839),
.B(n_204),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_840),
.B(n_205),
.Y(n_890)
);

BUFx2_ASAP7_75t_L g891 ( 
.A(n_840),
.Y(n_891)
);

AOI21x1_ASAP7_75t_L g892 ( 
.A1(n_822),
.A2(n_206),
.B(n_207),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_834),
.Y(n_893)
);

CKINVDCx11_ASAP7_75t_R g894 ( 
.A(n_828),
.Y(n_894)
);

A2O1A1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_797),
.A2(n_208),
.B(n_209),
.C(n_211),
.Y(n_895)
);

AO21x2_ASAP7_75t_L g896 ( 
.A1(n_825),
.A2(n_212),
.B(n_213),
.Y(n_896)
);

AOI222xp33_ASAP7_75t_L g897 ( 
.A1(n_843),
.A2(n_271),
.B1(n_216),
.B2(n_218),
.C1(n_219),
.C2(n_220),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_L g898 ( 
.A1(n_826),
.A2(n_214),
.B1(n_223),
.B2(n_224),
.Y(n_898)
);

AOI211xp5_ASAP7_75t_L g899 ( 
.A1(n_819),
.A2(n_225),
.B(n_226),
.C(n_228),
.Y(n_899)
);

BUFx2_ASAP7_75t_L g900 ( 
.A(n_834),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_842),
.B(n_229),
.Y(n_901)
);

AOI22xp33_ASAP7_75t_L g902 ( 
.A1(n_790),
.A2(n_230),
.B1(n_231),
.B2(n_233),
.Y(n_902)
);

AOI22xp5_ASAP7_75t_SL g903 ( 
.A1(n_788),
.A2(n_234),
.B1(n_236),
.B2(n_237),
.Y(n_903)
);

OR2x6_ASAP7_75t_L g904 ( 
.A(n_825),
.B(n_238),
.Y(n_904)
);

AOI22xp33_ASAP7_75t_L g905 ( 
.A1(n_818),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_905)
);

OR2x2_ASAP7_75t_L g906 ( 
.A(n_847),
.B(n_838),
.Y(n_906)
);

AOI22xp33_ASAP7_75t_L g907 ( 
.A1(n_851),
.A2(n_824),
.B1(n_818),
.B2(n_821),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_856),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_874),
.B(n_833),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_867),
.Y(n_910)
);

NOR2x1_ASAP7_75t_SL g911 ( 
.A(n_904),
.B(n_788),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_854),
.B(n_849),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_859),
.B(n_832),
.Y(n_913)
);

AND2x4_ASAP7_75t_L g914 ( 
.A(n_887),
.B(n_836),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_873),
.B(n_829),
.Y(n_915)
);

INVx2_ASAP7_75t_SL g916 ( 
.A(n_891),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_868),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_845),
.Y(n_918)
);

OAI221xp5_ASAP7_75t_L g919 ( 
.A1(n_884),
.A2(n_786),
.B1(n_798),
.B2(n_815),
.C(n_809),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_904),
.Y(n_920)
);

AND2x4_ASAP7_75t_L g921 ( 
.A(n_870),
.B(n_809),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_869),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_872),
.Y(n_923)
);

AND2x4_ASAP7_75t_L g924 ( 
.A(n_870),
.B(n_809),
.Y(n_924)
);

BUFx2_ASAP7_75t_SL g925 ( 
.A(n_889),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_865),
.B(n_788),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_875),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_853),
.B(n_824),
.Y(n_928)
);

AND2x4_ASAP7_75t_L g929 ( 
.A(n_886),
.B(n_781),
.Y(n_929)
);

AO31x2_ASAP7_75t_L g930 ( 
.A1(n_852),
.A2(n_821),
.A3(n_781),
.B(n_783),
.Y(n_930)
);

INVx2_ASAP7_75t_SL g931 ( 
.A(n_900),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_853),
.B(n_781),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_846),
.B(n_788),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_882),
.B(n_890),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_846),
.B(n_799),
.Y(n_935)
);

INVx2_ASAP7_75t_L g936 ( 
.A(n_846),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_846),
.Y(n_937)
);

BUFx3_ASAP7_75t_L g938 ( 
.A(n_894),
.Y(n_938)
);

INVx2_ASAP7_75t_SL g939 ( 
.A(n_885),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_904),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_896),
.Y(n_941)
);

INVx2_ASAP7_75t_SL g942 ( 
.A(n_877),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_848),
.B(n_815),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_896),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_848),
.B(n_815),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_858),
.Y(n_946)
);

OAI22xp33_ASAP7_75t_L g947 ( 
.A1(n_881),
.A2(n_799),
.B1(n_244),
.B2(n_245),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_892),
.Y(n_948)
);

OR2x6_ASAP7_75t_L g949 ( 
.A(n_861),
.B(n_243),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_902),
.B(n_246),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_850),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_848),
.B(n_270),
.Y(n_952)
);

AND2x4_ASAP7_75t_SL g953 ( 
.A(n_901),
.B(n_248),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_883),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_855),
.Y(n_955)
);

HB1xp67_ASAP7_75t_L g956 ( 
.A(n_857),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_902),
.B(n_250),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_860),
.B(n_251),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_912),
.B(n_860),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_917),
.Y(n_960)
);

AOI221xp5_ASAP7_75t_L g961 ( 
.A1(n_956),
.A2(n_876),
.B1(n_866),
.B2(n_864),
.C(n_862),
.Y(n_961)
);

HB1xp67_ASAP7_75t_L g962 ( 
.A(n_912),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_927),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_933),
.B(n_893),
.Y(n_964)
);

HB1xp67_ASAP7_75t_L g965 ( 
.A(n_918),
.Y(n_965)
);

NAND3xp33_ASAP7_75t_L g966 ( 
.A(n_955),
.B(n_897),
.C(n_880),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_933),
.B(n_880),
.Y(n_967)
);

OAI321xp33_ASAP7_75t_L g968 ( 
.A1(n_955),
.A2(n_876),
.A3(n_878),
.B1(n_879),
.B2(n_863),
.C(n_888),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_917),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_939),
.B(n_942),
.Y(n_970)
);

AOI22xp5_ASAP7_75t_L g971 ( 
.A1(n_950),
.A2(n_957),
.B1(n_949),
.B2(n_951),
.Y(n_971)
);

NAND3xp33_ASAP7_75t_L g972 ( 
.A(n_951),
.B(n_878),
.C(n_879),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_939),
.B(n_899),
.Y(n_973)
);

INVx2_ASAP7_75t_SL g974 ( 
.A(n_916),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_922),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_932),
.B(n_903),
.Y(n_976)
);

OR2x2_ASAP7_75t_L g977 ( 
.A(n_909),
.B(n_888),
.Y(n_977)
);

NOR2x1_ASAP7_75t_L g978 ( 
.A(n_925),
.B(n_871),
.Y(n_978)
);

AOI221xp5_ASAP7_75t_L g979 ( 
.A1(n_935),
.A2(n_898),
.B1(n_905),
.B2(n_895),
.C(n_256),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_921),
.B(n_905),
.Y(n_980)
);

INVx2_ASAP7_75t_SL g981 ( 
.A(n_916),
.Y(n_981)
);

AO21x2_ASAP7_75t_L g982 ( 
.A1(n_936),
.A2(n_252),
.B(n_253),
.Y(n_982)
);

OAI21x1_ASAP7_75t_L g983 ( 
.A1(n_946),
.A2(n_255),
.B(n_257),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_921),
.B(n_258),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_927),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_922),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_908),
.Y(n_987)
);

OAI221xp5_ASAP7_75t_L g988 ( 
.A1(n_949),
.A2(n_259),
.B1(n_260),
.B2(n_262),
.C(n_263),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_946),
.Y(n_989)
);

OAI211xp5_ASAP7_75t_L g990 ( 
.A1(n_950),
.A2(n_264),
.B(n_265),
.C(n_267),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_936),
.Y(n_991)
);

HB1xp67_ASAP7_75t_L g992 ( 
.A(n_965),
.Y(n_992)
);

AO21x1_ASAP7_75t_L g993 ( 
.A1(n_971),
.A2(n_935),
.B(n_957),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_960),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_960),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_991),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_991),
.Y(n_997)
);

AND2x2_ASAP7_75t_L g998 ( 
.A(n_962),
.B(n_931),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_969),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_969),
.B(n_910),
.Y(n_1000)
);

OR2x2_ASAP7_75t_L g1001 ( 
.A(n_974),
.B(n_908),
.Y(n_1001)
);

HB1xp67_ASAP7_75t_L g1002 ( 
.A(n_975),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_964),
.B(n_931),
.Y(n_1003)
);

INVx1_ASAP7_75t_SL g1004 ( 
.A(n_964),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_975),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_974),
.B(n_938),
.Y(n_1006)
);

INVx3_ASAP7_75t_L g1007 ( 
.A(n_989),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_991),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_989),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_986),
.B(n_987),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_986),
.B(n_910),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_987),
.B(n_915),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_981),
.B(n_915),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_989),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_981),
.B(n_970),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_959),
.B(n_913),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_996),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_992),
.B(n_959),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_994),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_1016),
.B(n_977),
.Y(n_1020)
);

INVx2_ASAP7_75t_SL g1021 ( 
.A(n_1001),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_993),
.A2(n_978),
.B(n_968),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_996),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_1004),
.B(n_925),
.Y(n_1024)
);

AOI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_993),
.A2(n_971),
.B1(n_966),
.B2(n_961),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_1012),
.B(n_1002),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_1001),
.B(n_977),
.Y(n_1027)
);

AOI22xp33_ASAP7_75t_L g1028 ( 
.A1(n_1006),
.A2(n_966),
.B1(n_972),
.B2(n_967),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_996),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_994),
.Y(n_1030)
);

INVx2_ASAP7_75t_SL g1031 ( 
.A(n_1015),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_995),
.Y(n_1032)
);

CKINVDCx8_ASAP7_75t_R g1033 ( 
.A(n_1022),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_1017),
.Y(n_1034)
);

OR2x2_ASAP7_75t_L g1035 ( 
.A(n_1027),
.B(n_1010),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_1019),
.Y(n_1036)
);

AND2x4_ASAP7_75t_L g1037 ( 
.A(n_1031),
.B(n_1015),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_1031),
.B(n_1021),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_1021),
.B(n_998),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_1030),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_1024),
.B(n_998),
.Y(n_1041)
);

INVxp67_ASAP7_75t_SL g1042 ( 
.A(n_1025),
.Y(n_1042)
);

AND2x2_ASAP7_75t_L g1043 ( 
.A(n_1018),
.B(n_1003),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_1032),
.Y(n_1044)
);

OAI22xp33_ASAP7_75t_L g1045 ( 
.A1(n_1033),
.A2(n_1042),
.B1(n_972),
.B2(n_973),
.Y(n_1045)
);

O2A1O1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_1033),
.A2(n_1028),
.B(n_988),
.C(n_990),
.Y(n_1046)
);

AOI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_1037),
.A2(n_1028),
.B1(n_976),
.B2(n_967),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_1043),
.B(n_1020),
.Y(n_1048)
);

INVxp33_ASAP7_75t_L g1049 ( 
.A(n_1037),
.Y(n_1049)
);

OAI32xp33_ASAP7_75t_L g1050 ( 
.A1(n_1038),
.A2(n_1026),
.A3(n_1007),
.B1(n_938),
.B2(n_1009),
.Y(n_1050)
);

OR2x2_ASAP7_75t_L g1051 ( 
.A(n_1035),
.B(n_1000),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_1040),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_1040),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1052),
.Y(n_1054)
);

INVx2_ASAP7_75t_SL g1055 ( 
.A(n_1053),
.Y(n_1055)
);

OAI32xp33_ASAP7_75t_L g1056 ( 
.A1(n_1049),
.A2(n_1038),
.A3(n_1035),
.B1(n_1039),
.B2(n_1036),
.Y(n_1056)
);

NAND2x1_ASAP7_75t_SL g1057 ( 
.A(n_1047),
.B(n_1037),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_1051),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1055),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1055),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1058),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1058),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_1054),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_1059),
.B(n_1043),
.Y(n_1064)
);

O2A1O1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_1061),
.A2(n_1045),
.B(n_1046),
.C(n_1056),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_SL g1066 ( 
.A(n_1062),
.B(n_978),
.Y(n_1066)
);

NOR3xp33_ASAP7_75t_L g1067 ( 
.A(n_1060),
.B(n_1050),
.C(n_1048),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1063),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1061),
.Y(n_1069)
);

NOR2x1_ASAP7_75t_R g1070 ( 
.A(n_1059),
.B(n_1057),
.Y(n_1070)
);

AOI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_1066),
.A2(n_1034),
.B1(n_979),
.B2(n_976),
.Y(n_1071)
);

OAI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_1065),
.A2(n_1044),
.B1(n_1039),
.B2(n_1041),
.Y(n_1072)
);

OAI22xp33_ASAP7_75t_L g1073 ( 
.A1(n_1069),
.A2(n_949),
.B1(n_1034),
.B2(n_934),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_1065),
.B(n_1041),
.Y(n_1074)
);

NOR4xp25_ASAP7_75t_L g1075 ( 
.A(n_1068),
.B(n_952),
.C(n_958),
.D(n_947),
.Y(n_1075)
);

AOI22xp33_ASAP7_75t_L g1076 ( 
.A1(n_1067),
.A2(n_949),
.B1(n_976),
.B2(n_937),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_1074),
.B(n_1070),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1072),
.Y(n_1078)
);

OA22x2_ASAP7_75t_L g1079 ( 
.A1(n_1071),
.A2(n_1064),
.B1(n_1003),
.B2(n_976),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_1075),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_1076),
.B(n_1009),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1073),
.Y(n_1082)
);

OAI322xp33_ASAP7_75t_L g1083 ( 
.A1(n_1074),
.A2(n_954),
.A3(n_948),
.B1(n_1009),
.B2(n_1014),
.C1(n_1011),
.C2(n_1005),
.Y(n_1083)
);

AND2x4_ASAP7_75t_L g1084 ( 
.A(n_1077),
.B(n_1007),
.Y(n_1084)
);

OAI221xp5_ASAP7_75t_L g1085 ( 
.A1(n_1080),
.A2(n_949),
.B1(n_948),
.B2(n_1017),
.C(n_1029),
.Y(n_1085)
);

OR2x2_ASAP7_75t_L g1086 ( 
.A(n_1078),
.B(n_1005),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_1079),
.B(n_1023),
.Y(n_1087)
);

AOI322xp5_ASAP7_75t_L g1088 ( 
.A1(n_1082),
.A2(n_1081),
.A3(n_1083),
.B1(n_907),
.B2(n_1023),
.C1(n_1029),
.C2(n_940),
.Y(n_1088)
);

NOR3xp33_ASAP7_75t_L g1089 ( 
.A(n_1080),
.B(n_983),
.C(n_919),
.Y(n_1089)
);

AOI211x1_ASAP7_75t_L g1090 ( 
.A1(n_1078),
.A2(n_1013),
.B(n_995),
.C(n_999),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1080),
.B(n_1007),
.Y(n_1091)
);

OAI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_1077),
.A2(n_984),
.B(n_1014),
.Y(n_1092)
);

NOR3xp33_ASAP7_75t_L g1093 ( 
.A(n_1080),
.B(n_983),
.C(n_943),
.Y(n_1093)
);

BUFx2_ASAP7_75t_L g1094 ( 
.A(n_1078),
.Y(n_1094)
);

NOR2x1_ASAP7_75t_L g1095 ( 
.A(n_1094),
.B(n_1007),
.Y(n_1095)
);

AOI22xp5_ASAP7_75t_L g1096 ( 
.A1(n_1087),
.A2(n_1089),
.B1(n_1093),
.B2(n_1085),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_1090),
.B(n_999),
.Y(n_1097)
);

INVx2_ASAP7_75t_SL g1098 ( 
.A(n_1086),
.Y(n_1098)
);

NOR3xp33_ASAP7_75t_SL g1099 ( 
.A(n_1091),
.B(n_945),
.C(n_926),
.Y(n_1099)
);

NOR3xp33_ASAP7_75t_L g1100 ( 
.A(n_1092),
.B(n_984),
.C(n_940),
.Y(n_1100)
);

NOR3xp33_ASAP7_75t_SL g1101 ( 
.A(n_1084),
.B(n_953),
.C(n_941),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_1084),
.A2(n_954),
.B(n_953),
.Y(n_1102)
);

OAI221xp5_ASAP7_75t_L g1103 ( 
.A1(n_1088),
.A2(n_989),
.B1(n_942),
.B2(n_937),
.C(n_920),
.Y(n_1103)
);

AOI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_1087),
.A2(n_982),
.B1(n_980),
.B2(n_920),
.Y(n_1104)
);

OAI22xp33_ASAP7_75t_L g1105 ( 
.A1(n_1094),
.A2(n_920),
.B1(n_1008),
.B2(n_997),
.Y(n_1105)
);

OA22x2_ASAP7_75t_L g1106 ( 
.A1(n_1094),
.A2(n_980),
.B1(n_932),
.B2(n_1008),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_1094),
.B(n_1008),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_1098),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_1103),
.A2(n_982),
.B1(n_941),
.B2(n_920),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_1096),
.Y(n_1110)
);

NOR4xp25_ASAP7_75t_L g1111 ( 
.A(n_1107),
.B(n_997),
.C(n_923),
.D(n_963),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_1101),
.Y(n_1112)
);

NOR2x1_ASAP7_75t_L g1113 ( 
.A(n_1095),
.B(n_982),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1106),
.Y(n_1114)
);

NOR2xp67_ASAP7_75t_L g1115 ( 
.A(n_1097),
.B(n_268),
.Y(n_1115)
);

CKINVDCx20_ASAP7_75t_R g1116 ( 
.A(n_1099),
.Y(n_1116)
);

CKINVDCx20_ASAP7_75t_R g1117 ( 
.A(n_1104),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_1102),
.Y(n_1118)
);

OAI22x1_ASAP7_75t_L g1119 ( 
.A1(n_1108),
.A2(n_1100),
.B1(n_1105),
.B2(n_924),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1114),
.Y(n_1120)
);

OAI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_1112),
.A2(n_997),
.B1(n_920),
.B2(n_985),
.Y(n_1121)
);

OAI221xp5_ASAP7_75t_L g1122 ( 
.A1(n_1115),
.A2(n_944),
.B1(n_963),
.B2(n_985),
.C(n_923),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1116),
.B(n_929),
.Y(n_1123)
);

OAI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1120),
.A2(n_1118),
.B(n_1110),
.Y(n_1124)
);

OAI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1123),
.A2(n_1117),
.B(n_1113),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_1119),
.Y(n_1126)
);

OA22x2_ASAP7_75t_L g1127 ( 
.A1(n_1121),
.A2(n_1109),
.B1(n_1111),
.B2(n_921),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_1126),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1124),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1129),
.A2(n_1125),
.B(n_1127),
.Y(n_1130)
);

NOR3xp33_ASAP7_75t_SL g1131 ( 
.A(n_1128),
.B(n_1122),
.C(n_269),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1128),
.Y(n_1132)
);

AOI22xp5_ASAP7_75t_R g1133 ( 
.A1(n_1130),
.A2(n_911),
.B1(n_921),
.B2(n_924),
.Y(n_1133)
);

OAI222xp33_ASAP7_75t_L g1134 ( 
.A1(n_1132),
.A2(n_944),
.B1(n_928),
.B2(n_906),
.C1(n_929),
.C2(n_924),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1133),
.Y(n_1135)
);

OAI211xp5_ASAP7_75t_L g1136 ( 
.A1(n_1134),
.A2(n_1131),
.B(n_928),
.C(n_911),
.Y(n_1136)
);

OAI221xp5_ASAP7_75t_R g1137 ( 
.A1(n_1135),
.A2(n_1136),
.B1(n_924),
.B2(n_930),
.C(n_929),
.Y(n_1137)
);

AOI211xp5_ASAP7_75t_L g1138 ( 
.A1(n_1137),
.A2(n_929),
.B(n_914),
.C(n_906),
.Y(n_1138)
);


endmodule