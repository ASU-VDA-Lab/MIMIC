module fake_jpeg_29278_n_38 (n_3, n_2, n_1, n_0, n_4, n_5, n_38);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_38;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g6 ( 
.A(n_4),
.B(n_3),
.Y(n_6)
);

BUFx24_ASAP7_75t_L g7 ( 
.A(n_1),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

INVx13_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_1),
.B(n_5),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_2),
.B(n_1),
.Y(n_12)
);

AOI22xp33_ASAP7_75t_SL g13 ( 
.A1(n_8),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_13)
);

AOI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_13),
.A2(n_19),
.B1(n_2),
.B2(n_3),
.Y(n_21)
);

OA22x2_ASAP7_75t_L g14 ( 
.A1(n_8),
.A2(n_7),
.B1(n_11),
.B2(n_9),
.Y(n_14)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_16),
.C(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_15),
.B(n_16),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_17),
.B(n_18),
.Y(n_24)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_21),
.A2(n_22),
.B(n_23),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_14),
.A2(n_6),
.B1(n_12),
.B2(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_24),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_26),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_22),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_14),
.Y(n_29)
);

OAI221xp5_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_30),
.B1(n_28),
.B2(n_25),
.C(n_19),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_14),
.C(n_18),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_32),
.A2(n_9),
.B(n_10),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_30),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_34),
.A2(n_35),
.B1(n_0),
.B2(n_23),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_0),
.C(n_28),
.Y(n_37)
);

BUFx24_ASAP7_75t_SL g38 ( 
.A(n_37),
.Y(n_38)
);


endmodule