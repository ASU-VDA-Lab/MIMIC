module fake_aes_10917_n_46 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_15, n_10, n_8, n_0, n_46);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_15;
input n_10;
input n_8;
input n_0;
output n_46;
wire n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_30;
wire n_26;
wire n_33;
wire n_16;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_42;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_43;
wire n_40;
wire n_29;
wire n_39;
AND2x4_ASAP7_75t_L g16 ( .A(n_10), .B(n_5), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_8), .Y(n_17) );
BUFx10_ASAP7_75t_L g18 ( .A(n_4), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_14), .B(n_4), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_13), .Y(n_20) );
AND2x2_ASAP7_75t_L g21 ( .A(n_3), .B(n_7), .Y(n_21) );
AND2x2_ASAP7_75t_L g22 ( .A(n_0), .B(n_1), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_6), .Y(n_23) );
INVx2_ASAP7_75t_L g24 ( .A(n_20), .Y(n_24) );
HB1xp67_ASAP7_75t_L g25 ( .A(n_22), .Y(n_25) );
AND2x2_ASAP7_75t_L g26 ( .A(n_18), .B(n_0), .Y(n_26) );
CKINVDCx5p33_ASAP7_75t_R g27 ( .A(n_18), .Y(n_27) );
INVx6_ASAP7_75t_L g28 ( .A(n_26), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_25), .Y(n_29) );
OAI21x1_ASAP7_75t_L g30 ( .A1(n_24), .A2(n_20), .B(n_23), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_30), .Y(n_31) );
NAND4xp25_ASAP7_75t_L g32 ( .A(n_29), .B(n_22), .C(n_19), .D(n_17), .Y(n_32) );
BUFx2_ASAP7_75t_L g33 ( .A(n_31), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_32), .Y(n_34) );
NAND2xp5_ASAP7_75t_L g35 ( .A(n_34), .B(n_25), .Y(n_35) );
AOI211x1_ASAP7_75t_L g36 ( .A1(n_33), .A2(n_21), .B(n_18), .C(n_28), .Y(n_36) );
INVx1_ASAP7_75t_L g37 ( .A(n_35), .Y(n_37) );
INVx1_ASAP7_75t_L g38 ( .A(n_36), .Y(n_38) );
AOI322xp5_ASAP7_75t_L g39 ( .A1(n_35), .A2(n_27), .A3(n_21), .B1(n_16), .B2(n_1), .C1(n_2), .C2(n_3), .Y(n_39) );
INVx1_ASAP7_75t_L g40 ( .A(n_37), .Y(n_40) );
INVx1_ASAP7_75t_L g41 ( .A(n_38), .Y(n_41) );
AND2x2_ASAP7_75t_SL g42 ( .A(n_39), .B(n_33), .Y(n_42) );
AOI22xp5_ASAP7_75t_L g43 ( .A1(n_42), .A2(n_28), .B1(n_16), .B2(n_30), .Y(n_43) );
INVx1_ASAP7_75t_L g44 ( .A(n_40), .Y(n_44) );
AOI22xp5_ASAP7_75t_SL g45 ( .A1(n_44), .A2(n_41), .B1(n_42), .B2(n_16), .Y(n_45) );
OA331x2_ASAP7_75t_L g46 ( .A1(n_45), .A2(n_43), .A3(n_2), .B1(n_11), .B2(n_12), .B3(n_15), .C1(n_9), .Y(n_46) );
endmodule