module fake_jpeg_28551_n_533 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_533);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_533;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_16),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_12),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_11),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_55),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_56),
.Y(n_128)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_31),
.Y(n_58)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_59),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_60),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_17),
.B(n_7),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_61),
.B(n_25),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g62 ( 
.A(n_21),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g111 ( 
.A(n_62),
.Y(n_111)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_63),
.Y(n_123)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_64),
.Y(n_113)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_65),
.Y(n_124)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_66),
.Y(n_154)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_67),
.Y(n_152)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_68),
.B(n_71),
.Y(n_119)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_69),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx3_ASAP7_75t_SL g136 ( 
.A(n_70),
.Y(n_136)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_72),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_74),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_75),
.Y(n_149)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_34),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_76),
.Y(n_137)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_80),
.Y(n_117)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_82),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_83),
.Y(n_147)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_84),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_85),
.Y(n_161)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_21),
.Y(n_86)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_86),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_87),
.Y(n_142)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_88),
.Y(n_155)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_37),
.Y(n_89)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_89),
.Y(n_133)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_90),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_91),
.Y(n_134)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_39),
.Y(n_92)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_92),
.Y(n_139)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_93),
.Y(n_143)
);

BUFx12_ASAP7_75t_L g94 ( 
.A(n_21),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_94),
.B(n_99),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_39),
.Y(n_95)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_36),
.Y(n_96)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_96),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_17),
.B(n_7),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_97),
.B(n_35),
.Y(n_148)
);

BUFx24_ASAP7_75t_L g98 ( 
.A(n_21),
.Y(n_98)
);

INVx2_ASAP7_75t_SL g160 ( 
.A(n_98),
.Y(n_160)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_24),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_36),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_100),
.Y(n_116)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_40),
.Y(n_101)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_101),
.Y(n_165)
);

INVx5_ASAP7_75t_SL g102 ( 
.A(n_18),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_102),
.B(n_108),
.Y(n_169)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_36),
.Y(n_103)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_103),
.Y(n_168)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_36),
.Y(n_104)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_104),
.Y(n_170)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_44),
.Y(n_105)
);

NAND2xp33_ASAP7_75t_SL g110 ( 
.A(n_105),
.B(n_106),
.Y(n_110)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

BUFx10_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_24),
.Y(n_108)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_54),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_109),
.B(n_28),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_102),
.A2(n_18),
.B1(n_19),
.B2(n_54),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_129),
.A2(n_150),
.B1(n_163),
.B2(n_164),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_61),
.A2(n_25),
.B1(n_53),
.B2(n_52),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_132),
.A2(n_146),
.B1(n_22),
.B2(n_33),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_144),
.B(n_148),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_76),
.A2(n_44),
.B1(n_19),
.B2(n_18),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_90),
.A2(n_19),
.B1(n_54),
.B2(n_44),
.Y(n_150)
);

OA22x2_ASAP7_75t_L g151 ( 
.A1(n_77),
.A2(n_43),
.B1(n_50),
.B2(n_47),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_151),
.A2(n_153),
.B1(n_173),
.B2(n_22),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_82),
.A2(n_73),
.B1(n_70),
.B2(n_78),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_87),
.B(n_42),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_158),
.B(n_167),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_94),
.B(n_35),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_162),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_55),
.B(n_42),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_75),
.A2(n_54),
.B1(n_28),
.B2(n_47),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_83),
.A2(n_28),
.B1(n_41),
.B2(n_50),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_91),
.B(n_53),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_172),
.Y(n_218)
);

OA22x2_ASAP7_75t_L g173 ( 
.A1(n_103),
.A2(n_41),
.B1(n_30),
.B2(n_45),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_119),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_174),
.B(n_185),
.Y(n_236)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_138),
.Y(n_175)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_175),
.Y(n_238)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_155),
.Y(n_176)
);

INVx13_ASAP7_75t_L g232 ( 
.A(n_176),
.Y(n_232)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_133),
.Y(n_178)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_178),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_179),
.A2(n_184),
.B1(n_129),
.B2(n_163),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_180),
.A2(n_181),
.B1(n_188),
.B2(n_211),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_153),
.A2(n_95),
.B1(n_104),
.B2(n_59),
.Y(n_181)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_128),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_182),
.Y(n_245)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_128),
.Y(n_183)
);

INVx6_ASAP7_75t_L g243 ( 
.A(n_183),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_151),
.A2(n_60),
.B1(n_56),
.B2(n_96),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_169),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_139),
.Y(n_186)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_186),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_161),
.Y(n_187)
);

INVx5_ASAP7_75t_L g246 ( 
.A(n_187),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_164),
.A2(n_72),
.B1(n_62),
.B2(n_86),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_143),
.Y(n_189)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_189),
.Y(n_248)
);

INVx13_ASAP7_75t_L g190 ( 
.A(n_149),
.Y(n_190)
);

BUFx12f_ASAP7_75t_L g252 ( 
.A(n_190),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_144),
.B(n_33),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_191),
.B(n_201),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_151),
.B(n_32),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_192),
.B(n_212),
.Y(n_233)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_168),
.Y(n_193)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_193),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_146),
.A2(n_45),
.B1(n_43),
.B2(n_30),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_194),
.A2(n_217),
.B1(n_226),
.B2(n_160),
.Y(n_241)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_122),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_195),
.Y(n_244)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_171),
.Y(n_196)
);

INVx8_ASAP7_75t_L g257 ( 
.A(n_196),
.Y(n_257)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_127),
.Y(n_198)
);

INVx5_ASAP7_75t_L g264 ( 
.A(n_198),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g263 ( 
.A(n_199),
.Y(n_263)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_140),
.Y(n_200)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_200),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_123),
.Y(n_201)
);

BUFx10_ASAP7_75t_L g202 ( 
.A(n_121),
.Y(n_202)
);

INVx13_ASAP7_75t_L g254 ( 
.A(n_202),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_130),
.B(n_52),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_203),
.B(n_208),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_135),
.A2(n_100),
.B1(n_28),
.B2(n_32),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_204),
.A2(n_209),
.B1(n_213),
.B2(n_214),
.Y(n_242)
);

BUFx12f_ASAP7_75t_L g205 ( 
.A(n_140),
.Y(n_205)
);

INVx13_ASAP7_75t_L g262 ( 
.A(n_205),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_112),
.Y(n_206)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_206),
.Y(n_265)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_170),
.Y(n_207)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_207),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_118),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_135),
.A2(n_28),
.B1(n_98),
.B2(n_51),
.Y(n_209)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_166),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_210),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_150),
.A2(n_51),
.B1(n_27),
.B2(n_9),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_173),
.B(n_9),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_110),
.A2(n_51),
.B1(n_27),
.B2(n_9),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_152),
.Y(n_214)
);

INVx3_ASAP7_75t_SL g215 ( 
.A(n_138),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_215),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_155),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_216),
.B(n_224),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_136),
.A2(n_27),
.B1(n_8),
.B2(n_10),
.Y(n_217)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_166),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_219),
.B(n_221),
.Y(n_256)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_117),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_114),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_222),
.B(n_223),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_173),
.B(n_159),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_124),
.B(n_27),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_157),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_225),
.B(n_137),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_136),
.A2(n_137),
.B1(n_147),
.B2(n_126),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_228),
.A2(n_253),
.B1(n_175),
.B2(n_200),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_220),
.A2(n_141),
.B(n_113),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_229),
.A2(n_241),
.B(n_268),
.Y(n_281)
);

AND2x2_ASAP7_75t_SL g231 ( 
.A(n_223),
.B(n_111),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_231),
.B(n_235),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_180),
.A2(n_154),
.B1(n_131),
.B2(n_115),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_234),
.A2(n_250),
.B1(n_142),
.B2(n_189),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_227),
.B(n_111),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_241),
.B(n_242),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_192),
.A2(n_212),
.B1(n_179),
.B2(n_194),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_227),
.A2(n_154),
.B1(n_134),
.B2(n_145),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_218),
.A2(n_160),
.B(n_116),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_259),
.A2(n_187),
.B(n_116),
.Y(n_282)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_261),
.Y(n_272)
);

NOR2x1_ASAP7_75t_R g268 ( 
.A(n_218),
.B(n_121),
.Y(n_268)
);

OAI21xp33_ASAP7_75t_L g293 ( 
.A1(n_268),
.A2(n_116),
.B(n_176),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_237),
.B(n_177),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_269),
.B(n_271),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_235),
.B(n_197),
.C(n_188),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_270),
.B(n_265),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_233),
.B(n_214),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_261),
.Y(n_273)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_273),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_275),
.B(n_277),
.Y(n_322)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_256),
.Y(n_276)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_276),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_230),
.B(n_228),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_236),
.B(n_222),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_278),
.B(n_283),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_279),
.B(n_290),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_256),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_280),
.B(n_289),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_281),
.A2(n_282),
.B(n_275),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_282),
.A2(n_302),
.B(n_252),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_233),
.B(n_178),
.Y(n_283)
);

OAI22x1_ASAP7_75t_SL g284 ( 
.A1(n_230),
.A2(n_211),
.B1(n_181),
.B2(n_215),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g318 ( 
.A1(n_284),
.A2(n_291),
.B1(n_267),
.B2(n_240),
.Y(n_318)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_248),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_285),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_234),
.A2(n_142),
.B1(n_186),
.B2(n_156),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_286),
.A2(n_287),
.B1(n_292),
.B2(n_296),
.Y(n_315)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_263),
.Y(n_288)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_288),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_249),
.B(n_198),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_260),
.B(n_207),
.Y(n_290)
);

OAI22xp33_ASAP7_75t_L g291 ( 
.A1(n_260),
.A2(n_219),
.B1(n_210),
.B2(n_208),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_242),
.A2(n_225),
.B1(n_193),
.B2(n_165),
.Y(n_292)
);

OAI21xp33_ASAP7_75t_L g311 ( 
.A1(n_293),
.A2(n_295),
.B(n_267),
.Y(n_311)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_239),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_294),
.B(n_298),
.Y(n_320)
);

HAxp5_ASAP7_75t_SL g295 ( 
.A(n_231),
.B(n_229),
.CON(n_295),
.SN(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_231),
.A2(n_196),
.B1(n_182),
.B2(n_183),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_253),
.A2(n_199),
.B1(n_205),
.B2(n_125),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_297),
.A2(n_299),
.B1(n_255),
.B2(n_263),
.Y(n_321)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_248),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_247),
.A2(n_120),
.B1(n_205),
.B2(n_13),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_244),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_300),
.B(n_301),
.Y(n_329)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_251),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_247),
.A2(n_202),
.B(n_121),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_274),
.B(n_259),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_303),
.B(n_308),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g350 ( 
.A1(n_304),
.A2(n_313),
.B(n_272),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_275),
.A2(n_265),
.B(n_255),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_306),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_275),
.A2(n_277),
.B(n_270),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_307),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_274),
.B(n_251),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_310),
.B(n_324),
.C(n_273),
.Y(n_337)
);

XNOR2x2_ASAP7_75t_SL g359 ( 
.A(n_311),
.B(n_202),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_278),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g361 ( 
.A(n_314),
.B(n_317),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_289),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_318),
.A2(n_272),
.B1(n_299),
.B2(n_302),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_284),
.A2(n_277),
.B1(n_287),
.B2(n_280),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_319),
.A2(n_321),
.B1(n_298),
.B2(n_285),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_283),
.B(n_266),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_300),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_325),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_269),
.B(n_244),
.Y(n_330)
);

CKINVDCx14_ASAP7_75t_R g363 ( 
.A(n_330),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_271),
.B(n_240),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_331),
.B(n_333),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_277),
.A2(n_266),
.B(n_258),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_332),
.B(n_238),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_290),
.B(n_258),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_329),
.Y(n_334)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_334),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_326),
.A2(n_284),
.B1(n_276),
.B2(n_296),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_335),
.A2(n_327),
.B1(n_331),
.B2(n_314),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_SL g374 ( 
.A(n_337),
.B(n_303),
.Y(n_374)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_329),
.Y(n_338)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_338),
.Y(n_389)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_320),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_339),
.B(n_341),
.Y(n_367)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_320),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_342),
.A2(n_351),
.B1(n_315),
.B2(n_326),
.Y(n_366)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_333),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_343),
.B(n_345),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_323),
.Y(n_344)
);

INVx4_ASAP7_75t_SL g386 ( 
.A(n_344),
.Y(n_386)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_312),
.Y(n_345)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_323),
.Y(n_348)
);

INVx2_ASAP7_75t_SL g384 ( 
.A(n_348),
.Y(n_384)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_312),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_349),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g385 ( 
.A1(n_350),
.A2(n_362),
.B(n_322),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_318),
.A2(n_281),
.B1(n_279),
.B2(n_292),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_L g352 ( 
.A1(n_319),
.A2(n_286),
.B1(n_297),
.B2(n_301),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_352),
.A2(n_353),
.B1(n_317),
.B2(n_305),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_316),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_355),
.Y(n_368)
);

CKINVDCx14_ASAP7_75t_R g387 ( 
.A(n_356),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_308),
.B(n_294),
.C(n_239),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_357),
.B(n_310),
.C(n_307),
.Y(n_373)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_316),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_358),
.B(n_360),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_359),
.A2(n_304),
.B(n_306),
.Y(n_364)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_327),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_313),
.A2(n_252),
.B(n_246),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_364),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_366),
.B(n_375),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_355),
.B(n_330),
.Y(n_370)
);

NAND3xp33_ASAP7_75t_L g418 ( 
.A(n_370),
.B(n_340),
.C(n_360),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_336),
.B(n_308),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_372),
.B(n_374),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_373),
.B(n_377),
.C(n_382),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_351),
.A2(n_322),
.B1(n_315),
.B2(n_321),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_376),
.A2(n_392),
.B1(n_342),
.B2(n_343),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_357),
.B(n_310),
.C(n_303),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_361),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_378),
.B(n_393),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_336),
.B(n_324),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_379),
.B(n_381),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_337),
.B(n_324),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_354),
.B(n_328),
.C(n_309),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_SL g383 ( 
.A(n_350),
.B(n_309),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_383),
.B(n_374),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_385),
.B(n_362),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_334),
.B(n_328),
.Y(n_388)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_388),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_363),
.B(n_361),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_390),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_347),
.B(n_325),
.Y(n_391)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_391),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_349),
.Y(n_393)
);

BUFx24_ASAP7_75t_SL g394 ( 
.A(n_358),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_394),
.B(n_338),
.Y(n_401)
);

INVx13_ASAP7_75t_L g400 ( 
.A(n_386),
.Y(n_400)
);

CKINVDCx14_ASAP7_75t_R g435 ( 
.A(n_400),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_401),
.B(n_419),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_368),
.B(n_341),
.Y(n_403)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_403),
.Y(n_446)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_367),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_406),
.B(n_410),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_369),
.B(n_339),
.Y(n_408)
);

CKINVDCx14_ASAP7_75t_R g443 ( 
.A(n_408),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_409),
.A2(n_416),
.B(n_288),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_369),
.B(n_340),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_389),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_411),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_412),
.A2(n_422),
.B1(n_375),
.B2(n_353),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_385),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_413),
.B(n_418),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_373),
.B(n_377),
.C(n_381),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_414),
.B(n_417),
.C(n_383),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_382),
.B(n_347),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_415),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_389),
.B(n_322),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_372),
.B(n_354),
.C(n_346),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_387),
.B(n_345),
.Y(n_419)
);

OA21x2_ASAP7_75t_SL g420 ( 
.A1(n_388),
.A2(n_359),
.B(n_346),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_420),
.A2(n_384),
.B1(n_246),
.B2(n_264),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_421),
.B(n_379),
.Y(n_427)
);

AOI22xp33_ASAP7_75t_L g422 ( 
.A1(n_386),
.A2(n_348),
.B1(n_344),
.B2(n_305),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_367),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_423),
.B(n_380),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_427),
.B(n_429),
.Y(n_460)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_428),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_396),
.A2(n_392),
.B1(n_322),
.B2(n_364),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_430),
.A2(n_404),
.B1(n_413),
.B2(n_410),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_431),
.A2(n_432),
.B1(n_438),
.B2(n_441),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_395),
.A2(n_366),
.B1(n_380),
.B2(n_371),
.Y(n_432)
);

MAJx2_ASAP7_75t_L g436 ( 
.A(n_417),
.B(n_371),
.C(n_332),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_SL g453 ( 
.A(n_436),
.B(n_408),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_398),
.B(n_365),
.C(n_384),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_437),
.B(n_440),
.C(n_444),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_395),
.A2(n_384),
.B1(n_243),
.B2(n_245),
.Y(n_438)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_439),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_402),
.B(n_238),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_412),
.A2(n_243),
.B1(n_245),
.B2(n_257),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_398),
.B(n_232),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_442),
.B(n_447),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_414),
.B(n_288),
.C(n_257),
.Y(n_444)
);

OR2x2_ASAP7_75t_L g448 ( 
.A(n_445),
.B(n_409),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_407),
.B(n_402),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_448),
.B(n_461),
.Y(n_476)
);

OR2x2_ASAP7_75t_L g449 ( 
.A(n_433),
.B(n_403),
.Y(n_449)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_449),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_428),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_452),
.B(n_459),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_453),
.B(n_465),
.C(n_429),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_454),
.B(n_457),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_426),
.A2(n_405),
.B1(n_397),
.B2(n_399),
.Y(n_456)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_456),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_432),
.A2(n_416),
.B1(n_404),
.B2(n_409),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_457),
.A2(n_466),
.B1(n_430),
.B2(n_443),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_426),
.A2(n_411),
.B1(n_416),
.B2(n_421),
.Y(n_459)
);

INVx1_ASAP7_75t_SL g461 ( 
.A(n_446),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_425),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_462),
.B(n_463),
.Y(n_480)
);

BUFx24_ASAP7_75t_SL g463 ( 
.A(n_424),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_437),
.B(n_407),
.C(n_400),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_431),
.A2(n_245),
.B1(n_264),
.B2(n_263),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_467),
.B(n_4),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_468),
.B(n_469),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_460),
.B(n_447),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_471),
.A2(n_262),
.B1(n_190),
.B2(n_11),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_455),
.A2(n_425),
.B1(n_445),
.B2(n_434),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_472),
.A2(n_461),
.B1(n_453),
.B2(n_455),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_449),
.B(n_444),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_474),
.B(n_475),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_458),
.A2(n_438),
.B1(n_441),
.B2(n_435),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_SL g477 ( 
.A1(n_448),
.A2(n_436),
.B(n_442),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_477),
.A2(n_6),
.B(n_14),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_464),
.B(n_440),
.C(n_427),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_478),
.B(n_481),
.C(n_6),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g479 ( 
.A(n_450),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_479),
.B(n_483),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_464),
.B(n_232),
.C(n_254),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_454),
.A2(n_263),
.B1(n_254),
.B2(n_14),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_484),
.B(n_485),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_469),
.B(n_465),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_482),
.A2(n_451),
.B1(n_466),
.B2(n_460),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_486),
.B(n_492),
.Y(n_508)
);

AOI22xp33_ASAP7_75t_SL g487 ( 
.A1(n_473),
.A2(n_252),
.B1(n_262),
.B2(n_202),
.Y(n_487)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_487),
.Y(n_501)
);

NOR2xp67_ASAP7_75t_L g488 ( 
.A(n_480),
.B(n_252),
.Y(n_488)
);

AOI21x1_ASAP7_75t_SL g510 ( 
.A1(n_488),
.A2(n_475),
.B(n_471),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_491),
.B(n_483),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_478),
.B(n_27),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_SL g494 ( 
.A1(n_476),
.A2(n_5),
.B(n_14),
.Y(n_494)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_494),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_L g495 ( 
.A1(n_467),
.A2(n_5),
.B(n_14),
.Y(n_495)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_495),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_SL g500 ( 
.A(n_496),
.B(n_497),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_498),
.B(n_11),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_489),
.B(n_476),
.Y(n_499)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_499),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_490),
.A2(n_472),
.B1(n_468),
.B2(n_498),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_503),
.B(n_509),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_493),
.B(n_481),
.C(n_470),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_506),
.B(n_507),
.Y(n_512)
);

INVxp33_ASAP7_75t_L g517 ( 
.A(n_510),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_L g511 ( 
.A1(n_504),
.A2(n_496),
.B(n_491),
.Y(n_511)
);

AO21x1_ASAP7_75t_L g522 ( 
.A1(n_511),
.A2(n_515),
.B(n_3),
.Y(n_522)
);

XNOR2x1_ASAP7_75t_L g513 ( 
.A(n_508),
.B(n_493),
.Y(n_513)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_513),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_SL g515 ( 
.A1(n_499),
.A2(n_501),
.B(n_502),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_SL g518 ( 
.A1(n_505),
.A2(n_487),
.B(n_494),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g519 ( 
.A1(n_518),
.A2(n_501),
.B(n_507),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_SL g526 ( 
.A1(n_519),
.A2(n_521),
.B(n_514),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_516),
.A2(n_477),
.B(n_500),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_522),
.B(n_523),
.Y(n_524)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_512),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_520),
.B(n_517),
.Y(n_525)
);

OAI21xp33_ASAP7_75t_L g527 ( 
.A1(n_525),
.A2(n_514),
.B(n_6),
.Y(n_527)
);

OAI311xp33_ASAP7_75t_L g528 ( 
.A1(n_526),
.A2(n_3),
.A3(n_13),
.B1(n_15),
.C1(n_0),
.Y(n_528)
);

A2O1A1Ixp33_ASAP7_75t_L g529 ( 
.A1(n_527),
.A2(n_528),
.B(n_524),
.C(n_1),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_SL g530 ( 
.A1(n_529),
.A2(n_1),
.B(n_2),
.Y(n_530)
);

AOI21x1_ASAP7_75t_L g531 ( 
.A1(n_530),
.A2(n_1),
.B(n_2),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_531),
.A2(n_1),
.B(n_2),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_532),
.B(n_2),
.Y(n_533)
);


endmodule