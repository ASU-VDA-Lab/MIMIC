module fake_netlist_6_3131_n_1902 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1902);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1902;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1348;
wire n_1209;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_268;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_297;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx2_ASAP7_75t_L g178 ( 
.A(n_107),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_108),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_142),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_118),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_16),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_117),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_3),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_32),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_103),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_45),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_68),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_62),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_13),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_93),
.Y(n_191)
);

BUFx2_ASAP7_75t_SL g192 ( 
.A(n_19),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_65),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_172),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_110),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_14),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_51),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_76),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_6),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_7),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_69),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_102),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_70),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_135),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_56),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_154),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_153),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_13),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_145),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_53),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_150),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_15),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_23),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_109),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_37),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_68),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_155),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_139),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_80),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_177),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_116),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_111),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_11),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_43),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_5),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_134),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_38),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_38),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_46),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_95),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_43),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_129),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_138),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_16),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_57),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_33),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_163),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_6),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_112),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_4),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_64),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_46),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_44),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_148),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_94),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_130),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_157),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_126),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_62),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_17),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_137),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_90),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_89),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_22),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_169),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_71),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_49),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_140),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_113),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_26),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_67),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_60),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_53),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_32),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_86),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_100),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_51),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_20),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_166),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_52),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_41),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_174),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_167),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_49),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_161),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_115),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_120),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_131),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_4),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_160),
.Y(n_280)
);

INVx2_ASAP7_75t_SL g281 ( 
.A(n_122),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_14),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_168),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_60),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_40),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_56),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_104),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_175),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_39),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_52),
.Y(n_290)
);

BUFx5_ASAP7_75t_L g291 ( 
.A(n_158),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_119),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_12),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_30),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_79),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_159),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_105),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_57),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_67),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_28),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_42),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_144),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_72),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_55),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_55),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_73),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_1),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_99),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_37),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_1),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_39),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_171),
.Y(n_312)
);

INVx2_ASAP7_75t_SL g313 ( 
.A(n_2),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_121),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_40),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_54),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_26),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_149),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_114),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_77),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_88),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_101),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_22),
.Y(n_323)
);

BUFx10_ASAP7_75t_L g324 ( 
.A(n_133),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_42),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_91),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_74),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_35),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_41),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_28),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_162),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_7),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_124),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_97),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_21),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_12),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_10),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_143),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_152),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_165),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_176),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_127),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_48),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_78),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_36),
.Y(n_345)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_123),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_24),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_54),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_65),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_47),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_164),
.Y(n_351)
);

BUFx10_ASAP7_75t_L g352 ( 
.A(n_31),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_87),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_61),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_59),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_181),
.Y(n_356)
);

BUFx2_ASAP7_75t_L g357 ( 
.A(n_210),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_193),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_183),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_R g360 ( 
.A(n_202),
.B(n_173),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_191),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_221),
.Y(n_362)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_224),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_193),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_224),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_193),
.Y(n_366)
);

OR2x2_ASAP7_75t_L g367 ( 
.A(n_187),
.B(n_0),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_193),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_193),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_299),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_288),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_194),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_299),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_198),
.Y(n_374)
);

INVxp67_ASAP7_75t_SL g375 ( 
.A(n_278),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_327),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_299),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_299),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_299),
.Y(n_379)
);

INVxp67_ASAP7_75t_SL g380 ( 
.A(n_278),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_237),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_352),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_315),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_315),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_237),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_247),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_315),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_203),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_315),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_315),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_207),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_316),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g393 ( 
.A(n_264),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_247),
.Y(n_394)
);

NOR2xp67_ASAP7_75t_L g395 ( 
.A(n_313),
.B(n_0),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_211),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_214),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_302),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_264),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_210),
.B(n_2),
.Y(n_400)
);

NOR2xp67_ASAP7_75t_L g401 ( 
.A(n_313),
.B(n_3),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_316),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_316),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_217),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_218),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_219),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_316),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_222),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_226),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_232),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_233),
.Y(n_411)
);

BUFx6f_ASAP7_75t_SL g412 ( 
.A(n_324),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_316),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_196),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_196),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_352),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_223),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_182),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_352),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_223),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_274),
.Y(n_421)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_324),
.Y(n_422)
);

INVxp33_ASAP7_75t_SL g423 ( 
.A(n_189),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_291),
.Y(n_424)
);

INVxp67_ASAP7_75t_SL g425 ( 
.A(n_339),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_239),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_274),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_281),
.B(n_5),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_284),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_284),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_190),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_248),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_289),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_255),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_256),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_289),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_187),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_258),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_188),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_188),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_208),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_208),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_291),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_259),
.Y(n_444)
);

INVxp33_ASAP7_75t_SL g445 ( 
.A(n_197),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_366),
.B(n_339),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_358),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_424),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_358),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_375),
.B(n_281),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_366),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_424),
.Y(n_452)
);

OAI21x1_ASAP7_75t_L g453 ( 
.A1(n_428),
.A2(n_206),
.B(n_178),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_364),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_364),
.Y(n_455)
);

BUFx2_ASAP7_75t_L g456 ( 
.A(n_381),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_368),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_400),
.B(n_234),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_368),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_443),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_380),
.B(n_425),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_369),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_369),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_370),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_443),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_370),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_373),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_373),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_363),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_377),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_377),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_378),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_423),
.B(n_445),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_378),
.Y(n_474)
);

AND2x2_ASAP7_75t_SL g475 ( 
.A(n_400),
.B(n_178),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_379),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_379),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_383),
.B(n_265),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_383),
.Y(n_479)
);

NOR2x1_ASAP7_75t_L g480 ( 
.A(n_384),
.B(n_206),
.Y(n_480)
);

BUFx2_ASAP7_75t_L g481 ( 
.A(n_385),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_384),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_387),
.Y(n_483)
);

BUFx8_ASAP7_75t_L g484 ( 
.A(n_412),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_387),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_389),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_357),
.B(n_234),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_357),
.B(n_286),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_389),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_390),
.B(n_269),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_390),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_392),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_392),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_402),
.B(n_272),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_402),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_403),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_422),
.B(n_324),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_403),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_407),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_407),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_399),
.Y(n_501)
);

INVx1_ASAP7_75t_SL g502 ( 
.A(n_386),
.Y(n_502)
);

AND2x4_ASAP7_75t_L g503 ( 
.A(n_413),
.B(n_179),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_418),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_413),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_414),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_414),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_415),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_422),
.B(n_199),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_415),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_367),
.A2(n_336),
.B1(n_317),
.B2(n_250),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_417),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_437),
.B(n_273),
.Y(n_513)
);

OAI21x1_ASAP7_75t_L g514 ( 
.A1(n_367),
.A2(n_180),
.B(n_179),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_417),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_420),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_431),
.B(n_326),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_420),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_421),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_421),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_427),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_427),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_429),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_475),
.B(n_356),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_473),
.B(n_359),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_473),
.B(n_361),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_SL g527 ( 
.A(n_469),
.B(n_394),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_446),
.Y(n_528)
);

OR2x6_ASAP7_75t_L g529 ( 
.A(n_461),
.B(n_192),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_460),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_446),
.B(n_180),
.Y(n_531)
);

INVx4_ASAP7_75t_L g532 ( 
.A(n_452),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_452),
.Y(n_533)
);

BUFx10_ASAP7_75t_L g534 ( 
.A(n_517),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_460),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_518),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_504),
.B(n_372),
.Y(n_537)
);

INVxp33_ASAP7_75t_L g538 ( 
.A(n_487),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_460),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_460),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_504),
.A2(n_405),
.B1(n_410),
.B2(n_408),
.Y(n_541)
);

CKINVDCx16_ASAP7_75t_R g542 ( 
.A(n_469),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_461),
.B(n_374),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_458),
.B(n_429),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_517),
.A2(n_398),
.B1(n_391),
.B2(n_396),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_452),
.Y(n_546)
);

INVxp33_ASAP7_75t_L g547 ( 
.A(n_487),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_446),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_518),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_466),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_475),
.B(n_388),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_518),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_484),
.B(n_397),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_466),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_487),
.Y(n_555)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_452),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_484),
.B(n_404),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_475),
.B(n_406),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_518),
.Y(n_559)
);

INVx1_ASAP7_75t_SL g560 ( 
.A(n_502),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_466),
.Y(n_561)
);

INVx4_ASAP7_75t_L g562 ( 
.A(n_452),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_484),
.B(n_409),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_466),
.Y(n_564)
);

AND2x2_ASAP7_75t_SL g565 ( 
.A(n_475),
.B(n_186),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_478),
.B(n_411),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_467),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_446),
.B(n_186),
.Y(n_568)
);

NAND3xp33_ASAP7_75t_L g569 ( 
.A(n_513),
.B(n_432),
.C(n_426),
.Y(n_569)
);

INVx5_ASAP7_75t_L g570 ( 
.A(n_452),
.Y(n_570)
);

INVxp67_ASAP7_75t_SL g571 ( 
.A(n_452),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_L g572 ( 
.A1(n_514),
.A2(n_395),
.B1(n_401),
.B2(n_286),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_520),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_467),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_467),
.Y(n_575)
);

NAND2xp33_ASAP7_75t_SL g576 ( 
.A(n_497),
.B(n_360),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_467),
.Y(n_577)
);

INVx4_ASAP7_75t_L g578 ( 
.A(n_452),
.Y(n_578)
);

OR2x6_ASAP7_75t_L g579 ( 
.A(n_497),
.B(n_192),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_472),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_520),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_478),
.B(n_434),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g583 ( 
.A(n_488),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_520),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_514),
.A2(n_260),
.B1(n_243),
.B2(n_290),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_490),
.B(n_435),
.Y(n_586)
);

AND3x2_ASAP7_75t_L g587 ( 
.A(n_501),
.B(n_416),
.C(n_382),
.Y(n_587)
);

INVx4_ASAP7_75t_L g588 ( 
.A(n_468),
.Y(n_588)
);

OR2x2_ASAP7_75t_L g589 ( 
.A(n_501),
.B(n_363),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_520),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_472),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_472),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_490),
.B(n_438),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_448),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_514),
.A2(n_458),
.B1(n_450),
.B2(n_488),
.Y(n_595)
);

BUFx10_ASAP7_75t_L g596 ( 
.A(n_446),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_455),
.Y(n_597)
);

NAND3xp33_ASAP7_75t_L g598 ( 
.A(n_513),
.B(n_444),
.C(n_419),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_484),
.B(n_365),
.Y(n_599)
);

BUFx2_ASAP7_75t_L g600 ( 
.A(n_488),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_484),
.B(n_365),
.Y(n_601)
);

INVx4_ASAP7_75t_L g602 ( 
.A(n_468),
.Y(n_602)
);

INVxp67_ASAP7_75t_SL g603 ( 
.A(n_494),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_472),
.Y(n_604)
);

BUFx6f_ASAP7_75t_L g605 ( 
.A(n_468),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_494),
.B(n_204),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_479),
.Y(n_607)
);

OAI22xp33_ASAP7_75t_SL g608 ( 
.A1(n_450),
.A2(n_393),
.B1(n_509),
.B2(n_201),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_479),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_446),
.B(n_220),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_479),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_458),
.A2(n_260),
.B1(n_290),
.B2(n_243),
.Y(n_612)
);

AND2x6_ASAP7_75t_L g613 ( 
.A(n_503),
.B(n_201),
.Y(n_613)
);

BUFx10_ASAP7_75t_L g614 ( 
.A(n_503),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_503),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_503),
.Y(n_616)
);

INVx2_ASAP7_75t_SL g617 ( 
.A(n_503),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_503),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_455),
.B(n_266),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_457),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_457),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_479),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_509),
.B(n_393),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_491),
.Y(n_624)
);

AND2x2_ASAP7_75t_SL g625 ( 
.A(n_456),
.B(n_209),
.Y(n_625)
);

BUFx2_ASAP7_75t_L g626 ( 
.A(n_456),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_495),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_484),
.B(n_275),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_448),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_523),
.B(n_412),
.Y(n_630)
);

NAND2xp33_ASAP7_75t_L g631 ( 
.A(n_480),
.B(n_195),
.Y(n_631)
);

INVx4_ASAP7_75t_L g632 ( 
.A(n_468),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_491),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_512),
.B(n_412),
.Y(n_634)
);

AND2x6_ASAP7_75t_L g635 ( 
.A(n_480),
.B(n_209),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_468),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_511),
.B(n_287),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_496),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_496),
.B(n_280),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_495),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_498),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g642 ( 
.A1(n_511),
.A2(n_300),
.B1(n_282),
.B2(n_279),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_523),
.B(n_362),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_498),
.B(n_447),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_447),
.B(n_295),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_453),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_447),
.B(n_449),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_502),
.B(n_292),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_449),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_512),
.B(n_430),
.Y(n_650)
);

BUFx10_ASAP7_75t_L g651 ( 
.A(n_512),
.Y(n_651)
);

NAND3xp33_ASAP7_75t_L g652 ( 
.A(n_516),
.B(n_212),
.C(n_200),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_506),
.B(n_308),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_495),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_516),
.B(n_430),
.Y(n_655)
);

INVx4_ASAP7_75t_L g656 ( 
.A(n_468),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_495),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_449),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_453),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_499),
.Y(n_660)
);

INVx1_ASAP7_75t_SL g661 ( 
.A(n_456),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_468),
.Y(n_662)
);

BUFx2_ASAP7_75t_L g663 ( 
.A(n_481),
.Y(n_663)
);

AND2x4_ASAP7_75t_SL g664 ( 
.A(n_516),
.B(n_371),
.Y(n_664)
);

AND2x4_ASAP7_75t_L g665 ( 
.A(n_453),
.B(n_230),
.Y(n_665)
);

NOR3xp33_ASAP7_75t_L g666 ( 
.A(n_481),
.B(n_332),
.C(n_227),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_454),
.Y(n_667)
);

OR2x2_ASAP7_75t_L g668 ( 
.A(n_481),
.B(n_437),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_454),
.B(n_346),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_454),
.Y(n_670)
);

OR2x6_ASAP7_75t_L g671 ( 
.A(n_519),
.B(n_225),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_468),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_459),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_523),
.B(n_376),
.Y(n_674)
);

OR2x6_ASAP7_75t_L g675 ( 
.A(n_519),
.B(n_225),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_519),
.B(n_213),
.Y(n_676)
);

NOR3xp33_ASAP7_75t_L g677 ( 
.A(n_576),
.B(n_216),
.C(n_215),
.Y(n_677)
);

INVx4_ASAP7_75t_SL g678 ( 
.A(n_613),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_603),
.B(n_448),
.Y(n_679)
);

INVx2_ASAP7_75t_SL g680 ( 
.A(n_664),
.Y(n_680)
);

OR2x2_ASAP7_75t_L g681 ( 
.A(n_668),
.B(n_439),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_649),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_543),
.B(n_448),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_649),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_528),
.Y(n_685)
);

OR2x2_ASAP7_75t_L g686 ( 
.A(n_668),
.B(n_589),
.Y(n_686)
);

OR2x2_ASAP7_75t_L g687 ( 
.A(n_589),
.B(n_439),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_565),
.B(n_448),
.Y(n_688)
);

INVxp67_ASAP7_75t_L g689 ( 
.A(n_623),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_664),
.Y(n_690)
);

AOI22xp5_ASAP7_75t_L g691 ( 
.A1(n_524),
.A2(n_314),
.B1(n_353),
.B2(n_351),
.Y(n_691)
);

INVxp33_ASAP7_75t_L g692 ( 
.A(n_626),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_565),
.B(n_195),
.Y(n_693)
);

INVxp67_ASAP7_75t_L g694 ( 
.A(n_643),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_658),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_544),
.B(n_440),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_595),
.B(n_195),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_544),
.Y(n_698)
);

NAND3xp33_ASAP7_75t_L g699 ( 
.A(n_555),
.B(n_240),
.C(n_236),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_538),
.B(n_241),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_606),
.B(n_465),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_658),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_538),
.B(n_242),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_670),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_547),
.B(n_319),
.Y(n_705)
);

AND2x4_ASAP7_75t_L g706 ( 
.A(n_528),
.B(n_440),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_670),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_547),
.B(n_551),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_558),
.B(n_249),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_R g710 ( 
.A(n_542),
.B(n_320),
.Y(n_710)
);

AOI22xp33_ASAP7_75t_L g711 ( 
.A1(n_585),
.A2(n_228),
.B1(n_348),
.B2(n_347),
.Y(n_711)
);

AND2x6_ASAP7_75t_SL g712 ( 
.A(n_579),
.B(n_228),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_617),
.B(n_195),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_583),
.B(n_254),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_L g715 ( 
.A1(n_665),
.A2(n_229),
.B1(n_348),
.B2(n_347),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_583),
.B(n_257),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_560),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_600),
.B(n_566),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_548),
.Y(n_719)
);

NOR3xp33_ASAP7_75t_L g720 ( 
.A(n_576),
.B(n_262),
.C(n_261),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_582),
.B(n_586),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_600),
.B(n_263),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_673),
.Y(n_723)
);

O2A1O1Ixp33_ASAP7_75t_L g724 ( 
.A1(n_608),
.A2(n_229),
.B(n_231),
.C(n_235),
.Y(n_724)
);

INVx4_ASAP7_75t_L g725 ( 
.A(n_548),
.Y(n_725)
);

BUFx6f_ASAP7_75t_L g726 ( 
.A(n_596),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_673),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_593),
.B(n_572),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_615),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_616),
.Y(n_730)
);

O2A1O1Ixp33_ASAP7_75t_L g731 ( 
.A1(n_610),
.A2(n_231),
.B(n_235),
.C(n_238),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_597),
.Y(n_732)
);

INVxp67_ASAP7_75t_L g733 ( 
.A(n_674),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_536),
.B(n_465),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_579),
.A2(n_344),
.B1(n_341),
.B2(n_338),
.Y(n_735)
);

NAND2xp33_ASAP7_75t_SL g736 ( 
.A(n_599),
.B(n_601),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_536),
.B(n_465),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_534),
.B(n_321),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_549),
.B(n_465),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_618),
.Y(n_740)
);

AND2x6_ASAP7_75t_SL g741 ( 
.A(n_579),
.B(n_238),
.Y(n_741)
);

NAND2xp33_ASAP7_75t_L g742 ( 
.A(n_613),
.B(n_291),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_549),
.Y(n_743)
);

OAI22xp33_ASAP7_75t_L g744 ( 
.A1(n_579),
.A2(n_283),
.B1(n_230),
.B2(n_244),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_552),
.B(n_465),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_552),
.B(n_515),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_559),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_534),
.B(n_529),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_559),
.B(n_515),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_529),
.B(n_267),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_534),
.B(n_322),
.Y(n_751)
);

OAI22xp33_ASAP7_75t_L g752 ( 
.A1(n_529),
.A2(n_283),
.B1(n_244),
.B2(n_245),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_573),
.B(n_515),
.Y(n_753)
);

INVx2_ASAP7_75t_SL g754 ( 
.A(n_626),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_597),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_573),
.B(n_515),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_581),
.B(n_515),
.Y(n_757)
);

INVx8_ASAP7_75t_L g758 ( 
.A(n_529),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_581),
.Y(n_759)
);

INVxp67_ASAP7_75t_L g760 ( 
.A(n_663),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_617),
.A2(n_331),
.B1(n_333),
.B2(n_334),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_651),
.B(n_195),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_624),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_624),
.Y(n_764)
);

INVx3_ASAP7_75t_L g765 ( 
.A(n_596),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_584),
.B(n_459),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_571),
.A2(n_462),
.B(n_459),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_665),
.A2(n_635),
.B1(n_613),
.B2(n_646),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_584),
.B(n_462),
.Y(n_769)
);

BUFx2_ASAP7_75t_R g770 ( 
.A(n_663),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_SL g771 ( 
.A1(n_625),
.A2(n_184),
.B1(n_185),
.B2(n_205),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_590),
.B(n_462),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_625),
.B(n_441),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_651),
.B(n_246),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_569),
.B(n_268),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_545),
.B(n_441),
.Y(n_776)
);

OAI22xp33_ASAP7_75t_L g777 ( 
.A1(n_671),
.A2(n_675),
.B1(n_598),
.B2(n_669),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_665),
.B(n_246),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_541),
.B(n_537),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_590),
.B(n_463),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_620),
.B(n_463),
.Y(n_781)
);

AND2x2_ASAP7_75t_SL g782 ( 
.A(n_531),
.B(n_245),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_651),
.B(n_442),
.Y(n_783)
);

AND2x6_ASAP7_75t_L g784 ( 
.A(n_531),
.B(n_251),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_525),
.B(n_270),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_614),
.B(n_246),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_650),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_633),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_633),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_646),
.A2(n_463),
.B(n_482),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_637),
.A2(n_277),
.B1(n_251),
.B2(n_342),
.Y(n_791)
);

INVx2_ASAP7_75t_SL g792 ( 
.A(n_531),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_650),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_659),
.A2(n_464),
.B(n_485),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_614),
.B(n_246),
.Y(n_795)
);

AND2x4_ASAP7_75t_L g796 ( 
.A(n_568),
.B(n_442),
.Y(n_796)
);

BUFx6f_ASAP7_75t_L g797 ( 
.A(n_596),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_655),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_638),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_638),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_621),
.B(n_464),
.Y(n_801)
);

INVxp67_ASAP7_75t_L g802 ( 
.A(n_527),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_614),
.B(n_246),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_526),
.B(n_271),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_648),
.B(n_285),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_L g806 ( 
.A(n_619),
.B(n_293),
.Y(n_806)
);

INVx8_ASAP7_75t_L g807 ( 
.A(n_613),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_641),
.B(n_464),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_676),
.B(n_521),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_641),
.B(n_474),
.Y(n_810)
);

BUFx3_ASAP7_75t_L g811 ( 
.A(n_613),
.Y(n_811)
);

AOI21xp5_ASAP7_75t_L g812 ( 
.A1(n_659),
.A2(n_485),
.B(n_474),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_655),
.Y(n_813)
);

AOI22xp5_ASAP7_75t_L g814 ( 
.A1(n_568),
.A2(n_563),
.B1(n_557),
.B2(n_553),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_667),
.B(n_474),
.Y(n_815)
);

INVx8_ASAP7_75t_L g816 ( 
.A(n_613),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_644),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_635),
.A2(n_304),
.B1(n_298),
.B2(n_328),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_L g819 ( 
.A1(n_635),
.A2(n_304),
.B1(n_298),
.B2(n_328),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_647),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_639),
.B(n_252),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_530),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_661),
.B(n_521),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_568),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_594),
.B(n_476),
.Y(n_825)
);

BUFx6f_ASAP7_75t_L g826 ( 
.A(n_546),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_594),
.Y(n_827)
);

INVx4_ASAP7_75t_L g828 ( 
.A(n_546),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_594),
.Y(n_829)
);

NAND2xp33_ASAP7_75t_L g830 ( 
.A(n_635),
.B(n_645),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_530),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_535),
.Y(n_832)
);

AOI22xp5_ASAP7_75t_L g833 ( 
.A1(n_652),
.A2(n_253),
.B1(n_252),
.B2(n_342),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_629),
.B(n_476),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_642),
.B(n_294),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_630),
.B(n_522),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_634),
.B(n_522),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_546),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_629),
.B(n_476),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_535),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_671),
.B(n_301),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_666),
.B(n_522),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_629),
.B(n_477),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_612),
.B(n_253),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_671),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_628),
.B(n_276),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_671),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_546),
.B(n_291),
.Y(n_848)
);

AOI21x1_ASAP7_75t_L g849 ( 
.A1(n_697),
.A2(n_653),
.B(n_540),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_694),
.B(n_675),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_721),
.B(n_809),
.Y(n_851)
);

NOR3xp33_ASAP7_75t_L g852 ( 
.A(n_771),
.B(n_277),
.C(n_276),
.Y(n_852)
);

O2A1O1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_693),
.A2(n_675),
.B(n_631),
.C(n_296),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_679),
.A2(n_683),
.B(n_688),
.Y(n_854)
);

A2O1A1Ixp33_ASAP7_75t_L g855 ( 
.A1(n_708),
.A2(n_318),
.B(n_312),
.C(n_306),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_817),
.B(n_533),
.Y(n_856)
);

OAI21xp33_ASAP7_75t_L g857 ( 
.A1(n_835),
.A2(n_675),
.B(n_307),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_728),
.A2(n_562),
.B(n_532),
.Y(n_858)
);

O2A1O1Ixp33_ASAP7_75t_SL g859 ( 
.A1(n_693),
.A2(n_296),
.B(n_297),
.C(n_340),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_697),
.A2(n_562),
.B(n_532),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_708),
.B(n_533),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_777),
.B(n_546),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_701),
.A2(n_562),
.B(n_532),
.Y(n_863)
);

INVx1_ASAP7_75t_SL g864 ( 
.A(n_717),
.Y(n_864)
);

OAI21xp5_ASAP7_75t_L g865 ( 
.A1(n_790),
.A2(n_533),
.B(n_539),
.Y(n_865)
);

INVx11_ASAP7_75t_L g866 ( 
.A(n_784),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_820),
.B(n_718),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_718),
.B(n_556),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_828),
.A2(n_578),
.B(n_556),
.Y(n_869)
);

OR2x4_ASAP7_75t_L g870 ( 
.A(n_835),
.B(n_587),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_682),
.Y(n_871)
);

INVx4_ASAP7_75t_L g872 ( 
.A(n_726),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_682),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_684),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_684),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_828),
.A2(n_578),
.B(n_556),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_765),
.A2(n_830),
.B(n_795),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_783),
.B(n_709),
.Y(n_878)
);

AOI22xp5_ASAP7_75t_L g879 ( 
.A1(n_709),
.A2(n_635),
.B1(n_578),
.B2(n_631),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_695),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_695),
.Y(n_881)
);

A2O1A1Ixp33_ASAP7_75t_L g882 ( 
.A1(n_715),
.A2(n_318),
.B(n_312),
.C(n_306),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_L g883 ( 
.A1(n_794),
.A2(n_540),
.B(n_539),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_702),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_765),
.A2(n_556),
.B(n_632),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_702),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_786),
.A2(n_556),
.B(n_632),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_836),
.B(n_635),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_837),
.B(n_550),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_704),
.Y(n_890)
);

INVx4_ASAP7_75t_L g891 ( 
.A(n_726),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_786),
.A2(n_656),
.B(n_602),
.Y(n_892)
);

AOI21x1_ASAP7_75t_L g893 ( 
.A1(n_778),
.A2(n_580),
.B(n_567),
.Y(n_893)
);

O2A1O1Ixp5_ASAP7_75t_L g894 ( 
.A1(n_795),
.A2(n_564),
.B(n_550),
.C(n_660),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_704),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_806),
.B(n_554),
.Y(n_896)
);

BUFx2_ASAP7_75t_L g897 ( 
.A(n_754),
.Y(n_897)
);

A2O1A1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_715),
.A2(n_303),
.B(n_297),
.C(n_340),
.Y(n_898)
);

AOI21xp5_ASAP7_75t_L g899 ( 
.A1(n_803),
.A2(n_838),
.B(n_826),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_733),
.B(n_310),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_823),
.B(n_433),
.Y(n_901)
);

AND2x2_ASAP7_75t_SL g902 ( 
.A(n_818),
.B(n_303),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_SL g903 ( 
.A(n_768),
.B(n_605),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_696),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_707),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_SL g906 ( 
.A(n_768),
.B(n_605),
.Y(n_906)
);

BUFx3_ASAP7_75t_L g907 ( 
.A(n_696),
.Y(n_907)
);

AND2x4_ASAP7_75t_L g908 ( 
.A(n_698),
.B(n_521),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_726),
.B(n_605),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_707),
.Y(n_910)
);

AOI22xp33_ASAP7_75t_L g911 ( 
.A1(n_711),
.A2(n_345),
.B1(n_291),
.B2(n_657),
.Y(n_911)
);

A2O1A1Ixp33_ASAP7_75t_L g912 ( 
.A1(n_711),
.A2(n_325),
.B(n_309),
.C(n_311),
.Y(n_912)
);

AOI21x1_ASAP7_75t_L g913 ( 
.A1(n_778),
.A2(n_592),
.B(n_554),
.Y(n_913)
);

AOI21xp33_ASAP7_75t_L g914 ( 
.A1(n_785),
.A2(n_329),
.B(n_355),
.Y(n_914)
);

AND2x6_ASAP7_75t_L g915 ( 
.A(n_811),
.B(n_605),
.Y(n_915)
);

OAI22xp5_ASAP7_75t_L g916 ( 
.A1(n_814),
.A2(n_689),
.B1(n_782),
.B2(n_824),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_723),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_686),
.B(n_773),
.Y(n_918)
);

AND2x4_ASAP7_75t_L g919 ( 
.A(n_845),
.B(n_433),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_776),
.B(n_436),
.Y(n_920)
);

INVx2_ASAP7_75t_SL g921 ( 
.A(n_681),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_802),
.B(n_305),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_723),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_803),
.A2(n_656),
.B(n_602),
.Y(n_924)
);

O2A1O1Ixp33_ASAP7_75t_L g925 ( 
.A1(n_744),
.A2(n_574),
.B(n_660),
.C(n_657),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_727),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_714),
.B(n_436),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_727),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_826),
.A2(n_588),
.B(n_602),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_806),
.B(n_561),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_826),
.A2(n_588),
.B(n_632),
.Y(n_931)
);

INVx3_ASAP7_75t_L g932 ( 
.A(n_725),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_826),
.A2(n_656),
.B(n_588),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_687),
.B(n_323),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_732),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_838),
.A2(n_570),
.B(n_662),
.Y(n_936)
);

NAND3xp33_ASAP7_75t_L g937 ( 
.A(n_785),
.B(n_350),
.C(n_330),
.Y(n_937)
);

NAND2xp33_ASAP7_75t_L g938 ( 
.A(n_726),
.B(n_291),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_838),
.A2(n_570),
.B(n_662),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_732),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_787),
.B(n_561),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_714),
.B(n_716),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_838),
.A2(n_570),
.B(n_662),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_793),
.B(n_564),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_755),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_755),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_SL g947 ( 
.A(n_770),
.B(n_335),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_763),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_797),
.A2(n_570),
.B(n_662),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_797),
.A2(n_792),
.B(n_737),
.Y(n_950)
);

O2A1O1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_724),
.A2(n_627),
.B(n_654),
.C(n_640),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_798),
.B(n_567),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_813),
.B(n_574),
.Y(n_953)
);

INVx3_ASAP7_75t_L g954 ( 
.A(n_725),
.Y(n_954)
);

INVx5_ASAP7_75t_L g955 ( 
.A(n_807),
.Y(n_955)
);

OAI21xp33_ASAP7_75t_L g956 ( 
.A1(n_804),
.A2(n_337),
.B(n_343),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_L g957 ( 
.A1(n_736),
.A2(n_604),
.B1(n_575),
.B2(n_654),
.Y(n_957)
);

INVx3_ASAP7_75t_L g958 ( 
.A(n_706),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_729),
.B(n_575),
.Y(n_959)
);

AOI21x1_ASAP7_75t_L g960 ( 
.A1(n_812),
.A2(n_577),
.B(n_580),
.Y(n_960)
);

OAI21xp5_ASAP7_75t_L g961 ( 
.A1(n_746),
.A2(n_592),
.B(n_604),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_716),
.B(n_349),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_730),
.B(n_740),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_763),
.B(n_577),
.Y(n_964)
);

INVx1_ASAP7_75t_SL g965 ( 
.A(n_692),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_764),
.B(n_591),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_797),
.A2(n_570),
.B(n_662),
.Y(n_967)
);

INVx3_ASAP7_75t_L g968 ( 
.A(n_706),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_797),
.A2(n_672),
.B(n_605),
.Y(n_969)
);

AOI22xp5_ASAP7_75t_L g970 ( 
.A1(n_782),
.A2(n_779),
.B1(n_685),
.B2(n_719),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_788),
.B(n_591),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_700),
.B(n_703),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_788),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_789),
.Y(n_974)
);

AOI33xp33_ASAP7_75t_L g975 ( 
.A1(n_842),
.A2(n_510),
.A3(n_354),
.B1(n_482),
.B2(n_485),
.B3(n_477),
.Y(n_975)
);

A2O1A1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_804),
.A2(n_510),
.B(n_640),
.C(n_607),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_700),
.B(n_607),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_748),
.B(n_636),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_789),
.B(n_799),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_799),
.B(n_609),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_800),
.Y(n_981)
);

INVx4_ASAP7_75t_L g982 ( 
.A(n_807),
.Y(n_982)
);

O2A1O1Ixp5_ASAP7_75t_L g983 ( 
.A1(n_713),
.A2(n_774),
.B(n_762),
.C(n_800),
.Y(n_983)
);

A2O1A1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_818),
.A2(n_510),
.B(n_609),
.C(n_627),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_743),
.Y(n_985)
);

OAI21xp5_ASAP7_75t_L g986 ( 
.A1(n_749),
.A2(n_622),
.B(n_611),
.Y(n_986)
);

O2A1O1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_752),
.A2(n_844),
.B(n_821),
.C(n_731),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_734),
.A2(n_672),
.B(n_636),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_703),
.B(n_796),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_760),
.B(n_611),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_827),
.B(n_636),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_796),
.B(n_622),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_747),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_722),
.B(n_510),
.Y(n_994)
);

A2O1A1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_819),
.A2(n_482),
.B(n_477),
.C(n_500),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_739),
.A2(n_672),
.B(n_636),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_745),
.A2(n_672),
.B(n_636),
.Y(n_997)
);

NOR2xp67_ASAP7_75t_L g998 ( 
.A(n_699),
.B(n_75),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_759),
.B(n_672),
.Y(n_999)
);

NAND2x1p5_ASAP7_75t_L g1000 ( 
.A(n_811),
.B(n_470),
.Y(n_1000)
);

INVx3_ASAP7_75t_L g1001 ( 
.A(n_829),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_722),
.B(n_500),
.Y(n_1002)
);

OR2x6_ASAP7_75t_L g1003 ( 
.A(n_758),
.B(n_680),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_822),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_822),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_753),
.A2(n_451),
.B(n_499),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_756),
.A2(n_451),
.B(n_499),
.Y(n_1007)
);

HB1xp67_ASAP7_75t_L g1008 ( 
.A(n_847),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_781),
.B(n_500),
.Y(n_1009)
);

INVx2_ASAP7_75t_SL g1010 ( 
.A(n_690),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_801),
.B(n_505),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_831),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_808),
.B(n_505),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_757),
.A2(n_451),
.B(n_499),
.Y(n_1014)
);

O2A1O1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_846),
.A2(n_505),
.B(n_470),
.C(n_483),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_766),
.A2(n_451),
.B(n_486),
.Y(n_1016)
);

AOI21x1_ASAP7_75t_L g1017 ( 
.A1(n_713),
.A2(n_489),
.B(n_470),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_691),
.B(n_775),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_769),
.A2(n_489),
.B(n_470),
.Y(n_1019)
);

AOI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_775),
.A2(n_291),
.B1(n_507),
.B2(n_506),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_810),
.B(n_489),
.Y(n_1021)
);

INVx4_ASAP7_75t_L g1022 ( 
.A(n_807),
.Y(n_1022)
);

O2A1O1Ixp5_ASAP7_75t_L g1023 ( 
.A1(n_805),
.A2(n_489),
.B(n_470),
.C(n_483),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_SL g1024 ( 
.A(n_758),
.B(n_291),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_831),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_805),
.B(n_493),
.Y(n_1026)
);

NOR2xp67_ASAP7_75t_L g1027 ( 
.A(n_735),
.B(n_128),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_832),
.B(n_493),
.Y(n_1028)
);

HB1xp67_ASAP7_75t_L g1029 ( 
.A(n_841),
.Y(n_1029)
);

HB1xp67_ASAP7_75t_L g1030 ( 
.A(n_841),
.Y(n_1030)
);

O2A1O1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_705),
.A2(n_493),
.B(n_489),
.C(n_486),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_816),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_832),
.B(n_493),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_840),
.Y(n_1034)
);

AND2x2_ASAP7_75t_SL g1035 ( 
.A(n_819),
.B(n_742),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_772),
.A2(n_483),
.B(n_486),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_780),
.A2(n_483),
.B(n_486),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_840),
.B(n_493),
.Y(n_1038)
);

A2O1A1Ixp33_ASAP7_75t_L g1039 ( 
.A1(n_750),
.A2(n_791),
.B(n_833),
.C(n_677),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_815),
.B(n_486),
.Y(n_1040)
);

O2A1O1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_972),
.A2(n_751),
.B(n_738),
.C(n_720),
.Y(n_1041)
);

NOR2xp33_ASAP7_75t_L g1042 ( 
.A(n_942),
.B(n_750),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_851),
.B(n_825),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_871),
.Y(n_1044)
);

O2A1O1Ixp33_ASAP7_75t_L g1045 ( 
.A1(n_972),
.A2(n_848),
.B(n_843),
.C(n_839),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_SL g1046 ( 
.A(n_878),
.B(n_761),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_867),
.B(n_712),
.Y(n_1047)
);

INVx2_ASAP7_75t_SL g1048 ( 
.A(n_897),
.Y(n_1048)
);

AOI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_1018),
.A2(n_784),
.B1(n_816),
.B2(n_848),
.Y(n_1049)
);

BUFx8_ASAP7_75t_L g1050 ( 
.A(n_921),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_871),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_900),
.B(n_918),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_918),
.B(n_710),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_927),
.B(n_834),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_900),
.B(n_741),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_SL g1056 ( 
.A(n_989),
.B(n_710),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_958),
.B(n_678),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_854),
.A2(n_816),
.B(n_767),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_945),
.Y(n_1059)
);

CKINVDCx20_ASAP7_75t_R g1060 ( 
.A(n_864),
.Y(n_1060)
);

INVx6_ASAP7_75t_L g1061 ( 
.A(n_1003),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_873),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_994),
.B(n_784),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_920),
.B(n_784),
.Y(n_1064)
);

INVx2_ASAP7_75t_SL g1065 ( 
.A(n_965),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_901),
.B(n_784),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_934),
.B(n_678),
.Y(n_1067)
);

BUFx6f_ASAP7_75t_L g1068 ( 
.A(n_904),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_1018),
.A2(n_483),
.B(n_678),
.C(n_507),
.Y(n_1069)
);

BUFx2_ASAP7_75t_L g1070 ( 
.A(n_1029),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_1035),
.A2(n_508),
.B1(n_507),
.B2(n_506),
.Y(n_1071)
);

O2A1O1Ixp5_ASAP7_75t_SL g1072 ( 
.A1(n_862),
.A2(n_8),
.B(n_9),
.C(n_10),
.Y(n_1072)
);

AOI221xp5_ASAP7_75t_L g1073 ( 
.A1(n_852),
.A2(n_508),
.B1(n_507),
.B2(n_506),
.C(n_15),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_945),
.Y(n_1074)
);

BUFx2_ASAP7_75t_L g1075 ( 
.A(n_1029),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_1035),
.A2(n_508),
.B1(n_507),
.B2(n_506),
.Y(n_1076)
);

BUFx12f_ASAP7_75t_L g1077 ( 
.A(n_1010),
.Y(n_1077)
);

OAI21xp33_ASAP7_75t_SL g1078 ( 
.A1(n_903),
.A2(n_906),
.B(n_970),
.Y(n_1078)
);

AO32x1_ASAP7_75t_L g1079 ( 
.A1(n_916),
.A2(n_917),
.A3(n_874),
.B1(n_875),
.B2(n_881),
.Y(n_1079)
);

OR2x6_ASAP7_75t_SL g1080 ( 
.A(n_937),
.B(n_8),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_877),
.A2(n_492),
.B(n_471),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_873),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_880),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_860),
.A2(n_492),
.B(n_471),
.Y(n_1084)
);

BUFx2_ASAP7_75t_L g1085 ( 
.A(n_1030),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_880),
.Y(n_1086)
);

INVx5_ASAP7_75t_L g1087 ( 
.A(n_1032),
.Y(n_1087)
);

AOI21xp5_ASAP7_75t_L g1088 ( 
.A1(n_858),
.A2(n_492),
.B(n_471),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_SL g1089 ( 
.A(n_958),
.B(n_508),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_973),
.Y(n_1090)
);

AOI21x1_ASAP7_75t_L g1091 ( 
.A1(n_909),
.A2(n_492),
.B(n_471),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_968),
.B(n_508),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_885),
.A2(n_492),
.B(n_471),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_977),
.B(n_508),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_902),
.A2(n_507),
.B1(n_506),
.B2(n_508),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_863),
.A2(n_492),
.B(n_471),
.Y(n_1096)
);

NOR3xp33_ASAP7_75t_SL g1097 ( 
.A(n_857),
.B(n_9),
.C(n_11),
.Y(n_1097)
);

O2A1O1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_914),
.A2(n_17),
.B(n_18),
.C(n_19),
.Y(n_1098)
);

OAI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_902),
.A2(n_507),
.B1(n_506),
.B2(n_508),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_962),
.B(n_507),
.Y(n_1100)
);

INVx6_ASAP7_75t_L g1101 ( 
.A(n_1003),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_977),
.B(n_506),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_889),
.B(n_492),
.Y(n_1103)
);

NOR2xp67_ASAP7_75t_L g1104 ( 
.A(n_1030),
.B(n_170),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_1003),
.Y(n_1105)
);

BUFx2_ASAP7_75t_L g1106 ( 
.A(n_904),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_886),
.Y(n_1107)
);

AO32x1_ASAP7_75t_L g1108 ( 
.A1(n_884),
.A2(n_18),
.A3(n_20),
.B1(n_21),
.B2(n_23),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_SL g1109 ( 
.A(n_872),
.B(n_156),
.Y(n_1109)
);

BUFx6f_ASAP7_75t_L g1110 ( 
.A(n_907),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1002),
.B(n_492),
.Y(n_1111)
);

OAI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_1039),
.A2(n_471),
.B1(n_25),
.B2(n_27),
.Y(n_1112)
);

OR2x2_ASAP7_75t_L g1113 ( 
.A(n_934),
.B(n_24),
.Y(n_1113)
);

INVxp67_ASAP7_75t_L g1114 ( 
.A(n_922),
.Y(n_1114)
);

NAND3xp33_ASAP7_75t_L g1115 ( 
.A(n_922),
.B(n_471),
.C(n_27),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_960),
.A2(n_151),
.B(n_147),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_973),
.B(n_146),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_850),
.B(n_25),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_974),
.B(n_141),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_974),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_868),
.A2(n_136),
.B(n_132),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_869),
.A2(n_125),
.B(n_106),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_1039),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_886),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_907),
.B(n_29),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_850),
.B(n_33),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_890),
.Y(n_1127)
);

BUFx2_ASAP7_75t_L g1128 ( 
.A(n_1008),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_908),
.B(n_34),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_890),
.Y(n_1130)
);

OA22x2_ASAP7_75t_L g1131 ( 
.A1(n_1008),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_956),
.B(n_44),
.Y(n_1132)
);

CKINVDCx16_ASAP7_75t_R g1133 ( 
.A(n_947),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_870),
.B(n_45),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_926),
.Y(n_1135)
);

INVx2_ASAP7_75t_SL g1136 ( 
.A(n_919),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_926),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_876),
.A2(n_98),
.B(n_96),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_872),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_SL g1140 ( 
.A(n_963),
.B(n_92),
.Y(n_1140)
);

O2A1O1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_855),
.A2(n_47),
.B(n_48),
.C(n_50),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_1032),
.Y(n_1142)
);

BUFx2_ASAP7_75t_L g1143 ( 
.A(n_919),
.Y(n_1143)
);

AOI22x1_ASAP7_75t_L g1144 ( 
.A1(n_928),
.A2(n_85),
.B1(n_84),
.B2(n_83),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_870),
.B(n_50),
.Y(n_1145)
);

OAI22xp5_ASAP7_75t_L g1146 ( 
.A1(n_882),
.A2(n_58),
.B1(n_59),
.B2(n_61),
.Y(n_1146)
);

AO32x1_ASAP7_75t_L g1147 ( 
.A1(n_895),
.A2(n_58),
.A3(n_63),
.B1(n_64),
.B2(n_66),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_892),
.A2(n_81),
.B(n_82),
.Y(n_1148)
);

BUFx2_ASAP7_75t_L g1149 ( 
.A(n_908),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_928),
.Y(n_1150)
);

AOI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_1027),
.A2(n_63),
.B1(n_66),
.B2(n_978),
.Y(n_1151)
);

HB1xp67_ASAP7_75t_L g1152 ( 
.A(n_985),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_882),
.A2(n_898),
.B1(n_888),
.B2(n_903),
.Y(n_1153)
);

NOR3xp33_ASAP7_75t_L g1154 ( 
.A(n_912),
.B(n_990),
.C(n_987),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_924),
.A2(n_1026),
.B(n_931),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_896),
.B(n_930),
.Y(n_1156)
);

INVx5_ASAP7_75t_L g1157 ( 
.A(n_1032),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_990),
.B(n_993),
.Y(n_1158)
);

INVx2_ASAP7_75t_SL g1159 ( 
.A(n_978),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_866),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_905),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_893),
.A2(n_913),
.B(n_883),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1034),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_1034),
.Y(n_1164)
);

AOI22x1_ASAP7_75t_L g1165 ( 
.A1(n_950),
.A2(n_910),
.B1(n_948),
.B2(n_946),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_L g1166 ( 
.A(n_1001),
.B(n_856),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_898),
.A2(n_906),
.B1(n_912),
.B2(n_855),
.Y(n_1167)
);

AOI22x1_ASAP7_75t_L g1168 ( 
.A1(n_923),
.A2(n_940),
.B1(n_935),
.B2(n_981),
.Y(n_1168)
);

BUFx3_ASAP7_75t_L g1169 ( 
.A(n_1032),
.Y(n_1169)
);

NOR2x1_ASAP7_75t_L g1170 ( 
.A(n_891),
.B(n_998),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_1001),
.B(n_932),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_929),
.A2(n_933),
.B(n_909),
.Y(n_1172)
);

NOR2xp67_ASAP7_75t_SL g1173 ( 
.A(n_955),
.B(n_932),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_SL g1174 ( 
.A1(n_911),
.A2(n_891),
.B1(n_879),
.B2(n_954),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_979),
.A2(n_861),
.B(n_899),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1013),
.B(n_1009),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_911),
.B(n_975),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1011),
.B(n_941),
.Y(n_1178)
);

AND2x4_ASAP7_75t_L g1179 ( 
.A(n_954),
.B(n_982),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_975),
.B(n_944),
.Y(n_1180)
);

O2A1O1Ixp33_ASAP7_75t_L g1181 ( 
.A1(n_862),
.A2(n_859),
.B(n_976),
.C(n_992),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_SL g1182 ( 
.A(n_955),
.B(n_1024),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_952),
.B(n_953),
.Y(n_1183)
);

OA22x2_ASAP7_75t_L g1184 ( 
.A1(n_957),
.A2(n_991),
.B1(n_1005),
.B2(n_1025),
.Y(n_1184)
);

CKINVDCx8_ASAP7_75t_R g1185 ( 
.A(n_915),
.Y(n_1185)
);

BUFx8_ASAP7_75t_L g1186 ( 
.A(n_915),
.Y(n_1186)
);

A2O1A1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_853),
.A2(n_983),
.B(n_951),
.C(n_1023),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_915),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1004),
.B(n_1012),
.Y(n_1189)
);

BUFx3_ASAP7_75t_L g1190 ( 
.A(n_915),
.Y(n_1190)
);

HB1xp67_ASAP7_75t_L g1191 ( 
.A(n_999),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_969),
.A2(n_887),
.B(n_997),
.Y(n_1192)
);

AOI21x1_ASAP7_75t_L g1193 ( 
.A1(n_849),
.A2(n_991),
.B(n_1017),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_SL g1194 ( 
.A(n_955),
.B(n_982),
.Y(n_1194)
);

AOI21xp33_ASAP7_75t_L g1195 ( 
.A1(n_959),
.A2(n_925),
.B(n_1040),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_988),
.A2(n_996),
.B(n_1021),
.Y(n_1196)
);

AOI21x1_ASAP7_75t_L g1197 ( 
.A1(n_964),
.A2(n_971),
.B(n_966),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_865),
.A2(n_980),
.B(n_955),
.Y(n_1198)
);

O2A1O1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_859),
.A2(n_976),
.B(n_995),
.C(n_938),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_984),
.A2(n_995),
.B1(n_1000),
.B2(n_1022),
.Y(n_1200)
);

OAI22x1_ASAP7_75t_L g1201 ( 
.A1(n_1052),
.A2(n_1020),
.B1(n_1000),
.B2(n_1022),
.Y(n_1201)
);

HB1xp67_ASAP7_75t_L g1202 ( 
.A(n_1065),
.Y(n_1202)
);

OAI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1046),
.A2(n_894),
.B(n_1037),
.Y(n_1203)
);

A2O1A1Ixp33_ASAP7_75t_L g1204 ( 
.A1(n_1042),
.A2(n_1031),
.B(n_1015),
.C(n_1036),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1158),
.B(n_984),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_L g1206 ( 
.A1(n_1162),
.A2(n_986),
.B(n_961),
.Y(n_1206)
);

OAI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1078),
.A2(n_1019),
.B(n_1016),
.Y(n_1207)
);

O2A1O1Ixp33_ASAP7_75t_SL g1208 ( 
.A1(n_1123),
.A2(n_1038),
.B(n_1033),
.C(n_1028),
.Y(n_1208)
);

OA21x2_ASAP7_75t_L g1209 ( 
.A1(n_1187),
.A2(n_1014),
.B(n_1007),
.Y(n_1209)
);

CKINVDCx11_ASAP7_75t_R g1210 ( 
.A(n_1060),
.Y(n_1210)
);

OA21x2_ASAP7_75t_L g1211 ( 
.A1(n_1175),
.A2(n_1006),
.B(n_949),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1114),
.B(n_915),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_SL g1213 ( 
.A(n_1047),
.B(n_967),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1043),
.B(n_1176),
.Y(n_1214)
);

AOI21xp33_ASAP7_75t_L g1215 ( 
.A1(n_1041),
.A2(n_936),
.B(n_939),
.Y(n_1215)
);

OAI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1154),
.A2(n_943),
.B(n_1176),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1043),
.B(n_1054),
.Y(n_1217)
);

INVx2_ASAP7_75t_SL g1218 ( 
.A(n_1050),
.Y(n_1218)
);

NAND2x1p5_ASAP7_75t_L g1219 ( 
.A(n_1087),
.B(n_1157),
.Y(n_1219)
);

HB1xp67_ASAP7_75t_L g1220 ( 
.A(n_1070),
.Y(n_1220)
);

AO32x2_ASAP7_75t_L g1221 ( 
.A1(n_1112),
.A2(n_1167),
.A3(n_1153),
.B1(n_1146),
.B2(n_1174),
.Y(n_1221)
);

BUFx6f_ASAP7_75t_L g1222 ( 
.A(n_1142),
.Y(n_1222)
);

AO31x2_ASAP7_75t_L g1223 ( 
.A1(n_1167),
.A2(n_1153),
.A3(n_1069),
.B(n_1200),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1163),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1054),
.B(n_1156),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1164),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1058),
.A2(n_1155),
.B(n_1198),
.Y(n_1227)
);

INVx2_ASAP7_75t_SL g1228 ( 
.A(n_1050),
.Y(n_1228)
);

O2A1O1Ixp33_ASAP7_75t_L g1229 ( 
.A1(n_1113),
.A2(n_1053),
.B(n_1112),
.C(n_1118),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1149),
.B(n_1129),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1161),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1156),
.A2(n_1172),
.B(n_1178),
.Y(n_1232)
);

AOI221xp5_ASAP7_75t_SL g1233 ( 
.A1(n_1132),
.A2(n_1098),
.B1(n_1055),
.B2(n_1126),
.C(n_1141),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_1133),
.Y(n_1234)
);

BUFx8_ASAP7_75t_L g1235 ( 
.A(n_1075),
.Y(n_1235)
);

AOI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1056),
.A2(n_1136),
.B1(n_1067),
.B2(n_1143),
.Y(n_1236)
);

BUFx2_ASAP7_75t_L g1237 ( 
.A(n_1085),
.Y(n_1237)
);

O2A1O1Ixp33_ASAP7_75t_SL g1238 ( 
.A1(n_1140),
.A2(n_1180),
.B(n_1057),
.C(n_1064),
.Y(n_1238)
);

A2O1A1Ixp33_ASAP7_75t_L g1239 ( 
.A1(n_1151),
.A2(n_1181),
.B(n_1177),
.C(n_1066),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1178),
.A2(n_1100),
.B(n_1183),
.Y(n_1240)
);

AO31x2_ASAP7_75t_L g1241 ( 
.A1(n_1200),
.A2(n_1071),
.A3(n_1076),
.B(n_1196),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1191),
.B(n_1152),
.Y(n_1242)
);

AND2x2_ASAP7_75t_SL g1243 ( 
.A(n_1109),
.B(n_1073),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1125),
.B(n_1128),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1044),
.Y(n_1245)
);

OR2x2_ASAP7_75t_L g1246 ( 
.A(n_1048),
.B(n_1106),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1094),
.A2(n_1102),
.B(n_1192),
.Y(n_1247)
);

CKINVDCx20_ASAP7_75t_R g1248 ( 
.A(n_1160),
.Y(n_1248)
);

O2A1O1Ixp33_ASAP7_75t_SL g1249 ( 
.A1(n_1063),
.A2(n_1119),
.B(n_1117),
.C(n_1182),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1051),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1094),
.A2(n_1102),
.B(n_1195),
.Y(n_1251)
);

AOI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1104),
.A2(n_1145),
.B1(n_1134),
.B2(n_1159),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1088),
.A2(n_1081),
.B(n_1096),
.Y(n_1253)
);

OAI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1193),
.A2(n_1084),
.B(n_1091),
.Y(n_1254)
);

OR2x2_ASAP7_75t_L g1255 ( 
.A(n_1068),
.B(n_1110),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1195),
.A2(n_1045),
.B(n_1063),
.Y(n_1256)
);

NAND3xp33_ASAP7_75t_L g1257 ( 
.A(n_1097),
.B(n_1115),
.C(n_1146),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1166),
.B(n_1189),
.Y(n_1258)
);

NOR4xp25_ASAP7_75t_L g1259 ( 
.A(n_1199),
.B(n_1080),
.C(n_1117),
.D(n_1119),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1111),
.A2(n_1103),
.B(n_1171),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1111),
.A2(n_1103),
.B(n_1049),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1109),
.A2(n_1184),
.B(n_1148),
.Y(n_1262)
);

NOR2xp67_ASAP7_75t_L g1263 ( 
.A(n_1077),
.B(n_1105),
.Y(n_1263)
);

NOR2xp67_ASAP7_75t_SL g1264 ( 
.A(n_1185),
.B(n_1157),
.Y(n_1264)
);

AO21x1_ASAP7_75t_L g1265 ( 
.A1(n_1121),
.A2(n_1071),
.B(n_1076),
.Y(n_1265)
);

INVx2_ASAP7_75t_SL g1266 ( 
.A(n_1061),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1184),
.A2(n_1179),
.B(n_1194),
.Y(n_1267)
);

BUFx6f_ASAP7_75t_L g1268 ( 
.A(n_1142),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_SL g1269 ( 
.A(n_1068),
.B(n_1110),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1062),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1093),
.A2(n_1165),
.B(n_1168),
.Y(n_1271)
);

INVxp67_ASAP7_75t_SL g1272 ( 
.A(n_1186),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1116),
.A2(n_1197),
.B(n_1138),
.Y(n_1273)
);

INVx3_ASAP7_75t_L g1274 ( 
.A(n_1179),
.Y(n_1274)
);

OAI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1170),
.A2(n_1092),
.B(n_1089),
.Y(n_1275)
);

NOR2xp67_ASAP7_75t_L g1276 ( 
.A(n_1087),
.B(n_1157),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1082),
.B(n_1107),
.Y(n_1277)
);

AO31x2_ASAP7_75t_L g1278 ( 
.A1(n_1095),
.A2(n_1099),
.A3(n_1079),
.B(n_1122),
.Y(n_1278)
);

BUFx12f_ASAP7_75t_L g1279 ( 
.A(n_1101),
.Y(n_1279)
);

INVx5_ASAP7_75t_L g1280 ( 
.A(n_1188),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1169),
.B(n_1087),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1095),
.A2(n_1099),
.B(n_1157),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_1083),
.B(n_1086),
.Y(n_1283)
);

AOI221xp5_ASAP7_75t_L g1284 ( 
.A1(n_1059),
.A2(n_1120),
.B1(n_1074),
.B2(n_1130),
.C(n_1150),
.Y(n_1284)
);

OA21x2_ASAP7_75t_L g1285 ( 
.A1(n_1090),
.A2(n_1135),
.B(n_1137),
.Y(n_1285)
);

A2O1A1Ixp33_ASAP7_75t_L g1286 ( 
.A1(n_1124),
.A2(n_1127),
.B(n_1190),
.C(n_1173),
.Y(n_1286)
);

AO31x2_ASAP7_75t_L g1287 ( 
.A1(n_1079),
.A2(n_1072),
.A3(n_1108),
.B(n_1147),
.Y(n_1287)
);

AOI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1131),
.A2(n_1079),
.B(n_1144),
.Y(n_1288)
);

AO31x2_ASAP7_75t_L g1289 ( 
.A1(n_1108),
.A2(n_1147),
.A3(n_1186),
.B(n_1188),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1087),
.A2(n_1139),
.B(n_1188),
.Y(n_1290)
);

O2A1O1Ixp33_ASAP7_75t_SL g1291 ( 
.A1(n_1147),
.A2(n_1018),
.B(n_1039),
.C(n_1123),
.Y(n_1291)
);

CKINVDCx6p67_ASAP7_75t_R g1292 ( 
.A(n_1060),
.Y(n_1292)
);

INVx3_ASAP7_75t_L g1293 ( 
.A(n_1179),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1058),
.A2(n_854),
.B(n_851),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1162),
.A2(n_1088),
.B(n_1081),
.Y(n_1295)
);

BUFx5_ASAP7_75t_L g1296 ( 
.A(n_1190),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1161),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1042),
.A2(n_851),
.B1(n_867),
.B2(n_972),
.Y(n_1298)
);

CKINVDCx6p67_ASAP7_75t_R g1299 ( 
.A(n_1060),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_1060),
.Y(n_1300)
);

O2A1O1Ixp33_ASAP7_75t_L g1301 ( 
.A1(n_1052),
.A2(n_694),
.B(n_733),
.C(n_942),
.Y(n_1301)
);

OR2x6_ASAP7_75t_L g1302 ( 
.A(n_1065),
.B(n_1048),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1162),
.A2(n_1088),
.B(n_1081),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1058),
.A2(n_854),
.B(n_851),
.Y(n_1304)
);

NOR2x1_ASAP7_75t_R g1305 ( 
.A(n_1077),
.B(n_717),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1058),
.A2(n_854),
.B(n_851),
.Y(n_1306)
);

BUFx8_ASAP7_75t_SL g1307 ( 
.A(n_1060),
.Y(n_1307)
);

INVx3_ASAP7_75t_L g1308 ( 
.A(n_1179),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1058),
.A2(n_854),
.B(n_851),
.Y(n_1309)
);

NAND3xp33_ASAP7_75t_L g1310 ( 
.A(n_1052),
.B(n_972),
.C(n_942),
.Y(n_1310)
);

AO31x2_ASAP7_75t_L g1311 ( 
.A1(n_1187),
.A2(n_1167),
.A3(n_1153),
.B(n_1069),
.Y(n_1311)
);

BUFx6f_ASAP7_75t_L g1312 ( 
.A(n_1142),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1058),
.A2(n_854),
.B(n_851),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_1065),
.Y(n_1314)
);

INVx2_ASAP7_75t_L g1315 ( 
.A(n_1044),
.Y(n_1315)
);

OAI21xp33_ASAP7_75t_L g1316 ( 
.A1(n_1052),
.A2(n_942),
.B(n_900),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1058),
.A2(n_854),
.B(n_851),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1058),
.A2(n_854),
.B(n_851),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_SL g1319 ( 
.A(n_1114),
.B(n_942),
.Y(n_1319)
);

A2O1A1Ixp33_ASAP7_75t_L g1320 ( 
.A1(n_1052),
.A2(n_972),
.B(n_942),
.C(n_851),
.Y(n_1320)
);

O2A1O1Ixp33_ASAP7_75t_L g1321 ( 
.A1(n_1052),
.A2(n_694),
.B(n_733),
.C(n_942),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1058),
.A2(n_854),
.B(n_851),
.Y(n_1322)
);

O2A1O1Ixp33_ASAP7_75t_SL g1323 ( 
.A1(n_1123),
.A2(n_1018),
.B(n_1039),
.C(n_693),
.Y(n_1323)
);

O2A1O1Ixp33_ASAP7_75t_L g1324 ( 
.A1(n_1052),
.A2(n_694),
.B(n_733),
.C(n_942),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1161),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1058),
.A2(n_854),
.B(n_851),
.Y(n_1326)
);

AO31x2_ASAP7_75t_L g1327 ( 
.A1(n_1187),
.A2(n_1167),
.A3(n_1153),
.B(n_1069),
.Y(n_1327)
);

O2A1O1Ixp33_ASAP7_75t_SL g1328 ( 
.A1(n_1123),
.A2(n_1018),
.B(n_1039),
.C(n_693),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_L g1329 ( 
.A(n_1052),
.B(n_851),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1162),
.A2(n_1088),
.B(n_1081),
.Y(n_1330)
);

NAND2xp5_ASAP7_75t_L g1331 ( 
.A(n_1052),
.B(n_851),
.Y(n_1331)
);

AOI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1198),
.A2(n_862),
.B(n_877),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1161),
.Y(n_1333)
);

INVxp67_ASAP7_75t_L g1334 ( 
.A(n_1065),
.Y(n_1334)
);

A2O1A1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1052),
.A2(n_972),
.B(n_942),
.C(n_851),
.Y(n_1335)
);

AO32x2_ASAP7_75t_L g1336 ( 
.A1(n_1112),
.A2(n_1167),
.A3(n_1153),
.B1(n_1146),
.B2(n_916),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1058),
.A2(n_854),
.B(n_851),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1052),
.B(n_694),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1162),
.A2(n_1088),
.B(n_1081),
.Y(n_1339)
);

OR2x2_ASAP7_75t_L g1340 ( 
.A(n_1065),
.B(n_686),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1052),
.B(n_851),
.Y(n_1341)
);

NAND2xp5_ASAP7_75t_L g1342 ( 
.A(n_1052),
.B(n_851),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_L g1343 ( 
.A(n_1052),
.B(n_694),
.Y(n_1343)
);

BUFx10_ASAP7_75t_L g1344 ( 
.A(n_1047),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1065),
.Y(n_1345)
);

INVxp67_ASAP7_75t_L g1346 ( 
.A(n_1065),
.Y(n_1346)
);

OAI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1046),
.A2(n_972),
.B(n_878),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1058),
.A2(n_854),
.B(n_851),
.Y(n_1348)
);

BUFx12f_ASAP7_75t_L g1349 ( 
.A(n_1077),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1058),
.A2(n_854),
.B(n_851),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_1052),
.B(n_851),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1162),
.A2(n_1088),
.B(n_1081),
.Y(n_1352)
);

AND2x4_ASAP7_75t_L g1353 ( 
.A(n_1068),
.B(n_904),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1042),
.A2(n_851),
.B1(n_867),
.B2(n_972),
.Y(n_1354)
);

NAND3xp33_ASAP7_75t_SL g1355 ( 
.A(n_1052),
.B(n_942),
.C(n_717),
.Y(n_1355)
);

AND2x4_ASAP7_75t_L g1356 ( 
.A(n_1068),
.B(n_904),
.Y(n_1356)
);

BUFx6f_ASAP7_75t_L g1357 ( 
.A(n_1142),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1052),
.B(n_851),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1058),
.A2(n_854),
.B(n_851),
.Y(n_1359)
);

OAI22xp33_ASAP7_75t_SL g1360 ( 
.A1(n_1329),
.A2(n_1341),
.B1(n_1331),
.B2(n_1358),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1310),
.A2(n_1243),
.B1(n_1316),
.B2(n_1257),
.Y(n_1361)
);

BUFx10_ASAP7_75t_L g1362 ( 
.A(n_1300),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1342),
.B(n_1351),
.Y(n_1363)
);

CKINVDCx20_ASAP7_75t_R g1364 ( 
.A(n_1307),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1298),
.A2(n_1354),
.B1(n_1347),
.B2(n_1338),
.Y(n_1365)
);

CKINVDCx11_ASAP7_75t_R g1366 ( 
.A(n_1292),
.Y(n_1366)
);

INVx6_ASAP7_75t_L g1367 ( 
.A(n_1235),
.Y(n_1367)
);

OAI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1214),
.A2(n_1343),
.B1(n_1225),
.B2(n_1217),
.Y(n_1368)
);

CKINVDCx6p67_ASAP7_75t_R g1369 ( 
.A(n_1299),
.Y(n_1369)
);

OAI21xp33_ASAP7_75t_L g1370 ( 
.A1(n_1320),
.A2(n_1335),
.B(n_1259),
.Y(n_1370)
);

BUFx4f_ASAP7_75t_SL g1371 ( 
.A(n_1248),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_1234),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1355),
.A2(n_1265),
.B1(n_1319),
.B2(n_1252),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1213),
.A2(n_1216),
.B1(n_1258),
.B2(n_1344),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1205),
.A2(n_1240),
.B1(n_1262),
.B2(n_1333),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1297),
.A2(n_1325),
.B1(n_1256),
.B2(n_1220),
.Y(n_1376)
);

BUFx8_ASAP7_75t_L g1377 ( 
.A(n_1349),
.Y(n_1377)
);

INVx6_ASAP7_75t_L g1378 ( 
.A(n_1235),
.Y(n_1378)
);

BUFx4_ASAP7_75t_SL g1379 ( 
.A(n_1302),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1237),
.A2(n_1236),
.B1(n_1232),
.B2(n_1242),
.Y(n_1380)
);

OAI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1301),
.A2(n_1321),
.B1(n_1324),
.B2(n_1340),
.Y(n_1381)
);

INVx2_ASAP7_75t_SL g1382 ( 
.A(n_1302),
.Y(n_1382)
);

BUFx3_ASAP7_75t_L g1383 ( 
.A(n_1279),
.Y(n_1383)
);

INVx4_ASAP7_75t_L g1384 ( 
.A(n_1280),
.Y(n_1384)
);

INVx1_ASAP7_75t_SL g1385 ( 
.A(n_1246),
.Y(n_1385)
);

INVx6_ASAP7_75t_L g1386 ( 
.A(n_1280),
.Y(n_1386)
);

OAI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1221),
.A2(n_1282),
.B1(n_1212),
.B2(n_1272),
.Y(n_1387)
);

BUFx2_ASAP7_75t_SL g1388 ( 
.A(n_1263),
.Y(n_1388)
);

OAI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1229),
.A2(n_1233),
.B(n_1239),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1230),
.A2(n_1224),
.B1(n_1226),
.B2(n_1270),
.Y(n_1390)
);

BUFx8_ASAP7_75t_L g1391 ( 
.A(n_1218),
.Y(n_1391)
);

CKINVDCx20_ASAP7_75t_R g1392 ( 
.A(n_1202),
.Y(n_1392)
);

BUFx12f_ASAP7_75t_L g1393 ( 
.A(n_1255),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1226),
.A2(n_1245),
.B1(n_1270),
.B2(n_1250),
.Y(n_1394)
);

CKINVDCx6p67_ASAP7_75t_R g1395 ( 
.A(n_1280),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1285),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1245),
.A2(n_1250),
.B1(n_1315),
.B2(n_1221),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_SL g1398 ( 
.A1(n_1221),
.A2(n_1336),
.B1(n_1345),
.B2(n_1314),
.Y(n_1398)
);

INVx4_ASAP7_75t_L g1399 ( 
.A(n_1281),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1283),
.A2(n_1336),
.B1(n_1284),
.B2(n_1251),
.Y(n_1400)
);

INVx8_ASAP7_75t_L g1401 ( 
.A(n_1281),
.Y(n_1401)
);

INVx4_ASAP7_75t_L g1402 ( 
.A(n_1219),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1285),
.Y(n_1403)
);

INVx2_ASAP7_75t_SL g1404 ( 
.A(n_1266),
.Y(n_1404)
);

CKINVDCx20_ASAP7_75t_R g1405 ( 
.A(n_1334),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1277),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1269),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1336),
.A2(n_1201),
.B1(n_1261),
.B2(n_1207),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_1228),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1222),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_L g1411 ( 
.A1(n_1267),
.A2(n_1260),
.B1(n_1356),
.B2(n_1353),
.Y(n_1411)
);

INVx11_ASAP7_75t_L g1412 ( 
.A(n_1305),
.Y(n_1412)
);

BUFx10_ASAP7_75t_L g1413 ( 
.A(n_1356),
.Y(n_1413)
);

INVx6_ASAP7_75t_L g1414 ( 
.A(n_1268),
.Y(n_1414)
);

AOI22xp5_ASAP7_75t_L g1415 ( 
.A1(n_1346),
.A2(n_1328),
.B1(n_1323),
.B2(n_1308),
.Y(n_1415)
);

OAI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1286),
.A2(n_1293),
.B1(n_1308),
.B2(n_1274),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1293),
.A2(n_1247),
.B1(n_1275),
.B2(n_1203),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1268),
.B(n_1357),
.Y(n_1418)
);

NAND2x1p5_ASAP7_75t_L g1419 ( 
.A(n_1264),
.B(n_1276),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1294),
.A2(n_1359),
.B1(n_1309),
.B2(n_1306),
.Y(n_1420)
);

BUFx3_ASAP7_75t_L g1421 ( 
.A(n_1312),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_L g1422 ( 
.A1(n_1304),
.A2(n_1322),
.B1(n_1318),
.B2(n_1350),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1204),
.A2(n_1348),
.B1(n_1337),
.B2(n_1326),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_L g1424 ( 
.A1(n_1313),
.A2(n_1317),
.B1(n_1215),
.B2(n_1209),
.Y(n_1424)
);

INVx2_ASAP7_75t_L g1425 ( 
.A(n_1296),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1311),
.Y(n_1426)
);

BUFx2_ASAP7_75t_L g1427 ( 
.A(n_1296),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1311),
.Y(n_1428)
);

INVx8_ASAP7_75t_L g1429 ( 
.A(n_1290),
.Y(n_1429)
);

CKINVDCx6p67_ASAP7_75t_R g1430 ( 
.A(n_1238),
.Y(n_1430)
);

BUFx4f_ASAP7_75t_SL g1431 ( 
.A(n_1249),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_SL g1432 ( 
.A1(n_1291),
.A2(n_1223),
.B1(n_1271),
.B2(n_1227),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1327),
.B(n_1223),
.Y(n_1433)
);

INVx4_ASAP7_75t_L g1434 ( 
.A(n_1211),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1211),
.A2(n_1206),
.B1(n_1223),
.B2(n_1253),
.Y(n_1435)
);

BUFx2_ASAP7_75t_SL g1436 ( 
.A(n_1208),
.Y(n_1436)
);

BUFx2_ASAP7_75t_L g1437 ( 
.A(n_1327),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1288),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1295),
.A2(n_1303),
.B1(n_1339),
.B2(n_1330),
.Y(n_1439)
);

INVx4_ASAP7_75t_L g1440 ( 
.A(n_1332),
.Y(n_1440)
);

CKINVDCx20_ASAP7_75t_R g1441 ( 
.A(n_1241),
.Y(n_1441)
);

BUFx4_ASAP7_75t_R g1442 ( 
.A(n_1241),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1289),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1254),
.Y(n_1444)
);

CKINVDCx11_ASAP7_75t_R g1445 ( 
.A(n_1241),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1352),
.A2(n_1273),
.B1(n_1289),
.B2(n_1287),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1289),
.A2(n_972),
.B1(n_1310),
.B2(n_1052),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1287),
.A2(n_972),
.B1(n_1310),
.B2(n_1052),
.Y(n_1448)
);

INVx2_ASAP7_75t_SL g1449 ( 
.A(n_1278),
.Y(n_1449)
);

INVx8_ASAP7_75t_L g1450 ( 
.A(n_1278),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1242),
.B(n_1340),
.Y(n_1451)
);

INVx6_ASAP7_75t_L g1452 ( 
.A(n_1235),
.Y(n_1452)
);

CKINVDCx11_ASAP7_75t_R g1453 ( 
.A(n_1210),
.Y(n_1453)
);

INVx1_ASAP7_75t_SL g1454 ( 
.A(n_1237),
.Y(n_1454)
);

INVx8_ASAP7_75t_L g1455 ( 
.A(n_1280),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1310),
.A2(n_972),
.B1(n_1052),
.B2(n_1243),
.Y(n_1456)
);

INVx2_ASAP7_75t_SL g1457 ( 
.A(n_1235),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_SL g1458 ( 
.A1(n_1243),
.A2(n_942),
.B1(n_771),
.B2(n_1052),
.Y(n_1458)
);

INVx8_ASAP7_75t_L g1459 ( 
.A(n_1280),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1310),
.A2(n_972),
.B1(n_1052),
.B2(n_1243),
.Y(n_1460)
);

CKINVDCx11_ASAP7_75t_R g1461 ( 
.A(n_1210),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1338),
.A2(n_1343),
.B1(n_1310),
.B2(n_1331),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_SL g1463 ( 
.A1(n_1243),
.A2(n_942),
.B1(n_771),
.B2(n_1052),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1310),
.A2(n_972),
.B1(n_1052),
.B2(n_1243),
.Y(n_1464)
);

BUFx8_ASAP7_75t_L g1465 ( 
.A(n_1349),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_SL g1466 ( 
.A1(n_1243),
.A2(n_942),
.B1(n_771),
.B2(n_1052),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_L g1467 ( 
.A1(n_1310),
.A2(n_972),
.B1(n_1052),
.B2(n_1243),
.Y(n_1467)
);

BUFx12f_ASAP7_75t_L g1468 ( 
.A(n_1210),
.Y(n_1468)
);

OAI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1310),
.A2(n_1329),
.B1(n_1341),
.B2(n_1331),
.Y(n_1469)
);

AOI22xp33_ASAP7_75t_L g1470 ( 
.A1(n_1310),
.A2(n_972),
.B1(n_1052),
.B2(n_1243),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1329),
.B(n_1331),
.Y(n_1471)
);

INVxp33_ASAP7_75t_L g1472 ( 
.A(n_1244),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1310),
.A2(n_972),
.B1(n_1052),
.B2(n_1243),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1310),
.A2(n_972),
.B1(n_1052),
.B2(n_1243),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1310),
.A2(n_972),
.B1(n_1052),
.B2(n_1243),
.Y(n_1475)
);

INVx3_ASAP7_75t_L g1476 ( 
.A(n_1274),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1230),
.B(n_1244),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1310),
.A2(n_972),
.B1(n_1052),
.B2(n_1243),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1231),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1231),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1310),
.A2(n_972),
.B1(n_1052),
.B2(n_1243),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1230),
.B(n_1244),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1363),
.B(n_1471),
.Y(n_1483)
);

AND2x2_ASAP7_75t_L g1484 ( 
.A(n_1437),
.B(n_1433),
.Y(n_1484)
);

BUFx2_ASAP7_75t_L g1485 ( 
.A(n_1443),
.Y(n_1485)
);

BUFx2_ASAP7_75t_L g1486 ( 
.A(n_1426),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1458),
.A2(n_1463),
.B1(n_1466),
.B2(n_1481),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1441),
.B(n_1428),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1385),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1368),
.B(n_1469),
.Y(n_1490)
);

INVx5_ASAP7_75t_L g1491 ( 
.A(n_1434),
.Y(n_1491)
);

HB1xp67_ASAP7_75t_L g1492 ( 
.A(n_1451),
.Y(n_1492)
);

OAI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1462),
.A2(n_1389),
.B1(n_1381),
.B2(n_1431),
.Y(n_1493)
);

INVx5_ASAP7_75t_L g1494 ( 
.A(n_1434),
.Y(n_1494)
);

OAI21xp5_ASAP7_75t_L g1495 ( 
.A1(n_1456),
.A2(n_1464),
.B(n_1460),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1396),
.Y(n_1496)
);

HB1xp67_ASAP7_75t_L g1497 ( 
.A(n_1407),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1403),
.Y(n_1498)
);

INVx3_ASAP7_75t_L g1499 ( 
.A(n_1440),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1398),
.B(n_1447),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1447),
.B(n_1445),
.Y(n_1501)
);

INVx2_ASAP7_75t_SL g1502 ( 
.A(n_1386),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1448),
.B(n_1438),
.Y(n_1503)
);

BUFx2_ASAP7_75t_L g1504 ( 
.A(n_1427),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1449),
.Y(n_1505)
);

OAI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1439),
.A2(n_1423),
.B(n_1424),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1408),
.B(n_1450),
.Y(n_1507)
);

OA21x2_ASAP7_75t_L g1508 ( 
.A1(n_1424),
.A2(n_1420),
.B(n_1422),
.Y(n_1508)
);

INVx3_ASAP7_75t_L g1509 ( 
.A(n_1440),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1442),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1444),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1442),
.Y(n_1512)
);

NOR2x1_ASAP7_75t_L g1513 ( 
.A(n_1368),
.B(n_1469),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1360),
.B(n_1456),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1408),
.B(n_1448),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1387),
.B(n_1376),
.Y(n_1516)
);

OR2x6_ASAP7_75t_L g1517 ( 
.A(n_1436),
.B(n_1429),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1387),
.B(n_1376),
.Y(n_1518)
);

OAI21x1_ASAP7_75t_L g1519 ( 
.A1(n_1439),
.A2(n_1422),
.B(n_1420),
.Y(n_1519)
);

OA21x2_ASAP7_75t_L g1520 ( 
.A1(n_1446),
.A2(n_1370),
.B(n_1435),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1479),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1480),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1397),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1397),
.B(n_1375),
.Y(n_1524)
);

INVx2_ASAP7_75t_SL g1525 ( 
.A(n_1386),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1446),
.Y(n_1526)
);

OAI21xp5_ASAP7_75t_L g1527 ( 
.A1(n_1460),
.A2(n_1475),
.B(n_1481),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1394),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1394),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1435),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1375),
.B(n_1472),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1406),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1472),
.B(n_1400),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1432),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1400),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1415),
.Y(n_1536)
);

OAI21x1_ASAP7_75t_L g1537 ( 
.A1(n_1417),
.A2(n_1411),
.B(n_1425),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1464),
.A2(n_1467),
.B1(n_1478),
.B2(n_1475),
.Y(n_1538)
);

INVxp67_ASAP7_75t_L g1539 ( 
.A(n_1477),
.Y(n_1539)
);

BUFx3_ASAP7_75t_L g1540 ( 
.A(n_1455),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1430),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1431),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1417),
.Y(n_1543)
);

INVx2_ASAP7_75t_SL g1544 ( 
.A(n_1386),
.Y(n_1544)
);

AND2x4_ASAP7_75t_L g1545 ( 
.A(n_1411),
.B(n_1476),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1390),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1454),
.Y(n_1547)
);

AO21x1_ASAP7_75t_SL g1548 ( 
.A1(n_1373),
.A2(n_1361),
.B(n_1365),
.Y(n_1548)
);

BUFx2_ASAP7_75t_L g1549 ( 
.A(n_1393),
.Y(n_1549)
);

OAI21x1_ASAP7_75t_L g1550 ( 
.A1(n_1416),
.A2(n_1374),
.B(n_1373),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1390),
.Y(n_1551)
);

BUFx3_ASAP7_75t_L g1552 ( 
.A(n_1455),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1410),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1374),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1429),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1429),
.Y(n_1556)
);

INVx1_ASAP7_75t_SL g1557 ( 
.A(n_1392),
.Y(n_1557)
);

AO21x2_ASAP7_75t_L g1558 ( 
.A1(n_1418),
.A2(n_1361),
.B(n_1478),
.Y(n_1558)
);

INVx5_ASAP7_75t_L g1559 ( 
.A(n_1455),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1482),
.B(n_1474),
.Y(n_1560)
);

OAI21xp5_ASAP7_75t_L g1561 ( 
.A1(n_1467),
.A2(n_1474),
.B(n_1473),
.Y(n_1561)
);

BUFx3_ASAP7_75t_L g1562 ( 
.A(n_1459),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1419),
.Y(n_1563)
);

INVx1_ASAP7_75t_SL g1564 ( 
.A(n_1405),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1380),
.Y(n_1565)
);

BUFx2_ASAP7_75t_L g1566 ( 
.A(n_1382),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1380),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1419),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_SL g1569 ( 
.A1(n_1367),
.A2(n_1452),
.B1(n_1378),
.B2(n_1473),
.Y(n_1569)
);

OR2x2_ASAP7_75t_L g1570 ( 
.A(n_1470),
.B(n_1369),
.Y(n_1570)
);

BUFx2_ASAP7_75t_L g1571 ( 
.A(n_1421),
.Y(n_1571)
);

AOI21xp5_ASAP7_75t_L g1572 ( 
.A1(n_1470),
.A2(n_1459),
.B(n_1384),
.Y(n_1572)
);

NOR2xp33_ASAP7_75t_L g1573 ( 
.A(n_1371),
.B(n_1372),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_SL g1574 ( 
.A(n_1377),
.Y(n_1574)
);

BUFx3_ASAP7_75t_L g1575 ( 
.A(n_1459),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1379),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1395),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1488),
.B(n_1413),
.Y(n_1578)
);

OAI21xp5_ASAP7_75t_L g1579 ( 
.A1(n_1513),
.A2(n_1404),
.B(n_1402),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1488),
.B(n_1510),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1498),
.Y(n_1581)
);

OA21x2_ASAP7_75t_L g1582 ( 
.A1(n_1506),
.A2(n_1457),
.B(n_1409),
.Y(n_1582)
);

A2O1A1Ixp33_ASAP7_75t_L g1583 ( 
.A1(n_1513),
.A2(n_1401),
.B(n_1388),
.C(n_1383),
.Y(n_1583)
);

NAND2x1_ASAP7_75t_L g1584 ( 
.A(n_1517),
.B(n_1452),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1492),
.B(n_1483),
.Y(n_1585)
);

INVx3_ASAP7_75t_L g1586 ( 
.A(n_1555),
.Y(n_1586)
);

AOI22xp5_ASAP7_75t_L g1587 ( 
.A1(n_1493),
.A2(n_1452),
.B1(n_1367),
.B2(n_1378),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1533),
.B(n_1413),
.Y(n_1588)
);

NOR2xp33_ASAP7_75t_L g1589 ( 
.A(n_1514),
.B(n_1399),
.Y(n_1589)
);

A2O1A1Ixp33_ASAP7_75t_L g1590 ( 
.A1(n_1487),
.A2(n_1401),
.B(n_1383),
.C(n_1364),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_SL g1591 ( 
.A(n_1490),
.B(n_1362),
.Y(n_1591)
);

INVx3_ASAP7_75t_L g1592 ( 
.A(n_1555),
.Y(n_1592)
);

OAI22xp5_ASAP7_75t_SL g1593 ( 
.A1(n_1569),
.A2(n_1378),
.B1(n_1367),
.B2(n_1468),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1533),
.B(n_1362),
.Y(n_1594)
);

AO32x2_ASAP7_75t_L g1595 ( 
.A1(n_1502),
.A2(n_1414),
.A3(n_1391),
.B1(n_1366),
.B2(n_1461),
.Y(n_1595)
);

INVx1_ASAP7_75t_SL g1596 ( 
.A(n_1489),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1512),
.B(n_1414),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1498),
.Y(n_1598)
);

AO32x2_ASAP7_75t_L g1599 ( 
.A1(n_1525),
.A2(n_1453),
.A3(n_1377),
.B1(n_1465),
.B2(n_1412),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_SL g1600 ( 
.A1(n_1495),
.A2(n_1371),
.B1(n_1465),
.B2(n_1527),
.Y(n_1600)
);

AO21x2_ASAP7_75t_L g1601 ( 
.A1(n_1519),
.A2(n_1561),
.B(n_1550),
.Y(n_1601)
);

OA21x2_ASAP7_75t_L g1602 ( 
.A1(n_1519),
.A2(n_1550),
.B(n_1537),
.Y(n_1602)
);

INVx4_ASAP7_75t_L g1603 ( 
.A(n_1517),
.Y(n_1603)
);

NAND2x1_ASAP7_75t_L g1604 ( 
.A(n_1517),
.B(n_1555),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_1504),
.Y(n_1605)
);

CKINVDCx5p33_ASAP7_75t_R g1606 ( 
.A(n_1574),
.Y(n_1606)
);

BUFx12f_ASAP7_75t_L g1607 ( 
.A(n_1549),
.Y(n_1607)
);

BUFx12f_ASAP7_75t_L g1608 ( 
.A(n_1549),
.Y(n_1608)
);

OAI21x1_ASAP7_75t_SL g1609 ( 
.A1(n_1572),
.A2(n_1538),
.B(n_1568),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1560),
.B(n_1531),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1560),
.B(n_1531),
.Y(n_1611)
);

HB1xp67_ASAP7_75t_L g1612 ( 
.A(n_1497),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1565),
.B(n_1567),
.Y(n_1613)
);

AND2x4_ASAP7_75t_SL g1614 ( 
.A(n_1517),
.B(n_1547),
.Y(n_1614)
);

NOR2xp33_ASAP7_75t_L g1615 ( 
.A(n_1570),
.B(n_1554),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1565),
.B(n_1567),
.Y(n_1616)
);

AO32x2_ASAP7_75t_L g1617 ( 
.A1(n_1525),
.A2(n_1544),
.A3(n_1503),
.B1(n_1485),
.B2(n_1486),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1484),
.B(n_1526),
.Y(n_1618)
);

NAND4xp25_ASAP7_75t_L g1619 ( 
.A(n_1539),
.B(n_1570),
.C(n_1532),
.D(n_1536),
.Y(n_1619)
);

O2A1O1Ixp33_ASAP7_75t_L g1620 ( 
.A1(n_1516),
.A2(n_1518),
.B(n_1541),
.C(n_1542),
.Y(n_1620)
);

NOR2xp33_ASAP7_75t_L g1621 ( 
.A(n_1558),
.B(n_1501),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1507),
.B(n_1530),
.Y(n_1622)
);

AOI21xp5_ASAP7_75t_SL g1623 ( 
.A1(n_1517),
.A2(n_1508),
.B(n_1562),
.Y(n_1623)
);

A2O1A1Ixp33_ASAP7_75t_L g1624 ( 
.A1(n_1516),
.A2(n_1518),
.B(n_1515),
.C(n_1524),
.Y(n_1624)
);

NOR4xp25_ASAP7_75t_SL g1625 ( 
.A(n_1541),
.B(n_1571),
.C(n_1566),
.D(n_1542),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_L g1626 ( 
.A(n_1558),
.B(n_1563),
.Y(n_1626)
);

AO21x2_ASAP7_75t_L g1627 ( 
.A1(n_1505),
.A2(n_1543),
.B(n_1534),
.Y(n_1627)
);

NOR2xp33_ASAP7_75t_L g1628 ( 
.A(n_1545),
.B(n_1535),
.Y(n_1628)
);

A2O1A1Ixp33_ASAP7_75t_L g1629 ( 
.A1(n_1524),
.A2(n_1500),
.B(n_1535),
.C(n_1548),
.Y(n_1629)
);

NOR2xp33_ASAP7_75t_L g1630 ( 
.A(n_1545),
.B(n_1546),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1521),
.B(n_1522),
.Y(n_1631)
);

OAI21x1_ASAP7_75t_L g1632 ( 
.A1(n_1499),
.A2(n_1509),
.B(n_1511),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1612),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1610),
.B(n_1521),
.Y(n_1634)
);

AND2x4_ASAP7_75t_L g1635 ( 
.A(n_1603),
.B(n_1491),
.Y(n_1635)
);

AOI22xp33_ASAP7_75t_L g1636 ( 
.A1(n_1600),
.A2(n_1548),
.B1(n_1545),
.B2(n_1546),
.Y(n_1636)
);

BUFx2_ASAP7_75t_L g1637 ( 
.A(n_1617),
.Y(n_1637)
);

OAI221xp5_ASAP7_75t_L g1638 ( 
.A1(n_1590),
.A2(n_1551),
.B1(n_1566),
.B2(n_1557),
.C(n_1529),
.Y(n_1638)
);

INVxp67_ASAP7_75t_SL g1639 ( 
.A(n_1626),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_L g1640 ( 
.A(n_1589),
.B(n_1564),
.Y(n_1640)
);

INVxp67_ASAP7_75t_L g1641 ( 
.A(n_1626),
.Y(n_1641)
);

AOI22xp33_ASAP7_75t_L g1642 ( 
.A1(n_1591),
.A2(n_1545),
.B1(n_1551),
.B2(n_1556),
.Y(n_1642)
);

AND2x4_ASAP7_75t_L g1643 ( 
.A(n_1603),
.B(n_1494),
.Y(n_1643)
);

OAI21xp5_ASAP7_75t_L g1644 ( 
.A1(n_1620),
.A2(n_1528),
.B(n_1529),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1581),
.Y(n_1645)
);

INVx3_ASAP7_75t_L g1646 ( 
.A(n_1632),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1631),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1581),
.Y(n_1648)
);

HB1xp67_ASAP7_75t_L g1649 ( 
.A(n_1627),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1598),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1622),
.B(n_1618),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1611),
.B(n_1522),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1618),
.B(n_1520),
.Y(n_1653)
);

CKINVDCx6p67_ASAP7_75t_R g1654 ( 
.A(n_1607),
.Y(n_1654)
);

NAND3xp33_ASAP7_75t_L g1655 ( 
.A(n_1624),
.B(n_1528),
.C(n_1508),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1615),
.B(n_1523),
.Y(n_1656)
);

HB1xp67_ASAP7_75t_L g1657 ( 
.A(n_1627),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1615),
.B(n_1523),
.Y(n_1658)
);

NOR2xp67_ASAP7_75t_SL g1659 ( 
.A(n_1623),
.B(n_1559),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1621),
.B(n_1496),
.Y(n_1660)
);

NOR2xp33_ASAP7_75t_L g1661 ( 
.A(n_1589),
.B(n_1596),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1651),
.B(n_1621),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1645),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1641),
.B(n_1630),
.Y(n_1664)
);

OAI211xp5_ASAP7_75t_L g1665 ( 
.A1(n_1644),
.A2(n_1624),
.B(n_1590),
.C(n_1629),
.Y(n_1665)
);

NAND3xp33_ASAP7_75t_L g1666 ( 
.A(n_1655),
.B(n_1629),
.C(n_1591),
.Y(n_1666)
);

AOI221xp5_ASAP7_75t_L g1667 ( 
.A1(n_1655),
.A2(n_1644),
.B1(n_1638),
.B2(n_1593),
.C(n_1656),
.Y(n_1667)
);

HB1xp67_ASAP7_75t_L g1668 ( 
.A(n_1633),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1645),
.Y(n_1669)
);

AOI21xp33_ASAP7_75t_L g1670 ( 
.A1(n_1638),
.A2(n_1601),
.B(n_1616),
.Y(n_1670)
);

HB1xp67_ASAP7_75t_L g1671 ( 
.A(n_1633),
.Y(n_1671)
);

OAI222xp33_ASAP7_75t_L g1672 ( 
.A1(n_1636),
.A2(n_1587),
.B1(n_1584),
.B2(n_1580),
.C1(n_1594),
.C2(n_1585),
.Y(n_1672)
);

AOI221xp5_ASAP7_75t_L g1673 ( 
.A1(n_1656),
.A2(n_1619),
.B1(n_1630),
.B2(n_1628),
.C(n_1609),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1648),
.Y(n_1674)
);

INVxp67_ASAP7_75t_L g1675 ( 
.A(n_1639),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1653),
.B(n_1617),
.Y(n_1676)
);

NAND3xp33_ASAP7_75t_SL g1677 ( 
.A(n_1661),
.B(n_1625),
.C(n_1579),
.Y(n_1677)
);

AND2x4_ASAP7_75t_L g1678 ( 
.A(n_1635),
.B(n_1586),
.Y(n_1678)
);

INVx3_ASAP7_75t_L g1679 ( 
.A(n_1646),
.Y(n_1679)
);

AND2x4_ASAP7_75t_L g1680 ( 
.A(n_1635),
.B(n_1592),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1641),
.B(n_1601),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1639),
.B(n_1605),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1648),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1653),
.B(n_1617),
.Y(n_1684)
);

OR2x2_ASAP7_75t_L g1685 ( 
.A(n_1660),
.B(n_1602),
.Y(n_1685)
);

NAND4xp25_ASAP7_75t_L g1686 ( 
.A(n_1640),
.B(n_1613),
.C(n_1583),
.D(n_1658),
.Y(n_1686)
);

BUFx3_ASAP7_75t_L g1687 ( 
.A(n_1654),
.Y(n_1687)
);

AOI33xp33_ASAP7_75t_L g1688 ( 
.A1(n_1642),
.A2(n_1577),
.A3(n_1588),
.B1(n_1578),
.B2(n_1553),
.B3(n_1597),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1650),
.Y(n_1689)
);

OR2x2_ASAP7_75t_L g1690 ( 
.A(n_1660),
.B(n_1602),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1676),
.B(n_1684),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1676),
.B(n_1637),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1684),
.B(n_1637),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1675),
.B(n_1658),
.Y(n_1694)
);

OR2x6_ASAP7_75t_L g1695 ( 
.A(n_1666),
.B(n_1604),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1674),
.Y(n_1696)
);

BUFx2_ASAP7_75t_L g1697 ( 
.A(n_1678),
.Y(n_1697)
);

INVx1_ASAP7_75t_SL g1698 ( 
.A(n_1682),
.Y(n_1698)
);

INVx1_ASAP7_75t_SL g1699 ( 
.A(n_1682),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1663),
.Y(n_1700)
);

NAND5xp2_ASAP7_75t_L g1701 ( 
.A(n_1667),
.B(n_1583),
.C(n_1573),
.D(n_1577),
.E(n_1599),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1685),
.B(n_1649),
.Y(n_1702)
);

BUFx2_ASAP7_75t_SL g1703 ( 
.A(n_1687),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1663),
.Y(n_1704)
);

NAND2xp67_ASAP7_75t_L g1705 ( 
.A(n_1687),
.B(n_1599),
.Y(n_1705)
);

INVx1_ASAP7_75t_SL g1706 ( 
.A(n_1668),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1674),
.Y(n_1707)
);

OR2x2_ASAP7_75t_L g1708 ( 
.A(n_1685),
.B(n_1649),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1675),
.B(n_1634),
.Y(n_1709)
);

HB1xp67_ASAP7_75t_L g1710 ( 
.A(n_1671),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1683),
.Y(n_1711)
);

INVx2_ASAP7_75t_SL g1712 ( 
.A(n_1679),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1683),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1663),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1689),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1689),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1662),
.B(n_1647),
.Y(n_1717)
);

INVx2_ASAP7_75t_L g1718 ( 
.A(n_1669),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1664),
.B(n_1634),
.Y(n_1719)
);

BUFx2_ASAP7_75t_L g1720 ( 
.A(n_1695),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1696),
.Y(n_1721)
);

NOR2x1_ASAP7_75t_L g1722 ( 
.A(n_1703),
.B(n_1687),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1696),
.Y(n_1723)
);

NAND3xp33_ASAP7_75t_L g1724 ( 
.A(n_1695),
.B(n_1667),
.C(n_1666),
.Y(n_1724)
);

NOR2xp33_ASAP7_75t_L g1725 ( 
.A(n_1705),
.B(n_1654),
.Y(n_1725)
);

INVx3_ASAP7_75t_L g1726 ( 
.A(n_1712),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1696),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1707),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1707),
.Y(n_1729)
);

INVx2_ASAP7_75t_SL g1730 ( 
.A(n_1697),
.Y(n_1730)
);

NOR2xp33_ASAP7_75t_SL g1731 ( 
.A(n_1703),
.B(n_1672),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1700),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1700),
.Y(n_1733)
);

INVx2_ASAP7_75t_SL g1734 ( 
.A(n_1697),
.Y(n_1734)
);

XNOR2x1_ASAP7_75t_L g1735 ( 
.A(n_1695),
.B(n_1606),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1698),
.B(n_1681),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1707),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1700),
.Y(n_1738)
);

NOR2x1_ASAP7_75t_L g1739 ( 
.A(n_1703),
.B(n_1677),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_SL g1740 ( 
.A(n_1694),
.B(n_1673),
.Y(n_1740)
);

AOI22xp33_ASAP7_75t_SL g1741 ( 
.A1(n_1695),
.A2(n_1665),
.B1(n_1607),
.B2(n_1608),
.Y(n_1741)
);

AND2x4_ASAP7_75t_L g1742 ( 
.A(n_1697),
.B(n_1679),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1700),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1710),
.Y(n_1744)
);

OAI21xp33_ASAP7_75t_L g1745 ( 
.A1(n_1701),
.A2(n_1665),
.B(n_1673),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1711),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1704),
.Y(n_1747)
);

HB1xp67_ASAP7_75t_L g1748 ( 
.A(n_1710),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1711),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1719),
.B(n_1694),
.Y(n_1750)
);

INVx2_ASAP7_75t_SL g1751 ( 
.A(n_1711),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1713),
.Y(n_1752)
);

INVx1_ASAP7_75t_SL g1753 ( 
.A(n_1706),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1713),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1691),
.B(n_1662),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1713),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1691),
.B(n_1678),
.Y(n_1757)
);

BUFx2_ASAP7_75t_L g1758 ( 
.A(n_1695),
.Y(n_1758)
);

AOI22xp5_ASAP7_75t_L g1759 ( 
.A1(n_1695),
.A2(n_1677),
.B1(n_1686),
.B2(n_1701),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1704),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1715),
.Y(n_1761)
);

AND2x2_ASAP7_75t_SL g1762 ( 
.A(n_1692),
.B(n_1688),
.Y(n_1762)
);

CKINVDCx16_ASAP7_75t_R g1763 ( 
.A(n_1731),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1755),
.B(n_1757),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1721),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1755),
.B(n_1695),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1753),
.B(n_1705),
.Y(n_1767)
);

NAND2x1p5_ASAP7_75t_L g1768 ( 
.A(n_1722),
.B(n_1659),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1757),
.B(n_1695),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1751),
.Y(n_1770)
);

INVx1_ASAP7_75t_SL g1771 ( 
.A(n_1735),
.Y(n_1771)
);

OR2x2_ASAP7_75t_L g1772 ( 
.A(n_1744),
.B(n_1698),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1721),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1723),
.Y(n_1774)
);

CKINVDCx16_ASAP7_75t_R g1775 ( 
.A(n_1739),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1723),
.Y(n_1776)
);

INVx1_ASAP7_75t_SL g1777 ( 
.A(n_1722),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1727),
.Y(n_1778)
);

AOI21xp5_ASAP7_75t_SL g1779 ( 
.A1(n_1724),
.A2(n_1606),
.B(n_1599),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1762),
.B(n_1691),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1727),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1751),
.Y(n_1782)
);

HB1xp67_ASAP7_75t_L g1783 ( 
.A(n_1748),
.Y(n_1783)
);

NOR2xp33_ASAP7_75t_L g1784 ( 
.A(n_1725),
.B(n_1654),
.Y(n_1784)
);

AND2x2_ASAP7_75t_SL g1785 ( 
.A(n_1762),
.B(n_1582),
.Y(n_1785)
);

AOI22x1_ASAP7_75t_L g1786 ( 
.A1(n_1724),
.A2(n_1576),
.B1(n_1608),
.B2(n_1706),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1762),
.B(n_1692),
.Y(n_1787)
);

CKINVDCx16_ASAP7_75t_R g1788 ( 
.A(n_1739),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1720),
.B(n_1692),
.Y(n_1789)
);

NAND2x1p5_ASAP7_75t_L g1790 ( 
.A(n_1759),
.B(n_1659),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1720),
.B(n_1693),
.Y(n_1791)
);

AO21x1_ASAP7_75t_L g1792 ( 
.A1(n_1740),
.A2(n_1693),
.B(n_1702),
.Y(n_1792)
);

NOR2xp33_ASAP7_75t_L g1793 ( 
.A(n_1745),
.B(n_1705),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1745),
.B(n_1719),
.Y(n_1794)
);

AOI21xp33_ASAP7_75t_SL g1795 ( 
.A1(n_1735),
.A2(n_1670),
.B(n_1599),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1750),
.B(n_1699),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1758),
.B(n_1693),
.Y(n_1797)
);

OR2x2_ASAP7_75t_L g1798 ( 
.A(n_1736),
.B(n_1699),
.Y(n_1798)
);

CKINVDCx16_ASAP7_75t_R g1799 ( 
.A(n_1763),
.Y(n_1799)
);

AOI221xp5_ASAP7_75t_L g1800 ( 
.A1(n_1795),
.A2(n_1779),
.B1(n_1793),
.B2(n_1787),
.C(n_1775),
.Y(n_1800)
);

AOI21xp5_ASAP7_75t_L g1801 ( 
.A1(n_1779),
.A2(n_1759),
.B(n_1741),
.Y(n_1801)
);

OAI21xp5_ASAP7_75t_L g1802 ( 
.A1(n_1771),
.A2(n_1758),
.B(n_1672),
.Y(n_1802)
);

NOR2xp33_ASAP7_75t_L g1803 ( 
.A(n_1794),
.B(n_1784),
.Y(n_1803)
);

AOI22xp5_ASAP7_75t_L g1804 ( 
.A1(n_1775),
.A2(n_1686),
.B1(n_1734),
.B2(n_1730),
.Y(n_1804)
);

OAI21xp33_ASAP7_75t_SL g1805 ( 
.A1(n_1787),
.A2(n_1734),
.B(n_1730),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1765),
.Y(n_1806)
);

OAI333xp33_ASAP7_75t_L g1807 ( 
.A1(n_1788),
.A2(n_1664),
.A3(n_1729),
.B1(n_1756),
.B2(n_1754),
.B3(n_1752),
.C1(n_1749),
.C2(n_1728),
.C3(n_1737),
.Y(n_1807)
);

XNOR2xp5_ASAP7_75t_L g1808 ( 
.A(n_1786),
.B(n_1578),
.Y(n_1808)
);

HB1xp67_ASAP7_75t_L g1809 ( 
.A(n_1783),
.Y(n_1809)
);

OAI21xp5_ASAP7_75t_L g1810 ( 
.A1(n_1786),
.A2(n_1670),
.B(n_1736),
.Y(n_1810)
);

AOI21xp5_ASAP7_75t_L g1811 ( 
.A1(n_1788),
.A2(n_1681),
.B(n_1709),
.Y(n_1811)
);

AOI22xp5_ASAP7_75t_L g1812 ( 
.A1(n_1763),
.A2(n_1628),
.B1(n_1709),
.B2(n_1643),
.Y(n_1812)
);

OR2x2_ASAP7_75t_L g1813 ( 
.A(n_1796),
.B(n_1652),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1764),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1780),
.B(n_1728),
.Y(n_1815)
);

AOI22xp5_ASAP7_75t_L g1816 ( 
.A1(n_1785),
.A2(n_1643),
.B1(n_1742),
.B2(n_1680),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1765),
.Y(n_1817)
);

OAI32xp33_ASAP7_75t_L g1818 ( 
.A1(n_1777),
.A2(n_1726),
.A3(n_1702),
.B1(n_1708),
.B2(n_1690),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1773),
.Y(n_1819)
);

AOI22xp5_ASAP7_75t_L g1820 ( 
.A1(n_1785),
.A2(n_1643),
.B1(n_1742),
.B2(n_1680),
.Y(n_1820)
);

OAI21xp5_ASAP7_75t_SL g1821 ( 
.A1(n_1790),
.A2(n_1742),
.B(n_1614),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1764),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1767),
.B(n_1717),
.Y(n_1823)
);

INVx1_ASAP7_75t_SL g1824 ( 
.A(n_1777),
.Y(n_1824)
);

AOI22xp5_ASAP7_75t_L g1825 ( 
.A1(n_1800),
.A2(n_1801),
.B1(n_1799),
.B2(n_1785),
.Y(n_1825)
);

BUFx2_ASAP7_75t_L g1826 ( 
.A(n_1805),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1809),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1806),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1824),
.B(n_1780),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1803),
.B(n_1795),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1817),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1819),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1814),
.Y(n_1833)
);

OAI22xp5_ASAP7_75t_L g1834 ( 
.A1(n_1802),
.A2(n_1790),
.B1(n_1768),
.B2(n_1772),
.Y(n_1834)
);

OAI22xp5_ASAP7_75t_L g1835 ( 
.A1(n_1802),
.A2(n_1790),
.B1(n_1768),
.B2(n_1772),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1815),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1815),
.Y(n_1837)
);

AOI322xp5_ASAP7_75t_SL g1838 ( 
.A1(n_1807),
.A2(n_1792),
.A3(n_1797),
.B1(n_1791),
.B2(n_1789),
.C1(n_1657),
.C2(n_1766),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1822),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1813),
.Y(n_1840)
);

INVxp67_ASAP7_75t_L g1841 ( 
.A(n_1804),
.Y(n_1841)
);

OAI31xp33_ASAP7_75t_L g1842 ( 
.A1(n_1821),
.A2(n_1768),
.A3(n_1796),
.B(n_1792),
.Y(n_1842)
);

NOR2xp33_ASAP7_75t_L g1843 ( 
.A(n_1808),
.B(n_1798),
.Y(n_1843)
);

INVxp67_ASAP7_75t_SL g1844 ( 
.A(n_1823),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1833),
.Y(n_1845)
);

AOI22xp5_ASAP7_75t_SL g1846 ( 
.A1(n_1826),
.A2(n_1810),
.B1(n_1791),
.B2(n_1797),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1833),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1843),
.B(n_1789),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1829),
.B(n_1769),
.Y(n_1849)
);

A2O1A1Ixp33_ASAP7_75t_L g1850 ( 
.A1(n_1842),
.A2(n_1825),
.B(n_1826),
.C(n_1843),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1827),
.B(n_1769),
.Y(n_1851)
);

AOI22xp5_ASAP7_75t_L g1852 ( 
.A1(n_1841),
.A2(n_1812),
.B1(n_1810),
.B2(n_1816),
.Y(n_1852)
);

NAND2xp33_ASAP7_75t_SL g1853 ( 
.A(n_1834),
.B(n_1798),
.Y(n_1853)
);

NOR3xp33_ASAP7_75t_L g1854 ( 
.A(n_1830),
.B(n_1818),
.C(n_1811),
.Y(n_1854)
);

AOI322xp5_ASAP7_75t_L g1855 ( 
.A1(n_1838),
.A2(n_1766),
.A3(n_1820),
.B1(n_1770),
.B2(n_1782),
.C1(n_1776),
.C2(n_1774),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1839),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1845),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1849),
.B(n_1844),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1856),
.Y(n_1859)
);

NAND3xp33_ASAP7_75t_SL g1860 ( 
.A(n_1850),
.B(n_1835),
.C(n_1838),
.Y(n_1860)
);

NAND4xp25_ASAP7_75t_L g1861 ( 
.A(n_1850),
.B(n_1837),
.C(n_1836),
.D(n_1839),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1847),
.B(n_1828),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1851),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1848),
.B(n_1840),
.Y(n_1864)
);

NOR2xp33_ASAP7_75t_L g1865 ( 
.A(n_1853),
.B(n_1831),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1846),
.Y(n_1866)
);

OAI21xp33_ASAP7_75t_SL g1867 ( 
.A1(n_1855),
.A2(n_1832),
.B(n_1782),
.Y(n_1867)
);

AOI21xp5_ASAP7_75t_L g1868 ( 
.A1(n_1860),
.A2(n_1854),
.B(n_1852),
.Y(n_1868)
);

AOI22xp5_ASAP7_75t_L g1869 ( 
.A1(n_1867),
.A2(n_1854),
.B1(n_1832),
.B2(n_1782),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1865),
.B(n_1770),
.Y(n_1870)
);

NOR2xp67_ASAP7_75t_L g1871 ( 
.A(n_1861),
.B(n_1770),
.Y(n_1871)
);

OAI22xp5_ASAP7_75t_L g1872 ( 
.A1(n_1866),
.A2(n_1863),
.B1(n_1864),
.B2(n_1858),
.Y(n_1872)
);

NAND4xp75_ASAP7_75t_L g1873 ( 
.A(n_1862),
.B(n_1781),
.C(n_1778),
.D(n_1776),
.Y(n_1873)
);

NAND4xp25_ASAP7_75t_SL g1874 ( 
.A(n_1862),
.B(n_1781),
.C(n_1778),
.D(n_1774),
.Y(n_1874)
);

OAI221xp5_ASAP7_75t_SL g1875 ( 
.A1(n_1868),
.A2(n_1859),
.B1(n_1857),
.B2(n_1773),
.C(n_1726),
.Y(n_1875)
);

AOI221x1_ASAP7_75t_L g1876 ( 
.A1(n_1872),
.A2(n_1726),
.B1(n_1761),
.B2(n_1756),
.C(n_1754),
.Y(n_1876)
);

OAI211xp5_ASAP7_75t_L g1877 ( 
.A1(n_1869),
.A2(n_1726),
.B(n_1760),
.C(n_1732),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1870),
.Y(n_1878)
);

OAI22xp33_ASAP7_75t_L g1879 ( 
.A1(n_1871),
.A2(n_1712),
.B1(n_1708),
.B2(n_1702),
.Y(n_1879)
);

AOI211xp5_ASAP7_75t_L g1880 ( 
.A1(n_1874),
.A2(n_1742),
.B(n_1737),
.C(n_1752),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1873),
.Y(n_1881)
);

NOR2x1_ASAP7_75t_L g1882 ( 
.A(n_1881),
.B(n_1878),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1879),
.B(n_1729),
.Y(n_1883)
);

INVx1_ASAP7_75t_SL g1884 ( 
.A(n_1875),
.Y(n_1884)
);

OR2x2_ASAP7_75t_L g1885 ( 
.A(n_1877),
.B(n_1746),
.Y(n_1885)
);

NOR2xp67_ASAP7_75t_L g1886 ( 
.A(n_1876),
.B(n_1746),
.Y(n_1886)
);

NAND3xp33_ASAP7_75t_L g1887 ( 
.A(n_1882),
.B(n_1880),
.C(n_1733),
.Y(n_1887)
);

NAND3xp33_ASAP7_75t_SL g1888 ( 
.A(n_1884),
.B(n_1595),
.C(n_1732),
.Y(n_1888)
);

AOI21xp33_ASAP7_75t_SL g1889 ( 
.A1(n_1885),
.A2(n_1761),
.B(n_1749),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1887),
.Y(n_1890)
);

OAI22xp5_ASAP7_75t_L g1891 ( 
.A1(n_1890),
.A2(n_1883),
.B1(n_1886),
.B2(n_1889),
.Y(n_1891)
);

XNOR2x1_ASAP7_75t_L g1892 ( 
.A(n_1891),
.B(n_1888),
.Y(n_1892)
);

OAI22xp5_ASAP7_75t_SL g1893 ( 
.A1(n_1891),
.A2(n_1760),
.B1(n_1747),
.B2(n_1743),
.Y(n_1893)
);

HB1xp67_ASAP7_75t_L g1894 ( 
.A(n_1892),
.Y(n_1894)
);

CKINVDCx20_ASAP7_75t_R g1895 ( 
.A(n_1893),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1895),
.Y(n_1896)
);

OAI21xp5_ASAP7_75t_L g1897 ( 
.A1(n_1894),
.A2(n_1738),
.B(n_1733),
.Y(n_1897)
);

AOI22xp33_ASAP7_75t_L g1898 ( 
.A1(n_1896),
.A2(n_1747),
.B1(n_1743),
.B2(n_1738),
.Y(n_1898)
);

OAI22xp5_ASAP7_75t_L g1899 ( 
.A1(n_1898),
.A2(n_1897),
.B1(n_1708),
.B2(n_1712),
.Y(n_1899)
);

OAI22xp33_ASAP7_75t_L g1900 ( 
.A1(n_1899),
.A2(n_1712),
.B1(n_1718),
.B2(n_1704),
.Y(n_1900)
);

AOI221xp5_ASAP7_75t_L g1901 ( 
.A1(n_1900),
.A2(n_1716),
.B1(n_1715),
.B2(n_1704),
.C(n_1714),
.Y(n_1901)
);

AOI211xp5_ASAP7_75t_L g1902 ( 
.A1(n_1901),
.A2(n_1575),
.B(n_1540),
.C(n_1552),
.Y(n_1902)
);


endmodule