module fake_jpeg_4560_n_320 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_320);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_320;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx4f_ASAP7_75t_SL g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_35),
.B(n_39),
.Y(n_50)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_22),
.B(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_38),
.A2(n_26),
.B1(n_31),
.B2(n_24),
.Y(n_69)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_43),
.Y(n_66)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_15),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_32),
.B1(n_22),
.B2(n_20),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_44),
.A2(n_36),
.B1(n_20),
.B2(n_29),
.Y(n_82)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_46),
.Y(n_80)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

BUFx2_ASAP7_75t_SL g87 ( 
.A(n_47),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_51),
.B(n_58),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_L g52 ( 
.A1(n_42),
.A2(n_33),
.B1(n_19),
.B2(n_28),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_52),
.A2(n_63),
.B1(n_17),
.B2(n_25),
.Y(n_83)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_59),
.Y(n_74)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_61),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_38),
.A2(n_32),
.B1(n_22),
.B2(n_20),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_65),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_37),
.B(n_32),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_37),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_71),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_64),
.A2(n_38),
.B1(n_39),
.B2(n_36),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_72),
.A2(n_56),
.B1(n_46),
.B2(n_36),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_75),
.Y(n_101)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_37),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_54),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_82),
.A2(n_57),
.B1(n_55),
.B2(n_53),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_83),
.A2(n_67),
.B1(n_27),
.B2(n_47),
.Y(n_100)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_88),
.Y(n_114)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_90),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_45),
.A2(n_39),
.B(n_35),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_91),
.B(n_35),
.C(n_41),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_74),
.A2(n_54),
.B1(n_67),
.B2(n_38),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_94),
.A2(n_100),
.B1(n_112),
.B2(n_120),
.Y(n_137)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_97),
.B(n_34),
.Y(n_142)
);

A2O1A1O1Ixp25_ASAP7_75t_L g98 ( 
.A1(n_89),
.A2(n_50),
.B(n_41),
.C(n_52),
.D(n_36),
.Y(n_98)
);

A2O1A1O1Ixp25_ASAP7_75t_L g123 ( 
.A1(n_98),
.A2(n_41),
.B(n_49),
.C(n_34),
.D(n_19),
.Y(n_123)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_99),
.B(n_103),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_102),
.A2(n_111),
.B1(n_75),
.B2(n_93),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_91),
.Y(n_103)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_39),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_113),
.Y(n_129)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

INVx4_ASAP7_75t_SL g108 ( 
.A(n_90),
.Y(n_108)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_110),
.A2(n_29),
.B(n_34),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_38),
.B1(n_56),
.B2(n_35),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_73),
.B(n_61),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_72),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_116),
.Y(n_136)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_119),
.Y(n_139)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_118),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_17),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_71),
.A2(n_41),
.B1(n_31),
.B2(n_17),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_121),
.A2(n_131),
.B1(n_146),
.B2(n_106),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_105),
.B(n_41),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_122),
.B(n_123),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_103),
.A2(n_27),
.B(n_26),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_124),
.A2(n_128),
.B(n_133),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_110),
.A2(n_27),
.B(n_26),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_116),
.A2(n_85),
.B1(n_79),
.B2(n_84),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_113),
.A2(n_29),
.B(n_31),
.Y(n_133)
);

AO22x1_ASAP7_75t_L g135 ( 
.A1(n_98),
.A2(n_102),
.B1(n_100),
.B2(n_115),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_135),
.A2(n_109),
.B1(n_34),
.B2(n_107),
.Y(n_162)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_120),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_140),
.B(n_106),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_99),
.A2(n_85),
.B1(n_24),
.B2(n_25),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_142),
.B(n_114),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_97),
.B(n_101),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_23),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_98),
.A2(n_79),
.B1(n_88),
.B2(n_34),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_144),
.A2(n_145),
.B1(n_30),
.B2(n_21),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_119),
.A2(n_34),
.B1(n_24),
.B2(n_25),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_111),
.A2(n_101),
.B1(n_117),
.B2(n_95),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_147),
.A2(n_28),
.B(n_21),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_149),
.B(n_150),
.Y(n_192)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_129),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_151),
.B(n_153),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_133),
.B(n_114),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_159),
.Y(n_180)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_154),
.A2(n_158),
.B1(n_162),
.B2(n_165),
.Y(n_177)
);

OAI21xp33_ASAP7_75t_SL g156 ( 
.A1(n_135),
.A2(n_104),
.B(n_108),
.Y(n_156)
);

FAx1_ASAP7_75t_SL g190 ( 
.A(n_156),
.B(n_166),
.CI(n_168),
.CON(n_190),
.SN(n_190)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_157),
.A2(n_124),
.B(n_145),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_135),
.A2(n_109),
.B1(n_118),
.B2(n_108),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_136),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_160),
.B(n_161),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_139),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_140),
.A2(n_30),
.B1(n_33),
.B2(n_21),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_164),
.A2(n_172),
.B(n_126),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_123),
.A2(n_19),
.B1(n_33),
.B2(n_21),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_136),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_167),
.B(n_142),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g169 ( 
.A(n_144),
.B(n_16),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_169),
.B(n_16),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_137),
.A2(n_70),
.B1(n_78),
.B2(n_33),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_170),
.A2(n_125),
.B1(n_130),
.B2(n_134),
.Y(n_187)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_134),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_171),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_139),
.B(n_1),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_146),
.Y(n_173)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_173),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g174 ( 
.A(n_121),
.Y(n_174)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_174),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_162),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_175),
.B(n_178),
.C(n_181),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_170),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_196),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_148),
.B(n_147),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_122),
.C(n_127),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g182 ( 
.A(n_171),
.Y(n_182)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_182),
.Y(n_209)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_184),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_150),
.B(n_122),
.C(n_127),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_185),
.B(n_186),
.C(n_188),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_128),
.C(n_123),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_187),
.A2(n_154),
.B1(n_157),
.B2(n_166),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_137),
.C(n_142),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_189),
.A2(n_194),
.B(n_152),
.Y(n_206)
);

AO21x1_ASAP7_75t_L g216 ( 
.A1(n_191),
.A2(n_197),
.B(n_179),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_155),
.A2(n_132),
.B(n_130),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_161),
.Y(n_196)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_149),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_167),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_160),
.B(n_125),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_23),
.C(n_77),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_188),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_195),
.A2(n_173),
.B1(n_174),
.B2(n_153),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_201),
.A2(n_208),
.B1(n_215),
.B2(n_217),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_213),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_204),
.Y(n_227)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_205),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_206),
.A2(n_225),
.B(n_190),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_178),
.B(n_165),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_207),
.B(n_221),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_177),
.A2(n_159),
.B1(n_168),
.B2(n_155),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_172),
.Y(n_210)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_210),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_R g211 ( 
.A(n_194),
.B(n_164),
.C(n_163),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_214),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_182),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_177),
.A2(n_126),
.B1(n_138),
.B2(n_70),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_218),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_176),
.A2(n_180),
.B1(n_192),
.B2(n_175),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_193),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_180),
.B(n_138),
.Y(n_220)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_220),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_181),
.B(n_77),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_222),
.B(n_199),
.C(n_191),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_182),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_223),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_185),
.B(n_28),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_1),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_189),
.A2(n_186),
.B(n_190),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_245),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_228),
.B(n_234),
.C(n_241),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_231),
.A2(n_209),
.B(n_215),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_205),
.A2(n_190),
.B1(n_200),
.B2(n_183),
.Y(n_233)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_233),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_183),
.C(n_62),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_225),
.A2(n_28),
.B1(n_30),
.B2(n_3),
.Y(n_235)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_235),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_202),
.A2(n_212),
.B1(n_216),
.B2(n_208),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_236),
.A2(n_211),
.B1(n_202),
.B2(n_206),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_219),
.B(n_1),
.C(n_2),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_224),
.B(n_15),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_242),
.B(n_246),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_219),
.C(n_207),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_14),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_210),
.B(n_2),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_244),
.B(n_222),
.Y(n_248)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_248),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g274 ( 
.A(n_250),
.B(n_245),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_246),
.B(n_220),
.Y(n_251)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_251),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_253),
.B(n_226),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_233),
.B(n_203),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_254),
.B(n_261),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_204),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_255),
.A2(n_256),
.B(n_237),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_238),
.B(n_209),
.C(n_214),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_260),
.C(n_263),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_13),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_231),
.B(n_11),
.Y(n_261)
);

FAx1_ASAP7_75t_SL g262 ( 
.A(n_236),
.B(n_232),
.CI(n_240),
.CON(n_262),
.SN(n_262)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_235),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_228),
.B(n_2),
.C(n_3),
.Y(n_263)
);

BUFx24_ASAP7_75t_SL g286 ( 
.A(n_264),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_257),
.A2(n_230),
.B1(n_232),
.B2(n_229),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_265),
.A2(n_263),
.B1(n_252),
.B2(n_237),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_266),
.A2(n_274),
.B(n_278),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_256),
.Y(n_269)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_269),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_243),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_270),
.B(n_271),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_262),
.B(n_227),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_259),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_272),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_252),
.C(n_254),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_275),
.C(n_253),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_234),
.C(n_241),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_277),
.A2(n_258),
.B1(n_250),
.B2(n_261),
.Y(n_279)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_279),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_4),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_268),
.B(n_247),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_282),
.B(n_280),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_284),
.C(n_285),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_273),
.B(n_260),
.C(n_3),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_274),
.A2(n_12),
.B1(n_3),
.B2(n_4),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_288),
.B(n_4),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_276),
.A2(n_272),
.B1(n_267),
.B2(n_275),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_283),
.C(n_284),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_267),
.B(n_276),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_291),
.A2(n_12),
.B(n_5),
.Y(n_295)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_294),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_297),
.Y(n_304)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_296),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_6),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_299),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_6),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_300),
.B(n_285),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_289),
.Y(n_301)
);

AO21x1_ASAP7_75t_L g309 ( 
.A1(n_301),
.A2(n_12),
.B(n_7),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_302),
.Y(n_311)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_301),
.Y(n_303)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_303),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_286),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_308),
.A2(n_309),
.B(n_294),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_310),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_292),
.Y(n_313)
);

MAJx2_ASAP7_75t_L g315 ( 
.A(n_313),
.B(n_305),
.C(n_306),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_312),
.B1(n_311),
.B2(n_304),
.Y(n_316)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g317 ( 
.A1(n_316),
.A2(n_314),
.B(n_304),
.C(n_9),
.D(n_10),
.Y(n_317)
);

OAI321xp33_ASAP7_75t_L g318 ( 
.A1(n_317),
.A2(n_6),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C(n_294),
.Y(n_318)
);

A2O1A1Ixp33_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_8),
.B(n_10),
.C(n_294),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_8),
.Y(n_320)
);


endmodule