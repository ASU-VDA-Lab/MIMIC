module real_jpeg_25204_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_1),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

INVx8_ASAP7_75t_SL g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_4),
.B(n_39),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_4),
.B(n_62),
.C(n_65),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_4),
.A2(n_26),
.B1(n_52),
.B2(n_53),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_4),
.B(n_55),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_4),
.A2(n_105),
.B1(n_165),
.B2(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_5),
.A2(n_65),
.B1(n_66),
.B2(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_5),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_5),
.A2(n_52),
.B1(n_53),
.B2(n_81),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_6),
.A2(n_25),
.B1(n_28),
.B2(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_6),
.A2(n_33),
.B1(n_34),
.B2(n_42),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_6),
.A2(n_42),
.B1(n_52),
.B2(n_53),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_6),
.A2(n_42),
.B1(n_65),
.B2(n_66),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_7),
.A2(n_33),
.B1(n_34),
.B2(n_46),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_7),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_7),
.A2(n_25),
.B1(n_38),
.B2(n_46),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_7),
.A2(n_46),
.B1(n_52),
.B2(n_53),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_7),
.A2(n_46),
.B1(n_65),
.B2(n_66),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_9),
.A2(n_33),
.B1(n_34),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_9),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_9),
.A2(n_57),
.B1(n_65),
.B2(n_66),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_9),
.A2(n_52),
.B1(n_53),
.B2(n_57),
.Y(n_190)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

NAND3xp33_ASAP7_75t_L g74 ( 
.A(n_10),
.B(n_32),
.C(n_33),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_11),
.A2(n_52),
.B1(n_53),
.B2(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_11),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_68),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_11),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_12),
.A2(n_52),
.B1(n_53),
.B2(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_12),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_12),
.A2(n_65),
.B1(n_66),
.B2(n_71),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_13),
.A2(n_65),
.B1(n_66),
.B2(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_13),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_15),
.Y(n_78)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_15),
.Y(n_85)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_15),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_128),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_126),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_101),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_20),
.B(n_101),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_72),
.C(n_90),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_21),
.B(n_211),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_43),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_22),
.B(n_44),
.C(n_58),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_29),
.B1(n_39),
.B2(n_40),
.Y(n_22)
);

OAI21xp33_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_26),
.B(n_27),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_26),
.B(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_26),
.B(n_64),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_26),
.B(n_172),
.Y(n_171)
);

HAxp5_ASAP7_75t_SL g182 ( 
.A(n_26),
.B(n_34),
.CON(n_182),
.SN(n_182)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_27),
.A2(n_31),
.B(n_34),
.C(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_29),
.Y(n_117)
);

AND2x2_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_36),
.Y(n_29)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_30),
.A2(n_41),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_L g36 ( 
.A1(n_31),
.A2(n_32),
.B1(n_37),
.B2(n_38),
.Y(n_36)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_33),
.A2(n_34),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

NOR3xp33_ASAP7_75t_L g183 ( 
.A(n_33),
.B(n_49),
.C(n_53),
.Y(n_183)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_58),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_47),
.B1(n_55),
.B2(n_56),
.Y(n_44)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_45),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_47),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_47),
.A2(n_55),
.B1(n_98),
.B2(n_182),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_51),
.Y(n_47)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_49),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_51)
);

O2A1O1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_50),
.A2(n_52),
.B(n_181),
.C(n_183),
.Y(n_180)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_51),
.A2(n_97),
.B1(n_99),
.B2(n_100),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_52),
.A2(n_53),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_53),
.B(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_55),
.B(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_56),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_67),
.B(n_69),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_59),
.B(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_59),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_59),
.A2(n_138),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_60),
.A2(n_64),
.B1(n_140),
.B2(n_153),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_60),
.A2(n_204),
.B(n_205),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_62),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

INVx3_ASAP7_75t_SL g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_70),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_64),
.A2(n_109),
.B(n_110),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_64),
.Y(n_138)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_66),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_67),
.B(n_138),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_70),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_72),
.B(n_90),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_75),
.B1(n_88),
.B2(n_89),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_73),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_73),
.B(n_88),
.Y(n_124)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_79),
.B1(n_82),
.B2(n_86),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_76),
.B(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_76),
.A2(n_82),
.B1(n_157),
.B2(n_159),
.Y(n_156)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_78),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_80),
.A2(n_85),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_82),
.B(n_93),
.Y(n_107)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_83),
.A2(n_105),
.B1(n_158),
.B2(n_165),
.Y(n_164)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_SL g145 ( 
.A(n_85),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_86),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_94),
.C(n_96),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_91),
.A2(n_94),
.B1(n_95),
.B2(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_91),
.Y(n_199)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_96),
.B(n_198),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_99),
.A2(n_121),
.B(n_122),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_113),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_112),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_108),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_106),
.B(n_107),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_105),
.A2(n_143),
.B(n_144),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_105),
.A2(n_107),
.B(n_147),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_124),
.B2(n_125),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_116),
.B(n_120),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_124),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_209),
.B(n_213),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_193),
.B(n_208),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_176),
.B(n_192),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_154),
.B(n_175),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_141),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_133),
.B(n_141),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_136),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_148),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_142),
.B(n_149),
.C(n_152),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_143),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_150),
.B1(n_151),
.B2(n_152),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_153),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_161),
.B(n_174),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_160),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_160),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_166),
.B(n_173),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_163),
.B(n_164),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_170),
.Y(n_166)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_191),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_177),
.B(n_191),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_186),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_187),
.C(n_188),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_184),
.B2(n_185),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_179),
.B(n_185),
.Y(n_202)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_190),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_195),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_200),
.B2(n_201),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_203),
.C(n_206),
.Y(n_212)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_206),
.B2(n_207),
.Y(n_201)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_202),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_203),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_212),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_210),
.B(n_212),
.Y(n_213)
);


endmodule