module fake_jpeg_12157_n_98 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_98);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_98;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g11 ( 
.A(n_9),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_0),
.B(n_7),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_13),
.B(n_2),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_28),
.B(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_14),
.B(n_5),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_29),
.B(n_32),
.Y(n_57)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_21),
.B(n_6),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_22),
.A2(n_3),
.B1(n_4),
.B2(n_19),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_33),
.A2(n_34),
.B1(n_40),
.B2(n_42),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_18),
.A2(n_3),
.B1(n_4),
.B2(n_20),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_17),
.B(n_26),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_28),
.Y(n_45)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_15),
.B(n_4),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_20),
.A2(n_12),
.B1(n_24),
.B2(n_23),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_24),
.A2(n_13),
.B1(n_16),
.B2(n_26),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_44),
.Y(n_58)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_45),
.B(n_51),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_30),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_52),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_42),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_37),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_40),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_55),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_27),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_41),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_SL g67 ( 
.A(n_61),
.B(n_58),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_35),
.B(n_38),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_57),
.Y(n_75)
);

MAJx2_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_45),
.C(n_62),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_63),
.B(n_75),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_59),
.A2(n_54),
.B(n_52),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_64),
.A2(n_66),
.B(n_49),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_58),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_67),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_59),
.A2(n_55),
.B(n_58),
.Y(n_66)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_72),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_74),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_72),
.C(n_56),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_71),
.A2(n_70),
.B1(n_64),
.B2(n_73),
.Y(n_81)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_81),
.B(n_75),
.Y(n_85)
);

NOR3xp33_ASAP7_75t_SL g89 ( 
.A(n_85),
.B(n_88),
.C(n_84),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_76),
.B(n_63),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_86),
.B(n_87),
.C(n_82),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_84),
.B(n_50),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_90),
.B(n_91),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_86),
.B(n_80),
.C(n_82),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_89),
.B(n_87),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_79),
.C(n_78),
.Y(n_94)
);

AOI31xp67_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_92),
.A3(n_93),
.B(n_47),
.Y(n_95)
);

BUFx24_ASAP7_75t_SL g96 ( 
.A(n_95),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_94),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_83),
.Y(n_98)
);


endmodule