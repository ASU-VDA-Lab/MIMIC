module real_jpeg_26410_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_173;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_200;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_133;
wire n_138;
wire n_25;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

INVx3_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_1),
.A2(n_35),
.B1(n_36),
.B2(n_56),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_1),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_1),
.A2(n_56),
.B1(n_64),
.B2(n_74),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_1),
.A2(n_28),
.B1(n_31),
.B2(n_56),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_1),
.A2(n_48),
.B1(n_51),
.B2(n_56),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_3),
.A2(n_48),
.B1(n_51),
.B2(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_3),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_31),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_4),
.A2(n_27),
.B1(n_64),
.B2(n_74),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_4),
.A2(n_27),
.B1(n_35),
.B2(n_36),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_4),
.A2(n_27),
.B1(n_48),
.B2(n_51),
.Y(n_184)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx8_ASAP7_75t_SL g63 ( 
.A(n_6),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_7),
.A2(n_35),
.B1(n_36),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_7),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_7),
.A2(n_46),
.B1(n_48),
.B2(n_51),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g71 ( 
.A(n_10),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_10),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_10),
.B(n_66),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_10),
.B(n_36),
.C(n_37),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_10),
.A2(n_28),
.B1(n_31),
.B2(n_71),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_10),
.B(n_40),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_10),
.A2(n_35),
.B1(n_36),
.B2(n_71),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_10),
.B(n_48),
.C(n_50),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_10),
.A2(n_81),
.B(n_172),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_11),
.A2(n_48),
.B1(n_51),
.B2(n_89),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_11),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_13),
.A2(n_48),
.B1(n_51),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_13),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_13),
.A2(n_35),
.B1(n_36),
.B2(n_85),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_14),
.A2(n_28),
.B1(n_31),
.B2(n_42),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_14),
.A2(n_35),
.B1(n_36),
.B2(n_42),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_14),
.A2(n_42),
.B1(n_48),
.B2(n_51),
.Y(n_171)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_15),
.Y(n_82)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_15),
.Y(n_87)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_15),
.Y(n_101)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_15),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_128),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_126),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_102),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_20),
.B(n_102),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_78),
.C(n_92),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_21),
.A2(n_22),
.B1(n_210),
.B2(n_211),
.Y(n_209)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_57),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_43),
.B2(n_44),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_25),
.B(n_43),
.C(n_57),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_32),
.B1(n_40),
.B2(n_41),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_26),
.Y(n_94)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_28),
.A2(n_31),
.B1(n_37),
.B2(n_38),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_28),
.A2(n_31),
.B1(n_61),
.B2(n_62),
.Y(n_66)
);

NAND2xp33_ASAP7_75t_SL g91 ( 
.A(n_28),
.B(n_61),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_28),
.B(n_134),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI32xp33_ASAP7_75t_L g90 ( 
.A1(n_31),
.A2(n_62),
.A3(n_64),
.B1(n_73),
.B2(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_32),
.B(n_96),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_33),
.A2(n_107),
.B(n_108),
.Y(n_106)
);

OAI21xp33_ASAP7_75t_L g148 ( 
.A1(n_33),
.A2(n_108),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_39),
.Y(n_33)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_34),
.A2(n_94),
.B(n_95),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_35),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_34)
);

OAI22xp33_ASAP7_75t_L g54 ( 
.A1(n_35),
.A2(n_36),
.B1(n_49),
.B2(n_50),
.Y(n_54)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_36),
.B(n_179),
.Y(n_178)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_40),
.B(n_96),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_41),
.Y(n_107)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_47),
.B(n_52),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_45),
.A2(n_47),
.B1(n_123),
.B2(n_124),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_47),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_47),
.A2(n_52),
.B(n_144),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_47),
.B(n_71),
.Y(n_191)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_47)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_48),
.B(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_51),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_53),
.B(n_55),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_53),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_53),
.A2(n_143),
.B1(n_145),
.B2(n_146),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_55),
.B(n_146),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_67),
.B(n_76),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_58),
.B(n_113),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_65),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_62),
.B2(n_64),
.Y(n_59)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_60),
.Y(n_75)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_65),
.A2(n_110),
.B(n_112),
.Y(n_109)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

OAI21xp33_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_71),
.B(n_72),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_71),
.B(n_120),
.Y(n_196)
);

INVxp33_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_78),
.B(n_92),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_90),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_90),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_83),
.B1(n_86),
.B2(n_88),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_80),
.A2(n_183),
.B1(n_185),
.B2(n_186),
.Y(n_182)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_81),
.A2(n_84),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_81),
.A2(n_117),
.B1(n_118),
.B2(n_120),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_81),
.B(n_141),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_81),
.A2(n_171),
.B(n_172),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_86),
.B(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_87),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_88),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_97),
.C(n_99),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_93),
.B(n_153),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_97),
.A2(n_98),
.B1(n_99),
.B2(n_154),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_99),
.Y(n_154)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_101),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_114),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_109),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_125),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_122),
.Y(n_115)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_123),
.A2(n_159),
.B(n_160),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_123),
.A2(n_160),
.B(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_208),
.B(n_213),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_161),
.B(n_207),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_150),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_131),
.B(n_150),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_142),
.C(n_147),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_132),
.B(n_203),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_133),
.B(n_135),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_135),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_137),
.B(n_140),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_139),
.A2(n_184),
.B(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_140),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_141),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_142),
.A2(n_147),
.B1(n_148),
.B2(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_142),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_145),
.Y(n_159)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_151),
.A2(n_152),
.B1(n_155),
.B2(n_156),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_151),
.B(n_157),
.C(n_158),
.Y(n_212)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_201),
.B(n_206),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_180),
.B(n_200),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_164),
.B(n_174),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_164),
.B(n_174),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_170),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_166),
.B(n_169),
.C(n_170),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_171),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_178),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_175),
.A2(n_176),
.B1(n_178),
.B2(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_178),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_189),
.B(n_199),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_187),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_182),
.B(n_187),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_194),
.B(n_198),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_191),
.B(n_192),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_197),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_205),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_202),
.B(n_205),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_212),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_212),
.Y(n_213)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);


endmodule