module real_jpeg_19441_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_344, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_344;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_0),
.A2(n_23),
.B1(n_25),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_0),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_0),
.A2(n_47),
.B1(n_48),
.B2(n_58),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_0),
.A2(n_41),
.B1(n_42),
.B2(n_58),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_0),
.A2(n_27),
.B1(n_29),
.B2(n_58),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_1),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_1),
.B(n_26),
.Y(n_153)
);

AOI21xp33_ASAP7_75t_L g174 ( 
.A1(n_1),
.A2(n_14),
.B(n_48),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_1),
.A2(n_41),
.B1(n_42),
.B2(n_123),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_1),
.A2(n_95),
.B1(n_132),
.B2(n_183),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_1),
.B(n_77),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_1),
.B(n_29),
.Y(n_209)
);

AOI21xp33_ASAP7_75t_L g213 ( 
.A1(n_1),
.A2(n_29),
.B(n_209),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_2),
.A2(n_23),
.B1(n_25),
.B2(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_2),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_2),
.A2(n_27),
.B1(n_29),
.B2(n_125),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_2),
.A2(n_41),
.B1(n_42),
.B2(n_125),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_2),
.A2(n_47),
.B1(n_48),
.B2(n_125),
.Y(n_183)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_4),
.A2(n_24),
.B1(n_41),
.B2(n_42),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_4),
.A2(n_24),
.B1(n_27),
.B2(n_29),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_4),
.A2(n_24),
.B1(n_47),
.B2(n_48),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_5),
.B(n_47),
.Y(n_96)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_5),
.Y(n_102)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_5),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_5),
.B(n_201),
.Y(n_200)
);

BUFx8_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_7),
.A2(n_23),
.B1(n_25),
.B2(n_56),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_7),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_7),
.A2(n_41),
.B1(n_42),
.B2(n_56),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_7),
.A2(n_47),
.B1(n_48),
.B2(n_56),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_7),
.A2(n_27),
.B1(n_29),
.B2(n_56),
.Y(n_274)
);

OAI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_8),
.A2(n_23),
.B1(n_25),
.B2(n_32),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_8),
.A2(n_27),
.B1(n_29),
.B2(n_32),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_8),
.A2(n_32),
.B1(n_47),
.B2(n_48),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_8),
.A2(n_32),
.B1(n_41),
.B2(n_42),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_9),
.A2(n_27),
.B1(n_29),
.B2(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_9),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_9),
.A2(n_23),
.B1(n_25),
.B2(n_118),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_9),
.A2(n_47),
.B1(n_48),
.B2(n_118),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_9),
.A2(n_41),
.B1(n_42),
.B2(n_118),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_11),
.A2(n_27),
.B1(n_29),
.B2(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_11),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_11),
.A2(n_47),
.B1(n_48),
.B2(n_120),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_11),
.A2(n_41),
.B1(n_42),
.B2(n_120),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_11),
.A2(n_23),
.B1(n_25),
.B2(n_120),
.Y(n_257)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_12),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_14),
.A2(n_41),
.B(n_45),
.C(n_46),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_14),
.B(n_41),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_14),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g49 ( 
.A(n_14),
.Y(n_49)
);

INVx11_ASAP7_75t_SL g44 ( 
.A(n_15),
.Y(n_44)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_20),
.C(n_341),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_83),
.B(n_339),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_35),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_20),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_30),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_21),
.A2(n_54),
.B(n_257),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_26),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_22),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_22),
.A2(n_26),
.B(n_33),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_23),
.Y(n_25)
);

O2A1O1Ixp33_ASAP7_75t_L g33 ( 
.A1(n_23),
.A2(n_26),
.B(n_28),
.C(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_28),
.Y(n_34)
);

HAxp5_ASAP7_75t_SL g122 ( 
.A(n_23),
.B(n_123),
.CON(n_122),
.SN(n_122)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_26),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_26),
.B(n_31),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_26),
.A2(n_33),
.B1(n_122),
.B2(n_124),
.Y(n_121)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_27),
.A2(n_34),
.B1(n_122),
.B2(n_129),
.Y(n_128)
);

AOI32xp33_ASAP7_75t_L g208 ( 
.A1(n_27),
.A2(n_41),
.A3(n_67),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_28),
.B(n_29),
.Y(n_129)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_29),
.A2(n_64),
.B(n_65),
.C(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_29),
.B(n_65),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_30),
.A2(n_55),
.B(n_59),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_33),
.Y(n_30)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_33),
.A2(n_80),
.B(n_81),
.Y(n_79)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_36),
.B(n_340),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_75),
.C(n_79),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_37),
.A2(n_38),
.B1(n_335),
.B2(n_337),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_52),
.C(n_60),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_39),
.A2(n_315),
.B1(n_316),
.B2(n_317),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_39),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_39),
.A2(n_60),
.B1(n_61),
.B2(n_315),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_46),
.B(n_50),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_40),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_40),
.A2(n_50),
.B(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_40),
.A2(n_46),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_40),
.A2(n_46),
.B1(n_178),
.B2(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_40),
.A2(n_46),
.B1(n_198),
.B2(n_216),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_40),
.A2(n_216),
.B(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_40),
.A2(n_46),
.B1(n_105),
.B2(n_249),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_40),
.A2(n_113),
.B(n_249),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_41),
.A2(n_42),
.B1(n_65),
.B2(n_67),
.Y(n_64)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_42),
.A2(n_49),
.B(n_123),
.C(n_174),
.Y(n_173)
);

NAND2xp33_ASAP7_75t_SL g210 ( 
.A(n_42),
.B(n_65),
.Y(n_210)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_46),
.A2(n_105),
.B(n_106),
.Y(n_104)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_46),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_46),
.B(n_123),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_47),
.B(n_187),
.Y(n_186)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_51),
.B(n_114),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_52),
.A2(n_53),
.B1(n_323),
.B2(n_324),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_57),
.B2(n_59),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_54),
.A2(n_59),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_54),
.A2(n_59),
.B1(n_137),
.B2(n_257),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_54),
.A2(n_82),
.B(n_303),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_57),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_69),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_63),
.A2(n_70),
.B(n_140),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_68),
.Y(n_63)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_64),
.A2(n_71),
.B1(n_117),
.B2(n_119),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_64),
.A2(n_71),
.B1(n_156),
.B2(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_64),
.B(n_74),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_64),
.A2(n_69),
.B(n_274),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_64),
.A2(n_71),
.B1(n_274),
.B2(n_295),
.Y(n_294)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_65),
.Y(n_67)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_68),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_70),
.B(n_73),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_70),
.A2(n_77),
.B(n_78),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_70),
.A2(n_77),
.B1(n_155),
.B2(n_157),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_70),
.A2(n_78),
.B(n_260),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_70),
.A2(n_260),
.B(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_75),
.A2(n_76),
.B1(n_79),
.B2(n_336),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_79),
.Y(n_336)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_332),
.B(n_338),
.Y(n_83)
);

OAI321xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_308),
.A3(n_327),
.B1(n_330),
.B2(n_331),
.C(n_344),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_287),
.B(n_307),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_265),
.B(n_286),
.Y(n_86)
);

O2A1O1Ixp33_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_158),
.B(n_240),
.C(n_264),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_142),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_89),
.B(n_142),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_126),
.B2(n_141),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_110),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_92),
.B(n_110),
.C(n_141),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_104),
.B2(n_109),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_93),
.B(n_109),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_97),
.B(n_98),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_95),
.A2(n_97),
.B1(n_131),
.B2(n_132),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_95),
.A2(n_102),
.B1(n_167),
.B2(n_183),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_95),
.A2(n_170),
.B(n_200),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_95),
.A2(n_102),
.B(n_282),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_96),
.B(n_152),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_96),
.A2(n_166),
.B1(n_168),
.B2(n_169),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_96),
.A2(n_99),
.B(n_201),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_103),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_102),
.B(n_123),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_103),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_104),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_106),
.B(n_231),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_108),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_107),
.B(n_114),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_115),
.C(n_121),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_111),
.A2(n_112),
.B1(n_115),
.B2(n_116),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_117),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_119),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_121),
.B(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_124),
.Y(n_136)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_133),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_127),
.B(n_134),
.C(n_139),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_130),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_130),
.Y(n_146)
);

OAI21x1_ASAP7_75t_SL g150 ( 
.A1(n_131),
.A2(n_132),
.B(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_132),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_138),
.B2(n_139),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_145),
.C(n_147),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_143),
.B(n_237),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_145),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_153),
.C(n_154),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_149),
.A2(n_150),
.B1(n_153),
.B2(n_227),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_151),
.B(n_200),
.Y(n_247)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_153),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_154),
.B(n_226),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_239),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_234),
.B(n_238),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_221),
.B(n_233),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_162),
.A2(n_203),
.B(n_220),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_163),
.A2(n_190),
.B(n_202),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_179),
.B(n_189),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_171),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_165),
.B(n_171),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_175),
.B2(n_176),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_173),
.B(n_175),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_184),
.B(n_188),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_182),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_191),
.B(n_192),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_199),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_197),
.C(n_199),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_201),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_204),
.B(n_205),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_211),
.B1(n_218),
.B2(n_219),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_206),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_207),
.B(n_208),
.Y(n_232)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_211),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_214),
.B1(n_215),
.B2(n_217),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_212),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_217),
.C(n_218),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_215),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_222),
.B(n_223),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_225),
.B1(n_228),
.B2(n_229),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_224),
.B(n_230),
.C(n_232),
.Y(n_235)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

XOR2x2_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_232),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_235),
.B(n_236),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_241),
.B(n_242),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_262),
.B2(n_263),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_250),
.B2(n_251),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_251),
.C(n_263),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_246),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_247),
.B(n_248),
.Y(n_271)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_254),
.B2(n_261),
.Y(n_251)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_252),
.Y(n_261)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_258),
.B2(n_259),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_255),
.B(n_259),
.C(n_261),
.Y(n_285)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_262),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_266),
.B(n_267),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_285),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_269),
.A2(n_270),
.B1(n_278),
.B2(n_279),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_279),
.C(n_285),
.Y(n_288)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_271),
.B(n_275),
.C(n_277),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_275),
.B1(n_276),
.B2(n_277),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_273),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_276),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_283),
.B2(n_284),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_280),
.A2(n_281),
.B1(n_302),
.B2(n_304),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_280),
.A2(n_298),
.B(n_302),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_283),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_283),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_288),
.B(n_289),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_305),
.B2(n_306),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_297),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_292),
.B(n_297),
.C(n_306),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_294),
.B(n_296),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_293),
.B(n_294),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_295),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_310),
.C(n_319),
.Y(n_309)
);

FAx1_ASAP7_75t_SL g329 ( 
.A(n_296),
.B(n_310),
.CI(n_319),
.CON(n_329),
.SN(n_329)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_299),
.B1(n_300),
.B2(n_301),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_302),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_305),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_320),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_309),
.B(n_320),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_312),
.B1(n_313),
.B2(n_314),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_311),
.A2(n_312),
.B1(n_322),
.B2(n_325),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_312),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_315),
.C(n_317),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_312),
.B(n_325),
.C(n_326),
.Y(n_333)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_317),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_326),
.Y(n_320)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_322),
.Y(n_325)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_328),
.B(n_329),
.Y(n_330)
);

BUFx24_ASAP7_75t_SL g342 ( 
.A(n_329),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_333),
.B(n_334),
.Y(n_338)
);

CKINVDCx14_ASAP7_75t_R g337 ( 
.A(n_335),
.Y(n_337)
);


endmodule