module fake_netlist_1_3214_n_30 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_30);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_30;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
AND2x2_ASAP7_75t_SL g13 ( .A(n_3), .B(n_8), .Y(n_13) );
AND2x6_ASAP7_75t_L g14 ( .A(n_7), .B(n_0), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_5), .B(n_11), .Y(n_15) );
INVx3_ASAP7_75t_L g16 ( .A(n_12), .Y(n_16) );
OAI22xp5_ASAP7_75t_SL g17 ( .A1(n_4), .A2(n_0), .B1(n_6), .B2(n_9), .Y(n_17) );
NAND2xp33_ASAP7_75t_R g18 ( .A(n_16), .B(n_10), .Y(n_18) );
INVx2_ASAP7_75t_L g19 ( .A(n_14), .Y(n_19) );
NAND2xp5_ASAP7_75t_SL g20 ( .A(n_19), .B(n_13), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_18), .B(n_14), .Y(n_21) );
NOR2xp33_ASAP7_75t_L g22 ( .A(n_21), .B(n_15), .Y(n_22) );
INVx1_ASAP7_75t_SL g23 ( .A(n_22), .Y(n_23) );
AND2x2_ASAP7_75t_L g24 ( .A(n_23), .B(n_20), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_24), .B(n_14), .Y(n_25) );
AOI21xp33_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_17), .B(n_1), .Y(n_26) );
OR2x6_ASAP7_75t_L g27 ( .A(n_26), .B(n_1), .Y(n_27) );
INVx2_ASAP7_75t_L g28 ( .A(n_27), .Y(n_28) );
CKINVDCx20_ASAP7_75t_R g29 ( .A(n_28), .Y(n_29) );
AOI21xp5_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_2), .B(n_28), .Y(n_30) );
endmodule