module real_jpeg_33628_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_657;
wire n_643;
wire n_656;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_669;
wire n_376;
wire n_354;
wire n_136;
wire n_679;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_666;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_685;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_680;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_678;
wire n_30;
wire n_328;
wire n_149;
wire n_620;
wire n_332;
wire n_366;
wire n_456;
wire n_578;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_682;
wire n_422;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_684;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_673;
wire n_631;
wire n_175;
wire n_338;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_470;
wire n_219;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_195;
wire n_110;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_615;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_670;
wire n_524;
wire n_589;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_638;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_316;
wire n_307;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_572;
wire n_155;
wire n_405;
wire n_412;
wire n_586;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_377;
wire n_616;
wire n_686;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_667;
wire n_330;
wire n_298;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_683;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_677;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_675;
wire n_179;
wire n_138;
wire n_662;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_358;
wire n_181;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_681;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_568;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_660;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g231 ( 
.A(n_0),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_0),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g619 ( 
.A(n_0),
.Y(n_619)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_1),
.A2(n_68),
.B1(n_383),
.B2(n_384),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_1),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_1),
.A2(n_383),
.B1(n_445),
.B2(n_450),
.Y(n_444)
);

AOI22xp33_ASAP7_75t_SL g568 ( 
.A1(n_1),
.A2(n_383),
.B1(n_569),
.B2(n_572),
.Y(n_568)
);

AOI22xp33_ASAP7_75t_SL g608 ( 
.A1(n_1),
.A2(n_383),
.B1(n_609),
.B2(n_615),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_3),
.A2(n_172),
.B1(n_274),
.B2(n_275),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_3),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_3),
.A2(n_274),
.B1(n_390),
.B2(n_392),
.Y(n_389)
);

AOI22xp33_ASAP7_75t_SL g547 ( 
.A1(n_3),
.A2(n_205),
.B1(n_274),
.B2(n_548),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_SL g589 ( 
.A1(n_3),
.A2(n_274),
.B1(n_590),
.B2(n_595),
.Y(n_589)
);

OAI22xp33_ASAP7_75t_R g56 ( 
.A1(n_4),
.A2(n_57),
.B1(n_61),
.B2(n_63),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_4),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_4),
.A2(n_63),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_4),
.A2(n_63),
.B1(n_158),
.B2(n_183),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_4),
.A2(n_63),
.B1(n_235),
.B2(n_237),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_5),
.A2(n_252),
.B1(n_256),
.B2(n_257),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_5),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_5),
.A2(n_214),
.B1(n_256),
.B2(n_397),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_5),
.A2(n_256),
.B1(n_431),
.B2(n_433),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_5),
.A2(n_256),
.B1(n_543),
.B2(n_544),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_6),
.B(n_372),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_6),
.Y(n_442)
);

NAND2xp33_ASAP7_75t_SL g475 ( 
.A(n_6),
.B(n_28),
.Y(n_475)
);

OAI32xp33_ASAP7_75t_L g521 ( 
.A1(n_6),
.A2(n_522),
.A3(n_524),
.B1(n_528),
.B2(n_534),
.Y(n_521)
);

OAI32xp33_ASAP7_75t_L g566 ( 
.A1(n_6),
.A2(n_522),
.A3(n_524),
.B1(n_528),
.B2(n_534),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_SL g574 ( 
.A1(n_6),
.A2(n_442),
.B1(n_575),
.B2(n_576),
.Y(n_574)
);

OAI21xp33_ASAP7_75t_L g654 ( 
.A1(n_6),
.A2(n_225),
.B(n_600),
.Y(n_654)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_7),
.A2(n_163),
.B1(n_164),
.B2(n_166),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_7),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_7),
.A2(n_163),
.B1(n_282),
.B2(n_285),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_7),
.A2(n_163),
.B1(n_408),
.B2(n_409),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_7),
.A2(n_163),
.B1(n_466),
.B2(n_470),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_8),
.A2(n_58),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_8),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_8),
.A2(n_170),
.B1(n_214),
.B2(n_216),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_8),
.A2(n_170),
.B1(n_300),
.B2(n_305),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_8),
.A2(n_170),
.B1(n_342),
.B2(n_345),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_9),
.Y(n_177)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_10),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_10),
.Y(n_131)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_11),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_11),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_11),
.Y(n_291)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_11),
.Y(n_614)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_12),
.Y(n_86)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_12),
.Y(n_96)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_12),
.Y(n_106)
);

CKINVDCx11_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_13),
.B(n_685),
.Y(n_684)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_14),
.A2(n_66),
.B1(n_67),
.B2(n_69),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_14),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_14),
.A2(n_66),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_14),
.A2(n_66),
.B1(n_205),
.B2(n_209),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_14),
.A2(n_66),
.B1(n_289),
.B2(n_292),
.Y(n_288)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_15),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_15),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_15),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_15),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_16),
.A2(n_20),
.B(n_23),
.Y(n_19)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_17),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_17),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_18),
.A2(n_145),
.B1(n_150),
.B2(n_151),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_18),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_18),
.A2(n_69),
.B1(n_150),
.B2(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_18),
.A2(n_150),
.B1(n_242),
.B2(n_245),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_18),
.A2(n_150),
.B1(n_356),
.B2(n_358),
.Y(n_355)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI21x1_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_73),
.B(n_684),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_64),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_26),
.B(n_686),
.Y(n_685)
);

OAI21xp33_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_43),
.B(n_56),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_27),
.A2(n_43),
.B1(n_56),
.B2(n_65),
.Y(n_64)
);

AO22x1_ASAP7_75t_L g161 ( 
.A1(n_27),
.A2(n_43),
.B1(n_162),
.B2(n_169),
.Y(n_161)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_27),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_27),
.A2(n_43),
.B1(n_65),
.B2(n_323),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_28),
.B(n_162),
.Y(n_259)
);

NAND2x1_ASAP7_75t_SL g271 ( 
.A(n_28),
.B(n_251),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_28),
.B(n_382),
.Y(n_381)
);

AO22x1_ASAP7_75t_L g417 ( 
.A1(n_28),
.A2(n_44),
.B1(n_273),
.B2(n_382),
.Y(n_417)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_34),
.B1(n_37),
.B2(n_39),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g137 ( 
.A(n_33),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_33),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_33),
.Y(n_159)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_34),
.Y(n_366)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_36),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_37),
.A2(n_135),
.B1(n_138),
.B2(n_141),
.Y(n_134)
);

INVx8_ASAP7_75t_L g215 ( 
.A(n_37),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx8_ASAP7_75t_L g394 ( 
.A(n_38),
.Y(n_394)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_43),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_44),
.B(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_44),
.B(n_273),
.Y(n_272)
);

OAI21xp33_ASAP7_75t_L g437 ( 
.A1(n_44),
.A2(n_371),
.B(n_438),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_49),
.B1(n_52),
.B2(n_54),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_47),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_48),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_48),
.Y(n_168)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_48),
.Y(n_255)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_59),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_60),
.Y(n_370)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_64),
.B(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_64),
.B(n_330),
.Y(n_683)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_64),
.Y(n_686)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_72),
.Y(n_258)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_72),
.Y(n_386)
);

OAI21x1_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_331),
.B(n_675),
.Y(n_73)
);

OR3x1_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_311),
.C(n_329),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_260),
.Y(n_75)
);

A2O1A1Ixp33_ASAP7_75t_L g678 ( 
.A1(n_76),
.A2(n_312),
.B(n_679),
.C(n_680),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_195),
.Y(n_76)
);

NOR3xp33_ASAP7_75t_L g680 ( 
.A(n_77),
.B(n_681),
.C(n_682),
.Y(n_680)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_178),
.Y(n_77)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_78),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_117),
.C(n_160),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_80),
.B(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_80),
.A2(n_117),
.B1(n_118),
.B2(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_80),
.Y(n_199)
);

OA21x2_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_97),
.B(n_112),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_81),
.A2(n_97),
.B1(n_112),
.B2(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_81),
.A2(n_97),
.B1(n_430),
.B2(n_435),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_81),
.B(n_430),
.Y(n_551)
);

INVx1_ASAP7_75t_SL g584 ( 
.A(n_81),
.Y(n_584)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_82),
.Y(n_240)
);

OAI22x1_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_87),
.B1(n_90),
.B2(n_94),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_89),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_89),
.Y(n_295)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_89),
.Y(n_348)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_89),
.Y(n_361)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_89),
.Y(n_469)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_90),
.Y(n_633)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_93),
.Y(n_236)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_93),
.Y(n_660)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_95),
.Y(n_625)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_96),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_97),
.B(n_644),
.Y(n_643)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_98),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_98),
.A2(n_204),
.B1(n_240),
.B2(n_241),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_98),
.A2(n_240),
.B1(n_241),
.B2(n_299),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_98),
.A2(n_240),
.B1(n_299),
.B2(n_407),
.Y(n_406)
);

OAI21xp33_ASAP7_75t_SL g546 ( 
.A1(n_98),
.A2(n_547),
.B(n_551),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_SL g567 ( 
.A1(n_98),
.A2(n_240),
.B1(n_547),
.B2(n_568),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_SL g583 ( 
.A1(n_98),
.A2(n_568),
.B1(n_584),
.B2(n_585),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_103),
.B1(n_107),
.B2(n_109),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_101),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_102),
.Y(n_539)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_106),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_109),
.Y(n_432)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_110),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_111),
.Y(n_211)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_111),
.Y(n_304)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_116),
.Y(n_244)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_144),
.B1(n_154),
.B2(n_156),
.Y(n_118)
);

AOI22x1_ASAP7_75t_L g443 ( 
.A1(n_119),
.A2(n_154),
.B1(n_444),
.B2(n_453),
.Y(n_443)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_120),
.A2(n_154),
.B1(n_156),
.B2(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_120),
.A2(n_144),
.B1(n_154),
.B2(n_213),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_120),
.A2(n_155),
.B1(n_213),
.B2(n_281),
.Y(n_280)
);

OAI21xp33_ASAP7_75t_SL g318 ( 
.A1(n_120),
.A2(n_182),
.B(n_319),
.Y(n_318)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_120),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_120),
.B(n_396),
.Y(n_463)
);

AND2x4_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_134),
.Y(n_120)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_121),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_125),
.B1(n_128),
.B2(n_132),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_126),
.Y(n_307)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_127),
.Y(n_133)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_127),
.Y(n_527)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_131),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_131),
.Y(n_533)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_137),
.Y(n_452)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_139),
.Y(n_138)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_148),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_149),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g284 ( 
.A(n_149),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_149),
.Y(n_449)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_153),
.Y(n_578)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_155),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_155),
.B(n_396),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_159),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_161),
.B(n_198),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_161),
.B(n_327),
.C(n_328),
.Y(n_326)
);

BUFx4f_ASAP7_75t_SL g164 ( 
.A(n_165),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_169),
.Y(n_189)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_175),
.Y(n_372)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_177),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_179),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_187),
.Y(n_179)
);

INVxp33_ASAP7_75t_L g316 ( 
.A(n_181),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_186),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_187),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_194),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_190),
.Y(n_323)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx11_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_221),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g682 ( 
.A(n_196),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_200),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_197),
.A2(n_200),
.B(n_222),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_197),
.B(n_309),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_SL g314 ( 
.A(n_199),
.B(n_315),
.C(n_316),
.Y(n_314)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_201),
.A2(n_202),
.B(n_212),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_201),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_212),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx4_ASAP7_75t_L g572 ( 
.A(n_207),
.Y(n_572)
);

INVx2_ASAP7_75t_SL g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_211),
.Y(n_408)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx8_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_220),
.Y(n_365)
);

INVxp67_ASAP7_75t_SL g681 ( 
.A(n_221),
.Y(n_681)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_222),
.B(n_310),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_238),
.B(n_249),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_223),
.A2(n_224),
.B1(n_249),
.B2(n_264),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_223),
.A2(n_224),
.B1(n_239),
.B2(n_499),
.Y(n_498)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_239),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_232),
.B(n_234),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_225),
.A2(n_234),
.B1(n_288),
.B2(n_296),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_225),
.A2(n_288),
.B1(n_402),
.B2(n_405),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_225),
.A2(n_341),
.B1(n_465),
.B2(n_471),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g588 ( 
.A1(n_225),
.A2(n_589),
.B(n_600),
.Y(n_588)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_226),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_226),
.A2(n_340),
.B1(n_349),
.B2(n_355),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_226),
.B(n_542),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_SL g606 ( 
.A1(n_226),
.A2(n_607),
.B1(n_618),
.B2(n_620),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx6_ASAP7_75t_L g357 ( 
.A(n_228),
.Y(n_357)
);

INVx4_ASAP7_75t_L g233 ( 
.A(n_229),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_231),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g540 ( 
.A1(n_232),
.A2(n_465),
.B(n_541),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_SL g652 ( 
.A1(n_232),
.A2(n_541),
.B(n_608),
.Y(n_652)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_236),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_239),
.Y(n_499)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_248),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_248),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_248),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_248),
.Y(n_638)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_249),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_259),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_250),
.B(n_381),
.Y(n_380)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_308),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_261),
.B(n_308),
.Y(n_679)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_265),
.C(n_267),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_262),
.B(n_484),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_266),
.B(n_268),
.Y(n_484)
);

INVxp67_ASAP7_75t_SL g267 ( 
.A(n_268),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_277),
.C(n_286),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_270),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_270),
.B(n_280),
.Y(n_492)
);

NAND2x1_ASAP7_75t_SL g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_271),
.B(n_437),
.Y(n_436)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

OAI21x1_ASAP7_75t_L g489 ( 
.A1(n_278),
.A2(n_490),
.B(n_492),
.Y(n_489)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_281),
.Y(n_416)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_284),
.Y(n_285)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_284),
.Y(n_397)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_286),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_298),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g419 ( 
.A(n_287),
.Y(n_419)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_291),
.Y(n_344)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_291),
.Y(n_594)
);

INVx4_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_295),
.Y(n_617)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_297),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_298),
.Y(n_420)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx4_ASAP7_75t_L g631 ( 
.A(n_304),
.Y(n_631)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVxp67_ASAP7_75t_SL g311 ( 
.A(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_326),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g677 ( 
.A(n_313),
.B(n_326),
.Y(n_677)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_317),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_314),
.B(n_322),
.C(n_324),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_318),
.A2(n_322),
.B1(n_324),
.B2(n_325),
.Y(n_317)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_318),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

OAI21x1_ASAP7_75t_L g461 ( 
.A1(n_320),
.A2(n_462),
.B(n_463),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

OAI22x1_ASAP7_75t_L g414 ( 
.A1(n_321),
.A2(n_388),
.B1(n_415),
.B2(n_416),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_321),
.B(n_442),
.Y(n_587)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_322),
.Y(n_325)
);

A2O1A1Ixp33_ASAP7_75t_L g676 ( 
.A1(n_329),
.A2(n_677),
.B(n_678),
.C(n_683),
.Y(n_676)
);

AND2x4_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_511),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_333),
.A2(n_480),
.B(n_505),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_421),
.C(n_454),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g513 ( 
.A1(n_335),
.A2(n_514),
.B(n_515),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_398),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_336),
.B(n_399),
.C(n_418),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_380),
.C(n_387),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

XNOR2x1_ASAP7_75t_L g423 ( 
.A(n_338),
.B(n_424),
.Y(n_423)
);

NOR2xp67_ASAP7_75t_SL g338 ( 
.A(n_339),
.B(n_362),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_339),
.B(n_362),
.Y(n_458)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_347),
.Y(n_470)
);

INVx4_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_349),
.B(n_542),
.Y(n_600)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_354),
.Y(n_404)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_354),
.Y(n_473)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_355),
.Y(n_405)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_357),
.Y(n_544)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_360),
.Y(n_543)
);

INVx4_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

AOI32xp33_ASAP7_75t_L g362 ( 
.A1(n_363),
.A2(n_366),
.A3(n_367),
.B1(n_371),
.B2(n_373),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx3_ASAP7_75t_SL g376 ( 
.A(n_365),
.Y(n_376)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx4_ASAP7_75t_SL g369 ( 
.A(n_370),
.Y(n_369)
);

NAND2xp33_ASAP7_75t_SL g373 ( 
.A(n_374),
.B(n_377),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g529 ( 
.A(n_376),
.Y(n_529)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

XNOR2x1_ASAP7_75t_L g424 ( 
.A(n_380),
.B(n_387),
.Y(n_424)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

OA21x2_ASAP7_75t_L g387 ( 
.A1(n_388),
.A2(n_389),
.B(n_395),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g573 ( 
.A1(n_388),
.A2(n_395),
.B(n_574),
.Y(n_573)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_389),
.Y(n_453)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_391),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx4_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_396),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_418),
.Y(n_398)
);

XNOR2x1_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_413),
.Y(n_399)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_400),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_406),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_401),
.B(n_406),
.Y(n_426)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_407),
.Y(n_435)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_411),
.Y(n_434)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

XNOR2x1_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_417),
.Y(n_413)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_414),
.Y(n_497)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_417),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_420),
.Y(n_418)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_421),
.Y(n_514)
);

MAJx2_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_425),
.C(n_427),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_422),
.A2(n_423),
.B1(n_477),
.B2(n_479),
.Y(n_476)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_425),
.A2(n_426),
.B1(n_428),
.B2(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_SL g478 ( 
.A(n_428),
.Y(n_478)
);

MAJx2_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_436),
.C(n_443),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_429),
.B(n_443),
.Y(n_457)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_430),
.Y(n_585)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g433 ( 
.A(n_434),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_436),
.B(n_457),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_442),
.Y(n_438)
);

INVx2_ASAP7_75t_SL g439 ( 
.A(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_442),
.B(n_535),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_442),
.B(n_628),
.Y(n_627)
);

OAI21xp33_ASAP7_75t_SL g644 ( 
.A1(n_442),
.A2(n_627),
.B(n_645),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_SL g651 ( 
.A(n_442),
.B(n_584),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_442),
.B(n_657),
.Y(n_656)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_444),
.Y(n_462)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

OR2x2_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_476),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_455),
.B(n_476),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_458),
.C(n_459),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_456),
.B(n_557),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_458),
.B(n_460),
.Y(n_557)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_464),
.C(n_474),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_461),
.B(n_554),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_464),
.A2(n_474),
.B1(n_475),
.B2(n_555),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_464),
.Y(n_555)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_467),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

BUFx12f_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_477),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_481),
.B(n_513),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_SL g481 ( 
.A1(n_482),
.A2(n_485),
.B(n_500),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_482),
.B(n_485),
.Y(n_510)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g509 ( 
.A(n_483),
.B(n_486),
.Y(n_509)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_494),
.C(n_498),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

XNOR2x1_ASAP7_75t_L g502 ( 
.A(n_488),
.B(n_503),
.Y(n_502)
);

XNOR2x1_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_493),
.Y(n_488)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_494),
.B(n_502),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_496),
.C(n_497),
.Y(n_494)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_498),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_501),
.B(n_504),
.Y(n_500)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_501),
.Y(n_508)
);

INVxp33_ASAP7_75t_SL g507 ( 
.A(n_504),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g505 ( 
.A1(n_506),
.A2(n_509),
.B(n_510),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_508),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_516),
.Y(n_511)
);

OAI21x1_ASAP7_75t_L g516 ( 
.A1(n_517),
.A2(n_558),
.B(n_673),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_518),
.B(n_556),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_519),
.B(n_674),
.Y(n_673)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_520),
.B(n_545),
.C(n_552),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_L g562 ( 
.A1(n_520),
.A2(n_545),
.B1(n_546),
.B2(n_563),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_520),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_521),
.B(n_540),
.Y(n_520)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVx4_ASAP7_75t_L g575 ( 
.A(n_523),
.Y(n_575)
);

BUFx2_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_529),
.B(n_530),
.Y(n_528)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

BUFx3_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_538),
.Y(n_647)
);

INVx5_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g565 ( 
.A(n_540),
.B(n_566),
.Y(n_565)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

INVx2_ASAP7_75t_SL g548 ( 
.A(n_549),
.Y(n_548)
);

INVx4_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_551),
.B(n_643),
.Y(n_642)
);

INVxp67_ASAP7_75t_L g552 ( 
.A(n_553),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_553),
.B(n_562),
.Y(n_561)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_556),
.Y(n_674)
);

AOI21x1_ASAP7_75t_L g558 ( 
.A1(n_559),
.A2(n_601),
.B(n_672),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_560),
.B(n_579),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_561),
.B(n_564),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_561),
.B(n_564),
.Y(n_672)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_565),
.B(n_567),
.C(n_573),
.Y(n_564)
);

XOR2xp5_ASAP7_75t_L g580 ( 
.A(n_565),
.B(n_581),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_L g581 ( 
.A(n_567),
.B(n_573),
.Y(n_581)
);

INVx2_ASAP7_75t_SL g569 ( 
.A(n_570),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_571),
.Y(n_570)
);

HB1xp67_ASAP7_75t_L g576 ( 
.A(n_577),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_578),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_580),
.B(n_582),
.Y(n_579)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_580),
.Y(n_670)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_582),
.Y(n_669)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_583),
.B(n_586),
.C(n_588),
.Y(n_582)
);

XNOR2xp5_ASAP7_75t_L g665 ( 
.A(n_583),
.B(n_587),
.Y(n_665)
);

HB1xp67_ASAP7_75t_L g586 ( 
.A(n_587),
.Y(n_586)
);

XOR2xp5_ASAP7_75t_L g664 ( 
.A(n_588),
.B(n_665),
.Y(n_664)
);

INVxp67_ASAP7_75t_L g620 ( 
.A(n_589),
.Y(n_620)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_591),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_591),
.B(n_624),
.Y(n_623)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_592),
.Y(n_591)
);

INVx4_ASAP7_75t_L g592 ( 
.A(n_593),
.Y(n_592)
);

INVx4_ASAP7_75t_L g593 ( 
.A(n_594),
.Y(n_593)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_594),
.Y(n_599)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_596),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_597),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_598),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_599),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_602),
.B(n_668),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_603),
.B(n_663),
.Y(n_602)
);

OAI21x1_ASAP7_75t_L g603 ( 
.A1(n_604),
.A2(n_648),
.B(n_662),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_605),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_606),
.B(n_621),
.Y(n_605)
);

OR2x2_ASAP7_75t_L g662 ( 
.A(n_606),
.B(n_621),
.Y(n_662)
);

INVxp67_ASAP7_75t_L g607 ( 
.A(n_608),
.Y(n_607)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_610),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_611),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_612),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_613),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_614),
.Y(n_613)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_616),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_617),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g618 ( 
.A(n_619),
.Y(n_618)
);

INVx5_ASAP7_75t_L g657 ( 
.A(n_619),
.Y(n_657)
);

XNOR2xp5_ASAP7_75t_L g621 ( 
.A(n_622),
.B(n_642),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_622),
.B(n_642),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_L g622 ( 
.A1(n_623),
.A2(n_626),
.B1(n_632),
.B2(n_634),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g624 ( 
.A(n_625),
.Y(n_624)
);

INVxp67_ASAP7_75t_L g626 ( 
.A(n_627),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_629),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_630),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_631),
.Y(n_630)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_633),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_635),
.B(n_639),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_636),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_637),
.Y(n_636)
);

HB1xp67_ASAP7_75t_L g637 ( 
.A(n_638),
.Y(n_637)
);

BUFx2_ASAP7_75t_L g639 ( 
.A(n_640),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_641),
.Y(n_640)
);

BUFx2_ASAP7_75t_L g645 ( 
.A(n_646),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_647),
.Y(n_646)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_649),
.Y(n_648)
);

OAI21xp5_ASAP7_75t_L g649 ( 
.A1(n_650),
.A2(n_653),
.B(n_661),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_651),
.B(n_652),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_651),
.B(n_652),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_654),
.B(n_655),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_SL g655 ( 
.A(n_656),
.B(n_658),
.Y(n_655)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_659),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_660),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_664),
.B(n_666),
.Y(n_663)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_664),
.Y(n_671)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_667),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_667),
.A2(n_669),
.B1(n_670),
.B2(n_671),
.Y(n_668)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_676),
.Y(n_675)
);


endmodule