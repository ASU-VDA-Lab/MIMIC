module fake_jpeg_29077_n_410 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_410);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_410;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx4f_ASAP7_75t_SL g23 ( 
.A(n_4),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_18),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_19),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_48),
.Y(n_114)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_49),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_26),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_50),
.B(n_58),
.Y(n_87)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_51),
.Y(n_91)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_52),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_54),
.Y(n_120)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_26),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_59),
.Y(n_130)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_60),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_26),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_61),
.B(n_68),
.Y(n_122)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_62),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_24),
.B(n_19),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_63),
.B(n_69),
.Y(n_110)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_64),
.Y(n_132)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_66),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_24),
.B(n_0),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_67),
.B(n_75),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_26),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_28),
.B(n_35),
.C(n_38),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

INVx3_ASAP7_75t_SL g116 ( 
.A(n_70),
.Y(n_116)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_31),
.B(n_19),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_74),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_26),
.B(n_0),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_32),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_32),
.Y(n_76)
);

CKINVDCx5p33_ASAP7_75t_R g107 ( 
.A(n_76),
.Y(n_107)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_40),
.Y(n_78)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_79),
.Y(n_99)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_31),
.B(n_37),
.Y(n_81)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_32),
.Y(n_82)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_85),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_37),
.B(n_18),
.Y(n_86)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_86),
.Y(n_124)
);

INVx5_ASAP7_75t_SL g89 ( 
.A(n_55),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_89),
.B(n_111),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_73),
.A2(n_47),
.B1(n_42),
.B2(n_43),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_97),
.A2(n_103),
.B1(n_105),
.B2(n_108),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_67),
.A2(n_22),
.B1(n_34),
.B2(n_36),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_54),
.A2(n_47),
.B1(n_43),
.B2(n_42),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_74),
.A2(n_34),
.B1(n_36),
.B2(n_41),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_117),
.B1(n_45),
.B2(n_84),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_57),
.A2(n_36),
.B1(n_34),
.B2(n_40),
.Y(n_108)
);

INVx4_ASAP7_75t_SL g111 ( 
.A(n_60),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_69),
.A2(n_41),
.B1(n_46),
.B2(n_30),
.Y(n_117)
);

OA22x2_ASAP7_75t_L g118 ( 
.A1(n_62),
.A2(n_42),
.B1(n_43),
.B2(n_47),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_118),
.A2(n_126),
.B1(n_129),
.B2(n_76),
.Y(n_151)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_71),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_125),
.B(n_128),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_80),
.A2(n_46),
.B1(n_25),
.B2(n_30),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_79),
.A2(n_25),
.B1(n_45),
.B2(n_32),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_61),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_134),
.B(n_143),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_110),
.B(n_77),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_151),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_137),
.A2(n_139),
.B1(n_116),
.B2(n_115),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_118),
.A2(n_85),
.B1(n_83),
.B2(n_53),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_90),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_140),
.Y(n_199)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_101),
.Y(n_141)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_141),
.Y(n_187)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_89),
.Y(n_142)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_142),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_94),
.B(n_82),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_87),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_147),
.Y(n_171)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_88),
.Y(n_145)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_145),
.Y(n_193)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_146),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_107),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_150),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_98),
.Y(n_149)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_149),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_75),
.Y(n_150)
);

A2O1A1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_133),
.A2(n_68),
.B(n_50),
.C(n_58),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_152),
.B(n_167),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_120),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_153),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_49),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_154),
.B(n_155),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_100),
.B(n_52),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_112),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_156),
.Y(n_177)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_95),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_158),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_111),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_102),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_160),
.Y(n_182)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_113),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_123),
.Y(n_162)
);

INVxp33_ASAP7_75t_L g198 ( 
.A(n_162),
.Y(n_198)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_96),
.Y(n_163)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_163),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_124),
.B(n_23),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_164),
.B(n_166),
.Y(n_190)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_95),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_165),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_126),
.B(n_23),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_119),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_114),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_168),
.A2(n_169),
.B1(n_170),
.B2(n_116),
.Y(n_183)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_127),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_99),
.Y(n_170)
);

OAI22x1_ASAP7_75t_L g172 ( 
.A1(n_138),
.A2(n_105),
.B1(n_97),
.B2(n_129),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_172),
.A2(n_151),
.B1(n_144),
.B2(n_156),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_138),
.A2(n_51),
.B1(n_56),
.B2(n_91),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_176),
.A2(n_192),
.B1(n_142),
.B2(n_136),
.Y(n_214)
);

OAI21xp33_ASAP7_75t_SL g180 ( 
.A1(n_134),
.A2(n_93),
.B(n_115),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_180),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_135),
.B(n_93),
.C(n_99),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_155),
.C(n_168),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_183),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_185),
.A2(n_197),
.B1(n_121),
.B2(n_149),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_154),
.A2(n_91),
.B1(n_104),
.B2(n_98),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_152),
.B(n_32),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_194),
.B(n_135),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_154),
.A2(n_104),
.B1(n_121),
.B2(n_130),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_200),
.A2(n_215),
.B1(n_172),
.B2(n_192),
.Y(n_235)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_193),
.Y(n_201)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_201),
.Y(n_238)
);

A2O1A1O1Ixp25_ASAP7_75t_L g237 ( 
.A1(n_202),
.A2(n_211),
.B(n_219),
.C(n_182),
.D(n_187),
.Y(n_237)
);

NOR2x1p5_ASAP7_75t_L g203 ( 
.A(n_173),
.B(n_143),
.Y(n_203)
);

AND2x2_ASAP7_75t_SL g233 ( 
.A(n_203),
.B(n_188),
.Y(n_233)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_193),
.Y(n_204)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_204),
.Y(n_243)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_195),
.Y(n_205)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_205),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_184),
.B(n_147),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_207),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_174),
.B(n_161),
.Y(n_207)
);

MAJx2_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_181),
.C(n_188),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_184),
.B(n_161),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_210),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_186),
.B(n_145),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_186),
.B(n_155),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_171),
.B(n_146),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_212),
.B(n_177),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_136),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_213),
.B(n_218),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_214),
.A2(n_197),
.B1(n_185),
.B2(n_220),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_172),
.A2(n_153),
.B1(n_131),
.B2(n_114),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_195),
.Y(n_216)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_216),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_173),
.A2(n_160),
.B(n_158),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_217),
.A2(n_188),
.B(n_178),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_173),
.B(n_140),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_171),
.B(n_141),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_174),
.B(n_163),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_221),
.B(n_222),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_177),
.B(n_159),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_224),
.A2(n_196),
.B1(n_199),
.B2(n_162),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_225),
.A2(n_239),
.B1(n_223),
.B2(n_218),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_212),
.B(n_190),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_226),
.B(n_23),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_244),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_219),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_230),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_211),
.C(n_208),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_233),
.B(n_217),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_234),
.A2(n_217),
.B(n_203),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_235),
.A2(n_206),
.B(n_202),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_200),
.A2(n_176),
.B1(n_190),
.B2(n_178),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_236),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_213),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_214),
.A2(n_182),
.B1(n_179),
.B2(n_191),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_215),
.A2(n_149),
.B1(n_175),
.B2(n_167),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_224),
.A2(n_175),
.B1(n_169),
.B2(n_191),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_201),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_203),
.A2(n_187),
.B1(n_130),
.B2(n_170),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_222),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_209),
.B(n_198),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_248),
.B(n_207),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_250),
.B(n_262),
.C(n_265),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_251),
.A2(n_275),
.B1(n_260),
.B2(n_242),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g291 ( 
.A(n_252),
.Y(n_291)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_254),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_255),
.A2(n_239),
.B1(n_225),
.B2(n_237),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_256),
.B(n_257),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_258),
.Y(n_281)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_238),
.Y(n_259)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_259),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_227),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_260),
.B(n_264),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_211),
.C(n_208),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_238),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_263),
.Y(n_295)
);

OAI32xp33_ASAP7_75t_L g264 ( 
.A1(n_247),
.A2(n_203),
.A3(n_210),
.B1(n_221),
.B2(n_223),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_233),
.B(n_234),
.C(n_247),
.Y(n_265)
);

NOR2x1_ASAP7_75t_L g266 ( 
.A(n_248),
.B(n_216),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_266),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_229),
.B(n_205),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_267),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_231),
.B(n_204),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_268),
.Y(n_289)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_243),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_269),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_229),
.B(n_199),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_270),
.B(n_277),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_233),
.B(n_189),
.C(n_165),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_246),
.C(n_249),
.Y(n_290)
);

XOR2x2_ASAP7_75t_L g273 ( 
.A(n_233),
.B(n_199),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_273),
.A2(n_274),
.B(n_275),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_235),
.A2(n_157),
.B(n_131),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_240),
.A2(n_132),
.B(n_196),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_276),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_230),
.A2(n_23),
.B(n_48),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_282),
.B(n_297),
.Y(n_321)
);

XOR2x1_ASAP7_75t_SL g283 ( 
.A(n_266),
.B(n_236),
.Y(n_283)
);

NAND2xp33_ASAP7_75t_SL g308 ( 
.A(n_283),
.B(n_253),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_261),
.A2(n_231),
.B1(n_228),
.B2(n_244),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_287),
.A2(n_288),
.B1(n_296),
.B2(n_269),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_261),
.A2(n_272),
.B1(n_258),
.B2(n_268),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_290),
.B(n_293),
.C(n_300),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_250),
.B(n_249),
.C(n_245),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_272),
.A2(n_243),
.B1(n_245),
.B2(n_241),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_251),
.A2(n_196),
.B1(n_65),
.B2(n_66),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_298),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_262),
.B(n_64),
.C(n_41),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_266),
.A2(n_70),
.B1(n_59),
.B2(n_3),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_303),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_279),
.B(n_265),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_305),
.B(n_310),
.C(n_314),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_291),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_306),
.B(n_307),
.Y(n_326)
);

CKINVDCx14_ASAP7_75t_R g307 ( 
.A(n_294),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_308),
.A2(n_325),
.B1(n_303),
.B2(n_302),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_286),
.B(n_271),
.C(n_273),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_286),
.B(n_256),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_311),
.B(n_319),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_283),
.A2(n_252),
.B(n_253),
.Y(n_312)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_312),
.Y(n_344)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_284),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_313),
.B(n_316),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_293),
.B(n_273),
.C(n_257),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_279),
.B(n_254),
.C(n_255),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_315),
.B(n_317),
.C(n_320),
.Y(n_337)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_284),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_287),
.B(n_264),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_288),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_318),
.B(n_324),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_282),
.B(n_270),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_290),
.B(n_267),
.C(n_274),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_322),
.A2(n_297),
.B1(n_281),
.B2(n_298),
.Y(n_334)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_296),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_285),
.A2(n_263),
.B1(n_259),
.B2(n_277),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_311),
.B(n_299),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_327),
.B(n_345),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_310),
.A2(n_280),
.B(n_300),
.Y(n_328)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_328),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_323),
.A2(n_281),
.B1(n_289),
.B2(n_280),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_329),
.A2(n_304),
.B1(n_23),
.B2(n_1),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_305),
.B(n_301),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_331),
.B(n_335),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_334),
.B(n_343),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_314),
.B(n_315),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_336),
.B(n_339),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_309),
.B(n_301),
.C(n_278),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_338),
.B(n_342),
.C(n_44),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_309),
.B(n_278),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_320),
.B(n_302),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_340),
.B(n_44),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_319),
.B(n_295),
.C(n_292),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_317),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_321),
.A2(n_12),
.B(n_16),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_344),
.A2(n_323),
.B(n_304),
.Y(n_346)
);

OR2x2_ASAP7_75t_L g371 ( 
.A(n_346),
.B(n_358),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_326),
.B(n_340),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_347),
.B(n_352),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_348),
.A2(n_332),
.B1(n_1),
.B2(n_2),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_342),
.B(n_12),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_333),
.B(n_12),
.Y(n_354)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_354),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_337),
.Y(n_355)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_355),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_357),
.B(n_360),
.Y(n_365)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_329),
.A2(n_10),
.B(n_17),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_337),
.A2(n_333),
.B(n_338),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_359),
.B(n_361),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_341),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_356),
.A2(n_334),
.B1(n_339),
.B2(n_331),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_362),
.B(n_368),
.Y(n_379)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_366),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_346),
.B(n_330),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_351),
.A2(n_335),
.B1(n_330),
.B2(n_6),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_369),
.B(n_357),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_355),
.A2(n_10),
.B(n_16),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_370),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_358),
.A2(n_10),
.B1(n_16),
.B2(n_6),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_373),
.B(n_353),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_363),
.B(n_350),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_374),
.B(n_376),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_364),
.B(n_349),
.C(n_353),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_375),
.B(n_378),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_377),
.B(n_383),
.Y(n_393)
);

INVx6_ASAP7_75t_L g378 ( 
.A(n_372),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_367),
.B(n_360),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_381),
.B(n_382),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_369),
.B(n_349),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_371),
.B(n_9),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_375),
.B(n_362),
.C(n_368),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_385),
.B(n_388),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_378),
.A2(n_371),
.B1(n_366),
.B2(n_365),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_387),
.B(n_389),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_379),
.B(n_368),
.C(n_377),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_379),
.Y(n_389)
);

OR2x2_ASAP7_75t_L g390 ( 
.A(n_384),
.B(n_373),
.Y(n_390)
);

OR2x2_ASAP7_75t_L g399 ( 
.A(n_390),
.B(n_8),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_380),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_391),
.B(n_13),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_394),
.A2(n_9),
.B(n_15),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_396),
.A2(n_397),
.B(n_400),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_386),
.B(n_8),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_399),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_391),
.A2(n_6),
.B(n_7),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_401),
.Y(n_405)
);

MAJx2_ASAP7_75t_L g404 ( 
.A(n_395),
.B(n_392),
.C(n_393),
.Y(n_404)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_404),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_402),
.A2(n_398),
.B(n_390),
.Y(n_407)
);

OAI321xp33_ASAP7_75t_L g408 ( 
.A1(n_407),
.A2(n_403),
.A3(n_405),
.B1(n_14),
.B2(n_44),
.C(n_1),
.Y(n_408)
);

AOI21x1_ASAP7_75t_L g409 ( 
.A1(n_408),
.A2(n_14),
.B(n_406),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_409),
.A2(n_1),
.B(n_2),
.Y(n_410)
);


endmodule