module real_jpeg_33593_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_553;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_546;
wire n_285;
wire n_172;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_545;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g157 ( 
.A(n_0),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_0),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_0),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_0),
.Y(n_315)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_0),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_1),
.B(n_62),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_1),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_1),
.B(n_242),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_1),
.B(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_1),
.B(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_1),
.B(n_431),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_1),
.B(n_434),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_1),
.Y(n_457)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_2),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_2),
.B(n_264),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_2),
.B(n_450),
.Y(n_449)
);

NAND2xp33_ASAP7_75t_SL g480 ( 
.A(n_2),
.B(n_481),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx11_ASAP7_75t_R g554 ( 
.A(n_3),
.Y(n_554)
);

INVx2_ASAP7_75t_R g50 ( 
.A(n_4),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_4),
.B(n_165),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_4),
.B(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_4),
.B(n_261),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_4),
.B(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_4),
.B(n_321),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_5),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_6),
.B(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_6),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_6),
.B(n_143),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_6),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_6),
.B(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_7),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_7),
.Y(n_101)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_8),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_8),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_9),
.B(n_35),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_9),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_9),
.B(n_80),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_9),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_9),
.B(n_130),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_9),
.B(n_130),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_9),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_9),
.B(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_9),
.B(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_10),
.B(n_203),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_10),
.B(n_264),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_10),
.B(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_10),
.Y(n_297)
);

AND2x2_ASAP7_75t_SL g448 ( 
.A(n_10),
.B(n_200),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_10),
.B(n_461),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_10),
.B(n_492),
.Y(n_491)
);

AOI21xp33_ASAP7_75t_L g18 ( 
.A1(n_11),
.A2(n_19),
.B(n_22),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_12),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_12),
.Y(n_145)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_12),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_13),
.Y(n_304)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_14),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_15),
.B(n_237),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_15),
.A2(n_126),
.B1(n_299),
.B2(n_301),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_15),
.B(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_15),
.B(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_15),
.B(n_360),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_15),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_15),
.B(n_484),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_15),
.B(n_497),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_16),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_16),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_16),
.Y(n_167)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_16),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_31),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_17),
.B(n_39),
.Y(n_38)
);

NAND2x1_ASAP7_75t_L g73 ( 
.A(n_17),
.B(n_74),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_17),
.B(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_17),
.B(n_119),
.Y(n_118)
);

AND2x2_ASAP7_75t_SL g121 ( 
.A(n_17),
.B(n_122),
.Y(n_121)
);

AND2x2_ASAP7_75t_SL g156 ( 
.A(n_17),
.B(n_157),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_17),
.B(n_169),
.Y(n_168)
);

BUFx4f_ASAP7_75t_SL g19 ( 
.A(n_20),
.Y(n_19)
);

BUFx12f_ASAP7_75t_SL g20 ( 
.A(n_21),
.Y(n_20)
);

A2O1A1Ixp33_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_251),
.B(n_534),
.C(n_555),
.Y(n_22)
);

NOR2xp67_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_170),
.Y(n_23)
);

OAI211xp5_ASAP7_75t_L g534 ( 
.A1(n_24),
.A2(n_535),
.B(n_538),
.C(n_553),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_107),
.Y(n_24)
);

NAND2xp33_ASAP7_75t_SL g540 ( 
.A(n_25),
.B(n_107),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_90),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_57),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_27),
.B(n_57),
.C(n_90),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_42),
.C(n_51),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_SL g92 ( 
.A(n_28),
.B(n_93),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_34),
.C(n_38),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_29),
.A2(n_30),
.B1(n_34),
.B2(n_115),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_29),
.B(n_117),
.C(n_121),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_29),
.A2(n_30),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_29),
.A2(n_30),
.B1(n_274),
.B2(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_30),
.B(n_274),
.C(n_277),
.Y(n_273)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_33),
.Y(n_161)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_33),
.Y(n_200)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_34),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g544 ( 
.A1(n_34),
.A2(n_115),
.B1(n_545),
.B2(n_546),
.Y(n_544)
);

BUFx4f_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_37),
.Y(n_120)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_38),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_38),
.A2(n_65),
.B1(n_72),
.B2(n_73),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_38),
.A2(n_65),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_38),
.A2(n_65),
.B1(n_263),
.B2(n_265),
.Y(n_262)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_40),
.Y(n_240)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_42),
.B(n_51),
.Y(n_93)
);

NOR2xp67_ASAP7_75t_SL g42 ( 
.A(n_43),
.B(n_50),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_49),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_50),
.B(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_50),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_52),
.B(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_52),
.B(n_96),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_52),
.B(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_55),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_56),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_56),
.Y(n_242)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_56),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_77),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_64),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_59),
.B(n_64),
.C(n_77),
.Y(n_551)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_63),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.C(n_72),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_65),
.B(n_260),
.C(n_263),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_66),
.B(n_121),
.C(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_68),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_68),
.B(n_142),
.Y(n_194)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_70),
.Y(n_328)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_72),
.A2(n_73),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_72),
.A2(n_73),
.B1(n_285),
.B2(n_286),
.Y(n_284)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_73),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_73),
.Y(n_550)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_75),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_76),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_83),
.B2(n_84),
.Y(n_77)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_78),
.Y(n_548)
);

INVxp67_ASAP7_75t_SL g78 ( 
.A(n_79),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_79),
.B(n_125),
.C(n_129),
.Y(n_124)
);

XOR2x2_ASAP7_75t_L g146 ( 
.A(n_79),
.B(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_82),
.Y(n_296)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_85),
.B(n_198),
.C(n_201),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g546 ( 
.A1(n_85),
.A2(n_86),
.B1(n_168),
.B2(n_191),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_85),
.B(n_548),
.C(n_549),
.Y(n_547)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_86),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_86),
.B(n_228),
.Y(n_227)
);

NOR3xp33_ASAP7_75t_SL g557 ( 
.A(n_86),
.B(n_115),
.C(n_168),
.Y(n_557)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_88),
.Y(n_98)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_94),
.C(n_105),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_109),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_105),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_99),
.C(n_102),
.Y(n_94)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_99),
.B(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_99),
.B(n_156),
.C(n_181),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_99),
.B(n_214),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_101),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_101),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_101),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_102),
.B(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_110),
.C(n_132),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_108),
.B(n_111),
.Y(n_206)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

MAJx2_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_116),
.C(n_124),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_112),
.B(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_116),
.B(n_124),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_117),
.A2(n_118),
.B1(n_121),
.B2(n_138),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_117),
.B(n_554),
.Y(n_553)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_121),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_121),
.B(n_232),
.Y(n_318)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_123),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_123),
.Y(n_432)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_123),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_125),
.A2(n_129),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_128),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_129),
.A2(n_148),
.B1(n_217),
.B2(n_344),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_132),
.A2(n_133),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_150),
.C(n_154),
.Y(n_133)
);

XNOR2x1_ASAP7_75t_SL g175 ( 
.A(n_134),
.B(n_176),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_139),
.C(n_146),
.Y(n_134)
);

XOR2x2_ASAP7_75t_L g248 ( 
.A(n_135),
.B(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

OA21x2_ASAP7_75t_L g436 ( 
.A1(n_138),
.A2(n_232),
.B(n_437),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_138),
.B(n_232),
.Y(n_437)
);

OAI21xp33_ASAP7_75t_L g468 ( 
.A1(n_138),
.A2(n_232),
.B(n_437),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_139),
.A2(n_140),
.B1(n_146),
.B2(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_145),
.Y(n_367)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_146),
.Y(n_250)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_148),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_154),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_163),
.C(n_168),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_155),
.B(n_190),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.C(n_159),
.Y(n_155)
);

XNOR2x1_ASAP7_75t_L g196 ( 
.A(n_156),
.B(n_158),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_156),
.B(n_181),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_156),
.B(n_429),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_156),
.B(n_430),
.Y(n_464)
);

INVx8_ASAP7_75t_L g506 ( 
.A(n_157),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_159),
.B(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g330 ( 
.A(n_159),
.B(n_331),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_159),
.B(n_331),
.C(n_336),
.Y(n_345)
);

OR2x2_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_162),
.Y(n_159)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_163),
.A2(n_164),
.B1(n_168),
.B2(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_167),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_168),
.B(n_180),
.C(n_183),
.Y(n_179)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_168),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_168),
.A2(n_183),
.B1(n_184),
.B2(n_191),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_207),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g535 ( 
.A1(n_171),
.A2(n_536),
.B(n_537),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_204),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_172),
.B(n_204),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_R g172 ( 
.A(n_173),
.B(n_175),
.C(n_177),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_173),
.B(n_175),
.Y(n_209)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_209),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_187),
.C(n_192),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_179),
.A2(n_188),
.B1(n_189),
.B2(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_179),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_180),
.B(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_181),
.B(n_267),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_181),
.B(n_267),
.Y(n_355)
);

BUFx2_ASAP7_75t_L g261 ( 
.A(n_182),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_182),
.Y(n_499)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx3_ASAP7_75t_SL g185 ( 
.A(n_186),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XNOR2x1_ASAP7_75t_L g245 ( 
.A(n_192),
.B(n_246),
.Y(n_245)
);

MAJx2_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_195),
.C(n_197),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_193),
.B(n_197),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_195),
.B(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_202),
.Y(n_228)
);

INVxp33_ASAP7_75t_SL g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g536 ( 
.A(n_208),
.B(n_210),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_245),
.C(n_248),
.Y(n_210)
);

XNOR2x1_ASAP7_75t_L g401 ( 
.A(n_211),
.B(n_402),
.Y(n_401)
);

MAJx2_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_229),
.C(n_243),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_212),
.B(n_393),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_215),
.C(n_226),
.Y(n_212)
);

XNOR2x1_ASAP7_75t_L g385 ( 
.A(n_213),
.B(n_386),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_215),
.A2(n_216),
.B1(n_226),
.B2(n_227),
.Y(n_386)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_221),
.C(n_222),
.Y(n_216)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_217),
.Y(n_344)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_222),
.Y(n_342)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_229),
.B(n_243),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_238),
.C(n_241),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_230),
.B(n_382),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_232),
.C(n_235),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_232),
.A2(n_233),
.B1(n_235),
.B2(n_236),
.Y(n_286)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_234),
.Y(n_494)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_SL g337 ( 
.A(n_237),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_238),
.A2(n_239),
.B1(n_241),
.B2(n_383),
.Y(n_382)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_241),
.Y(n_383)
);

XNOR2x1_ASAP7_75t_L g402 ( 
.A(n_245),
.B(n_248),
.Y(n_402)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_414),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_388),
.B(n_410),
.Y(n_253)
);

OAI21x1_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_370),
.B(n_387),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_346),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_256),
.B(n_346),
.Y(n_533)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_306),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_257),
.B(n_307),
.C(n_338),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_283),
.Y(n_257)
);

MAJx2_ASAP7_75t_L g374 ( 
.A(n_258),
.B(n_284),
.C(n_287),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_266),
.C(n_272),
.Y(n_258)
);

XOR2x2_ASAP7_75t_L g368 ( 
.A(n_259),
.B(n_369),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_262),
.Y(n_259)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_263),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_266),
.B(n_273),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_271),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

NOR2x1_ASAP7_75t_L g336 ( 
.A(n_271),
.B(n_337),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_271),
.B(n_432),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_271),
.B(n_509),
.Y(n_508)
);

HB1xp67_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_274),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_276),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_277),
.B(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_280),
.Y(n_446)
);

INVx5_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_282),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_287),
.Y(n_283)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_298),
.B2(n_305),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_295),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_290),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_292),
.Y(n_485)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx6_ASAP7_75t_L g435 ( 
.A(n_293),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_294),
.Y(n_512)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_295),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_297),
.B(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_298),
.Y(n_305)
);

MAJx2_ASAP7_75t_L g378 ( 
.A(n_298),
.B(n_379),
.C(n_380),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx5_ASAP7_75t_L g458 ( 
.A(n_300),
.Y(n_458)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

OA21x2_ASAP7_75t_SL g308 ( 
.A1(n_305),
.A2(n_309),
.B(n_313),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_338),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_316),
.C(n_329),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_308),
.B(n_329),
.Y(n_348)
);

INVx3_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

BUFx4f_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_SL g347 ( 
.A(n_316),
.B(n_348),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_319),
.C(n_324),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_317),
.A2(n_318),
.B1(n_425),
.B2(n_426),
.Y(n_424)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_319),
.A2(n_320),
.B1(n_324),
.B2(n_325),
.Y(n_426)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

XNOR2x2_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_336),
.Y(n_329)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx3_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx4_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

XOR2x2_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_345),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

MAJx2_ASAP7_75t_L g384 ( 
.A(n_340),
.B(n_341),
.C(n_345),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_343),
.Y(n_341)
);

MAJx2_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_349),
.C(n_368),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_347),
.B(n_418),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_350),
.B(n_368),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_355),
.C(n_356),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_352),
.B(n_422),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_355),
.A2(n_356),
.B1(n_357),
.B2(n_423),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_355),
.Y(n_423)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_363),
.C(n_365),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_358),
.A2(n_359),
.B1(n_363),
.B2(n_364),
.Y(n_472)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_SL g471 ( 
.A(n_365),
.B(n_472),
.Y(n_471)
);

INVx4_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_371),
.B(n_533),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

OR2x2_ASAP7_75t_L g387 ( 
.A(n_372),
.B(n_373),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_375),
.Y(n_373)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_374),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_385),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_376),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_384),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_381),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_378),
.B(n_396),
.C(n_397),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_381),
.Y(n_397)
);

INVxp67_ASAP7_75t_SL g396 ( 
.A(n_384),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_385),
.B(n_408),
.C(n_409),
.Y(n_407)
);

NAND3xp33_ASAP7_75t_SL g414 ( 
.A(n_388),
.B(n_415),
.C(n_532),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_389),
.A2(n_400),
.B1(n_403),
.B2(n_406),
.Y(n_388)
);

INVxp67_ASAP7_75t_SL g389 ( 
.A(n_390),
.Y(n_389)
);

NOR2xp67_ASAP7_75t_L g411 ( 
.A(n_390),
.B(n_401),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_390),
.B(n_401),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_394),
.C(n_398),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_392),
.B(n_398),
.Y(n_405)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_395),
.B(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_404),
.B(n_407),
.Y(n_412)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_411),
.A2(n_412),
.B(n_413),
.Y(n_410)
);

AO21x2_ASAP7_75t_L g415 ( 
.A1(n_416),
.A2(n_438),
.B(n_531),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_417),
.B(n_419),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_417),
.B(n_419),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_424),
.C(n_427),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_420),
.A2(n_421),
.B1(n_529),
.B2(n_530),
.Y(n_528)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_421),
.B(n_525),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_SL g525 ( 
.A(n_424),
.B(n_427),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_424),
.B(n_427),
.Y(n_530)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_433),
.C(n_436),
.Y(n_427)
);

XNOR2x1_ASAP7_75t_L g466 ( 
.A(n_428),
.B(n_467),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_433),
.A2(n_436),
.B1(n_468),
.B2(n_469),
.Y(n_467)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_433),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_439),
.A2(n_523),
.B(n_527),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_440),
.A2(n_474),
.B(n_522),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_465),
.Y(n_440)
);

NOR2x1_ASAP7_75t_L g522 ( 
.A(n_441),
.B(n_465),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_454),
.C(n_464),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_443),
.B(n_519),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_447),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_444),
.B(n_448),
.C(n_453),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_446),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_445),
.B(n_504),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_448),
.A2(n_449),
.B1(n_452),
.B2(n_453),
.Y(n_447)
);

CKINVDCx14_ASAP7_75t_R g452 ( 
.A(n_448),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_449),
.Y(n_453)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

AO22x1_ASAP7_75t_L g519 ( 
.A1(n_454),
.A2(n_455),
.B1(n_464),
.B2(n_520),
.Y(n_519)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_459),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_456),
.A2(n_459),
.B1(n_460),
.B2(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_456),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_458),
.Y(n_456)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx4_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_464),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_470),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_466),
.B(n_471),
.C(n_473),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_473),
.Y(n_470)
);

OAI21x1_ASAP7_75t_L g474 ( 
.A1(n_475),
.A2(n_516),
.B(n_521),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_476),
.A2(n_500),
.B(n_515),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_477),
.B(n_489),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_477),
.B(n_489),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_478),
.A2(n_479),
.B1(n_486),
.B2(n_487),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_SL g479 ( 
.A(n_480),
.B(n_483),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_480),
.B(n_483),
.C(n_486),
.Y(n_517)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_495),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_490),
.A2(n_491),
.B1(n_495),
.B2(n_496),
.Y(n_513)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx3_ASAP7_75t_SL g492 ( 
.A(n_493),
.Y(n_492)
);

INVx8_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

OAI21x1_ASAP7_75t_L g500 ( 
.A1(n_501),
.A2(n_507),
.B(n_514),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_503),
.Y(n_501)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVx5_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_508),
.B(n_513),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_508),
.B(n_513),
.Y(n_514)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_517),
.B(n_518),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_517),
.B(n_518),
.Y(n_521)
);

NOR2x1p5_ASAP7_75t_L g523 ( 
.A(n_524),
.B(n_526),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_526),
.B(n_528),
.Y(n_527)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

NOR3xp33_ASAP7_75t_L g538 ( 
.A(n_539),
.B(n_541),
.C(n_547),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_542),
.B(n_552),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_543),
.B(n_551),
.Y(n_542)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_544),
.B(n_547),
.Y(n_543)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_550),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_553),
.B(n_556),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_557),
.Y(n_556)
);


endmodule