module fake_jpeg_1225_n_126 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_29, n_12, n_8, n_15, n_7, n_126);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_126;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_23),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_25),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_11),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_50),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_1),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_49),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_1),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx8_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_51),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_37),
.C(n_43),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_59),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_47),
.A2(n_37),
.B1(n_43),
.B2(n_40),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_58),
.A2(n_62),
.B(n_31),
.Y(n_73)
);

NAND2x1p5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_40),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_33),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_60),
.B(n_32),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_50),
.B(n_41),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_61),
.B(n_41),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_51),
.A2(n_35),
.B1(n_34),
.B2(n_39),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_65),
.B(n_68),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_70),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_54),
.A2(n_39),
.B1(n_35),
.B2(n_34),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_67),
.A2(n_74),
.B1(n_62),
.B2(n_38),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_56),
.Y(n_68)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_69),
.Y(n_77)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_72),
.A2(n_73),
.B(n_59),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_57),
.B(n_44),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_75),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_10),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_73),
.A2(n_38),
.B1(n_4),
.B2(n_5),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_81),
.A2(n_82),
.B1(n_83),
.B2(n_86),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_71),
.A2(n_38),
.B1(n_5),
.B2(n_6),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_71),
.A2(n_38),
.B1(n_7),
.B2(n_8),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_67),
.A2(n_2),
.B(n_7),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_85),
.A2(n_87),
.B(n_82),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_70),
.A2(n_2),
.B1(n_8),
.B2(n_9),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_69),
.A2(n_9),
.B(n_10),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_88),
.B(n_90),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_89),
.A2(n_92),
.B(n_94),
.Y(n_103)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_80),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_20),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_11),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g92 ( 
.A(n_79),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_77),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_93),
.Y(n_107)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_95),
.B(n_98),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_87),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_97),
.A2(n_99),
.B(n_96),
.Y(n_108)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_83),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

NOR2xp67_ASAP7_75t_SL g104 ( 
.A(n_100),
.B(n_12),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_109),
.Y(n_114)
);

AOI21x1_ASAP7_75t_L g117 ( 
.A1(n_104),
.A2(n_108),
.B(n_110),
.Y(n_117)
);

OAI32xp33_ASAP7_75t_L g106 ( 
.A1(n_101),
.A2(n_88),
.A3(n_89),
.B1(n_96),
.B2(n_91),
.Y(n_106)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_106),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_101),
.B(n_30),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_24),
.C(n_13),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_26),
.C(n_14),
.Y(n_111)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_111),
.Y(n_115)
);

XOR2x1_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_12),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_107),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_103),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_118),
.A2(n_116),
.B1(n_117),
.B2(n_115),
.Y(n_122)
);

AOI321xp33_ASAP7_75t_L g119 ( 
.A1(n_114),
.A2(n_109),
.A3(n_102),
.B1(n_107),
.B2(n_112),
.C(n_27),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_119),
.B(n_120),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_15),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_123),
.A2(n_121),
.B(n_18),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_16),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_19),
.Y(n_126)
);


endmodule