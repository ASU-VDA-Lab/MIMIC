module real_jpeg_25498_n_16 (n_5, n_4, n_8, n_0, n_12, n_345, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_345;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_323;
wire n_176;
wire n_215;
wire n_166;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_1),
.A2(n_55),
.B1(n_56),
.B2(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_1),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_127),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_127),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_1),
.A2(n_47),
.B1(n_48),
.B2(n_127),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_2),
.A2(n_54),
.B1(n_55),
.B2(n_57),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_2),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_57),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_2),
.A2(n_47),
.B1(n_48),
.B2(n_57),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_2),
.A2(n_25),
.B1(n_26),
.B2(n_57),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_3),
.A2(n_69),
.B(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_3),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_3),
.B(n_60),
.Y(n_157)
);

OAI22xp33_ASAP7_75t_L g196 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_124),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_3),
.B(n_43),
.C(n_48),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_3),
.B(n_29),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_3),
.A2(n_98),
.B1(n_217),
.B2(n_224),
.Y(n_228)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_6),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_117),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_6),
.A2(n_47),
.B1(n_48),
.B2(n_117),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_6),
.A2(n_68),
.B1(n_69),
.B2(n_117),
.Y(n_261)
);

INVx8_ASAP7_75t_SL g63 ( 
.A(n_7),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_8),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_8),
.A2(n_55),
.B1(n_115),
.B2(n_135),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_115),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_8),
.A2(n_47),
.B1(n_48),
.B2(n_115),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_9),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_9),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_9),
.A2(n_47),
.B1(n_48),
.B2(n_67),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_9),
.A2(n_31),
.B1(n_32),
.B2(n_67),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_9),
.A2(n_25),
.B1(n_26),
.B2(n_67),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_10),
.A2(n_38),
.B1(n_55),
.B2(n_56),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_38),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_10),
.A2(n_38),
.B1(n_47),
.B2(n_48),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_12),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_12),
.A2(n_28),
.B1(n_55),
.B2(n_56),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_12),
.A2(n_28),
.B1(n_47),
.B2(n_48),
.Y(n_173)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_15),
.Y(n_101)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_15),
.Y(n_107)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_15),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_83),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_82),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_76),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_19),
.B(n_76),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_71),
.C(n_72),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_20),
.B(n_340),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_39),
.C(n_51),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_21),
.A2(n_22),
.B1(n_39),
.B2(n_324),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_34),
.Y(n_22)
);

OAI21xp33_ASAP7_75t_L g138 ( 
.A1(n_23),
.A2(n_113),
.B(n_116),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_29),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_24),
.A2(n_29),
.B(n_35),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_24),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_25),
.A2(n_26),
.B1(n_30),
.B2(n_33),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_25),
.A2(n_26),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g140 ( 
.A1(n_25),
.A2(n_62),
.B(n_123),
.C(n_141),
.Y(n_140)
);

HAxp5_ASAP7_75t_SL g169 ( 
.A(n_25),
.B(n_124),
.CON(n_169),
.SN(n_169)
);

INVx3_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

NAND3xp33_ASAP7_75t_L g141 ( 
.A(n_26),
.B(n_61),
.C(n_136),
.Y(n_141)
);

OAI32xp33_ASAP7_75t_L g168 ( 
.A1(n_26),
.A2(n_30),
.A3(n_32),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_29),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_29),
.A2(n_35),
.B1(n_160),
.B2(n_169),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_29),
.B(n_37),
.Y(n_265)
);

AO22x1_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_29)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_31),
.A2(n_32),
.B1(n_43),
.B2(n_45),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_31),
.B(n_33),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_32),
.B(n_199),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_34),
.A2(n_118),
.B(n_286),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_35),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_35),
.A2(n_322),
.B(n_323),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_39),
.A2(n_320),
.B1(n_321),
.B2(n_324),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_39),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_46),
.B(n_49),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_41),
.B(n_95),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_41),
.A2(n_50),
.B(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_41),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_41),
.A2(n_178),
.B(n_189),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_41),
.A2(n_177),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_41),
.A2(n_176),
.B1(n_177),
.B2(n_197),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_41),
.A2(n_177),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_41),
.A2(n_111),
.B(n_255),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_46),
.Y(n_41)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_43),
.A2(n_45),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_46),
.A2(n_93),
.B(n_94),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_46),
.B(n_96),
.Y(n_111)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_46),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_46),
.B(n_49),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_46),
.B(n_124),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_47),
.B(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_47),
.B(n_230),
.Y(n_229)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_SL g328 ( 
.A(n_51),
.B(n_329),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_58),
.B1(n_60),
.B2(n_66),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_53),
.A2(n_59),
.B(n_77),
.Y(n_317)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_56),
.A2(n_61),
.B1(n_62),
.B2(n_65),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_56),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_58),
.A2(n_66),
.B(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_58),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_58),
.A2(n_60),
.B1(n_126),
.B2(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_58),
.A2(n_60),
.B1(n_134),
.B2(n_261),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_58),
.A2(n_80),
.B(n_261),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_58),
.A2(n_74),
.B(n_305),
.Y(n_304)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_64),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_59),
.B(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_59),
.A2(n_120),
.B1(n_121),
.B2(n_125),
.Y(n_119)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

CKINVDCx5p33_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_70),
.B(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_71),
.A2(n_72),
.B1(n_73),
.B2(n_341),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_71),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_79),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_81),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_337),
.B(n_342),
.Y(n_83)
);

OAI321xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_313),
.A3(n_332),
.B1(n_335),
.B2(n_336),
.C(n_345),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_291),
.B(n_312),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_270),
.B(n_290),
.Y(n_86)
);

O2A1O1Ixp33_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_161),
.B(n_245),
.C(n_269),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_146),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_89),
.B(n_146),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_130),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_108),
.B1(n_128),
.B2(n_129),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_91),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_91),
.B(n_129),
.C(n_130),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_97),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_92),
.B(n_97),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_93),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_94),
.B(n_298),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_102),
.B(n_104),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_98),
.A2(n_104),
.B(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_98),
.A2(n_207),
.B(n_208),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_98),
.A2(n_214),
.B1(n_224),
.B2(n_225),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_98),
.A2(n_172),
.B(n_225),
.Y(n_278)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_99),
.A2(n_100),
.B1(n_103),
.B2(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_99),
.B(n_105),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_99),
.A2(n_213),
.B1(n_215),
.B2(n_216),
.Y(n_212)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_100),
.Y(n_154)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_101),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_SL g209 ( 
.A(n_107),
.Y(n_209)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_112),
.C(n_119),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_109),
.A2(n_110),
.B1(n_112),
.B2(n_149),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_114),
.B1(n_116),
.B2(n_118),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_113),
.A2(n_114),
.B1(n_118),
.B2(n_159),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_113),
.A2(n_264),
.B(n_265),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_113),
.A2(n_118),
.B1(n_286),
.B2(n_300),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_119),
.B(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_124),
.B(n_225),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_139),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_137),
.B2(n_138),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_133),
.B(n_137),
.C(n_139),
.Y(n_267)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_142),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_140),
.A2(n_142),
.B1(n_143),
.B2(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_140),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_145),
.A2(n_154),
.B(n_155),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_150),
.C(n_152),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_147),
.B(n_243),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_150),
.B(n_152),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_156),
.C(n_158),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_153),
.A2(n_156),
.B1(n_157),
.B2(n_183),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_153),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_155),
.B(n_208),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_182),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_240),
.B(n_244),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_191),
.B(n_239),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_179),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_166),
.B(n_179),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_174),
.C(n_175),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_167),
.B(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_168),
.B(n_171),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_171),
.Y(n_186)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_173),
.B(n_209),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_174),
.B(n_175),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_184),
.B2(n_185),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_180),
.B(n_187),
.C(n_190),
.Y(n_241)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_188),
.B2(n_190),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_186),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_189),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_234),
.B(n_238),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_210),
.B(n_233),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_200),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_194),
.B(n_200),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_195),
.B(n_198),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_198),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_206),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_202),
.B(n_205),
.C(n_206),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_204),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_207),
.Y(n_215)
);

AOI21xp33_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_220),
.B(n_232),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_219),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_212),
.B(n_219),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_227),
.B(n_231),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_222),
.B(n_223),
.Y(n_231)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_235),
.B(n_236),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_241),
.B(n_242),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_247),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_267),
.B2(n_268),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_257),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_257),
.C(n_268),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_253),
.B2(n_256),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_251),
.B(n_256),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_253),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_266),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_262),
.B2(n_263),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_260),
.B(n_262),
.C(n_266),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_263),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_265),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_267),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_271),
.B(n_272),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_289),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_279),
.B1(n_287),
.B2(n_288),
.Y(n_273)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_274),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_288),
.C(n_289),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_277),
.B2(n_278),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_276),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_276),
.B(n_277),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_277),
.A2(n_278),
.B1(n_304),
.B2(n_306),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_277),
.A2(n_306),
.B(n_307),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_279),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_280),
.B(n_283),
.C(n_284),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_283),
.B1(n_284),
.B2(n_285),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_292),
.B(n_293),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_294),
.A2(n_295),
.B1(n_310),
.B2(n_311),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_302),
.B1(n_308),
.B2(n_309),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_296),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_296),
.B(n_309),
.C(n_311),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_299),
.B(n_301),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_297),
.B(n_299),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_300),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_301),
.B(n_315),
.C(n_325),
.Y(n_314)
);

FAx1_ASAP7_75t_L g334 ( 
.A(n_301),
.B(n_315),
.CI(n_325),
.CON(n_334),
.SN(n_334)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_302),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_307),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_304),
.Y(n_306)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_310),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_326),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_314),
.B(n_326),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_316),
.A2(n_317),
.B1(n_318),
.B2(n_319),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_316),
.A2(n_317),
.B1(n_328),
.B2(n_330),
.Y(n_327)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_317),
.B(n_321),
.C(n_324),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_317),
.B(n_330),
.C(n_331),
.Y(n_338)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_321),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_331),
.Y(n_326)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_328),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_333),
.B(n_334),
.Y(n_335)
);

BUFx24_ASAP7_75t_SL g343 ( 
.A(n_334),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_338),
.B(n_339),
.Y(n_342)
);


endmodule