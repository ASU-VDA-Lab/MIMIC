module real_aes_366_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_453;
wire n_374;
wire n_379;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_547;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_552;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_488;
wire n_501;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_465;
wire n_473;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
INVx1_ASAP7_75t_L g178 ( .A(n_0), .Y(n_178) );
AO22x2_ASAP7_75t_L g92 ( .A1(n_1), .A2(n_51), .B1(n_89), .B2(n_93), .Y(n_92) );
AOI22xp5_ASAP7_75t_L g546 ( .A1(n_2), .A2(n_80), .B1(n_169), .B2(n_547), .Y(n_546) );
CKINVDCx20_ASAP7_75t_R g547 ( .A(n_2), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_3), .B(n_206), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_4), .B(n_221), .Y(n_314) );
INVx1_ASAP7_75t_L g191 ( .A(n_5), .Y(n_191) );
AO22x2_ASAP7_75t_L g88 ( .A1(n_6), .A2(n_16), .B1(n_89), .B2(n_90), .Y(n_88) );
AND2x2_ASAP7_75t_L g241 ( .A(n_7), .B(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g316 ( .A(n_8), .B(n_230), .Y(n_316) );
INVx2_ASAP7_75t_L g227 ( .A(n_9), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_10), .B(n_221), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g126 ( .A1(n_11), .A2(n_48), .B1(n_127), .B2(n_131), .Y(n_126) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_12), .B(n_206), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g161 ( .A1(n_13), .A2(n_49), .B1(n_162), .B2(n_165), .Y(n_161) );
AOI22xp33_ASAP7_75t_L g246 ( .A1(n_14), .A2(n_68), .B1(n_206), .B2(n_247), .Y(n_246) );
AOI22xp5_ASAP7_75t_L g172 ( .A1(n_15), .A2(n_64), .B1(n_173), .B2(n_174), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_15), .Y(n_173) );
OAI221xp5_ASAP7_75t_L g183 ( .A1(n_16), .A2(n_51), .B1(n_56), .B2(n_184), .C(n_186), .Y(n_183) );
OR2x2_ASAP7_75t_L g228 ( .A(n_17), .B(n_66), .Y(n_228) );
OA21x2_ASAP7_75t_L g231 ( .A1(n_17), .A2(n_66), .B(n_227), .Y(n_231) );
INVx3_ASAP7_75t_L g89 ( .A(n_18), .Y(n_89) );
AO21x2_ASAP7_75t_L g292 ( .A1(n_19), .A2(n_242), .B(n_293), .Y(n_292) );
AOI21xp5_ASAP7_75t_L g311 ( .A1(n_20), .A2(n_214), .B(n_312), .Y(n_311) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_21), .A2(n_80), .B1(n_168), .B2(n_169), .Y(n_79) );
INVx1_ASAP7_75t_L g168 ( .A(n_21), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_21), .B(n_221), .Y(n_286) );
INVx1_ASAP7_75t_SL g100 ( .A(n_22), .Y(n_100) );
AOI22xp33_ASAP7_75t_L g145 ( .A1(n_23), .A2(n_67), .B1(n_146), .B2(n_150), .Y(n_145) );
INVx1_ASAP7_75t_L g193 ( .A(n_24), .Y(n_193) );
AND2x2_ASAP7_75t_L g212 ( .A(n_24), .B(n_191), .Y(n_212) );
AND2x2_ASAP7_75t_L g215 ( .A(n_24), .B(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_25), .B(n_206), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_26), .B(n_221), .Y(n_265) );
AOI22xp5_ASAP7_75t_L g538 ( .A1(n_26), .A2(n_80), .B1(n_169), .B2(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_26), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_27), .B(n_206), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_28), .A2(n_214), .B(n_237), .Y(n_236) );
AOI22xp33_ASAP7_75t_L g138 ( .A1(n_29), .A2(n_72), .B1(n_139), .B2(n_142), .Y(n_138) );
AOI22xp5_ASAP7_75t_L g114 ( .A1(n_30), .A2(n_74), .B1(n_115), .B2(n_120), .Y(n_114) );
AOI22xp33_ASAP7_75t_L g153 ( .A1(n_31), .A2(n_53), .B1(n_154), .B2(n_158), .Y(n_153) );
AO22x2_ASAP7_75t_L g95 ( .A1(n_32), .A2(n_56), .B1(n_89), .B2(n_96), .Y(n_95) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_33), .B(n_223), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g294 ( .A(n_34), .B(n_206), .Y(n_294) );
INVx1_ASAP7_75t_L g209 ( .A(n_35), .Y(n_209) );
INVx1_ASAP7_75t_L g218 ( .A(n_35), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_36), .B(n_221), .Y(n_239) );
AND2x2_ASAP7_75t_L g260 ( .A(n_37), .B(n_225), .Y(n_260) );
INVx1_ASAP7_75t_L g101 ( .A(n_38), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_39), .B(n_223), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_40), .B(n_223), .Y(n_285) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_41), .B(n_206), .Y(n_240) );
AOI22xp33_ASAP7_75t_L g83 ( .A1(n_42), .A2(n_62), .B1(n_84), .B2(n_102), .Y(n_83) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_43), .B(n_206), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g283 ( .A1(n_44), .A2(n_214), .B(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g276 ( .A(n_45), .B(n_226), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_46), .B(n_223), .Y(n_266) );
INVx1_ASAP7_75t_L g556 ( .A(n_46), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_47), .B(n_223), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g251 ( .A1(n_50), .A2(n_69), .B1(n_214), .B2(n_252), .Y(n_251) );
INVxp33_ASAP7_75t_L g188 ( .A(n_51), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_52), .B(n_221), .Y(n_273) );
INVx1_ASAP7_75t_L g211 ( .A(n_54), .Y(n_211) );
INVx1_ASAP7_75t_L g216 ( .A(n_54), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_55), .B(n_223), .Y(n_313) );
INVxp67_ASAP7_75t_L g187 ( .A(n_56), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_57), .A2(n_214), .B(n_264), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_58), .A2(n_214), .B(n_219), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_59), .B(n_108), .Y(n_107) );
AOI21xp5_ASAP7_75t_L g295 ( .A1(n_60), .A2(n_214), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g288 ( .A(n_61), .B(n_226), .Y(n_288) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_63), .B(n_225), .Y(n_244) );
INVx1_ASAP7_75t_L g174 ( .A(n_64), .Y(n_174) );
AND2x2_ASAP7_75t_L g229 ( .A(n_65), .B(n_230), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_70), .A2(n_214), .B(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_71), .B(n_221), .Y(n_220) );
BUFx2_ASAP7_75t_L g275 ( .A(n_73), .Y(n_275) );
BUFx2_ASAP7_75t_SL g185 ( .A(n_75), .Y(n_185) );
OAI22xp5_ASAP7_75t_L g175 ( .A1(n_76), .A2(n_176), .B1(n_177), .B2(n_178), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_76), .Y(n_176) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_180), .B1(n_194), .B2(n_534), .C(n_537), .Y(n_77) );
XNOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_170), .Y(n_78) );
CKINVDCx16_ASAP7_75t_R g169 ( .A(n_80), .Y(n_169) );
HB1xp67_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
NOR2x1_ASAP7_75t_L g81 ( .A(n_82), .B(n_137), .Y(n_81) );
NAND4xp25_ASAP7_75t_L g82 ( .A(n_83), .B(n_107), .C(n_114), .D(n_126), .Y(n_82) );
BUFx2_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
BUFx6f_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
AND2x4_ASAP7_75t_L g86 ( .A(n_87), .B(n_94), .Y(n_86) );
AND2x2_ASAP7_75t_L g117 ( .A(n_87), .B(n_118), .Y(n_117) );
AND2x4_ASAP7_75t_L g160 ( .A(n_87), .B(n_144), .Y(n_160) );
AND2x4_ASAP7_75t_L g87 ( .A(n_88), .B(n_91), .Y(n_87) );
INVx1_ASAP7_75t_L g113 ( .A(n_88), .Y(n_113) );
AND2x2_ASAP7_75t_L g124 ( .A(n_88), .B(n_92), .Y(n_124) );
INVx1_ASAP7_75t_L g130 ( .A(n_88), .Y(n_130) );
INVx2_ASAP7_75t_L g90 ( .A(n_89), .Y(n_90) );
INVx1_ASAP7_75t_L g93 ( .A(n_89), .Y(n_93) );
INVx1_ASAP7_75t_L g96 ( .A(n_89), .Y(n_96) );
OAI22x1_ASAP7_75t_L g98 ( .A1(n_89), .A2(n_99), .B1(n_100), .B2(n_101), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_89), .Y(n_99) );
INVxp67_ASAP7_75t_L g105 ( .A(n_91), .Y(n_105) );
AND2x4_ASAP7_75t_L g112 ( .A(n_91), .B(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
AND2x2_ASAP7_75t_L g129 ( .A(n_92), .B(n_130), .Y(n_129) );
AND2x2_ASAP7_75t_L g149 ( .A(n_94), .B(n_129), .Y(n_149) );
AND2x2_ASAP7_75t_L g164 ( .A(n_94), .B(n_112), .Y(n_164) );
AND2x2_ASAP7_75t_L g94 ( .A(n_95), .B(n_97), .Y(n_94) );
AND2x2_ASAP7_75t_L g106 ( .A(n_95), .B(n_98), .Y(n_106) );
INVx2_ASAP7_75t_L g119 ( .A(n_95), .Y(n_119) );
BUFx2_ASAP7_75t_L g152 ( .A(n_95), .Y(n_152) );
AND2x4_ASAP7_75t_L g144 ( .A(n_97), .B(n_119), .Y(n_144) );
INVx2_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
AND2x2_ASAP7_75t_L g118 ( .A(n_98), .B(n_119), .Y(n_118) );
HB1xp67_ASAP7_75t_L g125 ( .A(n_98), .Y(n_125) );
INVx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
INVx6_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
AND2x4_ASAP7_75t_L g104 ( .A(n_105), .B(n_106), .Y(n_104) );
AND2x2_ASAP7_75t_L g111 ( .A(n_106), .B(n_112), .Y(n_111) );
AND2x4_ASAP7_75t_L g134 ( .A(n_106), .B(n_135), .Y(n_134) );
BUFx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx4_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
INVx6_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
AND2x4_ASAP7_75t_L g141 ( .A(n_112), .B(n_118), .Y(n_141) );
AND2x4_ASAP7_75t_L g157 ( .A(n_112), .B(n_144), .Y(n_157) );
BUFx6f_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
BUFx3_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AND2x2_ASAP7_75t_L g128 ( .A(n_118), .B(n_129), .Y(n_128) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx3_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx3_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_125), .Y(n_123) );
AND2x4_ASAP7_75t_L g143 ( .A(n_124), .B(n_144), .Y(n_143) );
AND2x4_ASAP7_75t_L g151 ( .A(n_124), .B(n_152), .Y(n_151) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
AND2x4_ASAP7_75t_L g167 ( .A(n_129), .B(n_144), .Y(n_167) );
HB1xp67_ASAP7_75t_L g136 ( .A(n_130), .Y(n_136) );
INVx3_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
BUFx2_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
NAND4xp25_ASAP7_75t_L g137 ( .A(n_138), .B(n_145), .C(n_153), .D(n_161), .Y(n_137) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx6_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
BUFx2_ASAP7_75t_SL g142 ( .A(n_143), .Y(n_142) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
BUFx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx4_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx8_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_SL g162 ( .A(n_163), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
INVx8_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
OAI22xp5_ASAP7_75t_SL g170 ( .A1(n_171), .A2(n_172), .B1(n_175), .B2(n_179), .Y(n_170) );
CKINVDCx20_ASAP7_75t_R g171 ( .A(n_172), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g179 ( .A(n_175), .Y(n_179) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx1_ASAP7_75t_SL g180 ( .A(n_181), .Y(n_180) );
CKINVDCx20_ASAP7_75t_R g181 ( .A(n_182), .Y(n_181) );
AND3x1_ASAP7_75t_SL g182 ( .A(n_183), .B(n_189), .C(n_192), .Y(n_182) );
INVxp67_ASAP7_75t_L g545 ( .A(n_183), .Y(n_545) );
CKINVDCx8_ASAP7_75t_R g184 ( .A(n_185), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g186 ( .A(n_187), .B(n_188), .Y(n_186) );
CKINVDCx16_ASAP7_75t_R g543 ( .A(n_189), .Y(n_543) );
AOI21xp33_ASAP7_75t_L g552 ( .A1(n_189), .A2(n_553), .B(n_554), .Y(n_552) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
AND2x2_ASAP7_75t_L g248 ( .A(n_190), .B(n_249), .Y(n_248) );
OR2x2_ASAP7_75t_SL g550 ( .A(n_190), .B(n_192), .Y(n_550) );
HB1xp67_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
AND2x2_ASAP7_75t_L g217 ( .A(n_191), .B(n_218), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_192), .B(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
NOR2x1p5_ASAP7_75t_L g253 ( .A(n_193), .B(n_254), .Y(n_253) );
HB1xp67_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AND2x4_ASAP7_75t_L g196 ( .A(n_197), .B(n_459), .Y(n_196) );
NOR2xp67_ASAP7_75t_L g197 ( .A(n_198), .B(n_378), .Y(n_197) );
NAND5xp2_ASAP7_75t_L g198 ( .A(n_199), .B(n_322), .C(n_332), .D(n_349), .E(n_365), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
OAI22xp5_ASAP7_75t_L g200 ( .A1(n_201), .A2(n_256), .B1(n_299), .B2(n_303), .Y(n_200) );
OR2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_232), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
AND2x4_ASAP7_75t_L g305 ( .A(n_203), .B(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g324 ( .A(n_203), .B(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g345 ( .A(n_203), .B(n_346), .Y(n_345) );
INVx4_ASAP7_75t_L g359 ( .A(n_203), .Y(n_359) );
AND2x2_ASAP7_75t_L g368 ( .A(n_203), .B(n_369), .Y(n_368) );
AND2x4_ASAP7_75t_SL g390 ( .A(n_203), .B(n_307), .Y(n_390) );
BUFx2_ASAP7_75t_L g433 ( .A(n_203), .Y(n_433) );
AND2x2_ASAP7_75t_L g448 ( .A(n_203), .B(n_233), .Y(n_448) );
OR2x2_ASAP7_75t_L g480 ( .A(n_203), .B(n_481), .Y(n_480) );
NOR4xp25_ASAP7_75t_L g529 ( .A(n_203), .B(n_530), .C(n_531), .D(n_532), .Y(n_529) );
OR2x6_ASAP7_75t_L g203 ( .A(n_204), .B(n_229), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_213), .B(n_225), .Y(n_204) );
AND2x4_ASAP7_75t_L g206 ( .A(n_207), .B(n_212), .Y(n_206) );
AND2x4_ASAP7_75t_L g207 ( .A(n_208), .B(n_210), .Y(n_207) );
AND2x6_ASAP7_75t_L g223 ( .A(n_208), .B(n_216), .Y(n_223) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
AND2x4_ASAP7_75t_L g221 ( .A(n_210), .B(n_218), .Y(n_221) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx5_ASAP7_75t_L g224 ( .A(n_212), .Y(n_224) );
AND2x6_ASAP7_75t_L g214 ( .A(n_215), .B(n_217), .Y(n_214) );
BUFx3_ASAP7_75t_L g250 ( .A(n_215), .Y(n_250) );
INVx2_ASAP7_75t_L g255 ( .A(n_216), .Y(n_255) );
AND2x4_ASAP7_75t_L g252 ( .A(n_217), .B(n_253), .Y(n_252) );
INVx2_ASAP7_75t_L g249 ( .A(n_218), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_222), .B(n_224), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_223), .B(n_275), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_224), .A2(n_238), .B(n_239), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_224), .A2(n_265), .B(n_266), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g272 ( .A1(n_224), .A2(n_273), .B(n_274), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_224), .A2(n_285), .B(n_286), .Y(n_284) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_224), .A2(n_297), .B(n_298), .Y(n_296) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_224), .A2(n_313), .B(n_314), .Y(n_312) );
AO21x2_ASAP7_75t_L g245 ( .A1(n_225), .A2(n_246), .B(n_251), .Y(n_245) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_225), .Y(n_309) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AND2x2_ASAP7_75t_SL g226 ( .A(n_227), .B(n_228), .Y(n_226) );
AND2x4_ASAP7_75t_L g267 ( .A(n_227), .B(n_228), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_230), .A2(n_270), .B(n_271), .Y(n_269) );
BUFx4f_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx3_ASAP7_75t_L g234 ( .A(n_231), .Y(n_234) );
AOI31xp33_ASAP7_75t_L g397 ( .A1(n_232), .A2(n_398), .A3(n_400), .B(n_402), .Y(n_397) );
INVx2_ASAP7_75t_SL g514 ( .A(n_232), .Y(n_514) );
OR2x2_ASAP7_75t_L g232 ( .A(n_233), .B(n_243), .Y(n_232) );
INVx2_ASAP7_75t_L g321 ( .A(n_233), .Y(n_321) );
AND2x2_ASAP7_75t_L g325 ( .A(n_233), .B(n_308), .Y(n_325) );
INVx2_ASAP7_75t_L g348 ( .A(n_233), .Y(n_348) );
AND2x2_ASAP7_75t_L g367 ( .A(n_233), .B(n_307), .Y(n_367) );
AO21x2_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B(n_241), .Y(n_233) );
INVx4_ASAP7_75t_L g242 ( .A(n_234), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_236), .B(n_240), .Y(n_235) );
INVx3_ASAP7_75t_L g281 ( .A(n_242), .Y(n_281) );
AND2x2_ASAP7_75t_L g319 ( .A(n_243), .B(n_320), .Y(n_319) );
BUFx3_ASAP7_75t_L g326 ( .A(n_243), .Y(n_326) );
INVx2_ASAP7_75t_L g344 ( .A(n_243), .Y(n_344) );
AND2x2_ASAP7_75t_L g399 ( .A(n_243), .B(n_359), .Y(n_399) );
AND2x4_ASAP7_75t_L g243 ( .A(n_244), .B(n_245), .Y(n_243) );
AND2x4_ASAP7_75t_L g370 ( .A(n_244), .B(n_245), .Y(n_370) );
INVx1_ASAP7_75t_L g536 ( .A(n_247), .Y(n_536) );
AND2x4_ASAP7_75t_L g247 ( .A(n_248), .B(n_250), .Y(n_247) );
HB1xp67_ASAP7_75t_L g553 ( .A(n_249), .Y(n_553) );
INVx1_ASAP7_75t_L g555 ( .A(n_250), .Y(n_555) );
INVx3_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_257), .B(n_289), .Y(n_256) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_258), .B(n_277), .Y(n_257) );
OR2x2_ASAP7_75t_L g299 ( .A(n_258), .B(n_300), .Y(n_299) );
INVx3_ASAP7_75t_L g451 ( .A(n_258), .Y(n_451) );
OR2x2_ASAP7_75t_L g499 ( .A(n_258), .B(n_500), .Y(n_499) );
NAND2x1_ASAP7_75t_L g258 ( .A(n_259), .B(n_268), .Y(n_258) );
OR2x2_ASAP7_75t_SL g290 ( .A(n_259), .B(n_291), .Y(n_290) );
INVx4_ASAP7_75t_L g329 ( .A(n_259), .Y(n_329) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_259), .Y(n_373) );
INVx2_ASAP7_75t_L g381 ( .A(n_259), .Y(n_381) );
OR2x2_ASAP7_75t_L g416 ( .A(n_259), .B(n_279), .Y(n_416) );
AND2x2_ASAP7_75t_L g528 ( .A(n_259), .B(n_383), .Y(n_528) );
AND2x2_ASAP7_75t_L g533 ( .A(n_259), .B(n_292), .Y(n_533) );
OR2x6_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_263), .B(n_267), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g293 ( .A1(n_267), .A2(n_294), .B(n_295), .Y(n_293) );
OR2x2_ASAP7_75t_L g291 ( .A(n_268), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g357 ( .A(n_268), .B(n_278), .Y(n_357) );
OR2x2_ASAP7_75t_L g364 ( .A(n_268), .B(n_329), .Y(n_364) );
NOR2x1_ASAP7_75t_SL g383 ( .A(n_268), .B(n_302), .Y(n_383) );
BUFx2_ASAP7_75t_L g415 ( .A(n_268), .Y(n_415) );
AND2x2_ASAP7_75t_L g424 ( .A(n_268), .B(n_329), .Y(n_424) );
AND2x2_ASAP7_75t_L g457 ( .A(n_268), .B(n_377), .Y(n_457) );
INVx2_ASAP7_75t_SL g466 ( .A(n_268), .Y(n_466) );
AND2x2_ASAP7_75t_L g469 ( .A(n_268), .B(n_279), .Y(n_469) );
OR2x6_ASAP7_75t_L g268 ( .A(n_269), .B(n_276), .Y(n_268) );
NAND3xp33_ASAP7_75t_L g464 ( .A(n_277), .B(n_334), .C(n_419), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_277), .B(n_381), .Y(n_484) );
INVxp67_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_278), .B(n_466), .Y(n_487) );
INVx2_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_279), .Y(n_331) );
AND2x2_ASAP7_75t_L g375 ( .A(n_279), .B(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g440 ( .A(n_279), .B(n_441), .Y(n_440) );
INVx3_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AO21x2_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_282), .B(n_288), .Y(n_280) );
AO21x1_ASAP7_75t_SL g302 ( .A1(n_281), .A2(n_282), .B(n_288), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_287), .Y(n_282) );
AND2x4_ASAP7_75t_L g335 ( .A(n_289), .B(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g471 ( .A(n_291), .B(n_416), .Y(n_471) );
AND2x2_ASAP7_75t_L g301 ( .A(n_292), .B(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g339 ( .A(n_292), .Y(n_339) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_292), .Y(n_356) );
INVx2_ASAP7_75t_L g377 ( .A(n_292), .Y(n_377) );
INVx1_ASAP7_75t_L g441 ( .A(n_292), .Y(n_441) );
INVx2_ASAP7_75t_L g523 ( .A(n_299), .Y(n_523) );
OR2x2_ASAP7_75t_L g387 ( .A(n_300), .B(n_364), .Y(n_387) );
INVx2_ASAP7_75t_SL g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g527 ( .A(n_301), .B(n_424), .Y(n_527) );
AND2x2_ASAP7_75t_L g420 ( .A(n_302), .B(n_377), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_317), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AOI22xp5_ASAP7_75t_L g511 ( .A1(n_305), .A2(n_434), .B1(n_451), .B2(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g347 ( .A(n_307), .Y(n_347) );
AND2x2_ASAP7_75t_L g401 ( .A(n_307), .B(n_321), .Y(n_401) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_307), .Y(n_428) );
INVx3_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_308), .Y(n_396) );
AOI21x1_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_310), .B(n_316), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_315), .Y(n_310) );
INVxp67_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_319), .B(n_433), .Y(n_432) );
OAI32xp33_ASAP7_75t_L g449 ( .A1(n_319), .A2(n_450), .A3(n_452), .B1(n_453), .B2(n_455), .Y(n_449) );
BUFx2_ASAP7_75t_L g334 ( .A(n_320), .Y(n_334) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g476 ( .A(n_321), .B(n_370), .Y(n_476) );
OR4x1_ASAP7_75t_L g322 ( .A(n_323), .B(n_326), .C(n_327), .D(n_330), .Y(n_322) );
OAI22xp5_ASAP7_75t_L g507 ( .A1(n_323), .A2(n_414), .B1(n_508), .B2(n_509), .Y(n_507) );
INVx2_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
HB1xp67_ASAP7_75t_L g516 ( .A(n_324), .Y(n_516) );
AND2x2_ASAP7_75t_L g358 ( .A(n_325), .B(n_359), .Y(n_358) );
BUFx2_ASAP7_75t_L g438 ( .A(n_325), .Y(n_438) );
INVx1_ASAP7_75t_L g454 ( .A(n_325), .Y(n_454) );
INVx1_ASAP7_75t_L g489 ( .A(n_325), .Y(n_489) );
OR2x2_ASAP7_75t_L g446 ( .A(n_326), .B(n_447), .Y(n_446) );
OR2x2_ASAP7_75t_L g490 ( .A(n_326), .B(n_491), .Y(n_490) );
OAI22xp5_ASAP7_75t_L g429 ( .A1(n_327), .A2(n_364), .B1(n_408), .B2(n_427), .Y(n_429) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g473 ( .A(n_328), .B(n_382), .Y(n_473) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
BUFx2_ASAP7_75t_L g340 ( .A(n_329), .Y(n_340) );
NOR2xp67_ASAP7_75t_L g355 ( .A(n_329), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g336 ( .A(n_330), .Y(n_336) );
NAND4xp25_ASAP7_75t_L g463 ( .A(n_330), .B(n_334), .C(n_415), .D(n_427), .Y(n_463) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g500 ( .A(n_331), .Y(n_500) );
AOI22xp5_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_335), .B1(n_337), .B2(n_341), .Y(n_332) );
OAI22xp33_ASAP7_75t_L g483 ( .A1(n_333), .A2(n_334), .B1(n_484), .B2(n_485), .Y(n_483) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVxp67_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
INVx3_ASAP7_75t_L g362 ( .A(n_339), .Y(n_362) );
AOI32xp33_ASAP7_75t_L g478 ( .A1(n_339), .A2(n_479), .A3(n_483), .B1(n_488), .B2(n_492), .Y(n_478) );
AND2x2_ASAP7_75t_L g341 ( .A(n_342), .B(n_345), .Y(n_341) );
NOR2xp67_ASAP7_75t_L g384 ( .A(n_342), .B(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g437 ( .A(n_342), .B(n_438), .Y(n_437) );
AOI221xp5_ASAP7_75t_L g461 ( .A1(n_342), .A2(n_350), .B1(n_462), .B2(n_467), .C(n_470), .Y(n_461) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OR2x2_ASAP7_75t_L g394 ( .A(n_343), .B(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g509 ( .A(n_343), .B(n_510), .Y(n_509) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_344), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g351 ( .A(n_346), .Y(n_351) );
AND2x2_ASAP7_75t_L g369 ( .A(n_346), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
INVx1_ASAP7_75t_SL g409 ( .A(n_347), .Y(n_409) );
INVx1_ASAP7_75t_L g393 ( .A(n_348), .Y(n_393) );
AOI22xp5_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_352), .B1(n_358), .B2(n_360), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OR2x2_ASAP7_75t_L g495 ( .A(n_351), .B(n_425), .Y(n_495) );
INVx1_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx2_ASAP7_75t_L g435 ( .A(n_354), .Y(n_435) );
AND2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_357), .Y(n_354) );
AND2x2_ASAP7_75t_L g366 ( .A(n_359), .B(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_359), .B(n_396), .Y(n_395) );
NAND2x1p5_ASAP7_75t_L g408 ( .A(n_359), .B(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_359), .B(n_401), .Y(n_522) );
AOI22xp33_ASAP7_75t_SL g519 ( .A1(n_360), .A2(n_520), .B1(n_521), .B2(n_523), .Y(n_519) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_362), .B(n_363), .Y(n_361) );
OR2x2_ASAP7_75t_L g402 ( .A(n_362), .B(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g412 ( .A(n_362), .B(n_413), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_362), .B(n_424), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_362), .B(n_466), .Y(n_465) );
AND2x4_ASAP7_75t_SL g467 ( .A(n_362), .B(n_468), .Y(n_467) );
INVx2_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
OR2x2_ASAP7_75t_L g443 ( .A(n_364), .B(n_444), .Y(n_443) );
OAI21xp5_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_368), .B(n_371), .Y(n_365) );
INVx1_ASAP7_75t_L g385 ( .A(n_367), .Y(n_385) );
AOI22xp5_ASAP7_75t_L g404 ( .A1(n_368), .A2(n_405), .B1(n_412), .B2(n_417), .Y(n_404) );
INVx3_ASAP7_75t_L g407 ( .A(n_370), .Y(n_407) );
INVx2_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
OR2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
OAI32xp33_ASAP7_75t_SL g462 ( .A1(n_373), .A2(n_433), .A3(n_463), .B1(n_464), .B2(n_465), .Y(n_462) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g382 ( .A(n_376), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NAND4xp25_ASAP7_75t_SL g378 ( .A(n_379), .B(n_404), .C(n_421), .D(n_436), .Y(n_378) );
AOI221xp5_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_384), .B1(n_386), .B2(n_388), .C(n_397), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
INVx2_ASAP7_75t_L g419 ( .A(n_381), .Y(n_419) );
AND2x2_ASAP7_75t_L g468 ( .A(n_381), .B(n_469), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_381), .B(n_420), .Y(n_506) );
AND2x2_ASAP7_75t_L g517 ( .A(n_381), .B(n_440), .Y(n_517) );
INVx2_ASAP7_75t_L g403 ( .A(n_383), .Y(n_403) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OAI21xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_391), .B(n_394), .Y(n_388) );
AND2x2_ASAP7_75t_L g520 ( .A(n_389), .B(n_391), .Y(n_520) );
INVx2_ASAP7_75t_SL g389 ( .A(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_390), .B(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g497 ( .A(n_395), .Y(n_497) );
INVx1_ASAP7_75t_L g482 ( .A(n_396), .Y(n_482) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_399), .B(n_454), .Y(n_453) );
NOR2x1_ASAP7_75t_L g411 ( .A(n_400), .B(n_407), .Y(n_411) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_SL g510 ( .A(n_401), .Y(n_510) );
INVx1_ASAP7_75t_L g492 ( .A(n_403), .Y(n_492) );
OR2x2_ASAP7_75t_L g508 ( .A(n_403), .B(n_419), .Y(n_508) );
NAND2xp33_ASAP7_75t_SL g405 ( .A(n_406), .B(n_410), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_408), .Y(n_406) );
INVx2_ASAP7_75t_L g425 ( .A(n_407), .Y(n_425) );
AND2x2_ASAP7_75t_L g430 ( .A(n_407), .B(n_420), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_407), .B(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g504 ( .A(n_408), .Y(n_504) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AOI22xp5_ASAP7_75t_L g493 ( .A1(n_413), .A2(n_494), .B1(n_496), .B2(n_498), .Y(n_493) );
INVx1_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
OR2x2_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
INVx1_ASAP7_75t_L g458 ( .A(n_416), .Y(n_458) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_419), .B(n_420), .Y(n_418) );
INVx1_ASAP7_75t_L g444 ( .A(n_420), .Y(n_444) );
AOI322xp5_ASAP7_75t_L g421 ( .A1(n_422), .A2(n_425), .A3(n_426), .B1(n_429), .B2(n_430), .C1(n_431), .C2(n_434), .Y(n_421) );
OAI21xp5_ASAP7_75t_SL g472 ( .A1(n_422), .A2(n_473), .B(n_474), .Y(n_472) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
AND2x2_ASAP7_75t_L g439 ( .A(n_424), .B(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g496 ( .A(n_425), .B(n_497), .Y(n_496) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_432), .B(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g452 ( .A(n_433), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_433), .B(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
AOI221xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_439), .B1(n_442), .B2(n_445), .C(n_449), .Y(n_436) );
AOI221xp5_ASAP7_75t_L g524 ( .A1(n_438), .A2(n_525), .B1(n_527), .B2(n_528), .C(n_529), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_440), .B(n_451), .Y(n_450) );
BUFx2_ASAP7_75t_L g491 ( .A(n_441), .Y(n_491) );
INVx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OAI21xp5_ASAP7_75t_L g515 ( .A1(n_445), .A2(n_516), .B(n_517), .Y(n_515) );
INVx1_ASAP7_75t_SL g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
NAND2xp33_ASAP7_75t_SL g525 ( .A(n_454), .B(n_526), .Y(n_525) );
INVx3_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AND2x4_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
NOR4xp75_ASAP7_75t_L g459 ( .A(n_460), .B(n_477), .C(n_501), .D(n_518), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_472), .Y(n_460) );
INVx1_ASAP7_75t_L g531 ( .A(n_469), .Y(n_531) );
INVx1_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g503 ( .A(n_476), .B(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g530 ( .A(n_476), .Y(n_530) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_478), .B(n_493), .Y(n_477) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
INVx1_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx2_ASAP7_75t_SL g526 ( .A(n_497), .Y(n_526) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
NAND3x1_ASAP7_75t_L g501 ( .A(n_502), .B(n_511), .C(n_515), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_505), .B(n_507), .Y(n_502) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVxp67_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_519), .B(n_524), .Y(n_518) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_535), .Y(n_534) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
OAI222xp33_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_540), .B1(n_546), .B2(n_548), .C1(n_551), .C2(n_556), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g540 ( .A(n_541), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_542), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
CKINVDCx20_ASAP7_75t_R g548 ( .A(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
CKINVDCx20_ASAP7_75t_R g551 ( .A(n_552), .Y(n_551) );
INVxp67_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
endmodule