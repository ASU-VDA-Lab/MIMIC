module fake_jpeg_28580_n_425 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_425);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_425;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_412;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx24_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx5_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g117 ( 
.A(n_50),
.Y(n_117)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_17),
.B(n_16),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_52),
.B(n_73),
.Y(n_101)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_53),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_57),
.Y(n_130)
);

BUFx8_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g135 ( 
.A(n_58),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_59),
.Y(n_122)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_61),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_19),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_76),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_64),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_65),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_66),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_67),
.Y(n_126)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_70),
.Y(n_137)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_72),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_17),
.B(n_15),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_74),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_18),
.B(n_15),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_77),
.Y(n_112)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_80),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_R g81 ( 
.A(n_19),
.B(n_15),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_81),
.B(n_14),
.Y(n_125)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

BUFx10_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_36),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_84),
.B(n_39),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_61),
.A2(n_36),
.B1(n_31),
.B2(n_28),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_85),
.A2(n_96),
.B1(n_118),
.B2(n_0),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_41),
.C(n_31),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_90),
.B(n_105),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_43),
.A2(n_26),
.B1(n_40),
.B2(n_18),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_83),
.A2(n_41),
.B1(n_37),
.B2(n_34),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_102),
.A2(n_56),
.B1(n_66),
.B2(n_64),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_72),
.B(n_40),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_108),
.B(n_114),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_58),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_48),
.A2(n_26),
.B1(n_38),
.B2(n_39),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_72),
.B(n_38),
.Y(n_119)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_119),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_63),
.A2(n_39),
.B1(n_20),
.B2(n_34),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_120),
.A2(n_39),
.B1(n_20),
.B2(n_67),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_58),
.Y(n_123)
);

NAND3xp33_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_125),
.C(n_127),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_47),
.B(n_37),
.Y(n_124)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_49),
.B(n_14),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_65),
.B(n_39),
.Y(n_131)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

BUFx2_ASAP7_75t_L g139 ( 
.A(n_130),
.Y(n_139)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_139),
.Y(n_197)
);

OA22x2_ASAP7_75t_L g140 ( 
.A1(n_102),
.A2(n_68),
.B1(n_19),
.B2(n_57),
.Y(n_140)
);

AO22x2_ASAP7_75t_L g190 ( 
.A1(n_140),
.A2(n_148),
.B1(n_169),
.B2(n_106),
.Y(n_190)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_134),
.Y(n_141)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_141),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_90),
.B(n_75),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_167),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_85),
.A2(n_70),
.B1(n_69),
.B2(n_54),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_144),
.A2(n_168),
.B1(n_132),
.B2(n_107),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_146),
.A2(n_133),
.B1(n_104),
.B2(n_122),
.Y(n_186)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_134),
.Y(n_147)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_147),
.Y(n_181)
);

OA22x2_ASAP7_75t_L g148 ( 
.A1(n_120),
.A2(n_19),
.B1(n_62),
.B2(n_59),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_89),
.Y(n_149)
);

INVx13_ASAP7_75t_L g187 ( 
.A(n_149),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_150),
.A2(n_163),
.B1(n_164),
.B2(n_166),
.Y(n_196)
);

OA22x2_ASAP7_75t_L g180 ( 
.A1(n_152),
.A2(n_165),
.B1(n_171),
.B2(n_133),
.Y(n_180)
);

INVx4_ASAP7_75t_SL g153 ( 
.A(n_130),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_155),
.Y(n_178)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_110),
.Y(n_155)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_89),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_156),
.B(n_158),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_157),
.Y(n_179)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_94),
.Y(n_158)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_93),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_160),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_113),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_161),
.B(n_162),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_109),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g163 ( 
.A(n_106),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_118),
.A2(n_115),
.B1(n_112),
.B2(n_132),
.Y(n_165)
);

INVx13_ASAP7_75t_L g166 ( 
.A(n_136),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_91),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_98),
.A2(n_20),
.B1(n_14),
.B2(n_2),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_99),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_111),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_170),
.B(n_173),
.Y(n_184)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_110),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_116),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_101),
.B(n_0),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_174),
.B(n_1),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_176),
.A2(n_190),
.B1(n_148),
.B2(n_135),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_180),
.A2(n_148),
.B1(n_140),
.B2(n_104),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_143),
.A2(n_86),
.B(n_121),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_183),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_92),
.C(n_129),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_186),
.A2(n_99),
.B1(n_100),
.B2(n_103),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_146),
.A2(n_137),
.B1(n_128),
.B2(n_88),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_188),
.A2(n_192),
.B1(n_97),
.B2(n_153),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_189),
.B(n_175),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_172),
.A2(n_88),
.B1(n_97),
.B2(n_128),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_140),
.A2(n_117),
.B(n_95),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_194),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_172),
.B(n_174),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_195),
.B(n_165),
.Y(n_199)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_185),
.Y(n_198)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_198),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_200),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_152),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_201),
.A2(n_192),
.B1(n_190),
.B2(n_196),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_177),
.B(n_154),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_202),
.B(n_207),
.Y(n_229)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_184),
.Y(n_203)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_203),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_205),
.A2(n_206),
.B1(n_211),
.B2(n_218),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_175),
.B(n_151),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_208),
.B(n_212),
.Y(n_239)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_184),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_209),
.Y(n_230)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_181),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_210),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_190),
.A2(n_180),
.B1(n_186),
.B2(n_194),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_141),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_183),
.B(n_159),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_189),
.C(n_145),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_190),
.A2(n_148),
.B1(n_140),
.B2(n_100),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_214),
.A2(n_216),
.B1(n_196),
.B2(n_190),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_193),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_193),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_190),
.A2(n_122),
.B1(n_103),
.B2(n_160),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_215),
.A2(n_192),
.B(n_182),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_219),
.A2(n_235),
.B(n_199),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_222),
.A2(n_223),
.B1(n_224),
.B2(n_232),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_214),
.A2(n_190),
.B1(n_180),
.B2(n_186),
.Y(n_224)
);

MAJx2_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_182),
.C(n_183),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_204),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_204),
.C(n_213),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_211),
.A2(n_180),
.B1(n_194),
.B2(n_176),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_228),
.A2(n_234),
.B1(n_201),
.B2(n_200),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_214),
.A2(n_180),
.B1(n_188),
.B2(n_176),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_233),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_218),
.A2(n_180),
.B1(n_188),
.B2(n_156),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_215),
.A2(n_178),
.B(n_179),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_207),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_236),
.B(n_203),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_178),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_237),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_240),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_232),
.A2(n_216),
.B1(n_201),
.B2(n_209),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_241),
.A2(n_245),
.B1(n_220),
.B2(n_228),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_242),
.A2(n_221),
.B(n_234),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_229),
.B(n_202),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_254),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_219),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_253),
.Y(n_265)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_238),
.Y(n_249)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_249),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_233),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_250),
.Y(n_279)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_238),
.Y(n_251)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_251),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_252),
.B(n_221),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_235),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_235),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_230),
.C(n_239),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_225),
.B(n_213),
.C(n_227),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_256),
.B(n_225),
.C(n_227),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_237),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_259),
.Y(n_276)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_226),
.Y(n_258)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_258),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_226),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_250),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_260),
.B(n_191),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_262),
.B(n_267),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_206),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_246),
.A2(n_241),
.B1(n_220),
.B2(n_228),
.Y(n_269)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_269),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_270),
.Y(n_284)
);

MAJx2_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_212),
.C(n_229),
.Y(n_271)
);

NAND5xp2_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_257),
.C(n_247),
.D(n_240),
.E(n_252),
.Y(n_283)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_249),
.Y(n_272)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_272),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_246),
.A2(n_220),
.B1(n_234),
.B2(n_223),
.Y(n_273)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_273),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_242),
.A2(n_222),
.B(n_223),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_274),
.A2(n_224),
.B(n_245),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_248),
.A2(n_239),
.B(n_230),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_275),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_278),
.B(n_255),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_248),
.B(n_208),
.Y(n_280)
);

NAND3xp33_ASAP7_75t_L g293 ( 
.A(n_280),
.B(n_279),
.C(n_277),
.Y(n_293)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_281),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_282),
.B(n_292),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_283),
.B(n_271),
.Y(n_307)
);

NOR3xp33_ASAP7_75t_L g285 ( 
.A(n_279),
.B(n_247),
.C(n_243),
.Y(n_285)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_285),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_280),
.A2(n_251),
.B1(n_231),
.B2(n_258),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_286),
.B(n_288),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_287),
.A2(n_270),
.B1(n_265),
.B2(n_266),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_260),
.A2(n_231),
.B1(n_259),
.B2(n_206),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_276),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_293),
.Y(n_306)
);

NOR3xp33_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_142),
.C(n_179),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_294),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_210),
.Y(n_295)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_295),
.Y(n_313)
);

OAI22x1_ASAP7_75t_L g297 ( 
.A1(n_274),
.A2(n_205),
.B1(n_252),
.B2(n_187),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_297),
.A2(n_303),
.B1(n_263),
.B2(n_261),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_264),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_298),
.B(n_302),
.Y(n_321)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_299),
.Y(n_318)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_261),
.Y(n_301)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_301),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_275),
.B(n_264),
.Y(n_302)
);

NAND3xp33_ASAP7_75t_L g303 ( 
.A(n_265),
.B(n_191),
.C(n_181),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_289),
.A2(n_273),
.B1(n_269),
.B2(n_268),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_305),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_307),
.B(n_166),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_308),
.B(n_312),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_291),
.B(n_262),
.C(n_278),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_310),
.B(n_322),
.C(n_301),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_289),
.A2(n_300),
.B1(n_297),
.B2(n_284),
.Y(n_312)
);

FAx1_ASAP7_75t_SL g314 ( 
.A(n_302),
.B(n_267),
.CI(n_262),
.CON(n_314),
.SN(n_314)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_314),
.B(n_325),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_284),
.A2(n_266),
.B(n_272),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_315),
.A2(n_320),
.B(n_327),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_291),
.B(n_271),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_316),
.B(n_164),
.Y(n_345)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_319),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_296),
.A2(n_263),
.B(n_267),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_296),
.B(n_197),
.C(n_198),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_281),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_300),
.A2(n_198),
.B1(n_149),
.B2(n_169),
.Y(n_326)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_326),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_295),
.A2(n_287),
.B(n_283),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_329),
.B(n_320),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_318),
.Y(n_330)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_330),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_310),
.B(n_290),
.C(n_197),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_332),
.B(n_335),
.C(n_338),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_316),
.B(n_290),
.C(n_197),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_323),
.B(n_173),
.Y(n_336)
);

CKINVDCx14_ASAP7_75t_R g361 ( 
.A(n_336),
.Y(n_361)
);

FAx1_ASAP7_75t_SL g337 ( 
.A(n_307),
.B(n_163),
.CI(n_157),
.CON(n_337),
.SN(n_337)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_337),
.B(n_340),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_314),
.B(n_185),
.C(n_155),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_317),
.B(n_163),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_339),
.B(n_344),
.Y(n_360)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_324),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_318),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_342),
.B(n_343),
.Y(n_352)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_324),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_327),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_345),
.B(n_348),
.Y(n_353)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_315),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_346),
.A2(n_349),
.B1(n_313),
.B2(n_306),
.Y(n_354)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_321),
.Y(n_349)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_354),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_329),
.B(n_314),
.C(n_304),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_355),
.B(n_357),
.C(n_359),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_328),
.A2(n_331),
.B1(n_305),
.B2(n_309),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_356),
.B(n_358),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_345),
.B(n_312),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_332),
.B(n_304),
.C(n_308),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_335),
.B(n_321),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_362),
.B(n_365),
.C(n_367),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_331),
.A2(n_311),
.B1(n_313),
.B2(n_322),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_364),
.B(n_366),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_338),
.B(n_311),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_334),
.A2(n_326),
.B1(n_185),
.B2(n_171),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_333),
.B(n_170),
.C(n_147),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_360),
.B(n_341),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_368),
.B(n_369),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_350),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_358),
.B(n_336),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_370),
.B(n_373),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_362),
.B(n_347),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_355),
.B(n_337),
.C(n_348),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_377),
.B(n_380),
.C(n_353),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_352),
.A2(n_117),
.B(n_136),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_378),
.A2(n_381),
.B(n_23),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_361),
.A2(n_139),
.B1(n_87),
.B2(n_126),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_379),
.B(n_371),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_351),
.B(n_126),
.C(n_116),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_365),
.A2(n_87),
.B(n_187),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_372),
.B(n_351),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_382),
.B(n_384),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_383),
.B(n_386),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_372),
.B(n_359),
.C(n_357),
.Y(n_384)
);

AOI322xp5_ASAP7_75t_L g385 ( 
.A1(n_369),
.A2(n_363),
.A3(n_367),
.B1(n_353),
.B2(n_187),
.C1(n_109),
.C2(n_135),
.Y(n_385)
);

HB1xp67_ASAP7_75t_SL g399 ( 
.A(n_385),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_376),
.B(n_109),
.C(n_23),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_376),
.B(n_23),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_387),
.B(n_388),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_374),
.B(n_2),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_389),
.B(n_392),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_375),
.B(n_2),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_393),
.B(n_3),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_391),
.A2(n_390),
.B(n_384),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_395),
.B(n_4),
.C(n_6),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_398),
.B(n_401),
.Y(n_404)
);

OAI21xp33_ASAP7_75t_L g400 ( 
.A1(n_382),
.A2(n_377),
.B(n_380),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_400),
.B(n_4),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_383),
.B(n_23),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_390),
.B(n_23),
.Y(n_402)
);

INVxp33_ASAP7_75t_L g406 ( 
.A(n_402),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_394),
.A2(n_4),
.B(n_5),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_405),
.B(n_410),
.C(n_6),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_407),
.B(n_408),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_396),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_409),
.B(n_411),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_399),
.A2(n_6),
.B(n_7),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_400),
.B(n_6),
.C(n_7),
.Y(n_411)
);

NOR3xp33_ASAP7_75t_L g412 ( 
.A(n_406),
.B(n_403),
.C(n_397),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_412),
.A2(n_413),
.B1(n_8),
.B2(n_10),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_404),
.A2(n_7),
.B(n_8),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_414),
.B(n_8),
.C(n_10),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_415),
.A2(n_8),
.B(n_9),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_417),
.Y(n_420)
);

NOR3xp33_ASAP7_75t_L g421 ( 
.A(n_418),
.B(n_419),
.C(n_416),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_421),
.B(n_420),
.C(n_12),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_SL g423 ( 
.A1(n_422),
.A2(n_11),
.B(n_12),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_423),
.B(n_11),
.Y(n_424)
);

O2A1O1Ixp33_ASAP7_75t_SL g425 ( 
.A1(n_424),
.A2(n_11),
.B(n_13),
.C(n_420),
.Y(n_425)
);


endmodule