module fake_jpeg_22864_n_249 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_249);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_249;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_24),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_31),
.Y(n_41)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx3_ASAP7_75t_SL g49 ( 
.A(n_32),
.Y(n_49)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_34),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_20),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_20),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_33),
.A2(n_20),
.B1(n_27),
.B2(n_26),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_39),
.A2(n_19),
.B(n_18),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_30),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_40),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_38),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_44),
.Y(n_71)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_46),
.Y(n_56)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_31),
.B(n_16),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_53),
.B(n_55),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_16),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_36),
.B1(n_27),
.B2(n_19),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_58),
.A2(n_54),
.B1(n_15),
.B2(n_23),
.Y(n_93)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_62),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_44),
.B(n_46),
.C(n_55),
.Y(n_60)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_60),
.A2(n_69),
.B(n_74),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g64 ( 
.A(n_47),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_66),
.Y(n_83)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_68),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_48),
.A2(n_27),
.B1(n_26),
.B2(n_29),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_70),
.A2(n_15),
.B1(n_23),
.B2(n_28),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_50),
.Y(n_72)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_73),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_48),
.A2(n_18),
.B1(n_28),
.B2(n_15),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_80),
.B(n_81),
.Y(n_107)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_45),
.C(n_32),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_88),
.C(n_72),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_57),
.B(n_42),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_90),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_69),
.A2(n_29),
.B1(n_43),
.B2(n_42),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_85),
.A2(n_93),
.B1(n_70),
.B2(n_91),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_71),
.A2(n_43),
.B1(n_32),
.B2(n_37),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_86),
.A2(n_87),
.B1(n_94),
.B2(n_49),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_71),
.A2(n_37),
.B1(n_35),
.B2(n_51),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_37),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_35),
.B(n_18),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_89),
.A2(n_28),
.B(n_23),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_34),
.Y(n_90)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_97),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_96),
.A2(n_101),
.B1(n_104),
.B2(n_108),
.Y(n_129)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_100),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_99),
.A2(n_88),
.B(n_50),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_83),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_85),
.A2(n_60),
.B1(n_65),
.B2(n_66),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_87),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_103),
.Y(n_125)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_106),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_81),
.B(n_25),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_112),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_91),
.A2(n_88),
.B1(n_93),
.B2(n_82),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_111),
.A2(n_49),
.B1(n_54),
.B2(n_64),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_78),
.B(n_25),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_61),
.Y(n_113)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_113),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_90),
.B(n_21),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_86),
.Y(n_122)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_115),
.Y(n_154)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

AND2x6_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_89),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_124),
.Y(n_152)
);

AOI22x1_ASAP7_75t_SL g121 ( 
.A1(n_99),
.A2(n_88),
.B1(n_50),
.B2(n_94),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_121),
.A2(n_99),
.B1(n_49),
.B2(n_64),
.Y(n_149)
);

NAND3xp33_ASAP7_75t_L g138 ( 
.A(n_122),
.B(n_135),
.C(n_100),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_76),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_128),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_21),
.Y(n_128)
);

CKINVDCx5p33_ASAP7_75t_R g130 ( 
.A(n_110),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_130),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_113),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_131),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_133),
.A2(n_63),
.B1(n_67),
.B2(n_61),
.Y(n_153)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_134),
.B(n_105),
.Y(n_137)
);

AND2x6_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_50),
.Y(n_135)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_137),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_138),
.A2(n_149),
.B1(n_151),
.B2(n_122),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_129),
.A2(n_103),
.B1(n_108),
.B2(n_111),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_139),
.A2(n_153),
.B1(n_117),
.B2(n_54),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_129),
.B(n_111),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_142),
.C(n_144),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_95),
.C(n_109),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_101),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_143),
.B(n_146),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_119),
.B(n_96),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_115),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_75),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_125),
.A2(n_108),
.B1(n_114),
.B2(n_76),
.Y(n_151)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_132),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_118),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_133),
.B(n_123),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_120),
.C(n_112),
.Y(n_170)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_157),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_136),
.A2(n_121),
.B1(n_124),
.B2(n_134),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_163),
.Y(n_192)
);

INVxp33_ASAP7_75t_L g160 ( 
.A(n_137),
.Y(n_160)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_160),
.Y(n_188)
);

NOR4xp25_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_136),
.C(n_131),
.D(n_143),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_161),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_162),
.Y(n_177)
);

NOR3xp33_ASAP7_75t_SL g163 ( 
.A(n_152),
.B(n_130),
.C(n_128),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_156),
.B(n_116),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_164),
.B(n_22),
.C(n_17),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_151),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_165),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_167),
.B(n_168),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_148),
.B(n_120),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_139),
.A2(n_117),
.B1(n_79),
.B2(n_92),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_173),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_172),
.C(n_140),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_142),
.B(n_141),
.C(n_144),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_152),
.A2(n_79),
.B1(n_92),
.B2(n_63),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_150),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_175),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_149),
.A2(n_61),
.B1(n_59),
.B2(n_22),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_176),
.A2(n_145),
.B(n_158),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_164),
.B(n_154),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_178),
.A2(n_17),
.B(n_2),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_179),
.B(n_191),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_181),
.A2(n_169),
.B1(n_167),
.B2(n_170),
.Y(n_196)
);

XOR2x2_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_34),
.Y(n_182)
);

XNOR2x1_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_17),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_68),
.C(n_22),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_185),
.B(n_186),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_166),
.B(n_172),
.C(n_173),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_184),
.B(n_171),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_195),
.Y(n_216)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_182),
.Y(n_194)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_194),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_188),
.B(n_160),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_196),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_183),
.A2(n_163),
.B1(n_174),
.B2(n_22),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_197),
.A2(n_200),
.B1(n_191),
.B2(n_177),
.Y(n_212)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_190),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_198),
.A2(n_201),
.B(n_204),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_189),
.B(n_13),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_203),
.A2(n_7),
.B(n_12),
.Y(n_218)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_190),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_181),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_205),
.A2(n_206),
.B(n_180),
.Y(n_211)
);

OAI21x1_ASAP7_75t_L g206 ( 
.A1(n_178),
.A2(n_7),
.B(n_12),
.Y(n_206)
);

NAND3xp33_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_180),
.C(n_192),
.Y(n_207)
);

MAJx2_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_194),
.C(n_8),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_186),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_1),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_202),
.B(n_179),
.C(n_185),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_213),
.Y(n_226)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_211),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_217),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_195),
.B(n_187),
.C(n_178),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_1),
.C(n_2),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_9),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_214),
.B(n_201),
.Y(n_219)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_219),
.Y(n_236)
);

NOR3xp33_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_9),
.C(n_3),
.Y(n_231)
);

MAJx2_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_6),
.C(n_11),
.Y(n_221)
);

AOI32xp33_ASAP7_75t_L g229 ( 
.A1(n_221),
.A2(n_210),
.A3(n_217),
.B1(n_216),
.B2(n_5),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_223),
.B(n_227),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_R g224 ( 
.A(n_207),
.B(n_6),
.C(n_3),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_224),
.A2(n_4),
.B1(n_5),
.B2(n_9),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_6),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_219),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_229),
.B(n_230),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_222),
.B(n_213),
.Y(n_230)
);

AOI31xp67_ASAP7_75t_L g241 ( 
.A1(n_231),
.A2(n_235),
.A3(n_10),
.B(n_11),
.Y(n_241)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_233),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_215),
.C(n_3),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_234),
.A2(n_228),
.B(n_225),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_232),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_239),
.Y(n_243)
);

OR2x2_ASAP7_75t_L g244 ( 
.A(n_241),
.B(n_231),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_236),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_244),
.Y(n_246)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_243),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_245),
.A2(n_240),
.B1(n_13),
.B2(n_2),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_247),
.A2(n_246),
.B(n_13),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_248),
.B(n_2),
.Y(n_249)
);


endmodule