module fake_jpeg_20662_n_135 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_135);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_30),
.Y(n_37)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_0),
.Y(n_30)
);

BUFx4f_ASAP7_75t_SL g31 ( 
.A(n_26),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_32),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_19),
.B(n_1),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_36),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_3),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_27),
.Y(n_42)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_35),
.A2(n_22),
.B1(n_21),
.B2(n_17),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_38),
.A2(n_39),
.B1(n_47),
.B2(n_20),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_13),
.B1(n_18),
.B2(n_27),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_42),
.B(n_23),
.Y(n_59)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_22),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_45),
.B(n_48),
.Y(n_64)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_29),
.A2(n_21),
.B1(n_20),
.B2(n_16),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_28),
.B(n_32),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_32),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_50),
.B(n_59),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_51),
.A2(n_53),
.B1(n_55),
.B2(n_41),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_47),
.A2(n_29),
.B1(n_30),
.B2(n_15),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_46),
.A2(n_13),
.B1(n_18),
.B2(n_14),
.Y(n_55)
);

NOR2x1_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_31),
.Y(n_57)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

NOR2x1_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_31),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_60),
.B(n_64),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_16),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_61),
.B(n_24),
.Y(n_77)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_62),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_43),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_66),
.B(n_72),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_41),
.C(n_37),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_33),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_71),
.A2(n_49),
.B1(n_56),
.B2(n_24),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_64),
.B(n_15),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_73),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_37),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_75),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_51),
.B(n_39),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_78),
.A2(n_60),
.B1(n_57),
.B2(n_25),
.Y(n_83)
);

NOR4xp25_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_60),
.C(n_57),
.D(n_53),
.Y(n_80)
);

AOI322xp5_ASAP7_75t_SL g100 ( 
.A1(n_80),
.A2(n_26),
.A3(n_33),
.B1(n_13),
.B2(n_18),
.C1(n_14),
.C2(n_12),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_70),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_82),
.B(n_83),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_65),
.A2(n_49),
.B(n_44),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_84),
.A2(n_79),
.B(n_76),
.Y(n_93)
);

OAI32xp33_ASAP7_75t_L g85 ( 
.A1(n_65),
.A2(n_72),
.A3(n_67),
.B1(n_75),
.B2(n_68),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_92),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_86),
.A2(n_89),
.B1(n_79),
.B2(n_63),
.Y(n_98)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_76),
.A2(n_49),
.B1(n_56),
.B2(n_25),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_93),
.A2(n_101),
.B(n_88),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_90),
.B(n_67),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_94),
.B(n_95),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_87),
.B(n_58),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_58),
.Y(n_97)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_98),
.A2(n_102),
.B1(n_40),
.B2(n_26),
.Y(n_108)
);

BUFx12f_ASAP7_75t_SL g106 ( 
.A(n_100),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_81),
.A2(n_69),
.B(n_52),
.Y(n_101)
);

NOR3xp33_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_84),
.C(n_85),
.Y(n_102)
);

AO21x1_ASAP7_75t_L g113 ( 
.A1(n_104),
.A2(n_99),
.B(n_98),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_96),
.A2(n_86),
.B1(n_92),
.B2(n_91),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_105),
.A2(n_108),
.B1(n_40),
.B2(n_52),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_26),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_110),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_93),
.A2(n_69),
.B(n_4),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_111),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_114),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_104),
.A2(n_103),
.B(n_94),
.Y(n_114)
);

AOI321xp33_ASAP7_75t_L g115 ( 
.A1(n_107),
.A2(n_103),
.A3(n_10),
.B1(n_11),
.B2(n_7),
.C(n_8),
.Y(n_115)
);

AOI31xp67_ASAP7_75t_L g120 ( 
.A1(n_115),
.A2(n_106),
.A3(n_111),
.B(n_8),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_118),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_112),
.A2(n_63),
.B1(n_6),
.B2(n_7),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_105),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_122),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_124),
.A2(n_112),
.B1(n_123),
.B2(n_120),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_121),
.A2(n_119),
.B(n_116),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_126),
.A2(n_106),
.B(n_115),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_128),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_109),
.C(n_52),
.Y(n_128)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_129),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_125),
.B(n_5),
.Y(n_130)
);

NAND3xp33_ASAP7_75t_L g133 ( 
.A(n_130),
.B(n_5),
.C(n_6),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_133),
.A2(n_131),
.B(n_8),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_132),
.Y(n_135)
);


endmodule