module fake_jpeg_3225_n_515 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_515);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_515;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_4),
.B(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_4),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

INVx8_ASAP7_75t_SL g47 ( 
.A(n_3),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_10),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_7),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_7),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_54),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx4_ASAP7_75t_SL g138 ( 
.A(n_55),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_21),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_56),
.B(n_71),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_28),
.B(n_15),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_57),
.B(n_76),
.Y(n_124)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_58),
.Y(n_166)
);

BUFx24_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g121 ( 
.A(n_59),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_18),
.Y(n_61)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_62),
.Y(n_149)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_63),
.Y(n_134)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_64),
.Y(n_118)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_65),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_66),
.Y(n_152)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_67),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_68),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_18),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_69),
.Y(n_133)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_70),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_47),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_72),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_73),
.Y(n_143)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_74),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_75),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_32),
.B(n_15),
.Y(n_76)
);

INVx2_ASAP7_75t_R g77 ( 
.A(n_47),
.Y(n_77)
);

INVx2_ASAP7_75t_R g157 ( 
.A(n_77),
.Y(n_157)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_78),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_80),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_28),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_82),
.B(n_91),
.Y(n_112)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_39),
.Y(n_83)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_35),
.Y(n_85)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_87),
.Y(n_137)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_88),
.Y(n_163)
);

INVx8_ASAP7_75t_SL g89 ( 
.A(n_30),
.Y(n_89)
);

INVx5_ASAP7_75t_SL g109 ( 
.A(n_89),
.Y(n_109)
);

NAND2x1_ASAP7_75t_L g90 ( 
.A(n_27),
.B(n_1),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_30),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_48),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_32),
.B(n_15),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_92),
.B(n_105),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_93),
.Y(n_154)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_27),
.Y(n_94)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_94),
.Y(n_156)
);

BUFx4f_ASAP7_75t_L g95 ( 
.A(n_37),
.Y(n_95)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_95),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_96),
.Y(n_145)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_97),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_98),
.Y(n_160)
);

INVx3_ASAP7_75t_SL g99 ( 
.A(n_39),
.Y(n_99)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_99),
.Y(n_162)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_37),
.Y(n_100)
);

INVx13_ASAP7_75t_L g127 ( 
.A(n_100),
.Y(n_127)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_102),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_51),
.Y(n_102)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_39),
.Y(n_103)
);

CKINVDCx9p33_ASAP7_75t_R g125 ( 
.A(n_103),
.Y(n_125)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_39),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g164 ( 
.A(n_104),
.Y(n_164)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_16),
.Y(n_105)
);

OAI21xp33_ASAP7_75t_L g180 ( 
.A1(n_110),
.A2(n_59),
.B(n_42),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_52),
.A2(n_40),
.B1(n_19),
.B2(n_51),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_128),
.A2(n_100),
.B1(n_45),
.B2(n_49),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_103),
.B(n_40),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_130),
.B(n_132),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_55),
.B(n_19),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_55),
.B(n_34),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_139),
.B(n_141),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_96),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_98),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_142),
.B(n_147),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_77),
.B(n_16),
.Y(n_144)
);

NAND3xp33_ASAP7_75t_L g189 ( 
.A(n_144),
.B(n_158),
.C(n_33),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_99),
.B(n_34),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_146),
.B(n_24),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_78),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_69),
.B(n_50),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_148),
.B(n_161),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_90),
.B(n_41),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_88),
.Y(n_161)
);

NAND2xp33_ASAP7_75t_SL g236 ( 
.A(n_167),
.B(n_211),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_121),
.A2(n_58),
.B1(n_95),
.B2(n_97),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_L g227 ( 
.A1(n_168),
.A2(n_177),
.B1(n_181),
.B2(n_151),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_135),
.A2(n_68),
.B1(n_75),
.B2(n_93),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_169),
.A2(n_170),
.B1(n_197),
.B2(n_200),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_124),
.B(n_112),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_171),
.B(n_185),
.Y(n_230)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_107),
.Y(n_172)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_172),
.Y(n_235)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_107),
.Y(n_173)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_173),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_138),
.Y(n_174)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_174),
.Y(n_244)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_121),
.Y(n_175)
);

INVx3_ASAP7_75t_SL g249 ( 
.A(n_175),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_162),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_176),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_157),
.A2(n_104),
.B1(n_36),
.B2(n_136),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_158),
.A2(n_80),
.B(n_73),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_178),
.B(n_184),
.Y(n_226)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_160),
.Y(n_179)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_179),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_180),
.B(n_208),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_157),
.A2(n_83),
.B1(n_42),
.B2(n_41),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_110),
.B(n_59),
.Y(n_182)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_182),
.Y(n_238)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_114),
.Y(n_183)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_183),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_125),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_126),
.Y(n_185)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_133),
.Y(n_186)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_186),
.Y(n_228)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_131),
.Y(n_187)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_187),
.Y(n_246)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_166),
.Y(n_188)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_188),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_189),
.B(n_201),
.Y(n_245)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_166),
.Y(n_190)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_190),
.Y(n_234)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_115),
.Y(n_192)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_192),
.Y(n_216)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_159),
.Y(n_193)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_193),
.Y(n_219)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_134),
.Y(n_194)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_194),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_153),
.B(n_43),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_195),
.B(n_209),
.Y(n_243)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_164),
.Y(n_196)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_196),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_154),
.A2(n_87),
.B1(n_86),
.B2(n_85),
.Y(n_197)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_114),
.Y(n_199)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_199),
.Y(n_232)
);

OAI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_163),
.A2(n_84),
.B1(n_81),
.B2(n_79),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_108),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_129),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_203),
.Y(n_239)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_106),
.Y(n_204)
);

INVx6_ASAP7_75t_L g223 ( 
.A(n_204),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_119),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_205),
.B(n_210),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_117),
.A2(n_66),
.B1(n_62),
.B2(n_60),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_207),
.A2(n_117),
.B1(n_184),
.B2(n_119),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_129),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_118),
.B(n_43),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_122),
.B(n_50),
.Y(n_210)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_140),
.Y(n_211)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_106),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_212),
.B(n_213),
.Y(n_250)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_133),
.Y(n_213)
);

INVx6_ASAP7_75t_SL g214 ( 
.A(n_138),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_214),
.B(n_215),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_150),
.B(n_49),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_200),
.A2(n_156),
.B1(n_155),
.B2(n_123),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_217),
.A2(n_168),
.B1(n_181),
.B2(n_120),
.Y(n_253)
);

FAx1_ASAP7_75t_SL g220 ( 
.A(n_180),
.B(n_165),
.CI(n_127),
.CON(n_220),
.SN(n_220)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_220),
.B(n_224),
.Y(n_256)
);

FAx1_ASAP7_75t_SL g224 ( 
.A(n_182),
.B(n_127),
.CI(n_109),
.CON(n_224),
.SN(n_224)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_227),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_237),
.A2(n_247),
.B1(n_205),
.B2(n_149),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_177),
.A2(n_109),
.B(n_163),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_242),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_198),
.A2(n_152),
.B1(n_149),
.B2(n_145),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_202),
.B(n_143),
.C(n_155),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_252),
.B(n_208),
.C(n_203),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_253),
.A2(n_284),
.B1(n_239),
.B2(n_231),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_206),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_254),
.B(n_261),
.Y(n_286)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_221),
.Y(n_255)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_255),
.Y(n_311)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_221),
.Y(n_257)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_257),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_258),
.B(n_274),
.C(n_276),
.Y(n_297)
);

INVx13_ASAP7_75t_L g259 ( 
.A(n_244),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_259),
.Y(n_287)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_241),
.Y(n_260)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_260),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_218),
.B(n_191),
.Y(n_261)
);

BUFx24_ASAP7_75t_L g262 ( 
.A(n_249),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_262),
.B(n_271),
.Y(n_293)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_232),
.Y(n_263)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_263),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_218),
.B(n_176),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_264),
.B(n_265),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_230),
.B(n_193),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_244),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_266),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_250),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_267),
.B(n_269),
.Y(n_309)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_223),
.Y(n_268)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_268),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_243),
.B(n_172),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_245),
.B(n_173),
.Y(n_270)
);

NOR2x1_ASAP7_75t_L g310 ( 
.A(n_270),
.B(n_278),
.Y(n_310)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_219),
.Y(n_272)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_272),
.Y(n_295)
);

INVx13_ASAP7_75t_L g273 ( 
.A(n_249),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_273),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_238),
.B(n_211),
.C(n_175),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_232),
.Y(n_275)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_275),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_238),
.B(n_188),
.C(n_143),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_236),
.B(n_219),
.Y(n_278)
);

INVx6_ASAP7_75t_L g279 ( 
.A(n_241),
.Y(n_279)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_279),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_234),
.B(n_174),
.Y(n_280)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_280),
.Y(n_305)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_225),
.Y(n_281)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_281),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_252),
.B(n_186),
.Y(n_282)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_282),
.Y(n_313)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_233),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_267),
.A2(n_226),
.B(n_240),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_289),
.A2(n_296),
.B(n_300),
.Y(n_334)
);

MAJx2_ASAP7_75t_L g292 ( 
.A(n_261),
.B(n_240),
.C(n_220),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_292),
.B(n_306),
.C(n_312),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_277),
.A2(n_283),
.B(n_242),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_283),
.A2(n_222),
.B1(n_240),
.B2(n_227),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_298),
.A2(n_300),
.B1(n_296),
.B2(n_315),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_277),
.A2(n_220),
.B(n_229),
.Y(n_300)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_303),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_256),
.A2(n_229),
.B(n_196),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_304),
.B(n_315),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_258),
.B(n_216),
.C(n_246),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_276),
.B(n_216),
.C(n_246),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_256),
.B(n_224),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_314),
.B(n_292),
.C(n_289),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_253),
.A2(n_233),
.B(n_228),
.Y(n_315)
);

INVx13_ASAP7_75t_L g316 ( 
.A(n_287),
.Y(n_316)
);

BUFx8_ASAP7_75t_L g356 ( 
.A(n_316),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_313),
.B(n_254),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_317),
.B(n_272),
.Y(n_365)
);

INVx13_ASAP7_75t_L g319 ( 
.A(n_287),
.Y(n_319)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_319),
.Y(n_373)
);

BUFx12f_ASAP7_75t_L g320 ( 
.A(n_290),
.Y(n_320)
);

INVx2_ASAP7_75t_SL g350 ( 
.A(n_320),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_305),
.B(n_255),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_322),
.B(n_323),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_313),
.B(n_235),
.Y(n_323)
);

INVx4_ASAP7_75t_L g324 ( 
.A(n_293),
.Y(n_324)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_324),
.Y(n_347)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_295),
.Y(n_325)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_325),
.Y(n_352)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_295),
.Y(n_326)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_326),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_286),
.B(n_257),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_327),
.B(n_333),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_286),
.B(n_309),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_328),
.B(n_329),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_307),
.Y(n_329)
);

MAJx2_ASAP7_75t_L g348 ( 
.A(n_330),
.B(n_297),
.C(n_312),
.Y(n_348)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_285),
.Y(n_331)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_331),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_332),
.A2(n_345),
.B1(n_297),
.B2(n_293),
.Y(n_349)
);

AND2x6_ASAP7_75t_L g333 ( 
.A(n_310),
.B(n_266),
.Y(n_333)
);

INVx13_ASAP7_75t_L g335 ( 
.A(n_299),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_335),
.Y(n_361)
);

BUFx2_ASAP7_75t_L g337 ( 
.A(n_305),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_337),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_310),
.B(n_235),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_338),
.B(n_340),
.Y(n_376)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_285),
.Y(n_339)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_339),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_306),
.B(n_251),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_311),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_341),
.B(n_342),
.Y(n_354)
);

BUFx5_ASAP7_75t_L g342 ( 
.A(n_304),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_291),
.B(n_263),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_343),
.B(n_344),
.Y(n_362)
);

AND2x6_ASAP7_75t_L g344 ( 
.A(n_314),
.B(n_274),
.Y(n_344)
);

CKINVDCx14_ASAP7_75t_R g345 ( 
.A(n_293),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_308),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_346),
.B(n_331),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_348),
.B(n_363),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_349),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_324),
.B(n_298),
.Y(n_355)
);

AOI21x1_ASAP7_75t_L g405 ( 
.A1(n_355),
.A2(n_259),
.B(n_262),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_318),
.B(n_291),
.C(n_308),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_357),
.B(n_377),
.C(n_326),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_332),
.A2(n_271),
.B1(n_222),
.B2(n_301),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_359),
.A2(n_321),
.B1(n_336),
.B2(n_339),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_SL g363 ( 
.A(n_330),
.B(n_318),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_337),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_364),
.B(n_320),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_365),
.B(n_224),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_327),
.A2(n_302),
.B1(n_301),
.B2(n_294),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_366),
.A2(n_367),
.B1(n_279),
.B2(n_319),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_336),
.A2(n_294),
.B1(n_302),
.B2(n_288),
.Y(n_367)
);

O2A1O1Ixp33_ASAP7_75t_L g370 ( 
.A1(n_334),
.A2(n_288),
.B(n_284),
.C(n_281),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_370),
.A2(n_342),
.B(n_335),
.Y(n_395)
);

AO22x1_ASAP7_75t_L g371 ( 
.A1(n_336),
.A2(n_275),
.B1(n_268),
.B2(n_260),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_371),
.B(n_321),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_343),
.B(n_275),
.Y(n_372)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_372),
.Y(n_381)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_374),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_317),
.B(n_228),
.C(n_251),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_378),
.A2(n_403),
.B1(n_367),
.B2(n_347),
.Y(n_408)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_379),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_382),
.B(n_385),
.C(n_391),
.Y(n_416)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_361),
.Y(n_383)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_383),
.Y(n_415)
);

AND2x2_ASAP7_75t_SL g411 ( 
.A(n_384),
.B(n_405),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_357),
.B(n_344),
.C(n_334),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_361),
.Y(n_386)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_386),
.Y(n_420)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_352),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_387),
.B(n_388),
.Y(n_406)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_353),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_355),
.A2(n_333),
.B(n_320),
.Y(n_389)
);

AOI21x1_ASAP7_75t_L g410 ( 
.A1(n_389),
.A2(n_355),
.B(n_362),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_368),
.B(n_325),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_390),
.B(n_392),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_348),
.B(n_225),
.C(n_231),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_358),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_366),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_393),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_394),
.B(n_350),
.Y(n_424)
);

OR2x2_ASAP7_75t_L g417 ( 
.A(n_395),
.B(n_399),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_368),
.B(n_372),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_396),
.B(n_397),
.Y(n_414)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_369),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_360),
.B(n_316),
.Y(n_399)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_354),
.Y(n_401)
);

NOR3xp33_ASAP7_75t_L g409 ( 
.A(n_401),
.B(n_402),
.C(n_351),
.Y(n_409)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_375),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_360),
.A2(n_152),
.B1(n_116),
.B2(n_137),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_404),
.B(n_262),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_408),
.A2(n_422),
.B1(n_424),
.B2(n_378),
.Y(n_437)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_409),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_410),
.A2(n_405),
.B(n_384),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_393),
.A2(n_359),
.B1(n_362),
.B2(n_371),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_418),
.A2(n_412),
.B1(n_424),
.B2(n_417),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_382),
.B(n_363),
.C(n_377),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_419),
.B(n_421),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_391),
.B(n_365),
.C(n_376),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_400),
.A2(n_370),
.B1(n_350),
.B2(n_356),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_398),
.B(n_350),
.C(n_373),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_423),
.B(n_427),
.C(n_395),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_380),
.B(n_356),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_425),
.B(n_426),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_385),
.B(n_356),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_398),
.B(n_223),
.C(n_137),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_428),
.B(n_390),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g429 ( 
.A(n_407),
.Y(n_429)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_429),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g455 ( 
.A(n_430),
.B(n_431),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_419),
.B(n_389),
.Y(n_431)
);

NOR2xp67_ASAP7_75t_SL g432 ( 
.A(n_416),
.B(n_399),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_432),
.A2(n_436),
.B(n_45),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_SL g433 ( 
.A(n_416),
.B(n_403),
.C(n_404),
.Y(n_433)
);

OR2x2_ASAP7_75t_L g456 ( 
.A(n_433),
.B(n_437),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_421),
.B(n_400),
.C(n_381),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_434),
.B(n_435),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_423),
.B(n_396),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_438),
.B(n_439),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_427),
.B(n_381),
.C(n_113),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_441),
.A2(n_446),
.B1(n_408),
.B2(n_411),
.Y(n_453)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_413),
.Y(n_444)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_444),
.Y(n_461)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_406),
.Y(n_445)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_445),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_422),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_417),
.A2(n_199),
.B1(n_183),
.B2(n_123),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_447),
.B(n_443),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_412),
.B(n_120),
.C(n_113),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_448),
.B(n_411),
.C(n_428),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_446),
.A2(n_418),
.B(n_424),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_450),
.A2(n_465),
.B(n_31),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_429),
.A2(n_411),
.B1(n_414),
.B2(n_415),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_451),
.B(n_454),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_452),
.B(n_111),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_453),
.Y(n_472)
);

FAx1_ASAP7_75t_SL g457 ( 
.A(n_434),
.B(n_420),
.CI(n_262),
.CON(n_457),
.SN(n_457)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_457),
.B(n_458),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_442),
.A2(n_213),
.B1(n_116),
.B2(n_212),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_440),
.B(n_204),
.C(n_273),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_460),
.B(n_464),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_462),
.A2(n_31),
.B(n_22),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_SL g464 ( 
.A(n_431),
.B(n_33),
.Y(n_464)
);

XOR2x2_ASAP7_75t_L g465 ( 
.A(n_438),
.B(n_430),
.Y(n_465)
);

OAI21xp5_ASAP7_75t_SL g467 ( 
.A1(n_456),
.A2(n_439),
.B(n_448),
.Y(n_467)
);

INVxp33_ASAP7_75t_SL g490 ( 
.A(n_467),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_455),
.B(n_111),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_468),
.B(n_471),
.Y(n_487)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_469),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_473),
.Y(n_493)
);

NOR2x1_ASAP7_75t_SL g474 ( 
.A(n_455),
.B(n_14),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_474),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_465),
.A2(n_456),
.B(n_459),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_475),
.A2(n_457),
.B1(n_458),
.B2(n_17),
.Y(n_489)
);

NAND3xp33_ASAP7_75t_L g478 ( 
.A(n_453),
.B(n_14),
.C(n_12),
.Y(n_478)
);

NOR3xp33_ASAP7_75t_L g486 ( 
.A(n_478),
.B(n_452),
.C(n_460),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_450),
.A2(n_106),
.B1(n_111),
.B2(n_22),
.Y(n_479)
);

AOI22xp33_ASAP7_75t_SL g488 ( 
.A1(n_479),
.A2(n_480),
.B1(n_481),
.B2(n_451),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_463),
.B(n_1),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_461),
.B(n_1),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_476),
.B(n_466),
.Y(n_482)
);

OR2x2_ASAP7_75t_L g501 ( 
.A(n_482),
.B(n_483),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_472),
.B(n_449),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_486),
.B(n_488),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_489),
.A2(n_491),
.B(n_17),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_478),
.B(n_457),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_477),
.B(n_17),
.C(n_3),
.Y(n_492)
);

NOR2xp67_ASAP7_75t_SL g498 ( 
.A(n_492),
.B(n_468),
.Y(n_498)
);

INVx6_ASAP7_75t_L g494 ( 
.A(n_490),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_494),
.B(n_498),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_493),
.B(n_480),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_495),
.A2(n_496),
.B(n_499),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_484),
.B(n_470),
.C(n_471),
.Y(n_496)
);

AOI21x1_ASAP7_75t_L g499 ( 
.A1(n_486),
.A2(n_17),
.B(n_4),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_500),
.B(n_2),
.Y(n_505)
);

A2O1A1Ixp33_ASAP7_75t_L g502 ( 
.A1(n_497),
.A2(n_485),
.B(n_487),
.C(n_8),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_L g507 ( 
.A1(n_502),
.A2(n_501),
.B(n_6),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_495),
.B(n_487),
.Y(n_503)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_503),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_505),
.B(n_506),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_507),
.A2(n_508),
.B1(n_504),
.B2(n_6),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_510),
.B(n_511),
.C(n_2),
.Y(n_512)
);

AOI21x1_ASAP7_75t_L g511 ( 
.A1(n_509),
.A2(n_2),
.B(n_8),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_512),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_513),
.B(n_11),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_514),
.B(n_11),
.Y(n_515)
);


endmodule