module real_jpeg_15410_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_470;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_0),
.A2(n_20),
.B(n_566),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_0),
.B(n_567),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_1),
.B(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_1),
.B(n_204),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_1),
.B(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_1),
.B(n_326),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_1),
.B(n_364),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_1),
.B(n_474),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_1),
.B(n_477),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_1),
.B(n_494),
.Y(n_493)
);

BUFx5_ASAP7_75t_L g168 ( 
.A(n_2),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_2),
.Y(n_250)
);

BUFx5_ASAP7_75t_L g297 ( 
.A(n_2),
.Y(n_297)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_2),
.Y(n_417)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_3),
.Y(n_567)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_4),
.Y(n_77)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_4),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g234 ( 
.A(n_4),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_5),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_5),
.B(n_35),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_5),
.B(n_88),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_5),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_5),
.B(n_236),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_5),
.B(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_5),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_5),
.B(n_168),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_6),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_6),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_6),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_6),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_6),
.B(n_154),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_6),
.B(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_6),
.B(n_257),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_6),
.A2(n_15),
.B1(n_295),
.B2(n_298),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g412 ( 
.A(n_6),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_7),
.B(n_62),
.Y(n_61)
);

INVxp33_ASAP7_75t_L g101 ( 
.A(n_7),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_7),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_7),
.B(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_7),
.B(n_199),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_7),
.B(n_306),
.Y(n_305)
);

AND2x4_ASAP7_75t_SL g323 ( 
.A(n_7),
.B(n_324),
.Y(n_323)
);

AND2x2_ASAP7_75t_SL g361 ( 
.A(n_7),
.B(n_168),
.Y(n_361)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_8),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_8),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_8),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_8),
.Y(n_313)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_8),
.Y(n_370)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_9),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g217 ( 
.A(n_9),
.Y(n_217)
);

BUFx4f_ASAP7_75t_L g254 ( 
.A(n_9),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_9),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_10),
.B(n_27),
.Y(n_26)
);

AND2x2_ASAP7_75t_SL g30 ( 
.A(n_10),
.B(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g44 ( 
.A(n_10),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_10),
.B(n_67),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_10),
.B(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_11),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_11),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_11),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_11),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_11),
.B(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_11),
.B(n_159),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_11),
.B(n_215),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_11),
.B(n_248),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_12),
.Y(n_96)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_12),
.Y(n_149)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_12),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_13),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g160 ( 
.A(n_13),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_13),
.Y(n_199)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_13),
.Y(n_321)
);

BUFx5_ASAP7_75t_L g508 ( 
.A(n_13),
.Y(n_508)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_14),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_14),
.B(n_59),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_14),
.B(n_240),
.Y(n_239)
);

AND2x2_ASAP7_75t_SL g262 ( 
.A(n_14),
.B(n_263),
.Y(n_262)
);

AND2x4_ASAP7_75t_SL g318 ( 
.A(n_14),
.B(n_319),
.Y(n_318)
);

AND2x4_ASAP7_75t_L g367 ( 
.A(n_14),
.B(n_368),
.Y(n_367)
);

AND2x4_ASAP7_75t_SL g420 ( 
.A(n_14),
.B(n_421),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_14),
.B(n_480),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_15),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_15),
.B(n_232),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_15),
.B(n_372),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_15),
.B(n_405),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_15),
.B(n_448),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_15),
.B(n_257),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_15),
.B(n_470),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_15),
.B(n_514),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_16),
.B(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_16),
.B(n_426),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_16),
.B(n_445),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_16),
.B(n_463),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_16),
.B(n_507),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_16),
.B(n_522),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_16),
.B(n_529),
.Y(n_528)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_17),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

BUFx8_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_18),
.Y(n_205)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_18),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_117),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_116),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_70),
.Y(n_22)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_23),
.B(n_70),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_51),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_38),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_30),
.C(n_34),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_26),
.A2(n_40),
.B1(n_45),
.B2(n_46),
.Y(n_39)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_26),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_26),
.A2(n_30),
.B1(n_45),
.B2(n_55),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_28),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_29),
.Y(n_301)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_30),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_30),
.B(n_61),
.C(n_65),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_30),
.A2(n_55),
.B1(n_65),
.B2(n_66),
.Y(n_111)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_33),
.Y(n_157)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_33),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_37),
.Y(n_202)
);

INVx4_ASAP7_75t_L g427 ( 
.A(n_37),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_47),
.Y(n_38)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_41),
.B(n_44),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OR2x2_ASAP7_75t_SL g106 ( 
.A(n_44),
.B(n_107),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_44),
.B(n_130),
.Y(n_129)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_56),
.C(n_60),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_52),
.A2(n_53),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_SL g115 ( 
.A(n_56),
.B(n_60),
.Y(n_115)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_61),
.B(n_111),
.Y(n_110)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_64),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_65),
.A2(n_66),
.B1(n_106),
.B2(n_127),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_66),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_SL g99 ( 
.A(n_66),
.B(n_100),
.C(n_106),
.Y(n_99)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_112),
.C(n_113),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_71),
.B(n_184),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_99),
.C(n_109),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_72),
.B(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_83),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_78),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_74),
.B(n_78),
.C(n_83),
.Y(n_112)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_82),
.Y(n_264)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_82),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_91),
.C(n_97),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_84),
.A2(n_85),
.B1(n_91),
.B2(n_92),
.Y(n_163)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g329 ( 
.A(n_90),
.Y(n_329)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g304 ( 
.A(n_96),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_97),
.B(n_163),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_99),
.B(n_110),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_100),
.B(n_177),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_105),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_106),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_106),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_106),
.B(n_128),
.C(n_133),
.Y(n_178)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_112),
.B(n_113),
.Y(n_184)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AOI21x1_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_284),
.B(n_561),
.Y(n_118)
);

NOR3x1_ASAP7_75t_SL g119 ( 
.A(n_120),
.B(n_185),
.C(n_278),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g561 ( 
.A1(n_120),
.A2(n_562),
.B(n_565),
.Y(n_561)
);

NOR2xp67_ASAP7_75t_R g120 ( 
.A(n_121),
.B(n_183),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_121),
.B(n_183),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_175),
.C(n_180),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_122),
.B(n_281),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_161),
.C(n_164),
.Y(n_122)
);

INVxp33_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_124),
.B(n_275),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_136),
.C(n_150),
.Y(n_124)
);

XNOR2x2_ASAP7_75t_SL g223 ( 
.A(n_125),
.B(n_224),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_126),
.B(n_133),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_128),
.A2(n_129),
.B1(n_167),
.B2(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

MAJx2_ASAP7_75t_L g166 ( 
.A(n_129),
.B(n_167),
.C(n_169),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_132),
.Y(n_422)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_136),
.B(n_150),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_141),
.C(n_145),
.Y(n_136)
);

XNOR2x1_ASAP7_75t_L g209 ( 
.A(n_137),
.B(n_145),
.Y(n_209)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx4_ASAP7_75t_L g366 ( 
.A(n_139),
.Y(n_366)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_140),
.Y(n_449)
);

XNOR2x1_ASAP7_75t_L g208 ( 
.A(n_141),
.B(n_209),
.Y(n_208)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_143),
.Y(n_324)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_151),
.B(n_153),
.C(n_158),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_158),
.Y(n_152)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_162),
.B(n_164),
.Y(n_275)
);

MAJx2_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_173),
.C(n_174),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_165),
.A2(n_166),
.B1(n_190),
.B2(n_192),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_166),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_167),
.B(n_211),
.C(n_213),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_167),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_167),
.A2(n_214),
.B1(n_222),
.B2(n_229),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_169),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_218)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_169),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_169),
.A2(n_219),
.B1(n_305),
.B2(n_356),
.Y(n_355)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_173),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_173),
.B(n_247),
.C(n_251),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_173),
.B(n_292),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g206 ( 
.A(n_174),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_174),
.A2(n_203),
.B1(n_206),
.B2(n_267),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_175),
.B(n_181),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.C(n_179),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_176),
.B(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_178),
.B(n_179),
.Y(n_273)
);

INVxp67_ASAP7_75t_SL g180 ( 
.A(n_181),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_268),
.Y(n_185)
);

NOR2x1_ASAP7_75t_L g563 ( 
.A(n_186),
.B(n_268),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_223),
.C(n_225),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_187),
.B(n_223),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_207),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_193),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_189),
.B(n_193),
.C(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_190),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_203),
.C(n_206),
.Y(n_193)
);

XNOR2x1_ASAP7_75t_L g265 ( 
.A(n_194),
.B(n_266),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_198),
.C(n_200),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_195),
.B(n_200),
.Y(n_244)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_198),
.B(n_244),
.Y(n_243)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_199),
.Y(n_237)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_203),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g212 ( 
.A(n_205),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_207),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.C(n_218),
.Y(n_207)
);

XNOR2x1_ASAP7_75t_L g339 ( 
.A(n_208),
.B(n_210),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_211),
.B(n_228),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_214),
.Y(n_229)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_217),
.Y(n_306)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_217),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_218),
.Y(n_338)
);

MAJx2_ASAP7_75t_L g302 ( 
.A(n_219),
.B(n_303),
.C(n_305),
.Y(n_302)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_225),
.B(n_383),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_245),
.C(n_265),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_226),
.B(n_336),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_230),
.C(n_243),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_227),
.B(n_230),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_235),
.C(n_238),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_231),
.A2(n_238),
.B1(n_239),
.B2(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_231),
.Y(n_380)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g378 ( 
.A(n_235),
.B(n_379),
.Y(n_378)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_238),
.B(n_444),
.C(n_447),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_238),
.A2(n_239),
.B1(n_444),
.B2(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx4_ASAP7_75t_L g465 ( 
.A(n_241),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_242),
.Y(n_373)
);

XNOR2x2_ASAP7_75t_L g348 ( 
.A(n_243),
.B(n_349),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_245),
.B(n_265),
.Y(n_336)
);

MAJx2_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_255),
.C(n_261),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_246),
.B(n_333),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_247),
.B(n_251),
.Y(n_292)
);

INVx6_ASAP7_75t_L g515 ( 
.A(n_248),
.Y(n_515)
);

INVx5_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_254),
.Y(n_478)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_256),
.B(n_262),
.Y(n_333)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_261),
.A2(n_262),
.B1(n_424),
.B2(n_425),
.Y(n_545)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_262),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_262),
.B(n_419),
.C(n_424),
.Y(n_418)
);

INVx2_ASAP7_75t_SL g263 ( 
.A(n_264),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_271),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_269),
.B(n_272),
.C(n_283),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_274),
.B1(n_276),
.B2(n_277),
.Y(n_271)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_272),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_274),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_277),
.Y(n_283)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g562 ( 
.A1(n_279),
.A2(n_563),
.B(n_564),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_282),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_280),
.B(n_282),
.Y(n_564)
);

AO21x2_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_388),
.B(n_558),
.Y(n_284)
);

NOR2xp67_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_381),
.Y(n_285)
);

AND2x2_ASAP7_75t_SL g286 ( 
.A(n_287),
.B(n_342),
.Y(n_286)
);

OR2x2_ASAP7_75t_L g559 ( 
.A(n_287),
.B(n_342),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_334),
.Y(n_287)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_288),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_307),
.C(n_330),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_290),
.B(n_346),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_293),
.C(n_302),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_291),
.B(n_429),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_293),
.A2(n_294),
.B1(n_302),
.B2(n_430),
.Y(n_429)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_294),
.A2(n_404),
.B(n_411),
.Y(n_403)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_297),
.Y(n_474)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_301),
.Y(n_446)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_302),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_303),
.B(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_305),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_308),
.A2(n_331),
.B1(n_332),
.B2(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_308),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_322),
.C(n_325),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_309),
.B(n_376),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_314),
.C(n_318),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_310),
.A2(n_318),
.B1(n_401),
.B2(n_402),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g402 ( 
.A(n_310),
.Y(n_402)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx6_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_314),
.B(n_400),
.Y(n_399)
);

INVx6_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_318),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_318),
.B(n_461),
.Y(n_460)
);

INVx6_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_322),
.A2(n_323),
.B1(n_325),
.B2(n_377),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_325),
.Y(n_377)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_335),
.A2(n_337),
.B1(n_340),
.B2(n_341),
.Y(n_334)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_335),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_337),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_337),
.Y(n_387)
);

XOR2x2_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_340),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_348),
.C(n_350),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_344),
.A2(n_345),
.B1(n_348),
.B2(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_348),
.Y(n_393)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_351),
.B(n_392),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_374),
.C(n_378),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_SL g396 ( 
.A(n_352),
.B(n_397),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_357),
.C(n_362),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

XNOR2x1_ASAP7_75t_L g452 ( 
.A(n_354),
.B(n_453),
.Y(n_452)
);

XNOR2x1_ASAP7_75t_L g453 ( 
.A(n_357),
.B(n_362),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_361),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_358),
.B(n_361),
.Y(n_451)
);

NOR2x1_ASAP7_75t_R g358 ( 
.A(n_359),
.B(n_360),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_367),
.C(n_371),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_363),
.B(n_439),
.Y(n_438)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_367),
.A2(n_371),
.B1(n_440),
.B2(n_441),
.Y(n_439)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_367),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_367),
.B(n_503),
.C(n_505),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_367),
.A2(n_441),
.B1(n_505),
.B2(n_506),
.Y(n_518)
);

INVx8_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_369),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_370),
.Y(n_524)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_371),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_375),
.B(n_378),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_L g558 ( 
.A1(n_381),
.A2(n_559),
.B(n_560),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_384),
.Y(n_381)
);

OR2x2_ASAP7_75t_L g560 ( 
.A(n_382),
.B(n_384),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_386),
.C(n_387),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_454),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_394),
.C(n_431),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_391),
.B(n_395),
.Y(n_557)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_398),
.C(n_428),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_396),
.B(n_433),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_398),
.B(n_428),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_403),
.C(n_418),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_399),
.B(n_403),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_401),
.B(n_462),
.C(n_466),
.Y(n_485)
);

INVx1_ASAP7_75t_SL g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_413),
.Y(n_411)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_417),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_418),
.B(n_436),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_SL g544 ( 
.A(n_419),
.B(n_545),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_423),
.Y(n_419)
);

XNOR2x1_ASAP7_75t_L g492 ( 
.A(n_420),
.B(n_423),
.Y(n_492)
);

CKINVDCx14_ASAP7_75t_R g512 ( 
.A(n_420),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_420),
.A2(n_512),
.B1(n_513),
.B2(n_526),
.Y(n_525)
);

INVx4_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

NOR2xp67_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_434),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_432),
.B(n_434),
.Y(n_556)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_437),
.C(n_452),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_435),
.B(n_554),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g554 ( 
.A(n_437),
.B(n_452),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_442),
.C(n_450),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_438),
.B(n_540),
.Y(n_539)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_443),
.B(n_451),
.Y(n_540)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_444),
.Y(n_488)
);

INVx4_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_447),
.B(n_487),
.Y(n_486)
);

INVx5_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

NAND3xp33_ASAP7_75t_L g454 ( 
.A(n_455),
.B(n_556),
.C(n_557),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_SL g455 ( 
.A1(n_456),
.A2(n_551),
.B(n_555),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_457),
.A2(n_536),
.B(n_550),
.Y(n_456)
);

OAI21x1_ASAP7_75t_L g457 ( 
.A1(n_458),
.A2(n_497),
.B(n_535),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_483),
.Y(n_458)
);

OR2x2_ASAP7_75t_L g535 ( 
.A(n_459),
.B(n_483),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_467),
.C(n_475),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_460),
.B(n_500),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_466),
.Y(n_461)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_467),
.A2(n_468),
.B1(n_475),
.B2(n_501),
.Y(n_500)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_473),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_SL g504 ( 
.A(n_469),
.B(n_473),
.Y(n_504)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_472),
.Y(n_531)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_475),
.Y(n_501)
);

AO22x1_ASAP7_75t_SL g475 ( 
.A1(n_476),
.A2(n_479),
.B1(n_481),
.B2(n_482),
.Y(n_475)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_476),
.Y(n_481)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_SL g482 ( 
.A(n_479),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_479),
.B(n_481),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_482),
.B(n_528),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_489),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_486),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_485),
.B(n_489),
.C(n_549),
.Y(n_548)
);

HB1xp67_ASAP7_75t_L g549 ( 
.A(n_486),
.Y(n_549)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_491),
.Y(n_489)
);

MAJx2_ASAP7_75t_L g547 ( 
.A(n_490),
.B(n_492),
.C(n_493),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_493),
.Y(n_491)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

AOI21x1_ASAP7_75t_L g497 ( 
.A1(n_498),
.A2(n_509),
.B(n_534),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_499),
.B(n_502),
.Y(n_498)
);

NOR2xp67_ASAP7_75t_SL g534 ( 
.A(n_499),
.B(n_502),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_503),
.A2(n_504),
.B1(n_517),
.B2(n_518),
.Y(n_516)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_510),
.A2(n_519),
.B(n_533),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_511),
.B(n_516),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_511),
.B(n_516),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_512),
.B(n_513),
.Y(n_511)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_513),
.Y(n_526)
);

INVx5_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_SL g519 ( 
.A1(n_520),
.A2(n_527),
.B(n_532),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_521),
.B(n_525),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_521),
.B(n_525),
.Y(n_532)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_524),
.Y(n_523)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_537),
.B(n_548),
.Y(n_536)
);

NOR2xp67_ASAP7_75t_SL g550 ( 
.A(n_537),
.B(n_548),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_538),
.A2(n_539),
.B1(n_541),
.B2(n_542),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_538),
.B(n_543),
.C(n_547),
.Y(n_552)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_543),
.A2(n_544),
.B1(n_546),
.B2(n_547),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

NOR2xp67_ASAP7_75t_L g551 ( 
.A(n_552),
.B(n_553),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_552),
.B(n_553),
.Y(n_555)
);


endmodule