module real_aes_2761_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_150;
wire n_147;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_481;
wire n_148;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_L g231 ( .A(n_0), .B(n_152), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_1), .B(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_2), .B(n_136), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_3), .B(n_154), .Y(n_509) );
INVx1_ASAP7_75t_L g143 ( .A(n_4), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_5), .B(n_136), .Y(n_135) );
NAND2xp33_ASAP7_75t_SL g222 ( .A(n_6), .B(n_142), .Y(n_222) );
INVx1_ASAP7_75t_L g203 ( .A(n_7), .Y(n_203) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_8), .Y(n_110) );
AND2x2_ASAP7_75t_L g130 ( .A(n_9), .B(n_131), .Y(n_130) );
XNOR2xp5_ASAP7_75t_L g121 ( .A(n_10), .B(n_122), .Y(n_121) );
AND2x2_ASAP7_75t_L g519 ( .A(n_10), .B(n_219), .Y(n_519) );
AND2x2_ASAP7_75t_L g511 ( .A(n_11), .B(n_193), .Y(n_511) );
INVx2_ASAP7_75t_L g132 ( .A(n_12), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_13), .B(n_154), .Y(n_528) );
XNOR2xp5_ASAP7_75t_L g480 ( .A(n_14), .B(n_481), .Y(n_480) );
CKINVDCx16_ASAP7_75t_R g112 ( .A(n_15), .Y(n_112) );
AOI221x1_ASAP7_75t_L g216 ( .A1(n_16), .A2(n_145), .B1(n_217), .B2(n_219), .C(n_221), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_17), .B(n_136), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_18), .B(n_136), .Y(n_542) );
INVx1_ASAP7_75t_L g114 ( .A(n_19), .Y(n_114) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_20), .A2(n_91), .B1(n_136), .B2(n_204), .Y(n_580) );
AOI21xp5_ASAP7_75t_L g144 ( .A1(n_21), .A2(n_145), .B(n_150), .Y(n_144) );
AOI221xp5_ASAP7_75t_SL g180 ( .A1(n_22), .A2(n_35), .B1(n_136), .B2(n_145), .C(n_181), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_23), .B(n_152), .Y(n_151) );
OR2x2_ASAP7_75t_L g133 ( .A(n_24), .B(n_90), .Y(n_133) );
OA21x2_ASAP7_75t_L g194 ( .A1(n_24), .A2(n_90), .B(n_132), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_25), .B(n_154), .Y(n_192) );
INVxp67_ASAP7_75t_L g215 ( .A(n_26), .Y(n_215) );
AND2x2_ASAP7_75t_L g176 ( .A(n_27), .B(n_166), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_28), .A2(n_145), .B(n_230), .Y(n_229) );
AO21x2_ASAP7_75t_L g523 ( .A1(n_29), .A2(n_219), .B(n_524), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_30), .B(n_154), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_31), .A2(n_145), .B(n_507), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_32), .B(n_154), .Y(n_537) );
AND2x2_ASAP7_75t_L g142 ( .A(n_33), .B(n_143), .Y(n_142) );
AND2x2_ASAP7_75t_L g146 ( .A(n_33), .B(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g211 ( .A(n_33), .Y(n_211) );
NOR3xp33_ASAP7_75t_L g108 ( .A(n_34), .B(n_109), .C(n_111), .Y(n_108) );
OR2x6_ASAP7_75t_L g470 ( .A(n_34), .B(n_471), .Y(n_470) );
XOR2xp5_ASAP7_75t_L g479 ( .A(n_36), .B(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_37), .B(n_136), .Y(n_510) );
AOI22xp5_ASAP7_75t_L g246 ( .A1(n_38), .A2(n_82), .B1(n_145), .B2(n_209), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_39), .B(n_154), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_40), .A2(n_74), .B1(n_461), .B2(n_462), .Y(n_460) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_40), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_41), .B(n_136), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_42), .B(n_152), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g795 ( .A(n_43), .Y(n_795) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_44), .A2(n_145), .B(n_515), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g473 ( .A(n_45), .B(n_474), .Y(n_473) );
AND2x2_ASAP7_75t_L g234 ( .A(n_46), .B(n_166), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_47), .B(n_152), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_48), .B(n_166), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_49), .B(n_136), .Y(n_525) );
OAI22xp5_ASAP7_75t_SL g458 ( .A1(n_50), .A2(n_459), .B1(n_460), .B2(n_463), .Y(n_458) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_50), .Y(n_463) );
INVx1_ASAP7_75t_L g139 ( .A(n_51), .Y(n_139) );
INVx1_ASAP7_75t_L g149 ( .A(n_51), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_52), .B(n_154), .Y(n_517) );
AND2x2_ASAP7_75t_L g553 ( .A(n_53), .B(n_166), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g175 ( .A(n_54), .B(n_136), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_55), .B(n_152), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_56), .B(n_152), .Y(n_536) );
AND2x2_ASAP7_75t_L g167 ( .A(n_57), .B(n_166), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_58), .B(n_136), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_59), .B(n_154), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_60), .B(n_136), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g534 ( .A1(n_61), .A2(n_145), .B(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_62), .B(n_152), .Y(n_163) );
AND2x2_ASAP7_75t_SL g195 ( .A(n_63), .B(n_131), .Y(n_195) );
AND2x2_ASAP7_75t_L g548 ( .A(n_64), .B(n_131), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g171 ( .A1(n_65), .A2(n_145), .B(n_172), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_66), .B(n_154), .Y(n_153) );
AND2x2_ASAP7_75t_SL g247 ( .A(n_67), .B(n_193), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_68), .B(n_152), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_69), .B(n_152), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_70), .A2(n_94), .B1(n_145), .B2(n_209), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_71), .B(n_154), .Y(n_545) );
INVx1_ASAP7_75t_L g141 ( .A(n_72), .Y(n_141) );
INVx1_ASAP7_75t_L g147 ( .A(n_72), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_73), .B(n_152), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g461 ( .A(n_74), .Y(n_461) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_75), .A2(n_145), .B(n_557), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_76), .A2(n_145), .B(n_499), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_77), .A2(n_145), .B(n_527), .Y(n_526) );
AND2x2_ASAP7_75t_L g539 ( .A(n_78), .B(n_131), .Y(n_539) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_79), .B(n_166), .Y(n_578) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_80), .B(n_136), .Y(n_164) );
AOI22xp5_ASAP7_75t_L g245 ( .A1(n_81), .A2(n_84), .B1(n_136), .B2(n_204), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_83), .B(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g472 ( .A(n_83), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_85), .B(n_152), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_86), .B(n_152), .Y(n_183) );
AND2x2_ASAP7_75t_L g502 ( .A(n_87), .B(n_193), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g799 ( .A(n_88), .Y(n_799) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_89), .A2(n_145), .B(n_161), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_92), .B(n_154), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_93), .A2(n_145), .B(n_544), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_95), .B(n_154), .Y(n_500) );
AOI22xp5_ASAP7_75t_L g481 ( .A1(n_96), .A2(n_103), .B1(n_482), .B2(n_483), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g482 ( .A(n_96), .Y(n_482) );
INVxp67_ASAP7_75t_L g218 ( .A(n_97), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_98), .B(n_136), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_99), .B(n_154), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_100), .A2(n_145), .B(n_190), .Y(n_189) );
BUFx2_ASAP7_75t_L g547 ( .A(n_101), .Y(n_547) );
BUFx2_ASAP7_75t_L g119 ( .A(n_102), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_102), .B(n_473), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_103), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_115), .B(n_798), .Y(n_104) );
BUFx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
BUFx8_ASAP7_75t_SL g800 ( .A(n_106), .Y(n_800) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
NAND2xp5_ASAP7_75t_SL g107 ( .A(n_108), .B(n_113), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_112), .B(n_469), .Y(n_468) );
AND2x6_ASAP7_75t_SL g488 ( .A(n_112), .B(n_470), .Y(n_488) );
OR2x6_ASAP7_75t_SL g790 ( .A(n_112), .B(n_469), .Y(n_790) );
OR2x2_ASAP7_75t_L g797 ( .A(n_112), .B(n_470), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_114), .B(n_472), .Y(n_471) );
OA22x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_120), .B1(n_477), .B2(n_478), .Y(n_115) );
CKINVDCx11_ASAP7_75t_R g116 ( .A(n_117), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI21xp5_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_464), .B(n_473), .Y(n_120) );
OAI22x1_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_124), .B1(n_457), .B2(n_458), .Y(n_122) );
OAI22x1_ASAP7_75t_L g792 ( .A1(n_123), .A2(n_485), .B1(n_790), .B2(n_793), .Y(n_792) );
INVx4_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OAI22xp5_ASAP7_75t_L g484 ( .A1(n_124), .A2(n_485), .B1(n_489), .B2(n_788), .Y(n_484) );
AND2x4_ASAP7_75t_L g124 ( .A(n_125), .B(n_368), .Y(n_124) );
NOR3xp33_ASAP7_75t_L g125 ( .A(n_126), .B(n_290), .C(n_340), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g126 ( .A(n_127), .B(n_257), .Y(n_126) );
AOI221xp5_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_177), .B1(n_196), .B2(n_239), .C(n_249), .Y(n_127) );
INVx1_ASAP7_75t_SL g339 ( .A(n_128), .Y(n_339) );
AND2x4_ASAP7_75t_SL g128 ( .A(n_129), .B(n_157), .Y(n_128) );
INVx2_ASAP7_75t_L g261 ( .A(n_129), .Y(n_261) );
OR2x2_ASAP7_75t_L g283 ( .A(n_129), .B(n_274), .Y(n_283) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_129), .Y(n_298) );
INVx5_ASAP7_75t_L g305 ( .A(n_129), .Y(n_305) );
AND2x4_ASAP7_75t_L g311 ( .A(n_129), .B(n_169), .Y(n_311) );
AND2x2_ASAP7_75t_SL g314 ( .A(n_129), .B(n_241), .Y(n_314) );
OR2x2_ASAP7_75t_L g323 ( .A(n_129), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g330 ( .A(n_129), .B(n_158), .Y(n_330) );
AND2x2_ASAP7_75t_L g431 ( .A(n_129), .B(n_168), .Y(n_431) );
OR2x6_ASAP7_75t_L g129 ( .A(n_130), .B(n_134), .Y(n_129) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_131), .Y(n_166) );
AND2x2_ASAP7_75t_SL g131 ( .A(n_132), .B(n_133), .Y(n_131) );
AND2x4_ASAP7_75t_L g156 ( .A(n_132), .B(n_133), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_144), .B(n_156), .Y(n_134) );
AND2x4_ASAP7_75t_L g136 ( .A(n_137), .B(n_142), .Y(n_136) );
INVx1_ASAP7_75t_L g223 ( .A(n_137), .Y(n_223) );
AND2x4_ASAP7_75t_L g137 ( .A(n_138), .B(n_140), .Y(n_137) );
AND2x6_ASAP7_75t_L g152 ( .A(n_138), .B(n_147), .Y(n_152) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x4_ASAP7_75t_L g154 ( .A(n_140), .B(n_149), .Y(n_154) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx5_ASAP7_75t_L g155 ( .A(n_142), .Y(n_155) );
AND2x2_ASAP7_75t_L g148 ( .A(n_143), .B(n_149), .Y(n_148) );
HB1xp67_ASAP7_75t_L g207 ( .A(n_143), .Y(n_207) );
AND2x6_ASAP7_75t_L g145 ( .A(n_146), .B(n_148), .Y(n_145) );
BUFx3_ASAP7_75t_L g208 ( .A(n_146), .Y(n_208) );
INVx2_ASAP7_75t_L g213 ( .A(n_147), .Y(n_213) );
AND2x4_ASAP7_75t_L g209 ( .A(n_148), .B(n_210), .Y(n_209) );
INVx2_ASAP7_75t_L g206 ( .A(n_149), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_153), .B(n_155), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_152), .B(n_547), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_155), .A2(n_162), .B(n_163), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_155), .A2(n_173), .B(n_174), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_155), .A2(n_182), .B(n_183), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_155), .A2(n_191), .B(n_192), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_155), .A2(n_231), .B(n_232), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_155), .A2(n_500), .B(n_501), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_155), .A2(n_508), .B(n_509), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_155), .A2(n_516), .B(n_517), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_155), .A2(n_528), .B(n_529), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_155), .A2(n_536), .B(n_537), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_155), .A2(n_545), .B(n_546), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_155), .A2(n_558), .B(n_559), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_156), .B(n_203), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g214 ( .A(n_156), .B(n_215), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_156), .B(n_218), .Y(n_217) );
NOR3xp33_ASAP7_75t_L g221 ( .A(n_156), .B(n_222), .C(n_223), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_156), .A2(n_525), .B(n_526), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g554 ( .A1(n_156), .A2(n_555), .B(n_556), .Y(n_554) );
INVx3_ASAP7_75t_SL g282 ( .A(n_157), .Y(n_282) );
AND2x2_ASAP7_75t_L g326 ( .A(n_157), .B(n_241), .Y(n_326) );
OAI21xp5_ASAP7_75t_L g329 ( .A1(n_157), .A2(n_330), .B(n_331), .Y(n_329) );
AND2x2_ASAP7_75t_L g367 ( .A(n_157), .B(n_305), .Y(n_367) );
AND2x4_ASAP7_75t_L g157 ( .A(n_158), .B(n_168), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_158), .B(n_169), .Y(n_248) );
OR2x2_ASAP7_75t_L g252 ( .A(n_158), .B(n_169), .Y(n_252) );
INVx1_ASAP7_75t_L g260 ( .A(n_158), .Y(n_260) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_158), .Y(n_272) );
INVx2_ASAP7_75t_L g280 ( .A(n_158), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_158), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g389 ( .A(n_158), .B(n_274), .Y(n_389) );
AND2x2_ASAP7_75t_L g404 ( .A(n_158), .B(n_241), .Y(n_404) );
AO21x2_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_165), .B(n_167), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_160), .B(n_164), .Y(n_159) );
AO21x2_ASAP7_75t_L g169 ( .A1(n_165), .A2(n_170), .B(n_176), .Y(n_169) );
AO21x2_ASAP7_75t_L g324 ( .A1(n_165), .A2(n_170), .B(n_176), .Y(n_324) );
AOI21x1_ASAP7_75t_L g504 ( .A1(n_165), .A2(n_505), .B(n_511), .Y(n_504) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_166), .Y(n_165) );
OA21x2_ASAP7_75t_L g179 ( .A1(n_166), .A2(n_180), .B(n_184), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_166), .A2(n_497), .B(n_498), .Y(n_496) );
AO21x2_ASAP7_75t_L g579 ( .A1(n_166), .A2(n_580), .B(n_581), .Y(n_579) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AND2x2_ASAP7_75t_L g273 ( .A(n_169), .B(n_274), .Y(n_273) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_169), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_171), .B(n_175), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_177), .B(n_397), .Y(n_396) );
NOR2x1p5_ASAP7_75t_L g177 ( .A(n_178), .B(n_185), .Y(n_177) );
BUFx3_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AND2x2_ASAP7_75t_L g225 ( .A(n_179), .B(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_179), .B(n_186), .Y(n_255) );
INVx1_ASAP7_75t_L g265 ( .A(n_179), .Y(n_265) );
INVx2_ASAP7_75t_L g288 ( .A(n_179), .Y(n_288) );
INVx2_ASAP7_75t_L g294 ( .A(n_179), .Y(n_294) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_179), .Y(n_364) );
OR2x2_ASAP7_75t_L g395 ( .A(n_179), .B(n_186), .Y(n_395) );
OR2x2_ASAP7_75t_L g411 ( .A(n_185), .B(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AND2x4_ASAP7_75t_SL g199 ( .A(n_186), .B(n_200), .Y(n_199) );
AND2x4_ASAP7_75t_L g237 ( .A(n_186), .B(n_238), .Y(n_237) );
OR2x2_ASAP7_75t_L g275 ( .A(n_186), .B(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g287 ( .A(n_186), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g300 ( .A(n_186), .B(n_266), .Y(n_300) );
OR2x2_ASAP7_75t_L g308 ( .A(n_186), .B(n_200), .Y(n_308) );
INVx2_ASAP7_75t_L g335 ( .A(n_186), .Y(n_335) );
INVx1_ASAP7_75t_L g353 ( .A(n_186), .Y(n_353) );
NOR2xp33_ASAP7_75t_R g386 ( .A(n_186), .B(n_226), .Y(n_386) );
OR2x6_ASAP7_75t_L g186 ( .A(n_187), .B(n_195), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B(n_193), .Y(n_187) );
INVx2_ASAP7_75t_SL g243 ( .A(n_193), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_193), .A2(n_542), .B(n_543), .Y(n_541) );
BUFx4f_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx3_ASAP7_75t_L g220 ( .A(n_194), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_197), .B(n_235), .Y(n_196) );
OAI22xp5_ASAP7_75t_L g277 ( .A1(n_197), .A2(n_278), .B1(n_281), .B2(n_284), .Y(n_277) );
OR2x2_ASAP7_75t_L g197 ( .A(n_198), .B(n_224), .Y(n_197) );
INVx1_ASAP7_75t_SL g198 ( .A(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g292 ( .A(n_199), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g327 ( .A(n_199), .B(n_328), .Y(n_327) );
AND2x4_ASAP7_75t_L g406 ( .A(n_199), .B(n_384), .Y(n_406) );
INVx3_ASAP7_75t_L g238 ( .A(n_200), .Y(n_238) );
AND2x4_ASAP7_75t_L g266 ( .A(n_200), .B(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_200), .B(n_226), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_200), .B(n_288), .Y(n_333) );
AND2x2_ASAP7_75t_L g338 ( .A(n_200), .B(n_335), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_200), .B(n_225), .Y(n_375) );
INVx1_ASAP7_75t_L g445 ( .A(n_200), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_200), .B(n_363), .Y(n_456) );
AND2x4_ASAP7_75t_L g200 ( .A(n_201), .B(n_216), .Y(n_200) );
AOI22xp5_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_204), .B1(n_209), .B2(n_214), .Y(n_201) );
AND2x4_ASAP7_75t_L g204 ( .A(n_205), .B(n_208), .Y(n_204) );
AND2x2_ASAP7_75t_L g205 ( .A(n_206), .B(n_207), .Y(n_205) );
NOR2x1p5_ASAP7_75t_L g210 ( .A(n_211), .B(n_212), .Y(n_210) );
INVx3_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx3_ASAP7_75t_L g532 ( .A(n_219), .Y(n_532) );
INVx4_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
AOI21x1_ASAP7_75t_L g227 ( .A1(n_220), .A2(n_228), .B(n_234), .Y(n_227) );
AO21x2_ASAP7_75t_L g512 ( .A1(n_220), .A2(n_513), .B(n_519), .Y(n_512) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g236 ( .A(n_226), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_226), .B(n_238), .Y(n_256) );
INVx2_ASAP7_75t_L g267 ( .A(n_226), .Y(n_267) );
AND2x2_ASAP7_75t_L g293 ( .A(n_226), .B(n_294), .Y(n_293) );
OR2x2_ASAP7_75t_L g309 ( .A(n_226), .B(n_288), .Y(n_309) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_226), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_226), .B(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g398 ( .A(n_226), .Y(n_398) );
INVx3_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_229), .B(n_233), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_236), .B(n_237), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_236), .B(n_265), .Y(n_276) );
AOI221x1_ASAP7_75t_SL g370 ( .A1(n_237), .A2(n_371), .B1(n_374), .B2(n_376), .C(n_380), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_237), .B(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g428 ( .A(n_237), .B(n_293), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_237), .B(n_450), .Y(n_449) );
OR2x2_ASAP7_75t_L g359 ( .A(n_238), .B(n_287), .Y(n_359) );
AND2x2_ASAP7_75t_L g397 ( .A(n_238), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_SL g239 ( .A(n_240), .Y(n_239) );
OR2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_248), .Y(n_240) );
AND2x2_ASAP7_75t_L g250 ( .A(n_241), .B(n_251), .Y(n_250) );
INVx2_ASAP7_75t_L g345 ( .A(n_241), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g350 ( .A(n_241), .B(n_261), .Y(n_350) );
AND2x4_ASAP7_75t_L g379 ( .A(n_241), .B(n_280), .Y(n_379) );
NAND2xp5_ASAP7_75t_SL g415 ( .A(n_241), .B(n_311), .Y(n_415) );
OR2x2_ASAP7_75t_L g433 ( .A(n_241), .B(n_364), .Y(n_433) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_241), .B(n_324), .Y(n_443) );
BUFx6f_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx2_ASAP7_75t_L g274 ( .A(n_242), .Y(n_274) );
AOI21x1_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_244), .B(n_247), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
INVx1_ASAP7_75t_L g299 ( .A(n_248), .Y(n_299) );
OAI22xp5_ASAP7_75t_L g306 ( .A1(n_248), .A2(n_307), .B1(n_310), .B2(n_312), .Y(n_306) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_253), .Y(n_249) );
INVx2_ASAP7_75t_L g262 ( .A(n_250), .Y(n_262) );
AND2x2_ASAP7_75t_L g401 ( .A(n_251), .B(n_261), .Y(n_401) );
AND2x2_ASAP7_75t_L g447 ( .A(n_251), .B(n_314), .Y(n_447) );
AND2x2_ASAP7_75t_L g452 ( .A(n_251), .B(n_303), .Y(n_452) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AOI32xp33_ASAP7_75t_L g421 ( .A1(n_253), .A2(n_323), .A3(n_403), .B1(n_422), .B2(n_424), .Y(n_421) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
OR2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
INVx1_ASAP7_75t_L g289 ( .A(n_256), .Y(n_289) );
AOI211xp5_ASAP7_75t_SL g257 ( .A1(n_258), .A2(n_263), .B(n_268), .C(n_277), .Y(n_257) );
OAI21xp5_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_261), .B(n_262), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_260), .B(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_261), .B(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g441 ( .A(n_261), .Y(n_441) );
AND2x2_ASAP7_75t_L g351 ( .A(n_263), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_SL g263 ( .A(n_264), .B(n_266), .Y(n_263) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_264), .Y(n_451) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVxp67_ASAP7_75t_SL g320 ( .A(n_265), .Y(n_320) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_265), .Y(n_420) );
INVx1_ASAP7_75t_L g317 ( .A(n_266), .Y(n_317) );
AND2x2_ASAP7_75t_L g383 ( .A(n_266), .B(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_266), .B(n_394), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_269), .B(n_275), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
OAI21xp33_ASAP7_75t_L g349 ( .A1(n_270), .A2(n_350), .B(n_351), .Y(n_349) );
AND2x2_ASAP7_75t_SL g270 ( .A(n_271), .B(n_273), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g279 ( .A(n_274), .B(n_280), .Y(n_279) );
BUFx2_ASAP7_75t_L g303 ( .A(n_274), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_279), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g410 ( .A(n_279), .Y(n_410) );
AND2x2_ASAP7_75t_L g440 ( .A(n_279), .B(n_441), .Y(n_440) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_280), .Y(n_417) );
OR2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_283), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_282), .B(n_430), .Y(n_429) );
INVx1_ASAP7_75t_SL g357 ( .A(n_283), .Y(n_357) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x4_ASAP7_75t_L g285 ( .A(n_286), .B(n_289), .Y(n_285) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g316 ( .A(n_287), .B(n_317), .Y(n_316) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_288), .Y(n_384) );
AND2x2_ASAP7_75t_L g393 ( .A(n_289), .B(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_313), .Y(n_290) );
AOI221xp5_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_295), .B1(n_300), .B2(n_301), .C(n_306), .Y(n_291) );
INVx1_ASAP7_75t_L g412 ( .A(n_293), .Y(n_412) );
INVxp33_ASAP7_75t_SL g444 ( .A(n_293), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g390 ( .A1(n_295), .A2(n_391), .B(n_399), .Y(n_390) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_SL g296 ( .A(n_297), .B(n_299), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_299), .B(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g312 ( .A(n_300), .Y(n_312) );
AND2x2_ASAP7_75t_L g347 ( .A(n_300), .B(n_348), .Y(n_347) );
AND2x2_ASAP7_75t_L g366 ( .A(n_300), .B(n_367), .Y(n_366) );
AOI22xp33_ASAP7_75t_SL g427 ( .A1(n_300), .A2(n_428), .B1(n_429), .B2(n_432), .Y(n_427) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OR2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
OR2x2_ASAP7_75t_L g322 ( .A(n_303), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_303), .B(n_311), .Y(n_361) );
AND2x4_ASAP7_75t_L g378 ( .A(n_305), .B(n_324), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_305), .B(n_379), .Y(n_425) );
AND2x2_ASAP7_75t_L g437 ( .A(n_305), .B(n_389), .Y(n_437) );
NAND2xp33_ASAP7_75t_L g422 ( .A(n_307), .B(n_423), .Y(n_422) );
OR2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
INVx1_ASAP7_75t_SL g365 ( .A(n_308), .Y(n_365) );
INVx1_ASAP7_75t_L g436 ( .A(n_309), .Y(n_436) );
INVx2_ASAP7_75t_SL g388 ( .A(n_311), .Y(n_388) );
AOI211xp5_ASAP7_75t_SL g313 ( .A1(n_314), .A2(n_315), .B(n_318), .C(n_336), .Y(n_313) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OAI211xp5_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_322), .B(n_325), .C(n_329), .Y(n_318) );
OR2x6_ASAP7_75t_SL g319 ( .A(n_320), .B(n_321), .Y(n_319) );
INVx1_ASAP7_75t_L g348 ( .A(n_320), .Y(n_348) );
INVx1_ASAP7_75t_SL g373 ( .A(n_323), .Y(n_373) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_323), .B(n_433), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_328), .B(n_338), .Y(n_337) );
INVx2_ASAP7_75t_SL g331 ( .A(n_332), .Y(n_331) );
OAI22xp33_ASAP7_75t_L g414 ( .A1(n_332), .A2(n_415), .B1(n_416), .B2(n_418), .Y(n_414) );
OR2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_337), .B(n_339), .Y(n_336) );
OAI211xp5_ASAP7_75t_SL g340 ( .A1(n_341), .A2(n_346), .B(n_349), .C(n_354), .Y(n_340) );
INVxp67_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_343), .B(n_345), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AOI221xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_358), .B1(n_360), .B2(n_362), .C(n_366), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_SL g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_365), .Y(n_362) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AOI222xp33_ASAP7_75t_L g446 ( .A1(n_365), .A2(n_447), .B1(n_448), .B2(n_452), .C1(n_453), .C2(n_455), .Y(n_446) );
INVx2_ASAP7_75t_L g381 ( .A(n_367), .Y(n_381) );
NOR3xp33_ASAP7_75t_L g368 ( .A(n_369), .B(n_407), .C(n_426), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_370), .B(n_390), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVxp67_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_378), .B(n_417), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_379), .B(n_441), .Y(n_454) );
OAI22xp33_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_382), .B1(n_385), .B2(n_387), .Y(n_380) );
INVx1_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
INVxp33_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_388), .B(n_410), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_392), .B(n_396), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_SL g394 ( .A(n_395), .Y(n_394) );
OAI22xp5_ASAP7_75t_L g399 ( .A1(n_396), .A2(n_400), .B1(n_402), .B2(n_405), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
BUFx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
CKINVDCx16_ASAP7_75t_R g405 ( .A(n_406), .Y(n_405) );
OAI211xp5_ASAP7_75t_SL g407 ( .A1(n_408), .A2(n_411), .B(n_413), .C(n_421), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVxp67_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
NAND3xp33_ASAP7_75t_L g426 ( .A(n_427), .B(n_434), .C(n_446), .Y(n_426) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OAI21xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_438), .B(n_445), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
AOI21xp5_ASAP7_75t_L g438 ( .A1(n_439), .A2(n_442), .B(n_444), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVxp33_ASAP7_75t_SL g457 ( .A(n_458), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_460), .Y(n_459) );
CKINVDCx11_ASAP7_75t_R g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_SL g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_SL g466 ( .A(n_467), .Y(n_466) );
BUFx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
BUFx3_ASAP7_75t_L g476 ( .A(n_468), .Y(n_476) );
CKINVDCx5p33_ASAP7_75t_R g469 ( .A(n_470), .Y(n_469) );
BUFx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
CKINVDCx20_ASAP7_75t_R g475 ( .A(n_476), .Y(n_475) );
AO221x1_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_484), .B1(n_791), .B2(n_792), .C(n_794), .Y(n_478) );
INVx1_ASAP7_75t_L g791 ( .A(n_479), .Y(n_791) );
CKINVDCx11_ASAP7_75t_R g485 ( .A(n_486), .Y(n_485) );
INVx3_ASAP7_75t_SL g486 ( .A(n_487), .Y(n_486) );
CKINVDCx5p33_ASAP7_75t_R g487 ( .A(n_488), .Y(n_487) );
INVx5_ASAP7_75t_L g793 ( .A(n_489), .Y(n_793) );
AND2x4_ASAP7_75t_L g489 ( .A(n_490), .B(n_692), .Y(n_489) );
NOR3xp33_ASAP7_75t_L g490 ( .A(n_491), .B(n_617), .C(n_653), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_492), .B(n_591), .Y(n_491) );
AOI211xp5_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_520), .B(n_549), .C(n_574), .Y(n_492) );
AND2x2_ASAP7_75t_L g682 ( .A(n_493), .B(n_551), .Y(n_682) );
AND2x2_ASAP7_75t_L g493 ( .A(n_494), .B(n_503), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_494), .B(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g715 ( .A(n_494), .B(n_597), .Y(n_715) );
AND2x2_ASAP7_75t_L g731 ( .A(n_494), .B(n_566), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_494), .B(n_741), .Y(n_740) );
NAND2x1p5_ASAP7_75t_L g764 ( .A(n_494), .B(n_765), .Y(n_764) );
INVx4_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AND2x4_ASAP7_75t_SL g561 ( .A(n_495), .B(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g586 ( .A(n_495), .Y(n_586) );
AND2x2_ASAP7_75t_L g633 ( .A(n_495), .B(n_576), .Y(n_633) );
AND2x2_ASAP7_75t_L g652 ( .A(n_495), .B(n_503), .Y(n_652) );
BUFx2_ASAP7_75t_L g657 ( .A(n_495), .Y(n_657) );
AND2x2_ASAP7_75t_L g701 ( .A(n_495), .B(n_512), .Y(n_701) );
AND2x4_ASAP7_75t_L g773 ( .A(n_495), .B(n_774), .Y(n_773) );
NOR2x1_ASAP7_75t_L g785 ( .A(n_495), .B(n_565), .Y(n_785) );
OR2x6_ASAP7_75t_L g495 ( .A(n_496), .B(n_502), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_503), .B(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g704 ( .A(n_503), .Y(n_704) );
BUFx2_ASAP7_75t_L g753 ( .A(n_503), .Y(n_753) );
INVx1_ASAP7_75t_L g775 ( .A(n_503), .Y(n_775) );
AND2x2_ASAP7_75t_L g503 ( .A(n_504), .B(n_512), .Y(n_503) );
INVx3_ASAP7_75t_L g562 ( .A(n_504), .Y(n_562) );
HB1xp67_ASAP7_75t_L g741 ( .A(n_504), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_510), .Y(n_505) );
INVx2_ASAP7_75t_L g565 ( .A(n_512), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_512), .B(n_562), .Y(n_566) );
INVx2_ASAP7_75t_L g641 ( .A(n_512), .Y(n_641) );
OR2x2_ASAP7_75t_L g648 ( .A(n_512), .B(n_597), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_518), .Y(n_513) );
AND2x2_ASAP7_75t_L g603 ( .A(n_520), .B(n_604), .Y(n_603) );
AND2x2_ASAP7_75t_L g637 ( .A(n_520), .B(n_600), .Y(n_637) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_530), .Y(n_520) );
AND2x2_ASAP7_75t_L g673 ( .A(n_521), .B(n_572), .Y(n_673) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g630 ( .A(n_522), .B(n_531), .Y(n_630) );
AND2x2_ASAP7_75t_L g749 ( .A(n_522), .B(n_540), .Y(n_749) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g571 ( .A(n_523), .Y(n_571) );
INVx1_ASAP7_75t_L g589 ( .A(n_523), .Y(n_589) );
AND2x2_ASAP7_75t_L g645 ( .A(n_523), .B(n_531), .Y(n_645) );
AND2x2_ASAP7_75t_L g650 ( .A(n_523), .B(n_552), .Y(n_650) );
OR2x2_ASAP7_75t_L g713 ( .A(n_523), .B(n_540), .Y(n_713) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_523), .Y(n_722) );
AND2x2_ASAP7_75t_L g551 ( .A(n_530), .B(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g590 ( .A(n_530), .Y(n_590) );
NOR2x1_ASAP7_75t_SL g530 ( .A(n_531), .B(n_540), .Y(n_530) );
AO21x1_ASAP7_75t_SL g531 ( .A1(n_532), .A2(n_533), .B(n_539), .Y(n_531) );
AO21x2_ASAP7_75t_L g573 ( .A1(n_532), .A2(n_533), .B(n_539), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_538), .Y(n_533) );
AND2x2_ASAP7_75t_L g568 ( .A(n_540), .B(n_569), .Y(n_568) );
INVx2_ASAP7_75t_SL g616 ( .A(n_540), .Y(n_616) );
NAND2x1_ASAP7_75t_L g626 ( .A(n_540), .B(n_552), .Y(n_626) );
OR2x2_ASAP7_75t_L g631 ( .A(n_540), .B(n_569), .Y(n_631) );
BUFx2_ASAP7_75t_L g687 ( .A(n_540), .Y(n_687) );
AND2x2_ASAP7_75t_L g723 ( .A(n_540), .B(n_602), .Y(n_723) );
AND2x2_ASAP7_75t_L g734 ( .A(n_540), .B(n_572), .Y(n_734) );
OR2x6_ASAP7_75t_L g540 ( .A(n_541), .B(n_548), .Y(n_540) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AOI22xp5_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_560), .B1(n_566), .B2(n_567), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g780 ( .A1(n_551), .A2(n_731), .B1(n_781), .B2(n_786), .Y(n_780) );
INVx4_ASAP7_75t_L g569 ( .A(n_552), .Y(n_569) );
INVx2_ASAP7_75t_L g600 ( .A(n_552), .Y(n_600) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_552), .Y(n_671) );
OR2x2_ASAP7_75t_L g686 ( .A(n_552), .B(n_572), .Y(n_686) );
OR2x2_ASAP7_75t_SL g712 ( .A(n_552), .B(n_713), .Y(n_712) );
OR2x6_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
AND2x2_ASAP7_75t_SL g560 ( .A(n_561), .B(n_563), .Y(n_560) );
INVx2_ASAP7_75t_SL g593 ( .A(n_561), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_561), .B(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g661 ( .A(n_561), .B(n_609), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_561), .B(n_699), .Y(n_698) );
INVx2_ASAP7_75t_L g583 ( .A(n_562), .Y(n_583) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_562), .Y(n_608) );
AND2x2_ASAP7_75t_L g664 ( .A(n_562), .B(n_641), .Y(n_664) );
INVx1_ASAP7_75t_L g774 ( .A(n_562), .Y(n_774) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_564), .B(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_564), .B(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g582 ( .A(n_565), .B(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_566), .B(n_715), .Y(n_714) );
AOI321xp33_ASAP7_75t_L g736 ( .A1(n_567), .A2(n_638), .A3(n_706), .B1(n_737), .B2(n_738), .C(n_742), .Y(n_736) );
AND2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_570), .Y(n_567) );
INVxp67_ASAP7_75t_SL g635 ( .A(n_568), .Y(n_635) );
AND2x2_ASAP7_75t_L g660 ( .A(n_568), .B(n_589), .Y(n_660) );
AND2x2_ASAP7_75t_L g735 ( .A(n_568), .B(n_645), .Y(n_735) );
INVx1_ASAP7_75t_L g604 ( .A(n_569), .Y(n_604) );
BUFx2_ASAP7_75t_L g614 ( .A(n_569), .Y(n_614) );
NOR2xp67_ASAP7_75t_L g721 ( .A(n_569), .B(n_722), .Y(n_721) );
INVx1_ASAP7_75t_SL g659 ( .A(n_570), .Y(n_659) );
AND2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
BUFx2_ASAP7_75t_L g666 ( .A(n_571), .Y(n_666) );
INVx2_ASAP7_75t_L g602 ( .A(n_572), .Y(n_602) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_572), .Y(n_625) );
INVx3_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AOI21xp33_ASAP7_75t_SL g574 ( .A1(n_575), .A2(n_584), .B(n_587), .Y(n_574) );
NOR2xp67_ASAP7_75t_L g718 ( .A(n_575), .B(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_582), .Y(n_576) );
INVx3_ASAP7_75t_L g609 ( .A(n_577), .Y(n_609) );
AND2x2_ASAP7_75t_L g640 ( .A(n_577), .B(n_641), .Y(n_640) );
AND2x4_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
AND2x4_ASAP7_75t_L g597 ( .A(n_578), .B(n_579), .Y(n_597) );
INVx1_ASAP7_75t_L g680 ( .A(n_582), .Y(n_680) );
INVx1_ASAP7_75t_SL g765 ( .A(n_583), .Y(n_765) );
INVxp33_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_SL g639 ( .A(n_586), .B(n_640), .Y(n_639) );
OR2x2_ASAP7_75t_L g691 ( .A(n_586), .B(n_648), .Y(n_691) );
OR2x2_ASAP7_75t_L g587 ( .A(n_588), .B(n_590), .Y(n_587) );
AND2x2_ASAP7_75t_L g695 ( .A(n_588), .B(n_696), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_588), .B(n_710), .Y(n_709) );
INVx3_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_589), .B(n_626), .Y(n_681) );
NOR4xp25_ASAP7_75t_L g776 ( .A(n_589), .B(n_620), .C(n_777), .D(n_778), .Y(n_776) );
OR2x2_ASAP7_75t_L g744 ( .A(n_590), .B(n_745), .Y(n_744) );
AOI221xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_598), .B1(n_603), .B2(n_605), .C(n_610), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
AND2x2_ASAP7_75t_L g619 ( .A(n_594), .B(n_620), .Y(n_619) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OR2x2_ASAP7_75t_L g656 ( .A(n_595), .B(n_657), .Y(n_656) );
INVx2_ASAP7_75t_L g676 ( .A(n_596), .Y(n_676) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
BUFx3_ASAP7_75t_L g699 ( .A(n_597), .Y(n_699) );
AND2x2_ASAP7_75t_L g706 ( .A(n_597), .B(n_707), .Y(n_706) );
INVxp67_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
OR2x2_ASAP7_75t_L g643 ( .A(n_600), .B(n_644), .Y(n_643) );
INVxp67_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_602), .B(n_616), .Y(n_615) );
INVxp67_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
OR2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_609), .Y(n_606) );
INVx2_ASAP7_75t_L g620 ( .A(n_607), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_607), .B(n_690), .Y(n_689) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g612 ( .A(n_609), .Y(n_612) );
OAI321xp33_ASAP7_75t_L g724 ( .A1(n_609), .A2(n_717), .A3(n_725), .B1(n_730), .B2(n_732), .C(n_736), .Y(n_724) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_611), .B(n_613), .Y(n_610) );
OR2x2_ASAP7_75t_L g679 ( .A(n_612), .B(n_680), .Y(n_679) );
OR2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
INVx1_ASAP7_75t_L g779 ( .A(n_615), .Y(n_779) );
NOR2xp33_ASAP7_75t_L g658 ( .A(n_616), .B(n_659), .Y(n_658) );
NAND2xp33_ASAP7_75t_SL g759 ( .A(n_616), .B(n_630), .Y(n_759) );
OAI211xp5_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_621), .B(n_632), .C(n_636), .Y(n_617) );
INVxp67_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
NOR2x1_ASAP7_75t_L g621 ( .A(n_622), .B(n_627), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OR2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_626), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g728 ( .A(n_625), .Y(n_728) );
INVx3_ASAP7_75t_L g667 ( .A(n_626), .Y(n_667) );
OR2x2_ASAP7_75t_L g770 ( .A(n_626), .B(n_644), .Y(n_770) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_628), .A2(n_712), .B1(n_714), .B2(n_716), .Y(n_711) );
OR2x2_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_SL g710 ( .A(n_631), .Y(n_710) );
OR2x2_ASAP7_75t_L g787 ( .A(n_631), .B(n_644), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
AOI21xp5_ASAP7_75t_SL g636 ( .A1(n_637), .A2(n_638), .B(n_642), .Y(n_636) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_640), .B(n_657), .Y(n_756) );
AND2x2_ASAP7_75t_L g762 ( .A(n_640), .B(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g707 ( .A(n_641), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_646), .B1(n_649), .B2(n_651), .Y(n_642) );
A2O1A1Ixp33_ASAP7_75t_L g688 ( .A1(n_644), .A2(n_687), .B(n_689), .C(n_691), .Y(n_688) );
INVx2_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_647), .B(n_717), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_647), .B(n_739), .Y(n_761) );
INVx2_ASAP7_75t_SL g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g733 ( .A(n_650), .B(n_734), .Y(n_733) );
INVx2_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
A2O1A1Ixp33_ASAP7_75t_L g683 ( .A1(n_652), .A2(n_684), .B(n_687), .C(n_688), .Y(n_683) );
NAND3xp33_ASAP7_75t_SL g653 ( .A(n_654), .B(n_668), .C(n_683), .Y(n_653) );
AOI222xp33_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_658), .B1(n_660), .B2(n_661), .C1(n_662), .C2(n_665), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx2_ASAP7_75t_L g717 ( .A(n_657), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_657), .B(n_690), .Y(n_743) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_SL g677 ( .A(n_664), .Y(n_677) );
AND2x2_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .Y(n_665) );
OR2x2_ASAP7_75t_L g782 ( .A(n_666), .B(n_699), .Y(n_782) );
AOI22xp5_ASAP7_75t_L g757 ( .A1(n_667), .A2(n_758), .B1(n_760), .B2(n_762), .Y(n_757) );
AOI221xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_674), .B1(n_678), .B2(n_681), .C(n_682), .Y(n_668) );
INVx2_ASAP7_75t_SL g669 ( .A(n_670), .Y(n_669) );
OR2x2_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .Y(n_670) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AOI21xp5_ASAP7_75t_SL g742 ( .A1(n_675), .A2(n_743), .B(n_744), .Y(n_742) );
OR2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_677), .Y(n_675) );
INVx2_ASAP7_75t_L g690 ( .A(n_676), .Y(n_690) );
AND2x2_ASAP7_75t_L g784 ( .A(n_676), .B(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx2_ASAP7_75t_L g768 ( .A(n_680), .Y(n_768) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
HB1xp67_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
OR2x2_ASAP7_75t_L g697 ( .A(n_686), .B(n_687), .Y(n_697) );
INVx1_ASAP7_75t_L g750 ( .A(n_686), .Y(n_750) );
NOR3xp33_ASAP7_75t_L g692 ( .A(n_693), .B(n_724), .C(n_746), .Y(n_692) );
OAI211xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_698), .B(n_700), .C(n_705), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
OAI21xp33_ASAP7_75t_L g700 ( .A1(n_695), .A2(n_701), .B(n_702), .Y(n_700) );
INVx1_ASAP7_75t_SL g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
AOI211xp5_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_708), .B(n_711), .C(n_718), .Y(n_705) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx2_ASAP7_75t_L g729 ( .A(n_712), .Y(n_729) );
INVxp67_ASAP7_75t_SL g754 ( .A(n_713), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_715), .B(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g777 ( .A(n_715), .Y(n_777) );
AND2x2_ASAP7_75t_L g767 ( .A(n_717), .B(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g737 ( .A(n_719), .Y(n_737) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
AND2x2_ASAP7_75t_L g720 ( .A(n_721), .B(n_723), .Y(n_720) );
INVx1_ASAP7_75t_L g745 ( .A(n_721), .Y(n_745) );
INVx2_ASAP7_75t_SL g725 ( .A(n_726), .Y(n_725) );
AND2x4_ASAP7_75t_L g726 ( .A(n_727), .B(n_729), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_SL g730 ( .A(n_731), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g732 ( .A(n_733), .B(n_735), .Y(n_732) );
AOI221xp5_ASAP7_75t_L g766 ( .A1(n_733), .A2(n_767), .B1(n_769), .B2(n_771), .C(n_776), .Y(n_766) );
OAI21xp33_ASAP7_75t_SL g781 ( .A1(n_738), .A2(n_782), .B(n_783), .Y(n_781) );
INVx2_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
NAND4xp25_ASAP7_75t_L g746 ( .A(n_747), .B(n_757), .C(n_766), .D(n_780), .Y(n_746) );
AOI22xp5_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_751), .B1(n_754), .B2(n_755), .Y(n_747) );
AND2x4_ASAP7_75t_L g748 ( .A(n_749), .B(n_750), .Y(n_748) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_SL g755 ( .A(n_756), .Y(n_755) );
INVxp67_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx2_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_772), .B(n_775), .Y(n_771) );
INVx2_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx2_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx1_ASAP7_75t_SL g788 ( .A(n_789), .Y(n_788) );
CKINVDCx11_ASAP7_75t_R g789 ( .A(n_790), .Y(n_789) );
NOR2xp33_ASAP7_75t_L g794 ( .A(n_795), .B(n_796), .Y(n_794) );
BUFx2_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
NOR2xp33_ASAP7_75t_L g798 ( .A(n_799), .B(n_800), .Y(n_798) );
endmodule