module fake_jpeg_4891_n_279 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_279);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_279;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_155;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx11_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_35),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_19),
.B(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_39),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_1),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_40),
.B(n_33),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

AND2x2_ASAP7_75t_SL g42 ( 
.A(n_37),
.B(n_26),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_42),
.A2(n_18),
.B1(n_36),
.B2(n_40),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_44),
.B(n_35),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_38),
.A2(n_16),
.B1(n_22),
.B2(n_27),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_46),
.A2(n_47),
.B1(n_48),
.B2(n_52),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_34),
.A2(n_27),
.B1(n_32),
.B2(n_16),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_34),
.A2(n_35),
.B1(n_38),
.B2(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_54),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_16),
.B1(n_22),
.B2(n_32),
.Y(n_52)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_57),
.Y(n_64)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx8_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_58),
.Y(n_70)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_59),
.B(n_33),
.Y(n_72)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

AO22x1_ASAP7_75t_SL g62 ( 
.A1(n_42),
.A2(n_26),
.B1(n_23),
.B2(n_18),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_62),
.A2(n_51),
.B1(n_43),
.B2(n_33),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_SL g107 ( 
.A(n_63),
.B(n_25),
.C(n_24),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_45),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_65),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_41),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_66),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_41),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_67),
.B(n_69),
.Y(n_92)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_75),
.Y(n_99)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_78),
.Y(n_101)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_53),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_80),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_57),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_44),
.B(n_39),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_30),
.Y(n_91)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

OAI21xp33_ASAP7_75t_L g97 ( 
.A1(n_86),
.A2(n_20),
.B(n_3),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_49),
.A2(n_35),
.B1(n_34),
.B2(n_40),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_87),
.A2(n_20),
.B1(n_40),
.B2(n_23),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_59),
.B(n_30),
.Y(n_88)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_88),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_69),
.A2(n_49),
.B1(n_55),
.B2(n_36),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_90),
.A2(n_106),
.B1(n_108),
.B2(n_70),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_107),
.Y(n_122)
);

FAx1_ASAP7_75t_SL g93 ( 
.A(n_84),
.B(n_23),
.CI(n_33),
.CON(n_93),
.SN(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_93),
.A2(n_85),
.B(n_67),
.C(n_66),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_97),
.B(n_100),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_79),
.A2(n_23),
.B(n_21),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_102),
.A2(n_29),
.B(n_68),
.Y(n_117)
);

AND2x2_ASAP7_75t_SL g103 ( 
.A(n_77),
.B(n_33),
.Y(n_103)
);

AND2x2_ASAP7_75t_SL g141 ( 
.A(n_103),
.B(n_25),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_74),
.A2(n_71),
.B1(n_65),
.B2(n_62),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_77),
.B(n_21),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_109),
.B(n_113),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_62),
.B(n_43),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_112),
.A2(n_114),
.B(n_64),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_77),
.B(n_21),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_21),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_115),
.B(n_118),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_116),
.A2(n_126),
.B1(n_131),
.B2(n_133),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_117),
.A2(n_119),
.B(n_120),
.Y(n_146)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_109),
.A2(n_68),
.B(n_61),
.Y(n_119)
);

AND2x4_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_24),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_104),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_121),
.Y(n_147)
);

INVx2_ASAP7_75t_SL g123 ( 
.A(n_94),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_123),
.B(n_127),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_110),
.Y(n_124)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_125),
.A2(n_129),
.B1(n_98),
.B2(n_25),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_108),
.A2(n_78),
.B1(n_75),
.B2(n_31),
.Y(n_126)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_89),
.Y(n_127)
);

AOI32xp33_ASAP7_75t_L g128 ( 
.A1(n_101),
.A2(n_31),
.A3(n_28),
.B1(n_17),
.B2(n_76),
.Y(n_128)
);

CKINVDCx12_ASAP7_75t_R g169 ( 
.A(n_128),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_76),
.Y(n_130)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_130),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_112),
.A2(n_28),
.B1(n_17),
.B2(n_31),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_96),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_132),
.B(n_134),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_112),
.A2(n_28),
.B1(n_81),
.B2(n_82),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_91),
.A2(n_25),
.B(n_24),
.Y(n_135)
);

MAJx2_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_102),
.C(n_93),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_92),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_136),
.Y(n_155)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_139),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_93),
.B(n_1),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_96),
.B(n_83),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_140),
.B(n_89),
.Y(n_143)
);

OA22x2_ASAP7_75t_L g150 ( 
.A1(n_141),
.A2(n_114),
.B1(n_107),
.B2(n_95),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_145),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_144),
.A2(n_122),
.B(n_142),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_126),
.Y(n_145)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_133),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_148),
.B(n_162),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_129),
.A2(n_106),
.B1(n_113),
.B2(n_95),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_149),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_150),
.A2(n_117),
.B(n_121),
.Y(n_179)
);

AND2x6_ASAP7_75t_L g153 ( 
.A(n_115),
.B(n_114),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_153),
.B(n_120),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_111),
.C(n_98),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_165),
.C(n_167),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_111),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_136),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_138),
.A2(n_25),
.B1(n_24),
.B2(n_73),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_125),
.A2(n_24),
.B1(n_73),
.B2(n_15),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_118),
.B(n_15),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_132),
.B(n_3),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_164),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_3),
.C(n_4),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_116),
.C(n_120),
.Y(n_167)
);

MAJx2_ASAP7_75t_L g170 ( 
.A(n_141),
.B(n_4),
.C(n_5),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_170),
.B(n_6),
.Y(n_188)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_123),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_171),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_182),
.Y(n_199)
);

A2O1A1O1Ixp25_ASAP7_75t_L g173 ( 
.A1(n_153),
.A2(n_120),
.B(n_122),
.C(n_119),
.D(n_135),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_173),
.B(n_188),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_175),
.B(n_178),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_163),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_177),
.B(n_192),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_157),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_179),
.A2(n_184),
.B(n_196),
.Y(n_217)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_168),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_180),
.B(n_185),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_167),
.B(n_122),
.C(n_131),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_149),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_146),
.A2(n_134),
.B(n_123),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_158),
.B(n_127),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_5),
.Y(n_186)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_186),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_148),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g201 ( 
.A(n_187),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_160),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_150),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_147),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_191),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_171),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_151),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_161),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_146),
.A2(n_6),
.B(n_7),
.Y(n_196)
);

NAND2x1_ASAP7_75t_L g197 ( 
.A(n_172),
.B(n_150),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_200),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_150),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_203),
.B(n_207),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_186),
.B(n_175),
.Y(n_205)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_205),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_174),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_190),
.Y(n_208)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_208),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_210),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_211),
.Y(n_221)
);

AOI21x1_ASAP7_75t_L g213 ( 
.A1(n_184),
.A2(n_144),
.B(n_170),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_196),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_178),
.B(n_154),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_214),
.B(n_181),
.Y(n_227)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_190),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_215),
.B(n_173),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_179),
.A2(n_156),
.B1(n_155),
.B2(n_169),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_216),
.B(n_182),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_212),
.Y(n_218)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_218),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_208),
.A2(n_189),
.B1(n_156),
.B2(n_180),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_220),
.A2(n_233),
.B1(n_198),
.B2(n_216),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_222),
.A2(n_228),
.B1(n_223),
.B2(n_231),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_200),
.B(n_183),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_223),
.B(n_227),
.C(n_231),
.Y(n_238)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_224),
.Y(n_235)
);

AOI21xp33_ASAP7_75t_L g225 ( 
.A1(n_197),
.A2(n_213),
.B(n_214),
.Y(n_225)
);

A2O1A1Ixp33_ASAP7_75t_L g242 ( 
.A1(n_225),
.A2(n_197),
.B(n_217),
.C(n_209),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_199),
.B(n_181),
.Y(n_231)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_232),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_215),
.A2(n_203),
.B1(n_210),
.B2(n_206),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_230),
.A2(n_217),
.B(n_206),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_234),
.A2(n_236),
.B(n_243),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_218),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_237),
.B(n_240),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_219),
.B(n_152),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_232),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_241),
.B(n_229),
.Y(n_250)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_242),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_226),
.A2(n_198),
.B(n_204),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_222),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_234),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_247),
.B(n_250),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_14),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_229),
.C(n_199),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_251),
.B(n_254),
.C(n_255),
.Y(n_262)
);

OAI321xp33_ASAP7_75t_L g253 ( 
.A1(n_236),
.A2(n_201),
.A3(n_221),
.B1(n_205),
.B2(n_195),
.C(n_202),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_253),
.A2(n_239),
.B1(n_235),
.B2(n_245),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_239),
.A2(n_209),
.B(n_202),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_176),
.C(n_165),
.Y(n_255)
);

NOR2x1_ASAP7_75t_L g256 ( 
.A(n_252),
.B(n_243),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_256),
.A2(n_249),
.B1(n_251),
.B2(n_10),
.Y(n_265)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_257),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_252),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_260),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_246),
.A2(n_242),
.B1(n_194),
.B2(n_166),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_248),
.A2(n_155),
.B1(n_188),
.B2(n_10),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_9),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_263),
.B(n_255),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_264),
.B(n_263),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_265),
.B(n_268),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_7),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_259),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_270),
.B(n_271),
.Y(n_274)
);

OAI21x1_ASAP7_75t_SL g272 ( 
.A1(n_267),
.A2(n_258),
.B(n_262),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_272),
.B(n_266),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_275),
.A2(n_269),
.B(n_273),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_276),
.B(n_274),
.Y(n_277)
);

OAI321xp33_ASAP7_75t_L g278 ( 
.A1(n_277),
.A2(n_9),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.C(n_256),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_12),
.Y(n_279)
);


endmodule