module fake_jpeg_13476_n_178 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_178);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_178;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g50 ( 
.A(n_29),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_26),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_6),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_11),
.B(n_23),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_16),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_48),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g66 ( 
.A(n_31),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_44),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_10),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_7),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_2),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_0),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_40),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_37),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_3),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_77),
.Y(n_88)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

BUFx4f_ASAP7_75t_SL g80 ( 
.A(n_68),
.Y(n_80)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_80),
.Y(n_97)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_0),
.Y(n_83)
);

BUFx8_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_76),
.A2(n_72),
.B1(n_52),
.B2(n_58),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_87),
.A2(n_89),
.B1(n_67),
.B2(n_3),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_81),
.A2(n_58),
.B1(n_68),
.B2(n_61),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_78),
.A2(n_50),
.B1(n_59),
.B2(n_62),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_93),
.A2(n_94),
.B1(n_96),
.B2(n_66),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g94 ( 
.A1(n_79),
.A2(n_69),
.B1(n_74),
.B2(n_73),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_60),
.B1(n_53),
.B2(n_65),
.Y(n_96)
);

BUFx12_ASAP7_75t_L g99 ( 
.A(n_80),
.Y(n_99)
);

BUFx4f_ASAP7_75t_SL g115 ( 
.A(n_99),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_95),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_100),
.A2(n_118),
.B1(n_104),
.B2(n_109),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_99),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_106),
.Y(n_128)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_103),
.B(n_110),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_92),
.A2(n_75),
.B1(n_66),
.B2(n_64),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_104),
.A2(n_114),
.B(n_8),
.Y(n_123)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_97),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_97),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_113),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_75),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

OA22x2_ASAP7_75t_L g109 ( 
.A1(n_89),
.A2(n_80),
.B1(n_64),
.B2(n_67),
.Y(n_109)
);

OAI32xp33_ASAP7_75t_L g138 ( 
.A1(n_109),
.A2(n_8),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_1),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_111),
.B(n_112),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_86),
.B(n_1),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_4),
.Y(n_113)
);

OR2x2_ASAP7_75t_SL g114 ( 
.A(n_98),
.B(n_4),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_90),
.B(n_5),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_116),
.B(n_119),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_91),
.A2(n_5),
.B(n_6),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_120),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_91),
.A2(n_28),
.B1(n_45),
.B2(n_43),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_85),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_7),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_123),
.A2(n_130),
.B(n_138),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_132),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_108),
.A2(n_27),
.B(n_41),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_131),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_25),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_113),
.B(n_46),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_135),
.B(n_139),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_115),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_30),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_39),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_9),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_140),
.B(n_141),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_115),
.B(n_12),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_114),
.B(n_38),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_142),
.B(n_35),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_136),
.A2(n_12),
.B(n_13),
.Y(n_143)
);

AO21x1_ASAP7_75t_L g164 ( 
.A1(n_143),
.A2(n_135),
.B(n_139),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_146),
.B(n_150),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_122),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_147),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_136),
.A2(n_14),
.B1(n_18),
.B2(n_22),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_121),
.Y(n_151)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_123),
.A2(n_33),
.B(n_34),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_152),
.A2(n_130),
.B(n_127),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_SL g153 ( 
.A(n_133),
.B(n_142),
.C(n_132),
.Y(n_153)
);

BUFx24_ASAP7_75t_SL g161 ( 
.A(n_153),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_128),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_125),
.C(n_129),
.Y(n_160)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_156),
.B(n_157),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_160),
.B(n_164),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_165),
.B(n_143),
.Y(n_170)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_159),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_167),
.A2(n_169),
.B1(n_170),
.B2(n_154),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_166),
.B(n_149),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_171),
.B(n_172),
.Y(n_173)
);

AOI321xp33_ASAP7_75t_L g172 ( 
.A1(n_168),
.A2(n_161),
.A3(n_144),
.B1(n_158),
.B2(n_163),
.C(n_164),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_173),
.B(n_170),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_174),
.B(n_157),
.C(n_158),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_175),
.A2(n_148),
.B(n_162),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_176),
.A2(n_138),
.B1(n_147),
.B2(n_150),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_145),
.Y(n_178)
);


endmodule