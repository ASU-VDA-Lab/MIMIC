module fake_jpeg_12925_n_460 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_460);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_460;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx24_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_11),
.B(n_8),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_40),
.B(n_9),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_47),
.B(n_83),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_48),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_9),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_54),
.B(n_84),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_55),
.Y(n_115)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_59),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_61),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_62),
.Y(n_108)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_65),
.Y(n_124)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_66),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_68),
.Y(n_130)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_70),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_17),
.Y(n_71)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_71),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_36),
.Y(n_74)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_74),
.Y(n_122)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_76),
.Y(n_127)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_80),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_79),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_81),
.B(n_82),
.Y(n_125)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_42),
.B(n_9),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_86),
.Y(n_94)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_16),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_88),
.Y(n_106)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_89),
.B(n_90),
.Y(n_126)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_49),
.B(n_19),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_99),
.B(n_129),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_63),
.A2(n_73),
.B1(n_81),
.B2(n_80),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_104),
.A2(n_119),
.B1(n_137),
.B2(n_20),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_57),
.A2(n_16),
.B1(n_37),
.B2(n_41),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_107),
.A2(n_110),
.B1(n_120),
.B2(n_123),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_49),
.A2(n_16),
.B1(n_37),
.B2(n_41),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_44),
.A2(n_37),
.B1(n_79),
.B2(n_74),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_60),
.A2(n_30),
.B1(n_38),
.B2(n_26),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_46),
.A2(n_61),
.B1(n_72),
.B2(n_50),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_53),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_51),
.A2(n_30),
.B1(n_38),
.B2(n_26),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_L g162 ( 
.A1(n_132),
.A2(n_35),
.B1(n_43),
.B2(n_20),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_60),
.B(n_18),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_135),
.B(n_27),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_56),
.A2(n_30),
.B1(n_38),
.B2(n_26),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_136),
.A2(n_69),
.B1(n_43),
.B2(n_35),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_55),
.A2(n_18),
.B1(n_39),
.B2(n_19),
.Y(n_137)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_143),
.Y(n_198)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_134),
.Y(n_144)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_144),
.Y(n_189)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_114),
.Y(n_145)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_145),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_126),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_146),
.B(n_158),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_147),
.A2(n_167),
.B(n_142),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_97),
.A2(n_20),
.B1(n_28),
.B2(n_31),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_32),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_149),
.B(n_150),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_32),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_117),
.Y(n_151)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_151),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_152),
.B(n_159),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_125),
.A2(n_58),
.B1(n_68),
.B2(n_67),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_153),
.A2(n_176),
.B1(n_128),
.B2(n_115),
.Y(n_205)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_96),
.Y(n_154)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_154),
.Y(n_192)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_140),
.Y(n_155)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_155),
.Y(n_214)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_122),
.Y(n_157)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_157),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_106),
.Y(n_158)
);

OAI21xp33_ASAP7_75t_L g159 ( 
.A1(n_121),
.A2(n_66),
.B(n_27),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_98),
.Y(n_160)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_160),
.Y(n_199)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_98),
.Y(n_161)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_161),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_162),
.A2(n_128),
.B1(n_92),
.B2(n_103),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_105),
.A2(n_76),
.B1(n_78),
.B2(n_45),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_164),
.Y(n_194)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_116),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_165),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_94),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_166),
.B(n_168),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_125),
.A2(n_28),
.B(n_31),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_102),
.B(n_39),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_169),
.B(n_170),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_105),
.B(n_77),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_141),
.Y(n_171)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_171),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_133),
.Y(n_172)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_172),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_127),
.B(n_65),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_174),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_132),
.B(n_43),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_93),
.Y(n_175)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_175),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_108),
.A2(n_62),
.B1(n_59),
.B2(n_89),
.Y(n_176)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_91),
.Y(n_177)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_177),
.Y(n_217)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_116),
.Y(n_178)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_178),
.Y(n_213)
);

AND2x4_ASAP7_75t_L g179 ( 
.A(n_124),
.B(n_70),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_179),
.A2(n_181),
.B(n_93),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_91),
.Y(n_180)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_180),
.Y(n_216)
);

AOI32xp33_ASAP7_75t_L g181 ( 
.A1(n_110),
.A2(n_31),
.A3(n_28),
.B1(n_35),
.B2(n_4),
.Y(n_181)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_118),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_182),
.A2(n_185),
.B1(n_186),
.B2(n_142),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_108),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_183),
.B(n_184),
.Y(n_208)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_109),
.Y(n_184)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_131),
.Y(n_185)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_118),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_152),
.A2(n_107),
.B1(n_120),
.B2(n_136),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_190),
.A2(n_205),
.B1(n_210),
.B2(n_179),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_191),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_196),
.A2(n_179),
.B(n_164),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_206),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_174),
.A2(n_115),
.B1(n_130),
.B2(n_109),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_149),
.B(n_130),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_211),
.B(n_215),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_150),
.B(n_139),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_220),
.A2(n_103),
.B1(n_112),
.B2(n_177),
.Y(n_247)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_217),
.Y(n_222)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_222),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_208),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_223),
.B(n_236),
.Y(n_258)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_188),
.Y(n_224)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_224),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_145),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_230),
.C(n_244),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_195),
.B(n_156),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_227),
.Y(n_252)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_188),
.Y(n_228)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_228),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_229),
.A2(n_219),
.B(n_212),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_197),
.B(n_170),
.C(n_179),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_208),
.Y(n_231)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_231),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_195),
.B(n_144),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_232),
.B(n_233),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_209),
.B(n_167),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_207),
.A2(n_163),
.B1(n_112),
.B2(n_92),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_234),
.A2(n_237),
.B1(n_239),
.B2(n_243),
.Y(n_268)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_199),
.Y(n_235)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_235),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_202),
.B(n_162),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_143),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_238),
.B(n_241),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_207),
.A2(n_170),
.B1(n_160),
.B2(n_161),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_209),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_187),
.A2(n_165),
.B1(n_178),
.B2(n_95),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_242),
.A2(n_100),
.B1(n_101),
.B2(n_131),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_207),
.A2(n_157),
.B1(n_151),
.B2(n_184),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_197),
.B(n_154),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_199),
.Y(n_245)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_245),
.Y(n_272)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_200),
.Y(n_246)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_246),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_247),
.A2(n_205),
.B1(n_210),
.B2(n_216),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_215),
.B(n_155),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_248),
.B(n_250),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_191),
.B(n_171),
.C(n_186),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_213),
.C(n_193),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_200),
.B(n_196),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_240),
.A2(n_194),
.B(n_220),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_253),
.A2(n_234),
.B(n_230),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_226),
.B(n_218),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_254),
.B(n_259),
.C(n_265),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_232),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_255),
.B(n_257),
.Y(n_303)
);

FAx1_ASAP7_75t_SL g257 ( 
.A(n_250),
.B(n_218),
.CI(n_194),
.CON(n_257),
.SN(n_257)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_244),
.B(n_203),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_225),
.B(n_203),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_266),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_267),
.A2(n_274),
.B1(n_277),
.B2(n_275),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_240),
.A2(n_216),
.B1(n_217),
.B2(n_180),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_276),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_271),
.B(n_239),
.C(n_245),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_231),
.A2(n_217),
.B1(n_213),
.B2(n_201),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_224),
.Y(n_275)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_275),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_236),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_228),
.Y(n_277)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_277),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_278),
.A2(n_229),
.B(n_273),
.Y(n_284)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_260),
.Y(n_280)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_280),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_264),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_281),
.B(n_299),
.Y(n_317)
);

OA21x2_ASAP7_75t_L g282 ( 
.A1(n_273),
.A2(n_237),
.B(n_243),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_282),
.B(n_257),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_255),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g329 ( 
.A(n_283),
.Y(n_329)
);

AO22x1_ASAP7_75t_L g326 ( 
.A1(n_284),
.A2(n_286),
.B1(n_289),
.B2(n_257),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_278),
.A2(n_221),
.B(n_249),
.Y(n_285)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_285),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_258),
.A2(n_223),
.B(n_241),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_256),
.B(n_225),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_292),
.B(n_295),
.C(n_300),
.Y(n_315)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_260),
.Y(n_293)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_293),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_256),
.B(n_233),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_SL g333 ( 
.A(n_294),
.B(n_302),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_276),
.A2(n_238),
.B1(n_248),
.B2(n_221),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_296),
.A2(n_297),
.B1(n_307),
.B2(n_268),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_258),
.A2(n_227),
.B1(n_235),
.B2(n_247),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_264),
.B(n_246),
.Y(n_298)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_298),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_274),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_254),
.B(n_201),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_259),
.B(n_193),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_268),
.A2(n_222),
.B1(n_212),
.B2(n_219),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_304),
.A2(n_267),
.B1(n_291),
.B2(n_251),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_269),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_305),
.B(n_252),
.Y(n_323)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_261),
.Y(n_306)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_306),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_271),
.B(n_214),
.C(n_204),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_309),
.C(n_279),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_265),
.B(n_214),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_282),
.Y(n_310)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_310),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_311),
.A2(n_336),
.B1(n_291),
.B2(n_272),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_289),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_312),
.B(n_325),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_314),
.A2(n_324),
.B1(n_270),
.B2(n_272),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_298),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_318),
.B(n_321),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_292),
.B(n_269),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_319),
.B(n_192),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_320),
.B(n_308),
.C(n_288),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_282),
.Y(n_321)
);

CKINVDCx14_ASAP7_75t_R g349 ( 
.A(n_323),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_286),
.A2(n_262),
.B1(n_257),
.B2(n_253),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_303),
.B(n_283),
.Y(n_325)
);

XNOR2x2_ASAP7_75t_SL g340 ( 
.A(n_326),
.B(n_302),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_284),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_330),
.B(n_332),
.Y(n_339)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_280),
.Y(n_331)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_331),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_295),
.B(n_262),
.Y(n_332)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_293),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_334),
.Y(n_350)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_290),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_335),
.B(n_222),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_311),
.A2(n_287),
.B1(n_285),
.B2(n_304),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_337),
.A2(n_351),
.B1(n_358),
.B2(n_321),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_317),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_338),
.B(n_348),
.Y(n_363)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_340),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_341),
.B(n_342),
.C(n_345),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_315),
.B(n_294),
.C(n_288),
.Y(n_342)
);

NOR3xp33_ASAP7_75t_SL g343 ( 
.A(n_336),
.B(n_252),
.C(n_301),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g362 ( 
.A(n_343),
.B(n_346),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_313),
.A2(n_287),
.B(n_296),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_344),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_315),
.B(n_309),
.C(n_300),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_319),
.B(n_320),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_333),
.B(n_297),
.C(n_279),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_347),
.B(n_345),
.C(n_342),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_329),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_324),
.B(n_192),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_352),
.B(n_322),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_353),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_SL g356 ( 
.A(n_333),
.B(n_263),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_SL g376 ( 
.A(n_356),
.B(n_361),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_310),
.A2(n_263),
.B1(n_261),
.B2(n_251),
.Y(n_358)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_359),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_350),
.B(n_318),
.Y(n_364)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_364),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_365),
.A2(n_353),
.B1(n_354),
.B2(n_355),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_337),
.A2(n_327),
.B1(n_326),
.B2(n_329),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_366),
.A2(n_367),
.B1(n_379),
.B2(n_381),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_354),
.A2(n_327),
.B1(n_326),
.B2(n_331),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_344),
.A2(n_334),
.B(n_322),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_369),
.A2(n_204),
.B(n_198),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_350),
.B(n_316),
.Y(n_373)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_373),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_374),
.B(n_383),
.Y(n_395)
);

INVx2_ASAP7_75t_SL g377 ( 
.A(n_360),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_377),
.Y(n_388)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_360),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_378),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_341),
.B(n_316),
.C(n_335),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_380),
.B(n_382),
.Y(n_385)
);

CKINVDCx14_ASAP7_75t_R g381 ( 
.A(n_357),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_358),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_SL g383 ( 
.A(n_356),
.B(n_328),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_384),
.A2(n_392),
.B1(n_400),
.B2(n_10),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_380),
.B(n_361),
.C(n_339),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_386),
.B(n_393),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_370),
.A2(n_355),
.B1(n_338),
.B2(n_349),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_390),
.A2(n_367),
.B1(n_372),
.B2(n_363),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_365),
.A2(n_347),
.B1(n_343),
.B2(n_340),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_371),
.B(n_348),
.C(n_359),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_362),
.A2(n_328),
.B1(n_189),
.B2(n_198),
.Y(n_394)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_394),
.Y(n_403)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_396),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g398 ( 
.A(n_371),
.B(n_189),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_398),
.B(n_401),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_366),
.A2(n_182),
.B1(n_139),
.B2(n_175),
.Y(n_399)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_399),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_375),
.A2(n_185),
.B1(n_95),
.B2(n_100),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_374),
.B(n_101),
.C(n_0),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_375),
.A2(n_10),
.B(n_1),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_402),
.B(n_377),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_393),
.B(n_369),
.C(n_376),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_404),
.B(n_408),
.Y(n_424)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_406),
.Y(n_429)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_407),
.Y(n_432)
);

OAI321xp33_ASAP7_75t_L g408 ( 
.A1(n_391),
.A2(n_363),
.A3(n_364),
.B1(n_373),
.B2(n_368),
.C(n_377),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_388),
.B(n_383),
.Y(n_409)
);

OR2x2_ASAP7_75t_L g419 ( 
.A(n_409),
.B(n_415),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_386),
.B(n_376),
.C(n_0),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_411),
.B(n_413),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_385),
.B(n_10),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_414),
.B(n_416),
.Y(n_431)
);

AOI22xp33_ASAP7_75t_SL g415 ( 
.A1(n_387),
.A2(n_384),
.B1(n_397),
.B2(n_400),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_390),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_395),
.B(n_0),
.C(n_1),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_418),
.B(n_411),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_405),
.A2(n_389),
.B1(n_387),
.B2(n_392),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_420),
.B(n_430),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_404),
.B(n_401),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_421),
.B(n_10),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_412),
.A2(n_395),
.B1(n_396),
.B2(n_402),
.Y(n_422)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_422),
.Y(n_433)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_423),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_410),
.A2(n_409),
.B(n_413),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_425),
.A2(n_406),
.B(n_5),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_412),
.A2(n_2),
.B(n_4),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_426),
.A2(n_11),
.B(n_12),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_417),
.B(n_2),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_427),
.B(n_6),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_403),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_424),
.B(n_418),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_435),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_436),
.A2(n_423),
.B(n_428),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g437 ( 
.A1(n_432),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_437),
.B(n_439),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_431),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_440),
.B(n_426),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_441),
.B(n_443),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_429),
.B(n_11),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_442),
.A2(n_422),
.B(n_419),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_445),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_447),
.A2(n_448),
.B(n_13),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_438),
.A2(n_419),
.B(n_14),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_450),
.A2(n_442),
.B(n_434),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_SL g455 ( 
.A1(n_451),
.A2(n_452),
.B(n_454),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_446),
.A2(n_433),
.B(n_434),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_453),
.B(n_444),
.C(n_449),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_456),
.A2(n_13),
.B(n_14),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_457),
.A2(n_455),
.B(n_13),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_458),
.A2(n_15),
.B(n_454),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_459),
.A2(n_15),
.B(n_443),
.Y(n_460)
);


endmodule