module fake_jpeg_9129_n_285 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_285);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_285;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_5),
.B(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_4),
.B(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVxp33_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_9),
.B(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_38),
.Y(n_47)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_24),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_41),
.B(n_16),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_21),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_27),
.Y(n_49)
);

BUFx2_ASAP7_75t_R g43 ( 
.A(n_42),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_43),
.B(n_46),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_44),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_45),
.B(n_36),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_41),
.B(n_33),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_36),
.A2(n_23),
.B1(n_31),
.B2(n_25),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_52),
.A2(n_26),
.B1(n_22),
.B2(n_19),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_29),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_57),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

BUFx4f_ASAP7_75t_SL g56 ( 
.A(n_42),
.Y(n_56)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_32),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_35),
.A2(n_23),
.B1(n_31),
.B2(n_25),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_60),
.A2(n_33),
.B1(n_18),
.B2(n_26),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_53),
.B(n_37),
.C(n_38),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_63),
.B(n_92),
.C(n_55),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_35),
.B1(n_36),
.B2(n_54),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_64),
.A2(n_76),
.B1(n_51),
.B2(n_59),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

INVxp67_ASAP7_75t_SL g112 ( 
.A(n_66),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_47),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_69),
.Y(n_93)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_47),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_53),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_75),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_31),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_72),
.B(n_80),
.Y(n_105)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_43),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_54),
.A2(n_48),
.B1(n_58),
.B2(n_57),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_77),
.B(n_81),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_43),
.A2(n_33),
.B1(n_18),
.B2(n_16),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_78),
.A2(n_84),
.B1(n_91),
.B2(n_37),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_44),
.B(n_25),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_45),
.B(n_34),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_86),
.B(n_89),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_87),
.Y(n_96)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_51),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_52),
.B(n_34),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_54),
.A2(n_37),
.B1(n_38),
.B2(n_23),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_90),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_48),
.A2(n_22),
.B1(n_19),
.B2(n_42),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_49),
.B(n_40),
.Y(n_92)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_110),
.Y(n_121)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_86),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_98),
.B(n_103),
.Y(n_134)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_101),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_102),
.A2(n_65),
.B1(n_75),
.B2(n_74),
.Y(n_125)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_70),
.Y(n_103)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_71),
.A2(n_51),
.B1(n_56),
.B2(n_34),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_104),
.A2(n_107),
.B1(n_85),
.B2(n_55),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g106 ( 
.A(n_68),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_106),
.B(n_111),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_108),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_109),
.B(n_40),
.Y(n_139)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_24),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_69),
.B(n_59),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_89),
.Y(n_120)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_114),
.B(n_93),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_92),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_117),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_87),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_82),
.Y(n_118)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_118),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_74),
.A2(n_17),
.B1(n_20),
.B2(n_29),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_119),
.A2(n_62),
.B1(n_82),
.B2(n_85),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_120),
.A2(n_127),
.B(n_132),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_122),
.B(n_135),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_105),
.B(n_63),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_138),
.Y(n_156)
);

OAI21xp33_ASAP7_75t_L g124 ( 
.A1(n_116),
.A2(n_72),
.B(n_65),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_124),
.A2(n_125),
.B(n_143),
.Y(n_149)
);

AOI22x1_ASAP7_75t_SL g127 ( 
.A1(n_102),
.A2(n_79),
.B1(n_109),
.B2(n_113),
.Y(n_127)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_133),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_131),
.A2(n_145),
.B1(n_122),
.B2(n_100),
.Y(n_169)
);

AOI21xp33_ASAP7_75t_L g132 ( 
.A1(n_105),
.A2(n_79),
.B(n_83),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_101),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g136 ( 
.A(n_118),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_146),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_88),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_137),
.B(n_141),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_79),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_139),
.B(n_107),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_116),
.A2(n_81),
.B(n_77),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_140),
.A2(n_40),
.B(n_39),
.Y(n_175)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_104),
.Y(n_141)
);

OAI21xp33_ASAP7_75t_L g143 ( 
.A1(n_115),
.A2(n_14),
.B(n_12),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_144),
.A2(n_128),
.B1(n_140),
.B2(n_119),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_97),
.A2(n_61),
.B1(n_40),
.B2(n_39),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_104),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_110),
.A2(n_13),
.B1(n_15),
.B2(n_14),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_148),
.A2(n_93),
.B(n_28),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_121),
.Y(n_150)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_150),
.Y(n_184)
);

O2A1O1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_141),
.A2(n_146),
.B(n_120),
.C(n_129),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_151),
.A2(n_160),
.B(n_162),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_152),
.A2(n_164),
.B1(n_174),
.B2(n_131),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_128),
.A2(n_117),
.B1(n_96),
.B2(n_98),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_153),
.A2(n_169),
.B1(n_133),
.B2(n_126),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_155),
.B(n_157),
.C(n_130),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_114),
.C(n_94),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g159 ( 
.A(n_136),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_159),
.Y(n_181)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_134),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_172),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_136),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_127),
.A2(n_94),
.B1(n_108),
.B2(n_95),
.Y(n_164)
);

INVx13_ASAP7_75t_L g166 ( 
.A(n_136),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_166),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_134),
.B(n_113),
.Y(n_167)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_167),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_125),
.A2(n_111),
.B(n_95),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_168),
.A2(n_175),
.B(n_138),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_106),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_171),
.Y(n_195)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_135),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_104),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_177),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_144),
.A2(n_104),
.B1(n_100),
.B2(n_61),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_142),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_176),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_147),
.B(n_29),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_145),
.Y(n_178)
);

NOR3xp33_ASAP7_75t_L g190 ( 
.A(n_178),
.B(n_112),
.C(n_61),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_139),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_186),
.C(n_187),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_182),
.A2(n_170),
.B1(n_178),
.B2(n_172),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_183),
.A2(n_167),
.B(n_163),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_139),
.C(n_126),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_188),
.A2(n_191),
.B1(n_199),
.B2(n_200),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_157),
.C(n_165),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_189),
.B(n_192),
.C(n_149),
.Y(n_206)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_190),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_164),
.A2(n_66),
.B1(n_20),
.B2(n_17),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_155),
.B(n_39),
.C(n_28),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_158),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_193),
.B(n_177),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_159),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_194),
.B(n_201),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_151),
.A2(n_20),
.B1(n_17),
.B2(n_39),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_174),
.A2(n_20),
.B1(n_27),
.B2(n_2),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_159),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_185),
.B(n_161),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_203),
.B(n_210),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_205),
.A2(n_212),
.B1(n_219),
.B2(n_199),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_206),
.B(n_211),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_168),
.C(n_175),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_213),
.Y(n_229)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_185),
.Y(n_210)
);

A2O1A1O1Ixp25_ASAP7_75t_L g211 ( 
.A1(n_183),
.A2(n_149),
.B(n_170),
.C(n_154),
.D(n_173),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_182),
.A2(n_152),
.B1(n_150),
.B2(n_154),
.Y(n_212)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_214),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_181),
.B(n_201),
.Y(n_215)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_215),
.Y(n_234)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_202),
.Y(n_216)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_216),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_196),
.B(n_163),
.Y(n_217)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_217),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_202),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_218),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_196),
.A2(n_169),
.B1(n_153),
.B2(n_162),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_181),
.B(n_159),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_220),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_188),
.A2(n_166),
.B1(n_160),
.B2(n_27),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_222),
.A2(n_193),
.B1(n_184),
.B2(n_195),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_179),
.B(n_166),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_223),
.B(n_204),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_225),
.A2(n_227),
.B1(n_205),
.B2(n_213),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_207),
.A2(n_180),
.B1(n_191),
.B2(n_184),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_228),
.A2(n_231),
.B1(n_207),
.B2(n_222),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_230),
.B(n_238),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_212),
.A2(n_200),
.B1(n_189),
.B2(n_180),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_219),
.A2(n_197),
.B1(n_194),
.B2(n_192),
.Y(n_233)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_233),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_204),
.B(n_208),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_229),
.B(n_187),
.C(n_206),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_250),
.C(n_252),
.Y(n_260)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_242),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_236),
.B(n_209),
.Y(n_243)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_243),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_244),
.A2(n_230),
.B1(n_1),
.B2(n_2),
.Y(n_258)
);

AOI21xp33_ASAP7_75t_SL g245 ( 
.A1(n_232),
.A2(n_229),
.B(n_223),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_245),
.A2(n_246),
.B(n_237),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_234),
.A2(n_210),
.B(n_221),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_214),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_249),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_216),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_211),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_225),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_252),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_198),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_248),
.A2(n_228),
.B1(n_231),
.B2(n_235),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_253),
.B(n_258),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_254),
.A2(n_255),
.B(n_261),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_244),
.A2(n_227),
.B(n_224),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_250),
.A2(n_8),
.B(n_14),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_8),
.C(n_13),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_8),
.C(n_13),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_263),
.B(n_240),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_259),
.B(n_241),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_264),
.B(n_265),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_266),
.B(n_267),
.C(n_15),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_7),
.C(n_11),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_257),
.B(n_7),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_5),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_256),
.A2(n_7),
.B(n_11),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_271),
.A2(n_262),
.B1(n_258),
.B2(n_9),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_265),
.B(n_260),
.C(n_253),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_272),
.A2(n_275),
.B(n_276),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_274),
.A2(n_268),
.B(n_269),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_278),
.B(n_279),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_272),
.A2(n_10),
.B(n_6),
.Y(n_279)
);

NOR2xp67_ASAP7_75t_SL g281 ( 
.A(n_277),
.B(n_273),
.Y(n_281)
);

OAI321xp33_ASAP7_75t_L g282 ( 
.A1(n_281),
.A2(n_280),
.A3(n_6),
.B1(n_3),
.B2(n_1),
.C(n_0),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_282),
.B(n_1),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_6),
.C(n_3),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_284),
.Y(n_285)
);


endmodule