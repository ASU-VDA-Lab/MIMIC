module real_jpeg_19600_n_17 (n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_337, n_11, n_14, n_336, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_337;
input n_11;
input n_14;
input n_336;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_0),
.A2(n_46),
.B1(n_48),
.B2(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_0),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_0),
.A2(n_69),
.B1(n_70),
.B2(n_116),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_0),
.A2(n_35),
.B1(n_36),
.B2(n_116),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_0),
.A2(n_26),
.B1(n_27),
.B2(n_116),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_1),
.A2(n_69),
.B1(n_70),
.B2(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_1),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_1),
.A2(n_46),
.B1(n_48),
.B2(n_121),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_1),
.A2(n_35),
.B1(n_36),
.B2(n_121),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_1),
.A2(n_26),
.B1(n_27),
.B2(n_121),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_2),
.A2(n_26),
.B1(n_27),
.B2(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_2),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_2),
.A2(n_69),
.B1(n_70),
.B2(n_83),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_2),
.A2(n_46),
.B1(n_48),
.B2(n_83),
.Y(n_214)
);

OAI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_2),
.A2(n_35),
.B1(n_36),
.B2(n_83),
.Y(n_257)
);

A2O1A1O1Ixp25_ASAP7_75t_L g100 ( 
.A1(n_3),
.A2(n_48),
.B(n_65),
.C(n_101),
.D(n_102),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_3),
.B(n_48),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_3),
.B(n_45),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_3),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_3),
.A2(n_122),
.B(n_124),
.Y(n_144)
);

A2O1A1O1Ixp25_ASAP7_75t_L g157 ( 
.A1(n_3),
.A2(n_35),
.B(n_42),
.C(n_158),
.D(n_159),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_3),
.B(n_35),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_3),
.B(n_39),
.Y(n_184)
);

AOI21xp33_ASAP7_75t_L g202 ( 
.A1(n_3),
.A2(n_36),
.B(n_203),
.Y(n_202)
);

OAI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_3),
.A2(n_26),
.B1(n_27),
.B2(n_139),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_4),
.A2(n_35),
.B1(n_36),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_4),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_4),
.A2(n_46),
.B1(n_48),
.B2(n_51),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_4),
.A2(n_51),
.B1(n_69),
.B2(n_70),
.Y(n_249)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_6),
.A2(n_26),
.B1(n_27),
.B2(n_29),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_6),
.A2(n_29),
.B1(n_35),
.B2(n_36),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_6),
.A2(n_29),
.B1(n_69),
.B2(n_70),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_6),
.A2(n_29),
.B1(n_46),
.B2(n_48),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_7),
.A2(n_26),
.B1(n_27),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_7),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_7),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_7),
.A2(n_38),
.B1(n_69),
.B2(n_70),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_7),
.A2(n_38),
.B1(n_46),
.B2(n_48),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_8),
.A2(n_26),
.B1(n_27),
.B2(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_8),
.A2(n_62),
.B1(n_69),
.B2(n_70),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_8),
.A2(n_46),
.B1(n_48),
.B2(n_62),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_8),
.A2(n_35),
.B1(n_36),
.B2(n_62),
.Y(n_276)
);

BUFx10_ASAP7_75t_L g69 ( 
.A(n_9),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_10),
.A2(n_46),
.B1(n_48),
.B2(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_10),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_10),
.A2(n_69),
.B1(n_70),
.B2(n_104),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_10),
.A2(n_35),
.B1(n_36),
.B2(n_104),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_10),
.A2(n_26),
.B1(n_27),
.B2(n_104),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_11),
.B(n_70),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_11),
.B(n_125),
.Y(n_124)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_11),
.Y(n_133)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_11),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_11),
.A2(n_123),
.B1(n_169),
.B2(n_186),
.Y(n_185)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_14),
.A2(n_32),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_15),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_91),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_89),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_75),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_20),
.B(n_75),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_52),
.B1(n_53),
.B2(n_74),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_21),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_40),
.B2(n_41),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B1(n_37),
.B2(n_39),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_25),
.A2(n_31),
.B1(n_34),
.B2(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

A2O1A1Ixp33_ASAP7_75t_L g31 ( 
.A1(n_27),
.A2(n_32),
.B(n_33),
.C(n_34),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_32),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g201 ( 
.A1(n_27),
.A2(n_32),
.B(n_139),
.C(n_202),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_30),
.A2(n_220),
.B(n_221),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_30),
.B(n_223),
.Y(n_232)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_31),
.A2(n_34),
.B1(n_61),
.B2(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_31),
.A2(n_34),
.B1(n_231),
.B2(n_260),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_31),
.A2(n_222),
.B(n_260),
.Y(n_278)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_32),
.Y(n_203)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

OAI21xp33_ASAP7_75t_L g230 ( 
.A1(n_34),
.A2(n_231),
.B(n_232),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_34),
.A2(n_82),
.B(n_232),
.Y(n_302)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

O2A1O1Ixp33_ASAP7_75t_SL g42 ( 
.A1(n_36),
.A2(n_43),
.B(n_44),
.C(n_45),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_43),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_39),
.B(n_223),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_45),
.B(n_49),
.Y(n_41)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_42),
.B(n_182),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_42),
.A2(n_45),
.B1(n_257),
.B2(n_276),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_42),
.A2(n_45),
.B1(n_88),
.B2(n_276),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_43),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_45)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_43),
.B(n_48),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_44),
.A2(n_46),
.B1(n_165),
.B2(n_166),
.Y(n_164)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

O2A1O1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_46),
.A2(n_66),
.B(n_67),
.C(n_68),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_66),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_50),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_55)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_59),
.C(n_63),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_54),
.A2(n_55),
.B1(n_63),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_56),
.A2(n_57),
.B1(n_58),
.B2(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_56),
.A2(n_58),
.B1(n_180),
.B2(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_56),
.A2(n_217),
.B(n_235),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_58),
.B(n_160),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_58),
.A2(n_180),
.B(n_181),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_58),
.A2(n_181),
.B(n_256),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_59),
.A2(n_60),
.B1(n_78),
.B2(n_79),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_63),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_63),
.A2(n_80),
.B1(n_85),
.B2(n_86),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_64),
.A2(n_72),
.B(n_73),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_64),
.A2(n_72),
.B1(n_115),
.B2(n_156),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_64),
.A2(n_156),
.B(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_64),
.A2(n_72),
.B1(n_214),
.B2(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_64),
.A2(n_72),
.B1(n_242),
.B2(n_251),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_64),
.A2(n_72),
.B1(n_251),
.B2(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_65),
.B(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_65),
.A2(n_68),
.B1(n_292),
.B2(n_293),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_66),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_68)
);

CKINVDCx9p33_ASAP7_75t_R g71 ( 
.A(n_66),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_66),
.B(n_70),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_67),
.A2(n_69),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_68),
.Y(n_72)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_70),
.B(n_146),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_72),
.A2(n_115),
.B(n_117),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_72),
.B(n_139),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_72),
.A2(n_117),
.B(n_214),
.Y(n_213)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_73),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_81),
.C(n_84),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_76),
.A2(n_77),
.B1(n_81),
.B2(n_321),
.Y(n_327)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_81),
.C(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_81),
.A2(n_321),
.B1(n_322),
.B2(n_323),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_81),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_84),
.B(n_327),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

OAI321xp33_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_318),
.A3(n_328),
.B1(n_333),
.B2(n_334),
.C(n_336),
.Y(n_91)
);

AOI321xp33_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_268),
.A3(n_306),
.B1(n_312),
.B2(n_317),
.C(n_337),
.Y(n_92)
);

NOR3xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_225),
.C(n_264),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_195),
.B(n_224),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_174),
.B(n_194),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_150),
.B(n_173),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_126),
.B(n_149),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_109),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_99),
.B(n_109),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_105),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_100),
.A2(n_105),
.B1(n_106),
.B2(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_100),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_101),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_102),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_119),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_111),
.B(n_114),
.C(n_119),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_122),
.B(n_124),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_120),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_122),
.A2(n_133),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_122),
.A2(n_133),
.B1(n_207),
.B2(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_122),
.A2(n_133),
.B1(n_240),
.B2(n_249),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_122),
.A2(n_141),
.B(n_249),
.Y(n_281)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_123),
.A2(n_129),
.B1(n_131),
.B2(n_132),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_123),
.B(n_125),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_136),
.B(n_148),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_134),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_128),
.B(n_134),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_130),
.A2(n_141),
.B(n_142),
.Y(n_140)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_143),
.B(n_147),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_138),
.B(n_140),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_141),
.Y(n_146)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_141),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_142),
.A2(n_168),
.B(n_170),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_145),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_151),
.B(n_152),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_163),
.B2(n_172),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_157),
.B1(n_161),
.B2(n_162),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_155),
.Y(n_162)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_157),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_157),
.B(n_162),
.C(n_172),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_158),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_159),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_160),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_163),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_167),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_167),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_175),
.B(n_176),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_188),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_177),
.B(n_190),
.C(n_192),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_183),
.B2(n_187),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_178),
.B(n_184),
.C(n_185),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_183),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_186),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_192),
.B2(n_193),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_189),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_190),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_197),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_196),
.B(n_197),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_211),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_208),
.B1(n_209),
.B2(n_210),
.Y(n_198)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_199),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_199),
.B(n_210),
.C(n_211),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_201),
.B1(n_204),
.B2(n_205),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_200),
.B(n_205),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_208),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_219),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_215),
.B1(n_216),
.B2(n_218),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_213),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_218),
.C(n_219),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

AOI21xp33_ASAP7_75t_L g313 ( 
.A1(n_226),
.A2(n_314),
.B(n_315),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_244),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_227),
.B(n_244),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_238),
.C(n_243),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_228),
.B(n_267),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_237),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_233),
.B1(n_234),
.B2(n_236),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_230),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_233),
.B(n_236),
.C(n_237),
.Y(n_262)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_238),
.B(n_243),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_239),
.B(n_241),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_262),
.B2(n_263),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_252),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_247),
.B(n_252),
.C(n_263),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_250),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_250),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_253),
.B(n_258),
.C(n_261),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_255),
.A2(n_258),
.B1(n_259),
.B2(n_261),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_255),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_262),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_265),
.B(n_266),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_286),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_269),
.B(n_286),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_279),
.C(n_285),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_270),
.A2(n_271),
.B1(n_279),
.B2(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_272),
.B(n_275),
.C(n_277),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_277),
.B2(n_278),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_275),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_279),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_282),
.B2(n_284),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_280),
.A2(n_281),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_280),
.A2(n_298),
.B(n_302),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_282),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_282),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_283),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_285),
.B(n_310),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_304),
.B2(n_305),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_296),
.B2(n_297),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_289),
.B(n_297),
.C(n_305),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_290),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_294),
.B(n_295),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_291),
.B(n_294),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_295),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_295),
.A2(n_320),
.B1(n_324),
.B2(n_332),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_297),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_299),
.B1(n_300),
.B2(n_303),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_300),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_302),
.Y(n_301)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_304),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_307),
.A2(n_313),
.B(n_316),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_308),
.B(n_309),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_326),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_319),
.B(n_326),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_324),
.C(n_325),
.Y(n_319)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_320),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_323),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_331),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_329),
.B(n_330),
.Y(n_333)
);


endmodule