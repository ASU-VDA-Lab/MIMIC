module fake_jpeg_16412_n_93 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_93);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_93;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_22;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

INVx13_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_SL g16 ( 
.A(n_1),
.B(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g23 ( 
.A(n_22),
.Y(n_23)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_24),
.B(n_28),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_17),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_29),
.Y(n_35)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_16),
.B(n_0),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_30),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_19),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_16),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_13),
.Y(n_33)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_33),
.B(n_48),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_26),
.A2(n_20),
.B1(n_18),
.B2(n_15),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_37),
.A2(n_49),
.B1(n_15),
.B2(n_14),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_22),
.C(n_17),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_42),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_27),
.B(n_22),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_SL g58 ( 
.A(n_41),
.B(n_47),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_20),
.Y(n_42)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_24),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_46),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_28),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_20),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_32),
.B(n_21),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_29),
.A2(n_18),
.B1(n_15),
.B2(n_1),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_25),
.A2(n_14),
.B1(n_13),
.B2(n_19),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_50),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_59),
.B1(n_36),
.B2(n_37),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_1),
.B(n_21),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_53),
.B(n_55),
.C(n_61),
.Y(n_67)
);

NAND2x1_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_21),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_2),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_33),
.Y(n_64)
);

AO22x2_ASAP7_75t_L g57 ( 
.A1(n_48),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_57),
.A2(n_38),
.B1(n_36),
.B2(n_35),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_47),
.B1(n_49),
.B2(n_38),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_57),
.B1(n_54),
.B2(n_58),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_6),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_64),
.B(n_66),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_40),
.Y(n_65)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_63),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_72),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_69),
.A2(n_70),
.B1(n_71),
.B2(n_57),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_55),
.A2(n_43),
.B1(n_9),
.B2(n_11),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_62),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_58),
.C(n_61),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_78),
.C(n_76),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_80),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_SL g76 ( 
.A(n_71),
.B(n_57),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_76),
.A2(n_81),
.B(n_78),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_53),
.C(n_62),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_72),
.A2(n_68),
.B(n_67),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_82),
.B(n_83),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_67),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_85),
.Y(n_90)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_86),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_86),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_89),
.B(n_74),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_91),
.A2(n_92),
.B1(n_88),
.B2(n_90),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);


endmodule