module real_aes_11154_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_400;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_417;
wire n_323;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_552;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1250;
wire n_1284;
wire n_1095;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_789;
wire n_738;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_837;
wire n_829;
wire n_1030;
wire n_375;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_264;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_665;
wire n_991;
wire n_667;
wire n_580;
wire n_1004;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_678;
wire n_415;
wire n_564;
wire n_638;
wire n_510;
wire n_550;
wire n_966;
wire n_333;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1182;
wire n_872;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_354;
wire n_265;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_639;
wire n_1186;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1223;
wire n_405;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_769;
wire n_434;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_714;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1033;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_546;
wire n_1010;
wire n_1015;
wire n_863;
wire n_1226;
wire n_525;
wire n_644;
wire n_1150;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1156;
wire n_988;
wire n_921;
wire n_1176;
wire n_640;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_857;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_886;
wire n_767;
wire n_889;
wire n_379;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_269;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_698;
wire n_371;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_272;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_703;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_0), .A2(n_221), .B1(n_594), .B2(n_614), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_0), .A2(n_221), .B1(n_394), .B2(n_568), .Y(n_733) );
OAI22xp5_ASAP7_75t_L g939 ( .A1(n_1), .A2(n_19), .B1(n_543), .B2(n_893), .Y(n_939) );
OAI22xp5_ASAP7_75t_L g945 ( .A1(n_1), .A2(n_234), .B1(n_335), .B2(n_551), .Y(n_945) );
AO221x1_ASAP7_75t_L g1054 ( .A1(n_2), .A2(n_150), .B1(n_1007), .B2(n_1055), .C(n_1057), .Y(n_1054) );
INVx1_ASAP7_75t_L g452 ( .A(n_3), .Y(n_452) );
INVxp67_ASAP7_75t_SL g769 ( .A(n_4), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g786 ( .A1(n_4), .A2(n_22), .B1(n_575), .B2(n_787), .Y(n_786) );
OAI22xp5_ASAP7_75t_L g546 ( .A1(n_5), .A2(n_171), .B1(n_547), .B2(n_551), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_5), .A2(n_171), .B1(n_505), .B2(n_587), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g1297 ( .A1(n_6), .A2(n_108), .B1(n_575), .B2(n_576), .Y(n_1297) );
AOI22xp33_ASAP7_75t_L g1305 ( .A1(n_6), .A2(n_108), .B1(n_413), .B2(n_505), .Y(n_1305) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_7), .Y(n_262) );
INVx1_ASAP7_75t_L g404 ( .A(n_7), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_8), .A2(n_93), .B1(n_416), .B2(n_418), .Y(n_987) );
AOI22xp33_ASAP7_75t_L g1000 ( .A1(n_8), .A2(n_93), .B1(n_378), .B2(n_1001), .Y(n_1000) );
AOI22xp33_ASAP7_75t_SL g825 ( .A1(n_9), .A2(n_205), .B1(n_483), .B2(n_602), .Y(n_825) );
AOI22xp33_ASAP7_75t_SL g833 ( .A1(n_9), .A2(n_205), .B1(n_588), .B2(n_730), .Y(n_833) );
AOI22xp5_ASAP7_75t_L g1036 ( .A1(n_10), .A2(n_115), .B1(n_1007), .B2(n_1031), .Y(n_1036) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_11), .A2(n_36), .B1(n_580), .B2(n_689), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_11), .A2(n_36), .B1(n_501), .B2(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g658 ( .A(n_12), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_13), .A2(n_202), .B1(n_568), .B2(n_571), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_13), .A2(n_202), .B1(n_583), .B2(n_584), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_14), .A2(n_177), .B1(n_483), .B2(n_602), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_14), .A2(n_177), .B1(n_588), .B2(n_794), .Y(n_793) );
AO22x2_ASAP7_75t_L g438 ( .A1(n_15), .A2(n_439), .B1(n_519), .B2(n_520), .Y(n_438) );
INVx1_ASAP7_75t_L g519 ( .A(n_15), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g377 ( .A1(n_16), .A2(n_129), .B1(n_378), .B2(n_382), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_16), .A2(n_129), .B1(n_416), .B2(n_418), .Y(n_415) );
CKINVDCx5p33_ASAP7_75t_R g890 ( .A(n_17), .Y(n_890) );
INVx1_ASAP7_75t_L g760 ( .A(n_18), .Y(n_760) );
INVx1_ASAP7_75t_L g932 ( .A(n_19), .Y(n_932) );
AOI22xp33_ASAP7_75t_SL g484 ( .A1(n_20), .A2(n_243), .B1(n_485), .B2(n_486), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_20), .A2(n_243), .B1(n_499), .B2(n_501), .Y(n_498) );
AO221x2_ASAP7_75t_L g1175 ( .A1(n_21), .A2(n_168), .B1(n_1055), .B2(n_1176), .C(n_1178), .Y(n_1175) );
AOI222xp33_ASAP7_75t_L g1214 ( .A1(n_21), .A2(n_1215), .B1(n_1270), .B2(n_1272), .C1(n_1310), .C2(n_1312), .Y(n_1214) );
AO22x2_ASAP7_75t_L g1215 ( .A1(n_21), .A2(n_1216), .B1(n_1217), .B2(n_1269), .Y(n_1215) );
INVxp67_ASAP7_75t_SL g1216 ( .A(n_21), .Y(n_1216) );
INVx1_ASAP7_75t_L g768 ( .A(n_22), .Y(n_768) );
INVx1_ASAP7_75t_L g804 ( .A(n_23), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_23), .A2(n_125), .B1(n_605), .B2(n_774), .Y(n_830) );
XNOR2xp5_ASAP7_75t_L g899 ( .A(n_24), .B(n_900), .Y(n_899) );
INVxp67_ASAP7_75t_SL g358 ( .A(n_25), .Y(n_358) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_25), .A2(n_198), .B1(n_428), .B2(n_430), .Y(n_427) );
INVx2_ASAP7_75t_L g284 ( .A(n_26), .Y(n_284) );
INVx1_ASAP7_75t_L g755 ( .A(n_27), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_28), .A2(n_215), .B1(n_602), .B2(n_608), .Y(n_607) );
INVxp67_ASAP7_75t_SL g642 ( .A(n_28), .Y(n_642) );
INVx1_ASAP7_75t_L g970 ( .A(n_29), .Y(n_970) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_29), .A2(n_113), .B1(n_411), .B2(n_986), .Y(n_985) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_30), .A2(n_184), .B1(n_451), .B2(n_623), .Y(n_622) );
OAI211xp5_ASAP7_75t_SL g626 ( .A1(n_30), .A2(n_474), .B(n_627), .C(n_630), .Y(n_626) );
BUFx2_ASAP7_75t_L g329 ( .A(n_31), .Y(n_329) );
BUFx2_ASAP7_75t_L g370 ( .A(n_31), .Y(n_370) );
INVx1_ASAP7_75t_L g402 ( .A(n_31), .Y(n_402) );
INVx1_ASAP7_75t_L g963 ( .A(n_32), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g990 ( .A1(n_32), .A2(n_99), .B1(n_480), .B2(n_991), .Y(n_990) );
AOI22xp33_ASAP7_75t_SL g729 ( .A1(n_33), .A2(n_106), .B1(n_730), .B2(n_731), .Y(n_729) );
INVxp67_ASAP7_75t_L g741 ( .A(n_33), .Y(n_741) );
INVx1_ASAP7_75t_L g978 ( .A(n_34), .Y(n_978) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_34), .A2(n_45), .B1(n_416), .B2(n_984), .Y(n_983) );
INVx1_ASAP7_75t_L g661 ( .A(n_35), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_35), .A2(n_97), .B1(n_571), .B2(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g665 ( .A(n_37), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g670 ( .A1(n_37), .A2(n_143), .B1(n_354), .B2(n_671), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_38), .A2(n_176), .B1(n_571), .B2(n_605), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_38), .A2(n_176), .B1(n_613), .B2(n_614), .Y(n_612) );
INVxp67_ASAP7_75t_SL g293 ( .A(n_39), .Y(n_293) );
OAI22xp5_ASAP7_75t_L g350 ( .A1(n_39), .A2(n_121), .B1(n_351), .B2(n_354), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_40), .A2(n_51), .B1(n_575), .B2(n_684), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_40), .A2(n_51), .B1(n_621), .B2(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g943 ( .A(n_41), .Y(n_943) );
AO22x2_ASAP7_75t_L g952 ( .A1(n_42), .A2(n_953), .B1(n_954), .B2(n_1003), .Y(n_952) );
INVx1_ASAP7_75t_L g1003 ( .A(n_42), .Y(n_1003) );
AOI22xp33_ASAP7_75t_L g1252 ( .A1(n_43), .A2(n_59), .B1(n_1250), .B2(n_1253), .Y(n_1252) );
INVxp67_ASAP7_75t_SL g1261 ( .A(n_43), .Y(n_1261) );
INVxp33_ASAP7_75t_L g1291 ( .A(n_44), .Y(n_1291) );
AOI22xp33_ASAP7_75t_L g1300 ( .A1(n_44), .A2(n_157), .B1(n_564), .B2(n_686), .Y(n_1300) );
INVx1_ASAP7_75t_L g972 ( .A(n_45), .Y(n_972) );
INVx1_ASAP7_75t_L g808 ( .A(n_46), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_46), .A2(n_230), .B1(n_483), .B2(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g759 ( .A(n_47), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g789 ( .A1(n_47), .A2(n_194), .B1(n_681), .B2(n_774), .Y(n_789) );
INVx1_ASAP7_75t_L g1058 ( .A(n_48), .Y(n_1058) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_49), .A2(n_241), .B1(n_505), .B2(n_588), .Y(n_883) );
OAI22xp5_ASAP7_75t_L g895 ( .A1(n_49), .A2(n_178), .B1(n_335), .B2(n_551), .Y(n_895) );
INVx1_ASAP7_75t_L g445 ( .A(n_50), .Y(n_445) );
XNOR2xp5_ASAP7_75t_L g523 ( .A(n_52), .B(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g962 ( .A(n_53), .Y(n_962) );
AOI22xp33_ASAP7_75t_SL g992 ( .A1(n_53), .A2(n_68), .B1(n_993), .B2(n_995), .Y(n_992) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_54), .A2(n_222), .B1(n_451), .B2(n_613), .Y(n_728) );
INVxp33_ASAP7_75t_L g743 ( .A(n_54), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_55), .A2(n_212), .B1(n_568), .B2(n_571), .Y(n_609) );
INVx1_ASAP7_75t_L g637 ( .A(n_55), .Y(n_637) );
AOI22xp33_ASAP7_75t_SL g1236 ( .A1(n_56), .A2(n_109), .B1(n_394), .B2(n_1237), .Y(n_1236) );
AOI22xp33_ASAP7_75t_L g1249 ( .A1(n_56), .A2(n_109), .B1(n_1250), .B2(n_1251), .Y(n_1249) );
INVxp33_ASAP7_75t_L g1285 ( .A(n_57), .Y(n_1285) );
AOI22xp33_ASAP7_75t_L g1307 ( .A1(n_57), .A2(n_91), .B1(n_501), .B2(n_613), .Y(n_1307) );
INVx1_ASAP7_75t_L g863 ( .A(n_58), .Y(n_863) );
OAI22xp5_ASAP7_75t_L g885 ( .A1(n_58), .A2(n_178), .B1(n_538), .B2(n_543), .Y(n_885) );
INVxp33_ASAP7_75t_L g1268 ( .A(n_59), .Y(n_1268) );
INVx1_ASAP7_75t_L g1059 ( .A(n_60), .Y(n_1059) );
INVx1_ASAP7_75t_L g942 ( .A(n_61), .Y(n_942) );
INVx1_ASAP7_75t_L g533 ( .A(n_62), .Y(n_533) );
INVx1_ASAP7_75t_L g536 ( .A(n_63), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g574 ( .A1(n_63), .A2(n_123), .B1(n_575), .B2(n_576), .Y(n_574) );
INVx1_ASAP7_75t_L g913 ( .A(n_64), .Y(n_913) );
INVxp67_ASAP7_75t_SL g1226 ( .A(n_65), .Y(n_1226) );
AOI22xp33_ASAP7_75t_SL g1241 ( .A1(n_65), .A2(n_107), .B1(n_1237), .B2(n_1242), .Y(n_1241) );
INVx1_ASAP7_75t_L g1282 ( .A(n_66), .Y(n_1282) );
INVxp67_ASAP7_75t_SL g674 ( .A(n_67), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_67), .A2(n_144), .B1(n_411), .B2(n_699), .Y(n_698) );
OAI222xp33_ASAP7_75t_L g957 ( .A1(n_68), .A2(n_154), .B1(n_238), .B2(n_765), .C1(n_766), .C2(n_958), .Y(n_957) );
INVx1_ASAP7_75t_L g822 ( .A(n_69), .Y(n_822) );
AOI22xp33_ASAP7_75t_SL g836 ( .A1(n_69), .A2(n_81), .B1(n_721), .B2(n_730), .Y(n_836) );
INVx1_ASAP7_75t_L g857 ( .A(n_70), .Y(n_857) );
OAI22xp5_ASAP7_75t_L g891 ( .A1(n_70), .A2(n_165), .B1(n_892), .B2(n_893), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_71), .A2(n_147), .B1(n_605), .B2(n_774), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_71), .A2(n_147), .B1(n_594), .B2(n_614), .Y(n_832) );
OAI22xp5_ASAP7_75t_L g812 ( .A1(n_72), .A2(n_102), .B1(n_766), .B2(n_813), .Y(n_812) );
OAI22xp5_ASAP7_75t_L g817 ( .A1(n_72), .A2(n_102), .B1(n_354), .B2(n_559), .Y(n_817) );
INVx1_ASAP7_75t_L g778 ( .A(n_73), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_73), .A2(n_96), .B1(n_721), .B2(n_730), .Y(n_798) );
INVx1_ASAP7_75t_L g918 ( .A(n_74), .Y(n_918) );
OAI211xp5_ASAP7_75t_SL g946 ( .A1(n_74), .A2(n_474), .B(n_553), .C(n_947), .Y(n_946) );
AOI22xp5_ASAP7_75t_L g1020 ( .A1(n_75), .A2(n_117), .B1(n_1021), .B2(n_1027), .Y(n_1020) );
AO221x1_ASAP7_75t_L g1038 ( .A1(n_76), .A2(n_118), .B1(n_1007), .B2(n_1031), .C(n_1039), .Y(n_1038) );
INVx1_ASAP7_75t_L g1181 ( .A(n_77), .Y(n_1181) );
AOI22xp33_ASAP7_75t_L g1255 ( .A1(n_78), .A2(n_112), .B1(n_1256), .B2(n_1257), .Y(n_1255) );
INVxp33_ASAP7_75t_SL g1265 ( .A(n_78), .Y(n_1265) );
INVxp67_ASAP7_75t_SL g446 ( .A(n_79), .Y(n_446) );
AOI22xp33_ASAP7_75t_SL g491 ( .A1(n_79), .A2(n_197), .B1(n_480), .B2(n_492), .Y(n_491) );
INVxp33_ASAP7_75t_SL g656 ( .A(n_80), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_80), .A2(n_162), .B1(n_575), .B2(n_576), .Y(n_679) );
INVx1_ASAP7_75t_L g820 ( .A(n_81), .Y(n_820) );
INVx1_ASAP7_75t_L g712 ( .A(n_82), .Y(n_712) );
OAI22xp5_ASAP7_75t_L g737 ( .A1(n_82), .A2(n_89), .B1(n_671), .B2(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g645 ( .A(n_83), .Y(n_645) );
INVx1_ASAP7_75t_L g327 ( .A(n_84), .Y(n_327) );
INVxp33_ASAP7_75t_SL g460 ( .A(n_85), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_85), .A2(n_188), .B1(n_515), .B2(n_516), .Y(n_514) );
INVx1_ASAP7_75t_L g448 ( .A(n_86), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_86), .A2(n_181), .B1(n_486), .B2(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g632 ( .A(n_87), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_88), .A2(n_191), .B1(n_480), .B2(n_481), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_88), .A2(n_191), .B1(n_503), .B2(n_506), .Y(n_502) );
INVx1_ASAP7_75t_L g713 ( .A(n_89), .Y(n_713) );
AO221x1_ASAP7_75t_L g1044 ( .A1(n_90), .A2(n_159), .B1(n_1007), .B2(n_1031), .C(n_1045), .Y(n_1044) );
INVx1_ASAP7_75t_L g1281 ( .A(n_91), .Y(n_1281) );
INVx1_ASAP7_75t_L g882 ( .A(n_92), .Y(n_882) );
OAI211xp5_ASAP7_75t_SL g896 ( .A1(n_92), .A2(n_474), .B(n_553), .C(n_897), .Y(n_896) );
OAI22xp5_ASAP7_75t_L g764 ( .A1(n_94), .A2(n_186), .B1(n_765), .B2(n_766), .Y(n_764) );
OAI22xp5_ASAP7_75t_L g775 ( .A1(n_94), .A2(n_186), .B1(n_354), .B2(n_671), .Y(n_775) );
INVx1_ASAP7_75t_L g907 ( .A(n_95), .Y(n_907) );
INVxp67_ASAP7_75t_L g780 ( .A(n_96), .Y(n_780) );
INVxp33_ASAP7_75t_SL g655 ( .A(n_97), .Y(n_655) );
INVxp67_ASAP7_75t_SL g309 ( .A(n_98), .Y(n_309) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_98), .A2(n_236), .B1(n_396), .B2(n_398), .Y(n_395) );
INVx1_ASAP7_75t_L g966 ( .A(n_99), .Y(n_966) );
INVx1_ASAP7_75t_L g936 ( .A(n_100), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_101), .A2(n_138), .B1(n_620), .B2(n_621), .Y(n_619) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_101), .A2(n_138), .B1(n_547), .B2(n_551), .Y(n_625) );
AOI22xp33_ASAP7_75t_L g988 ( .A1(n_103), .A2(n_131), .B1(n_515), .B2(n_986), .Y(n_988) );
AOI22xp33_ASAP7_75t_L g996 ( .A1(n_103), .A2(n_131), .B1(n_386), .B2(n_997), .Y(n_996) );
INVxp67_ASAP7_75t_SL g854 ( .A(n_104), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_104), .A2(n_185), .B1(n_588), .B2(n_620), .Y(n_875) );
AOI22xp33_ASAP7_75t_L g1070 ( .A1(n_105), .A2(n_209), .B1(n_1007), .B2(n_1031), .Y(n_1070) );
INVxp33_ASAP7_75t_L g740 ( .A(n_106), .Y(n_740) );
INVxp33_ASAP7_75t_SL g1220 ( .A(n_107), .Y(n_1220) );
INVx1_ASAP7_75t_L g917 ( .A(n_110), .Y(n_917) );
OAI22xp33_ASAP7_75t_SL g948 ( .A1(n_110), .A2(n_145), .B1(n_263), .B2(n_547), .Y(n_948) );
AO22x2_ASAP7_75t_L g704 ( .A1(n_111), .A2(n_705), .B1(n_744), .B2(n_745), .Y(n_704) );
INVx1_ASAP7_75t_L g744 ( .A(n_111), .Y(n_744) );
INVxp67_ASAP7_75t_SL g1266 ( .A(n_112), .Y(n_1266) );
INVx1_ASAP7_75t_L g969 ( .A(n_113), .Y(n_969) );
INVx1_ASAP7_75t_L g254 ( .A(n_114), .Y(n_254) );
INVx1_ASAP7_75t_L g819 ( .A(n_116), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_116), .A2(n_201), .B1(n_594), .B2(n_797), .Y(n_835) );
INVx1_ASAP7_75t_L g1040 ( .A(n_119), .Y(n_1040) );
OAI22xp5_ASAP7_75t_L g633 ( .A1(n_120), .A2(n_184), .B1(n_263), .B2(n_335), .Y(n_633) );
OAI22xp33_ASAP7_75t_L g644 ( .A1(n_120), .A2(n_212), .B1(n_538), .B2(n_543), .Y(n_644) );
INVxp67_ASAP7_75t_SL g301 ( .A(n_121), .Y(n_301) );
OAI22xp5_ASAP7_75t_L g1272 ( .A1(n_122), .A2(n_1273), .B1(n_1274), .B2(n_1309), .Y(n_1272) );
CKINVDCx5p33_ASAP7_75t_R g1309 ( .A(n_122), .Y(n_1309) );
INVxp67_ASAP7_75t_SL g535 ( .A(n_123), .Y(n_535) );
INVx1_ASAP7_75t_L g715 ( .A(n_124), .Y(n_715) );
INVx1_ASAP7_75t_L g811 ( .A(n_125), .Y(n_811) );
AOI22xp5_ASAP7_75t_L g1030 ( .A1(n_126), .A2(n_173), .B1(n_1007), .B2(n_1031), .Y(n_1030) );
AOI22xp5_ASAP7_75t_L g1071 ( .A1(n_127), .A2(n_248), .B1(n_1021), .B2(n_1027), .Y(n_1071) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_128), .A2(n_155), .B1(n_386), .B2(n_388), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_128), .A2(n_155), .B1(n_411), .B2(n_413), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_130), .A2(n_133), .B1(n_720), .B2(n_721), .Y(n_719) );
AOI22xp33_ASAP7_75t_SL g732 ( .A1(n_130), .A2(n_133), .B1(n_483), .B2(n_602), .Y(n_732) );
XOR2xp5_ASAP7_75t_L g838 ( .A(n_132), .B(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g1179 ( .A(n_134), .Y(n_1179) );
INVxp33_ASAP7_75t_SL g708 ( .A(n_135), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_135), .A2(n_148), .B1(n_394), .B2(n_605), .Y(n_724) );
INVx1_ASAP7_75t_L g1286 ( .A(n_136), .Y(n_1286) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_137), .A2(n_142), .B1(n_602), .B2(n_603), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_137), .A2(n_142), .B1(n_505), .B2(n_616), .Y(n_615) );
OAI22xp33_ASAP7_75t_L g537 ( .A1(n_139), .A2(n_182), .B1(n_538), .B2(n_543), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_139), .A2(n_211), .B1(n_579), .B2(n_580), .Y(n_578) );
INVxp33_ASAP7_75t_L g1279 ( .A(n_140), .Y(n_1279) );
AOI22xp33_ASAP7_75t_L g1308 ( .A1(n_140), .A2(n_153), .B1(n_505), .B2(n_621), .Y(n_1308) );
INVx1_ASAP7_75t_L g910 ( .A(n_141), .Y(n_910) );
INVx1_ASAP7_75t_L g664 ( .A(n_143), .Y(n_664) );
INVxp33_ASAP7_75t_L g673 ( .A(n_144), .Y(n_673) );
INVx1_ASAP7_75t_L g921 ( .A(n_145), .Y(n_921) );
INVx1_ASAP7_75t_L g1283 ( .A(n_146), .Y(n_1283) );
INVxp67_ASAP7_75t_SL g711 ( .A(n_148), .Y(n_711) );
INVxp33_ASAP7_75t_SL g716 ( .A(n_149), .Y(n_716) );
AOI22xp33_ASAP7_75t_SL g723 ( .A1(n_149), .A2(n_172), .B1(n_483), .B2(n_602), .Y(n_723) );
INVx1_ASAP7_75t_L g931 ( .A(n_151), .Y(n_931) );
OAI22xp33_ASAP7_75t_L g938 ( .A1(n_151), .A2(n_170), .B1(n_538), .B2(n_892), .Y(n_938) );
INVx1_ASAP7_75t_L g849 ( .A(n_152), .Y(n_849) );
INVxp33_ASAP7_75t_L g1278 ( .A(n_153), .Y(n_1278) );
INVx1_ASAP7_75t_L g974 ( .A(n_154), .Y(n_974) );
INVxp33_ASAP7_75t_SL g1221 ( .A(n_156), .Y(n_1221) );
AOI22xp33_ASAP7_75t_SL g1238 ( .A1(n_156), .A2(n_190), .B1(n_1234), .B2(n_1239), .Y(n_1238) );
INVxp33_ASAP7_75t_L g1293 ( .A(n_157), .Y(n_1293) );
AOI22xp33_ASAP7_75t_L g1298 ( .A1(n_158), .A2(n_214), .B1(n_571), .B2(n_681), .Y(n_1298) );
AOI22xp33_ASAP7_75t_L g1303 ( .A1(n_158), .A2(n_214), .B1(n_614), .B2(n_1304), .Y(n_1303) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_160), .Y(n_256) );
AND3x2_ASAP7_75t_L g1011 ( .A(n_160), .B(n_254), .C(n_1012), .Y(n_1011) );
NAND2xp5_ASAP7_75t_L g1026 ( .A(n_160), .B(n_254), .Y(n_1026) );
INVxp33_ASAP7_75t_SL g317 ( .A(n_161), .Y(n_317) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_161), .A2(n_225), .B1(n_378), .B2(n_393), .Y(n_392) );
INVxp33_ASAP7_75t_SL g659 ( .A(n_162), .Y(n_659) );
INVxp33_ASAP7_75t_SL g676 ( .A(n_163), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g697 ( .A1(n_163), .A2(n_216), .B1(n_501), .B2(n_693), .Y(n_697) );
INVx1_ASAP7_75t_L g531 ( .A(n_164), .Y(n_531) );
INVx1_ASAP7_75t_L g860 ( .A(n_165), .Y(n_860) );
INVxp33_ASAP7_75t_L g1294 ( .A(n_166), .Y(n_1294) );
AOI22xp33_ASAP7_75t_L g1301 ( .A1(n_166), .A2(n_169), .B1(n_568), .B2(n_571), .Y(n_1301) );
INVx2_ASAP7_75t_L g267 ( .A(n_167), .Y(n_267) );
INVx1_ASAP7_75t_L g1289 ( .A(n_169), .Y(n_1289) );
INVx1_ASAP7_75t_L g934 ( .A(n_170), .Y(n_934) );
INVxp33_ASAP7_75t_SL g709 ( .A(n_172), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_174), .A2(n_193), .B1(n_564), .B2(n_565), .Y(n_563) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_174), .A2(n_193), .B1(n_505), .B2(n_587), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g1233 ( .A1(n_175), .A2(n_203), .B1(n_1234), .B2(n_1235), .Y(n_1233) );
AOI22xp33_ASAP7_75t_L g1245 ( .A1(n_175), .A2(n_203), .B1(n_1246), .B2(n_1247), .Y(n_1245) );
INVx1_ASAP7_75t_L g1012 ( .A(n_179), .Y(n_1012) );
OAI211xp5_ASAP7_75t_L g552 ( .A1(n_180), .A2(n_474), .B(n_553), .C(n_557), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_180), .A2(n_246), .B1(n_584), .B2(n_594), .Y(n_593) );
INVxp33_ASAP7_75t_SL g442 ( .A(n_181), .Y(n_442) );
OAI22xp5_ASAP7_75t_L g560 ( .A1(n_182), .A2(n_246), .B1(n_263), .B2(n_335), .Y(n_560) );
INVxp67_ASAP7_75t_SL g340 ( .A(n_183), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_183), .A2(n_218), .B1(n_421), .B2(n_424), .Y(n_420) );
INVxp67_ASAP7_75t_SL g851 ( .A(n_185), .Y(n_851) );
INVx1_ASAP7_75t_L g846 ( .A(n_187), .Y(n_846) );
INVxp33_ASAP7_75t_SL g461 ( .A(n_188), .Y(n_461) );
CKINVDCx5p33_ASAP7_75t_R g806 ( .A(n_189), .Y(n_806) );
INVxp33_ASAP7_75t_L g1224 ( .A(n_190), .Y(n_1224) );
INVx1_ASAP7_75t_L g269 ( .A(n_192), .Y(n_269) );
INVx2_ASAP7_75t_L g338 ( .A(n_192), .Y(n_338) );
INVx1_ASAP7_75t_L g763 ( .A(n_194), .Y(n_763) );
INVx1_ASAP7_75t_L g772 ( .A(n_195), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g796 ( .A1(n_195), .A2(n_240), .B1(n_583), .B2(n_797), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_196), .A2(n_223), .B1(n_341), .B2(n_681), .Y(n_784) );
AOI22xp33_ASAP7_75t_L g791 ( .A1(n_196), .A2(n_223), .B1(n_291), .B2(n_792), .Y(n_791) );
INVxp33_ASAP7_75t_SL g443 ( .A(n_197), .Y(n_443) );
INVxp33_ASAP7_75t_SL g364 ( .A(n_198), .Y(n_364) );
AO22x2_ASAP7_75t_L g276 ( .A1(n_199), .A2(n_277), .B1(n_435), .B2(n_436), .Y(n_276) );
CKINVDCx14_ASAP7_75t_R g435 ( .A(n_199), .Y(n_435) );
XNOR2xp5_ASAP7_75t_L g800 ( .A(n_200), .B(n_801), .Y(n_800) );
AOI22xp5_ASAP7_75t_L g1035 ( .A1(n_200), .A2(n_210), .B1(n_1021), .B2(n_1027), .Y(n_1035) );
INVx1_ASAP7_75t_L g816 ( .A(n_201), .Y(n_816) );
INVx1_ASAP7_75t_L g1046 ( .A(n_204), .Y(n_1046) );
INVx1_ASAP7_75t_L g865 ( .A(n_206), .Y(n_865) );
CKINVDCx5p33_ASAP7_75t_R g965 ( .A(n_207), .Y(n_965) );
INVx1_ASAP7_75t_L g879 ( .A(n_208), .Y(n_879) );
OAI22xp33_ASAP7_75t_SL g898 ( .A1(n_208), .A2(n_241), .B1(n_263), .B2(n_547), .Y(n_898) );
INVx1_ASAP7_75t_L g528 ( .A(n_211), .Y(n_528) );
INVx1_ASAP7_75t_L g306 ( .A(n_213), .Y(n_306) );
INVx1_ASAP7_75t_L g643 ( .A(n_215), .Y(n_643) );
INVxp67_ASAP7_75t_SL g669 ( .A(n_216), .Y(n_669) );
INVx1_ASAP7_75t_L g1010 ( .A(n_217), .Y(n_1010) );
NAND2xp5_ASAP7_75t_L g1029 ( .A(n_217), .B(n_1024), .Y(n_1029) );
INVxp33_ASAP7_75t_SL g332 ( .A(n_218), .Y(n_332) );
INVx1_ASAP7_75t_L g454 ( .A(n_219), .Y(n_454) );
XOR2x2_ASAP7_75t_L g651 ( .A(n_220), .B(n_652), .Y(n_651) );
INVxp67_ASAP7_75t_SL g736 ( .A(n_222), .Y(n_736) );
INVx1_ASAP7_75t_L g905 ( .A(n_224), .Y(n_905) );
INVx1_ASAP7_75t_L g290 ( .A(n_225), .Y(n_290) );
INVx1_ASAP7_75t_L g631 ( .A(n_226), .Y(n_631) );
INVx1_ASAP7_75t_L g1223 ( .A(n_227), .Y(n_1223) );
INVx1_ASAP7_75t_L g1227 ( .A(n_228), .Y(n_1227) );
OAI22xp5_ASAP7_75t_L g1263 ( .A1(n_228), .A2(n_239), .B1(n_559), .B2(n_738), .Y(n_1263) );
CKINVDCx5p33_ASAP7_75t_R g889 ( .A(n_229), .Y(n_889) );
INVx1_ASAP7_75t_L g809 ( .A(n_230), .Y(n_809) );
AO22x1_ASAP7_75t_L g1063 ( .A1(n_231), .A2(n_235), .B1(n_1031), .B2(n_1064), .Y(n_1063) );
INVx2_ASAP7_75t_L g266 ( .A(n_232), .Y(n_266) );
AO22x1_ASAP7_75t_L g1065 ( .A1(n_233), .A2(n_242), .B1(n_1021), .B2(n_1027), .Y(n_1065) );
INVx1_ASAP7_75t_L g922 ( .A(n_234), .Y(n_922) );
INVxp67_ASAP7_75t_SL g321 ( .A(n_236), .Y(n_321) );
INVxp33_ASAP7_75t_SL g473 ( .A(n_237), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_237), .A2(n_247), .B1(n_511), .B2(n_513), .Y(n_510) );
INVx1_ASAP7_75t_L g975 ( .A(n_238), .Y(n_975) );
INVx1_ASAP7_75t_L g1228 ( .A(n_239), .Y(n_1228) );
INVxp33_ASAP7_75t_L g777 ( .A(n_240), .Y(n_777) );
BUFx3_ASAP7_75t_L g287 ( .A(n_244), .Y(n_287) );
INVx1_ASAP7_75t_L g315 ( .A(n_244), .Y(n_315) );
BUFx3_ASAP7_75t_L g288 ( .A(n_245), .Y(n_288) );
INVx1_ASAP7_75t_L g324 ( .A(n_245), .Y(n_324) );
INVx1_ASAP7_75t_L g468 ( .A(n_247), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_270), .B(n_1004), .Y(n_249) );
BUFx3_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x4_ASAP7_75t_L g251 ( .A(n_252), .B(n_257), .Y(n_251) );
AND2x4_ASAP7_75t_L g1271 ( .A(n_252), .B(n_258), .Y(n_1271) );
NOR2xp33_ASAP7_75t_SL g252 ( .A(n_253), .B(n_255), .Y(n_252) );
INVx1_ASAP7_75t_SL g1311 ( .A(n_253), .Y(n_1311) );
NAND2xp5_ASAP7_75t_L g1316 ( .A(n_253), .B(n_255), .Y(n_1316) );
HB1xp67_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g1310 ( .A(n_255), .B(n_1311), .Y(n_1310) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_259), .B(n_263), .Y(n_258) );
INVxp67_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
OR2x2_ASAP7_75t_L g369 ( .A(n_260), .B(n_370), .Y(n_369) );
OR2x6_ASAP7_75t_L g476 ( .A(n_260), .B(n_370), .Y(n_476) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g376 ( .A(n_261), .B(n_269), .Y(n_376) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
OR2x2_ASAP7_75t_L g843 ( .A(n_262), .B(n_337), .Y(n_843) );
INVx8_ASAP7_75t_L g333 ( .A(n_263), .Y(n_333) );
OR2x6_ASAP7_75t_L g263 ( .A(n_264), .B(n_268), .Y(n_263) );
OR2x6_ASAP7_75t_L g335 ( .A(n_264), .B(n_336), .Y(n_335) );
BUFx6f_ASAP7_75t_L g845 ( .A(n_264), .Y(n_845) );
HB1xp67_ASAP7_75t_L g862 ( .A(n_264), .Y(n_862) );
INVx2_ASAP7_75t_SL g927 ( .A(n_264), .Y(n_927) );
BUFx6f_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
INVx1_ASAP7_75t_L g344 ( .A(n_266), .Y(n_344) );
INVx1_ASAP7_75t_L g356 ( .A(n_266), .Y(n_356) );
INVx2_ASAP7_75t_L g361 ( .A(n_266), .Y(n_361) );
AND2x4_ASAP7_75t_L g368 ( .A(n_266), .B(n_345), .Y(n_368) );
AND2x2_ASAP7_75t_L g381 ( .A(n_266), .B(n_267), .Y(n_381) );
INVx2_ASAP7_75t_L g345 ( .A(n_267), .Y(n_345) );
INVx1_ASAP7_75t_L g353 ( .A(n_267), .Y(n_353) );
INVx1_ASAP7_75t_L g363 ( .A(n_267), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_267), .B(n_361), .Y(n_550) );
INVx1_ASAP7_75t_L g556 ( .A(n_267), .Y(n_556) );
AND2x4_ASAP7_75t_L g352 ( .A(n_268), .B(n_353), .Y(n_352) );
INVx2_ASAP7_75t_SL g268 ( .A(n_269), .Y(n_268) );
OR2x2_ASAP7_75t_L g354 ( .A(n_269), .B(n_355), .Y(n_354) );
OR2x2_ASAP7_75t_L g738 ( .A(n_269), .B(n_355), .Y(n_738) );
OAI22xp33_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_272), .B1(n_747), .B2(n_748), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AOI22xp5_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_274), .B1(n_648), .B2(n_649), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AO22x1_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_522), .B1(n_646), .B2(n_647), .Y(n_274) );
INVx1_ASAP7_75t_L g646 ( .A(n_275), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g275 ( .A1(n_276), .A2(n_437), .B1(n_438), .B2(n_521), .Y(n_275) );
INVx1_ASAP7_75t_L g521 ( .A(n_276), .Y(n_521) );
INVx1_ASAP7_75t_L g436 ( .A(n_277), .Y(n_436) );
AOI211x1_ASAP7_75t_SL g277 ( .A1(n_278), .A2(n_325), .B(n_330), .C(n_371), .Y(n_277) );
NAND4xp25_ASAP7_75t_SL g278 ( .A(n_279), .B(n_289), .C(n_305), .D(n_316), .Y(n_278) );
NAND3xp33_ASAP7_75t_SL g526 ( .A(n_279), .B(n_527), .C(n_534), .Y(n_526) );
NAND3xp33_ASAP7_75t_SL g635 ( .A(n_279), .B(n_636), .C(n_641), .Y(n_635) );
NAND4xp25_ASAP7_75t_L g653 ( .A(n_279), .B(n_654), .C(n_657), .D(n_660), .Y(n_653) );
NAND4xp25_ASAP7_75t_L g706 ( .A(n_279), .B(n_707), .C(n_710), .D(n_714), .Y(n_706) );
NAND2xp5_ASAP7_75t_SL g886 ( .A(n_279), .B(n_887), .Y(n_886) );
NAND2xp5_ASAP7_75t_SL g940 ( .A(n_279), .B(n_941), .Y(n_940) );
CKINVDCx8_ASAP7_75t_R g279 ( .A(n_280), .Y(n_279) );
INVx5_ASAP7_75t_L g456 ( .A(n_280), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g956 ( .A(n_280), .B(n_957), .Y(n_956) );
AOI221xp5_ASAP7_75t_L g1290 ( .A1(n_280), .A2(n_307), .B1(n_310), .B2(n_1286), .C(n_1291), .Y(n_1290) );
AND2x4_ASAP7_75t_L g280 ( .A(n_281), .B(n_285), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x6_ASAP7_75t_L g322 ( .A(n_282), .B(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g539 ( .A(n_282), .Y(n_539) );
AND2x2_ASAP7_75t_L g762 ( .A(n_282), .B(n_614), .Y(n_762) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x6_ASAP7_75t_L g302 ( .A(n_283), .B(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_284), .Y(n_296) );
INVx1_ASAP7_75t_L g312 ( .A(n_284), .Y(n_312) );
AND2x2_ASAP7_75t_L g409 ( .A(n_284), .B(n_327), .Y(n_409) );
INVx2_ASAP7_75t_L g434 ( .A(n_284), .Y(n_434) );
INVx1_ASAP7_75t_L g292 ( .A(n_285), .Y(n_292) );
INVx2_ASAP7_75t_L g419 ( .A(n_285), .Y(n_419) );
BUFx6f_ASAP7_75t_L g614 ( .A(n_285), .Y(n_614) );
BUFx6f_ASAP7_75t_L g663 ( .A(n_285), .Y(n_663) );
BUFx6f_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_286), .Y(n_426) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
INVx2_ASAP7_75t_L g304 ( .A(n_287), .Y(n_304) );
AND2x4_ASAP7_75t_L g323 ( .A(n_287), .B(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g300 ( .A(n_288), .Y(n_300) );
AND2x4_ASAP7_75t_L g314 ( .A(n_288), .B(n_315), .Y(n_314) );
AOI222xp33_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_291), .B1(n_293), .B2(n_294), .C1(n_301), .C2(n_302), .Y(n_289) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
BUFx4f_ASAP7_75t_L g453 ( .A(n_294), .Y(n_453) );
AOI222xp33_ASAP7_75t_L g1225 ( .A1(n_294), .A2(n_302), .B1(n_513), .B2(n_1226), .C1(n_1227), .C2(n_1228), .Y(n_1225) );
AND2x4_ASAP7_75t_L g294 ( .A(n_295), .B(n_297), .Y(n_294) );
AND2x4_ASAP7_75t_L g307 ( .A(n_295), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_SL g532 ( .A(n_295), .B(n_297), .Y(n_532) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g640 ( .A(n_298), .Y(n_640) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x4_ASAP7_75t_L g308 ( .A(n_300), .B(n_304), .Y(n_308) );
AOI222xp33_ASAP7_75t_L g447 ( .A1(n_302), .A2(n_448), .B1(n_449), .B2(n_452), .C1(n_453), .C2(n_454), .Y(n_447) );
AOI222xp33_ASAP7_75t_L g527 ( .A1(n_302), .A2(n_528), .B1(n_529), .B2(n_531), .C1(n_532), .C2(n_533), .Y(n_527) );
AOI222xp33_ASAP7_75t_L g636 ( .A1(n_302), .A2(n_631), .B1(n_632), .B2(n_637), .C1(n_638), .C2(n_639), .Y(n_636) );
AOI222xp33_ASAP7_75t_L g660 ( .A1(n_302), .A2(n_532), .B1(n_661), .B2(n_662), .C1(n_664), .C2(n_665), .Y(n_660) );
AOI222xp33_ASAP7_75t_L g710 ( .A1(n_302), .A2(n_424), .B1(n_532), .B2(n_711), .C1(n_712), .C2(n_713), .Y(n_710) );
INVx3_ASAP7_75t_L g766 ( .A(n_302), .Y(n_766) );
AOI222xp33_ASAP7_75t_L g887 ( .A1(n_302), .A2(n_639), .B1(n_865), .B2(n_888), .C1(n_889), .C2(n_890), .Y(n_887) );
AOI222xp33_ASAP7_75t_L g941 ( .A1(n_302), .A2(n_418), .B1(n_639), .B2(n_936), .C1(n_942), .C2(n_943), .Y(n_941) );
AOI222xp33_ASAP7_75t_L g1288 ( .A1(n_302), .A2(n_532), .B1(n_662), .B2(n_1282), .C1(n_1283), .C2(n_1289), .Y(n_1288) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AOI22xp33_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_307), .B1(n_309), .B2(n_310), .Y(n_305) );
AOI22xp5_ASAP7_75t_L g331 ( .A1(n_306), .A2(n_332), .B1(n_333), .B2(n_334), .Y(n_331) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_307), .A2(n_310), .B1(n_445), .B2(n_446), .Y(n_444) );
INVx4_ASAP7_75t_L g543 ( .A(n_307), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_307), .A2(n_310), .B1(n_658), .B2(n_659), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g714 ( .A1(n_307), .A2(n_310), .B1(n_715), .B2(n_716), .Y(n_714) );
AOI22xp5_ASAP7_75t_SL g758 ( .A1(n_307), .A2(n_318), .B1(n_759), .B2(n_760), .Y(n_758) );
AOI22xp5_ASAP7_75t_SL g803 ( .A1(n_307), .A2(n_804), .B1(n_805), .B2(n_806), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g964 ( .A1(n_307), .A2(n_310), .B1(n_965), .B2(n_966), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g1222 ( .A1(n_307), .A2(n_310), .B1(n_1223), .B2(n_1224), .Y(n_1222) );
INVx6_ASAP7_75t_L g320 ( .A(n_308), .Y(n_320) );
BUFx2_ASAP7_75t_L g583 ( .A(n_308), .Y(n_583) );
INVx2_ASAP7_75t_L g595 ( .A(n_308), .Y(n_595) );
AOI22xp5_ASAP7_75t_L g534 ( .A1(n_310), .A2(n_322), .B1(n_535), .B2(n_536), .Y(n_534) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_310), .A2(n_322), .B1(n_642), .B2(n_643), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g767 ( .A1(n_310), .A2(n_322), .B1(n_768), .B2(n_769), .Y(n_767) );
AOI22xp5_ASAP7_75t_L g807 ( .A1(n_310), .A2(n_322), .B1(n_808), .B2(n_809), .Y(n_807) );
INVx4_ASAP7_75t_L g893 ( .A(n_310), .Y(n_893) );
AND2x6_ASAP7_75t_L g310 ( .A(n_311), .B(n_313), .Y(n_310) );
AND2x4_ASAP7_75t_L g318 ( .A(n_311), .B(n_319), .Y(n_318) );
AND2x4_ASAP7_75t_L g805 ( .A(n_311), .B(n_319), .Y(n_805) );
INVx1_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g639 ( .A(n_312), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g414 ( .A(n_313), .Y(n_414) );
INVx1_ASAP7_75t_L g431 ( .A(n_313), .Y(n_431) );
INVx2_ASAP7_75t_L g507 ( .A(n_313), .Y(n_507) );
BUFx6f_ASAP7_75t_L g621 ( .A(n_313), .Y(n_621) );
BUFx6f_ASAP7_75t_L g721 ( .A(n_313), .Y(n_721) );
INVx1_ASAP7_75t_L g1248 ( .A(n_313), .Y(n_1248) );
BUFx6f_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
BUFx6f_ASAP7_75t_L g588 ( .A(n_314), .Y(n_588) );
INVx1_ASAP7_75t_L g617 ( .A(n_314), .Y(n_617) );
INVx2_ASAP7_75t_L g702 ( .A(n_314), .Y(n_702) );
INVx1_ASAP7_75t_L g1258 ( .A(n_314), .Y(n_1258) );
INVx1_ASAP7_75t_L g541 ( .A(n_315), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_318), .B1(n_321), .B2(n_322), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_318), .A2(n_322), .B1(n_442), .B2(n_443), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_318), .A2(n_322), .B1(n_655), .B2(n_656), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_318), .A2(n_322), .B1(n_708), .B2(n_709), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g1219 ( .A1(n_318), .A2(n_322), .B1(n_1220), .B2(n_1221), .Y(n_1219) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx2_ASAP7_75t_L g417 ( .A(n_320), .Y(n_417) );
INVx2_ASAP7_75t_SL g423 ( .A(n_320), .Y(n_423) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_320), .Y(n_500) );
HB1xp67_ASAP7_75t_L g512 ( .A(n_320), .Y(n_512) );
INVx1_ASAP7_75t_L g623 ( .A(n_320), .Y(n_623) );
INVx1_ASAP7_75t_L g792 ( .A(n_320), .Y(n_792) );
CKINVDCx6p67_ASAP7_75t_R g892 ( .A(n_322), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g961 ( .A1(n_322), .A2(n_805), .B1(n_962), .B2(n_963), .Y(n_961) );
AOI22xp5_ASAP7_75t_L g1292 ( .A1(n_322), .A2(n_805), .B1(n_1293), .B2(n_1294), .Y(n_1292) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_323), .Y(n_412) );
INVx2_ASAP7_75t_SL g429 ( .A(n_323), .Y(n_429) );
BUFx6f_ASAP7_75t_L g505 ( .A(n_323), .Y(n_505) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_323), .Y(n_515) );
BUFx6f_ASAP7_75t_L g620 ( .A(n_323), .Y(n_620) );
BUFx2_ASAP7_75t_L g695 ( .A(n_323), .Y(n_695) );
BUFx6f_ASAP7_75t_L g720 ( .A(n_323), .Y(n_720) );
BUFx3_ASAP7_75t_L g730 ( .A(n_323), .Y(n_730) );
INVx1_ASAP7_75t_L g542 ( .A(n_324), .Y(n_542) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_325), .Y(n_457) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_325), .A2(n_475), .B1(n_653), .B2(n_666), .C(n_677), .Y(n_652) );
INVx1_ASAP7_75t_L g1230 ( .A(n_325), .Y(n_1230) );
AOI221x1_ASAP7_75t_L g1275 ( .A1(n_325), .A2(n_475), .B1(n_1276), .B2(n_1287), .C(n_1295), .Y(n_1275) );
AND2x4_ASAP7_75t_L g325 ( .A(n_326), .B(n_328), .Y(n_325) );
AND2x4_ASAP7_75t_L g544 ( .A(n_326), .B(n_328), .Y(n_544) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AND2x4_ASAP7_75t_L g433 ( .A(n_327), .B(n_434), .Y(n_433) );
BUFx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx2_ASAP7_75t_L g375 ( .A(n_329), .Y(n_375) );
OR2x6_ASAP7_75t_L g842 ( .A(n_329), .B(n_843), .Y(n_842) );
AOI31xp33_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_339), .A3(n_357), .B(n_369), .Y(n_330) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_333), .A2(n_334), .B1(n_445), .B2(n_473), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g675 ( .A1(n_333), .A2(n_334), .B1(n_658), .B2(n_676), .Y(n_675) );
AOI22xp33_ASAP7_75t_SL g742 ( .A1(n_333), .A2(n_334), .B1(n_715), .B2(n_743), .Y(n_742) );
AOI22xp33_ASAP7_75t_SL g776 ( .A1(n_333), .A2(n_359), .B1(n_777), .B2(n_778), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_333), .A2(n_359), .B1(n_819), .B2(n_820), .Y(n_818) );
AOI22xp33_ASAP7_75t_L g977 ( .A1(n_333), .A2(n_965), .B1(n_978), .B2(n_979), .Y(n_977) );
AOI22xp33_ASAP7_75t_SL g1267 ( .A1(n_333), .A2(n_334), .B1(n_1223), .B2(n_1268), .Y(n_1267) );
AOI22xp33_ASAP7_75t_L g1284 ( .A1(n_333), .A2(n_334), .B1(n_1285), .B2(n_1286), .Y(n_1284) );
AOI22xp33_ASAP7_75t_SL g779 ( .A1(n_334), .A2(n_365), .B1(n_760), .B2(n_780), .Y(n_779) );
AOI22xp33_ASAP7_75t_L g821 ( .A1(n_334), .A2(n_365), .B1(n_806), .B2(n_822), .Y(n_821) );
INVx5_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx4_ASAP7_75t_L g979 ( .A(n_335), .Y(n_979) );
AND2x4_ASAP7_75t_L g359 ( .A(n_336), .B(n_360), .Y(n_359) );
AND2x4_ASAP7_75t_L g365 ( .A(n_336), .B(n_366), .Y(n_365) );
AND2x4_ASAP7_75t_L g462 ( .A(n_336), .B(n_366), .Y(n_462) );
INVx1_ASAP7_75t_L g548 ( .A(n_336), .Y(n_548) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g349 ( .A(n_338), .Y(n_349) );
AOI211xp5_ASAP7_75t_L g339 ( .A1(n_340), .A2(n_341), .B(n_346), .C(n_350), .Y(n_339) );
INVx2_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x4_ASAP7_75t_L g346 ( .A(n_343), .B(n_347), .Y(n_346) );
BUFx6f_ASAP7_75t_L g384 ( .A(n_343), .Y(n_384) );
BUFx6f_ASAP7_75t_L g394 ( .A(n_343), .Y(n_394) );
BUFx2_ASAP7_75t_L g471 ( .A(n_343), .Y(n_471) );
BUFx3_ASAP7_75t_L g572 ( .A(n_343), .Y(n_572) );
BUFx3_ASAP7_75t_L g774 ( .A(n_343), .Y(n_774) );
AND2x4_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
CKINVDCx11_ASAP7_75t_R g474 ( .A(n_346), .Y(n_474) );
AOI211xp5_ASAP7_75t_L g667 ( .A1(n_346), .A2(n_668), .B(n_669), .C(n_670), .Y(n_667) );
AOI211xp5_ASAP7_75t_L g735 ( .A1(n_346), .A2(n_393), .B(n_736), .C(n_737), .Y(n_735) );
AOI211xp5_ASAP7_75t_L g771 ( .A1(n_346), .A2(n_772), .B(n_773), .C(n_775), .Y(n_771) );
AOI211xp5_ASAP7_75t_L g815 ( .A1(n_346), .A2(n_382), .B(n_816), .C(n_817), .Y(n_815) );
AOI211xp5_ASAP7_75t_L g1260 ( .A1(n_346), .A2(n_1261), .B(n_1262), .C(n_1263), .Y(n_1260) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVxp67_ASAP7_75t_L g467 ( .A(n_348), .Y(n_467) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
NAND2x1p5_ASAP7_75t_L g403 ( .A(n_349), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g464 ( .A(n_351), .Y(n_464) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g559 ( .A(n_352), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_352), .A2(n_465), .B1(n_631), .B2(n_632), .Y(n_630) );
INVx2_ASAP7_75t_L g671 ( .A(n_352), .Y(n_671) );
AOI22xp5_ASAP7_75t_L g897 ( .A1(n_352), .A2(n_465), .B1(n_889), .B2(n_890), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_352), .A2(n_465), .B1(n_942), .B2(n_943), .Y(n_947) );
INVx1_ASAP7_75t_L g466 ( .A(n_355), .Y(n_466) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g555 ( .A(n_356), .B(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g848 ( .A(n_356), .B(n_556), .Y(n_848) );
AOI22xp5_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_359), .B1(n_364), .B2(n_365), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_359), .A2(n_460), .B1(n_461), .B2(n_462), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_359), .A2(n_462), .B1(n_673), .B2(n_674), .Y(n_672) );
AOI22xp33_ASAP7_75t_SL g739 ( .A1(n_359), .A2(n_462), .B1(n_740), .B2(n_741), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g968 ( .A1(n_359), .A2(n_365), .B1(n_969), .B2(n_970), .Y(n_968) );
AOI22xp33_ASAP7_75t_SL g1264 ( .A1(n_359), .A2(n_462), .B1(n_1265), .B2(n_1266), .Y(n_1264) );
AOI22xp33_ASAP7_75t_L g1277 ( .A1(n_359), .A2(n_462), .B1(n_1278), .B2(n_1279), .Y(n_1277) );
INVx1_ASAP7_75t_L g387 ( .A(n_360), .Y(n_387) );
INVx1_ASAP7_75t_L g397 ( .A(n_360), .Y(n_397) );
BUFx2_ASAP7_75t_L g480 ( .A(n_360), .Y(n_480) );
BUFx6f_ASAP7_75t_L g575 ( .A(n_360), .Y(n_575) );
BUFx6f_ASAP7_75t_L g602 ( .A(n_360), .Y(n_602) );
BUFx6f_ASAP7_75t_L g829 ( .A(n_360), .Y(n_829) );
AND2x4_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx5_ASAP7_75t_SL g551 ( .A(n_365), .Y(n_551) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
HB1xp67_ASAP7_75t_L g788 ( .A(n_367), .Y(n_788) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx3_ASAP7_75t_L g391 ( .A(n_368), .Y(n_391) );
BUFx6f_ASAP7_75t_L g483 ( .A(n_368), .Y(n_483) );
INVx1_ASAP7_75t_L g687 ( .A(n_368), .Y(n_687) );
AOI31xp33_ASAP7_75t_L g734 ( .A1(n_369), .A2(n_735), .A3(n_739), .B(n_742), .Y(n_734) );
AOI31xp33_ASAP7_75t_L g770 ( .A1(n_369), .A2(n_771), .A3(n_776), .B(n_779), .Y(n_770) );
AOI31xp33_ASAP7_75t_L g814 ( .A1(n_369), .A2(n_815), .A3(n_818), .B(n_821), .Y(n_814) );
AOI31xp33_ASAP7_75t_L g1259 ( .A1(n_369), .A2(n_1260), .A3(n_1264), .B(n_1267), .Y(n_1259) );
AND2x4_ASAP7_75t_L g432 ( .A(n_370), .B(n_433), .Y(n_432) );
AND2x4_ASAP7_75t_L g518 ( .A(n_370), .B(n_433), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_372), .B(n_405), .Y(n_371) );
AOI33xp33_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_377), .A3(n_385), .B1(n_392), .B2(n_395), .B3(n_399), .Y(n_372) );
BUFx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AND2x4_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
OR2x6_ASAP7_75t_L g407 ( .A(n_375), .B(n_408), .Y(n_407) );
AND2x4_ASAP7_75t_L g489 ( .A(n_375), .B(n_376), .Y(n_489) );
OR2x2_ASAP7_75t_L g590 ( .A(n_375), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g725 ( .A(n_375), .B(n_726), .Y(n_725) );
OR2x2_ASAP7_75t_L g903 ( .A(n_375), .B(n_408), .Y(n_903) );
BUFx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g496 ( .A(n_379), .Y(n_496) );
INVx1_ASAP7_75t_L g690 ( .A(n_379), .Y(n_690) );
BUFx3_ASAP7_75t_L g1237 ( .A(n_379), .Y(n_1237) );
INVx2_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g485 ( .A(n_380), .Y(n_485) );
INVx2_ASAP7_75t_SL g994 ( .A(n_380), .Y(n_994) );
INVx3_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
BUFx6f_ASAP7_75t_L g570 ( .A(n_381), .Y(n_570) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g580 ( .A(n_383), .Y(n_580) );
INVx2_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
HB1xp67_ASAP7_75t_L g995 ( .A(n_384), .Y(n_995) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx2_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g398 ( .A(n_389), .Y(n_398) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx2_ASAP7_75t_L g566 ( .A(n_390), .Y(n_566) );
INVx1_ASAP7_75t_L g855 ( .A(n_390), .Y(n_855) );
INVx3_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
BUFx6f_ASAP7_75t_L g577 ( .A(n_391), .Y(n_577) );
INVx3_ASAP7_75t_L g859 ( .A(n_391), .Y(n_859) );
BUFx6f_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_SL g1243 ( .A(n_394), .Y(n_1243) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g564 ( .A(n_397), .Y(n_564) );
NAND3xp33_ASAP7_75t_L g490 ( .A(n_399), .B(n_491), .C(n_494), .Y(n_490) );
NAND3xp33_ASAP7_75t_L g573 ( .A(n_399), .B(n_574), .C(n_578), .Y(n_573) );
NAND3xp33_ASAP7_75t_L g678 ( .A(n_399), .B(n_679), .C(n_680), .Y(n_678) );
AOI33xp33_ASAP7_75t_L g989 ( .A1(n_399), .A2(n_489), .A3(n_990), .B1(n_992), .B2(n_996), .B3(n_1000), .Y(n_989) );
AOI33xp33_ASAP7_75t_L g1232 ( .A1(n_399), .A2(n_487), .A3(n_1233), .B1(n_1236), .B2(n_1238), .B3(n_1241), .Y(n_1232) );
INVx5_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx6_ASAP7_75t_L g610 ( .A(n_400), .Y(n_610) );
OR2x6_ASAP7_75t_L g400 ( .A(n_401), .B(n_403), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g726 ( .A(n_403), .Y(n_726) );
AOI33xp33_ASAP7_75t_L g405 ( .A1(n_406), .A2(n_410), .A3(n_415), .B1(n_420), .B2(n_427), .B3(n_432), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
CKINVDCx5p33_ASAP7_75t_R g508 ( .A(n_407), .Y(n_508) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g591 ( .A(n_409), .Y(n_591) );
BUFx4f_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g906 ( .A(n_412), .Y(n_906) );
BUFx2_ASAP7_75t_L g1256 ( .A(n_412), .Y(n_1256) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
BUFx6f_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx3_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g451 ( .A(n_419), .Y(n_451) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
BUFx4f_ASAP7_75t_L g501 ( .A(n_426), .Y(n_501) );
BUFx3_ASAP7_75t_L g513 ( .A(n_426), .Y(n_513) );
INVx1_ASAP7_75t_L g530 ( .A(n_426), .Y(n_530) );
INVx2_ASAP7_75t_SL g585 ( .A(n_426), .Y(n_585) );
BUFx6f_ASAP7_75t_L g797 ( .A(n_426), .Y(n_797) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_SL g794 ( .A(n_429), .Y(n_794) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
NAND3xp33_ASAP7_75t_L g592 ( .A(n_432), .B(n_593), .C(n_596), .Y(n_592) );
NAND3xp33_ASAP7_75t_L g618 ( .A(n_432), .B(n_619), .C(n_622), .Y(n_618) );
NAND3xp33_ASAP7_75t_L g696 ( .A(n_432), .B(n_697), .C(n_698), .Y(n_696) );
AOI33xp33_ASAP7_75t_L g727 ( .A1(n_432), .A2(n_489), .A3(n_728), .B1(n_729), .B2(n_732), .B3(n_733), .Y(n_727) );
NAND3xp33_ASAP7_75t_L g795 ( .A(n_432), .B(n_796), .C(n_798), .Y(n_795) );
NAND3xp33_ASAP7_75t_L g834 ( .A(n_432), .B(n_835), .C(n_836), .Y(n_834) );
INVx1_ASAP7_75t_L g923 ( .A(n_432), .Y(n_923) );
NAND3xp33_ASAP7_75t_L g1306 ( .A(n_432), .B(n_1307), .C(n_1308), .Y(n_1306) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g520 ( .A(n_439), .Y(n_520) );
AOI221x1_ASAP7_75t_L g439 ( .A1(n_440), .A2(n_457), .B1(n_458), .B2(n_475), .C(n_477), .Y(n_439) );
NAND4xp25_ASAP7_75t_L g440 ( .A(n_441), .B(n_444), .C(n_447), .D(n_455), .Y(n_440) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
AOI222xp33_ASAP7_75t_L g463 ( .A1(n_452), .A2(n_454), .B1(n_464), .B2(n_465), .C1(n_468), .C2(n_469), .Y(n_463) );
BUFx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NAND4xp25_ASAP7_75t_L g757 ( .A(n_456), .B(n_758), .C(n_761), .D(n_767), .Y(n_757) );
NAND4xp25_ASAP7_75t_L g802 ( .A(n_456), .B(n_803), .C(n_807), .D(n_810), .Y(n_802) );
NAND4xp25_ASAP7_75t_L g1218 ( .A(n_456), .B(n_1219), .C(n_1222), .D(n_1225), .Y(n_1218) );
AOI221x1_ASAP7_75t_L g954 ( .A1(n_457), .A2(n_475), .B1(n_955), .B2(n_967), .C(n_980), .Y(n_954) );
NAND4xp25_ASAP7_75t_SL g458 ( .A(n_459), .B(n_463), .C(n_472), .D(n_474), .Y(n_458) );
AOI222xp33_ASAP7_75t_L g971 ( .A1(n_464), .A2(n_972), .B1(n_973), .B2(n_974), .C1(n_975), .C2(n_976), .Y(n_971) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_465), .A2(n_531), .B1(n_533), .B2(n_558), .Y(n_557) );
AND2x4_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
AND2x4_ASAP7_75t_L g976 ( .A(n_466), .B(n_467), .Y(n_976) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g486 ( .A(n_470), .Y(n_486) );
INVx1_ASAP7_75t_L g973 ( .A(n_470), .Y(n_973) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
AOI222xp33_ASAP7_75t_L g1280 ( .A1(n_471), .A2(n_558), .B1(n_976), .B2(n_1281), .C1(n_1282), .C2(n_1283), .Y(n_1280) );
NAND4xp25_ASAP7_75t_SL g967 ( .A(n_474), .B(n_968), .C(n_971), .D(n_977), .Y(n_967) );
NAND4xp25_ASAP7_75t_L g1276 ( .A(n_474), .B(n_1277), .C(n_1280), .D(n_1284), .Y(n_1276) );
OAI31xp33_ASAP7_75t_L g545 ( .A1(n_475), .A2(n_546), .A3(n_552), .B(n_560), .Y(n_545) );
OAI31xp33_ASAP7_75t_SL g624 ( .A1(n_475), .A2(n_625), .A3(n_626), .B(n_633), .Y(n_624) );
OAI31xp33_ASAP7_75t_SL g894 ( .A1(n_475), .A2(n_895), .A3(n_896), .B(n_898), .Y(n_894) );
OAI31xp33_ASAP7_75t_SL g944 ( .A1(n_475), .A2(n_945), .A3(n_946), .B(n_948), .Y(n_944) );
CKINVDCx16_ASAP7_75t_R g475 ( .A(n_476), .Y(n_475) );
NAND4xp25_ASAP7_75t_L g477 ( .A(n_478), .B(n_490), .C(n_497), .D(n_509), .Y(n_477) );
NAND3xp33_ASAP7_75t_L g478 ( .A(n_479), .B(n_484), .C(n_487), .Y(n_478) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_SL g482 ( .A(n_483), .Y(n_482) );
INVx4_ASAP7_75t_L g493 ( .A(n_483), .Y(n_493) );
INVx2_ASAP7_75t_SL g1240 ( .A(n_483), .Y(n_1240) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
NAND3xp33_ASAP7_75t_L g562 ( .A(n_489), .B(n_563), .C(n_567), .Y(n_562) );
NAND3xp33_ASAP7_75t_L g600 ( .A(n_489), .B(n_601), .C(n_604), .Y(n_600) );
NAND3xp33_ASAP7_75t_L g682 ( .A(n_489), .B(n_683), .C(n_688), .Y(n_682) );
NAND3xp33_ASAP7_75t_L g782 ( .A(n_489), .B(n_783), .C(n_784), .Y(n_782) );
NAND3xp33_ASAP7_75t_L g824 ( .A(n_489), .B(n_825), .C(n_826), .Y(n_824) );
NAND3xp33_ASAP7_75t_L g1296 ( .A(n_489), .B(n_1297), .C(n_1298), .Y(n_1296) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
NAND3xp33_ASAP7_75t_L g497 ( .A(n_498), .B(n_502), .C(n_508), .Y(n_497) );
INVx4_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g693 ( .A(n_500), .Y(n_693) );
INVx1_ASAP7_75t_L g1304 ( .A(n_500), .Y(n_1304) );
INVx2_ASAP7_75t_SL g503 ( .A(n_504), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g516 ( .A(n_507), .Y(n_516) );
OAI22xp5_ASAP7_75t_L g919 ( .A1(n_507), .A2(n_920), .B1(n_921), .B2(n_922), .Y(n_919) );
AOI33xp33_ASAP7_75t_L g1244 ( .A1(n_508), .A2(n_518), .A3(n_1245), .B1(n_1249), .B2(n_1252), .B3(n_1255), .Y(n_1244) );
NAND3xp33_ASAP7_75t_L g509 ( .A(n_510), .B(n_514), .C(n_517), .Y(n_509) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
BUFx4f_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx4_ASAP7_75t_L g876 ( .A(n_518), .Y(n_876) );
BUFx4f_ASAP7_75t_L g982 ( .A(n_518), .Y(n_982) );
INVx2_ASAP7_75t_L g647 ( .A(n_522), .Y(n_647) );
XOR2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_597), .Y(n_522) );
NAND3x1_ASAP7_75t_L g524 ( .A(n_525), .B(n_545), .C(n_561), .Y(n_524) );
OAI21xp5_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_537), .B(n_544), .Y(n_525) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g638 ( .A(n_530), .Y(n_638) );
OR2x2_ASAP7_75t_L g538 ( .A(n_539), .B(n_540), .Y(n_538) );
INVx2_ASAP7_75t_L g870 ( .A(n_540), .Y(n_870) );
INVx1_ASAP7_75t_L g912 ( .A(n_540), .Y(n_912) );
OR2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
AND2x2_ASAP7_75t_L g874 ( .A(n_541), .B(n_542), .Y(n_874) );
OAI21xp5_ASAP7_75t_SL g634 ( .A1(n_544), .A2(n_635), .B(n_644), .Y(n_634) );
AOI211x1_ASAP7_75t_L g705 ( .A1(n_544), .A2(n_706), .B(n_717), .C(n_734), .Y(n_705) );
AOI211xp5_ASAP7_75t_L g756 ( .A1(n_544), .A2(n_757), .B(n_770), .C(n_781), .Y(n_756) );
AOI211xp5_ASAP7_75t_L g801 ( .A1(n_544), .A2(n_802), .B(n_814), .C(n_823), .Y(n_801) );
OAI31xp33_ASAP7_75t_SL g884 ( .A1(n_544), .A2(n_885), .A3(n_886), .B(n_891), .Y(n_884) );
OAI31xp33_ASAP7_75t_L g937 ( .A1(n_544), .A2(n_938), .A3(n_939), .B(n_940), .Y(n_937) );
OR2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
BUFx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g853 ( .A(n_550), .Y(n_853) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
BUFx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g629 ( .A(n_555), .Y(n_629) );
INVx2_ASAP7_75t_L g864 ( .A(n_555), .Y(n_864) );
INVx3_ASAP7_75t_L g935 ( .A(n_555), .Y(n_935) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND4x1_ASAP7_75t_L g561 ( .A(n_562), .B(n_573), .C(n_581), .D(n_592), .Y(n_561) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
INVx2_ASAP7_75t_SL g568 ( .A(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g605 ( .A(n_569), .Y(n_605) );
INVx2_ASAP7_75t_L g681 ( .A(n_569), .Y(n_681) );
INVx3_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
BUFx2_ASAP7_75t_L g579 ( .A(n_570), .Y(n_579) );
HB1xp67_ASAP7_75t_L g668 ( .A(n_571), .Y(n_668) );
BUFx6f_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g1002 ( .A(n_572), .Y(n_1002) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g603 ( .A(n_577), .Y(n_603) );
INVx2_ASAP7_75t_L g608 ( .A(n_577), .Y(n_608) );
NAND3xp33_ASAP7_75t_L g581 ( .A(n_582), .B(n_586), .C(n_589), .Y(n_581) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g888 ( .A(n_585), .Y(n_888) );
INVx1_ASAP7_75t_L g984 ( .A(n_585), .Y(n_984) );
BUFx6f_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g908 ( .A(n_588), .Y(n_908) );
NAND3xp33_ASAP7_75t_L g611 ( .A(n_589), .B(n_612), .C(n_615), .Y(n_611) );
NAND3xp33_ASAP7_75t_L g691 ( .A(n_589), .B(n_692), .C(n_694), .Y(n_691) );
AOI33xp33_ASAP7_75t_L g718 ( .A1(n_589), .A2(n_719), .A3(n_722), .B1(n_723), .B2(n_724), .B3(n_725), .Y(n_718) );
NAND3xp33_ASAP7_75t_L g790 ( .A(n_589), .B(n_791), .C(n_793), .Y(n_790) );
NAND3xp33_ASAP7_75t_L g831 ( .A(n_589), .B(n_832), .C(n_833), .Y(n_831) );
AOI33xp33_ASAP7_75t_L g981 ( .A1(n_589), .A2(n_982), .A3(n_983), .B1(n_985), .B2(n_987), .B3(n_988), .Y(n_981) );
NAND3xp33_ASAP7_75t_L g1302 ( .A(n_589), .B(n_1303), .C(n_1305), .Y(n_1302) );
INVx3_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OAI22xp5_ASAP7_75t_SL g867 ( .A1(n_590), .A2(n_868), .B1(n_876), .B2(n_877), .Y(n_867) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_SL g613 ( .A(n_595), .Y(n_613) );
XOR2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_645), .Y(n_597) );
NAND3xp33_ASAP7_75t_L g598 ( .A(n_599), .B(n_624), .C(n_634), .Y(n_598) );
AND4x1_ASAP7_75t_L g599 ( .A(n_600), .B(n_606), .C(n_611), .D(n_618), .Y(n_599) );
BUFx3_ASAP7_75t_L g1234 ( .A(n_602), .Y(n_1234) );
NAND3xp33_ASAP7_75t_L g606 ( .A(n_607), .B(n_609), .C(n_610), .Y(n_606) );
HB1xp67_ASAP7_75t_L g1235 ( .A(n_608), .Y(n_1235) );
BUFx2_ASAP7_75t_L g1250 ( .A(n_613), .Y(n_1250) );
HB1xp67_ASAP7_75t_L g1251 ( .A(n_614), .Y(n_1251) );
INVx2_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g765 ( .A(n_639), .Y(n_765) );
INVx1_ASAP7_75t_L g813 ( .A(n_639), .Y(n_813) );
OAI22xp33_ASAP7_75t_L g1045 ( .A1(n_645), .A2(n_1041), .B1(n_1043), .B2(n_1046), .Y(n_1045) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_703), .B1(n_704), .B2(n_746), .Y(n_650) );
INVx1_ASAP7_75t_L g746 ( .A(n_651), .Y(n_746) );
BUFx6f_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NAND3xp33_ASAP7_75t_L g666 ( .A(n_667), .B(n_672), .C(n_675), .Y(n_666) );
NAND4xp25_ASAP7_75t_L g677 ( .A(n_678), .B(n_682), .C(n_691), .D(n_696), .Y(n_677) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g991 ( .A(n_685), .Y(n_991) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g999 ( .A(n_687), .Y(n_999) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx2_ASAP7_75t_SL g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g986 ( .A(n_700), .Y(n_986) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
BUFx2_ASAP7_75t_L g731 ( .A(n_701), .Y(n_731) );
INVx2_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx2_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g745 ( .A(n_705), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_718), .B(n_727), .Y(n_717) );
INVx1_ASAP7_75t_L g920 ( .A(n_720), .Y(n_920) );
NAND3xp33_ASAP7_75t_L g785 ( .A(n_725), .B(n_786), .C(n_789), .Y(n_785) );
NAND3xp33_ASAP7_75t_L g827 ( .A(n_725), .B(n_828), .C(n_830), .Y(n_827) );
INVx1_ASAP7_75t_L g866 ( .A(n_725), .Y(n_866) );
NAND3xp33_ASAP7_75t_L g1299 ( .A(n_725), .B(n_1300), .C(n_1301), .Y(n_1299) );
BUFx3_ASAP7_75t_L g1246 ( .A(n_730), .Y(n_1246) );
OAI22xp5_ASAP7_75t_L g1039 ( .A1(n_744), .A2(n_1040), .B1(n_1041), .B2(n_1043), .Y(n_1039) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_750), .B1(n_951), .B2(n_952), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
XOR2x2_ASAP7_75t_L g751 ( .A(n_752), .B(n_837), .Y(n_751) );
OAI22xp5_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_754), .B1(n_799), .B2(n_800), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
XNOR2xp5_ASAP7_75t_L g754 ( .A(n_755), .B(n_756), .Y(n_754) );
AOI21xp5_ASAP7_75t_L g761 ( .A1(n_762), .A2(n_763), .B(n_764), .Y(n_761) );
AOI21xp5_ASAP7_75t_L g810 ( .A1(n_762), .A2(n_811), .B(n_812), .Y(n_810) );
BUFx2_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
NAND4xp25_ASAP7_75t_L g781 ( .A(n_782), .B(n_785), .C(n_790), .D(n_795), .Y(n_781) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g1254 ( .A(n_797), .Y(n_1254) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
NAND4xp25_ASAP7_75t_L g823 ( .A(n_824), .B(n_827), .C(n_831), .D(n_834), .Y(n_823) );
OAI22xp5_ASAP7_75t_L g837 ( .A1(n_838), .A2(n_899), .B1(n_949), .B2(n_950), .Y(n_837) );
INVx1_ASAP7_75t_L g949 ( .A(n_838), .Y(n_949) );
NAND3xp33_ASAP7_75t_L g839 ( .A(n_840), .B(n_884), .C(n_894), .Y(n_839) );
NOR2xp33_ASAP7_75t_L g840 ( .A(n_841), .B(n_867), .Y(n_840) );
OAI33xp33_ASAP7_75t_L g841 ( .A1(n_842), .A2(n_844), .A3(n_850), .B1(n_856), .B2(n_861), .B3(n_866), .Y(n_841) );
OAI33xp33_ASAP7_75t_L g924 ( .A1(n_842), .A2(n_866), .A3(n_925), .B1(n_928), .B2(n_929), .B3(n_933), .Y(n_924) );
OAI22xp33_ASAP7_75t_L g844 ( .A1(n_845), .A2(n_846), .B1(n_847), .B2(n_849), .Y(n_844) );
OAI221xp5_ASAP7_75t_L g868 ( .A1(n_846), .A2(n_849), .B1(n_869), .B2(n_871), .C(n_875), .Y(n_868) );
OAI22xp33_ASAP7_75t_L g925 ( .A1(n_847), .A2(n_910), .B1(n_913), .B2(n_926), .Y(n_925) );
BUFx6f_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
OAI22xp33_ASAP7_75t_SL g850 ( .A1(n_851), .A2(n_852), .B1(n_854), .B2(n_855), .Y(n_850) );
OAI22xp5_ASAP7_75t_L g856 ( .A1(n_852), .A2(n_857), .B1(n_858), .B2(n_860), .Y(n_856) );
OAI22xp33_ASAP7_75t_L g928 ( .A1(n_852), .A2(n_858), .B1(n_905), .B2(n_907), .Y(n_928) );
INVx2_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g930 ( .A(n_853), .Y(n_930) );
OAI22xp33_ASAP7_75t_L g929 ( .A1(n_858), .A2(n_930), .B1(n_931), .B2(n_932), .Y(n_929) );
INVx2_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
OAI22xp33_ASAP7_75t_L g861 ( .A1(n_862), .A2(n_863), .B1(n_864), .B2(n_865), .Y(n_861) );
INVx2_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
INVx2_ASAP7_75t_L g878 ( .A(n_870), .Y(n_878) );
INVx2_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
INVx1_ASAP7_75t_L g872 ( .A(n_873), .Y(n_872) );
INVx1_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
BUFx2_ASAP7_75t_L g881 ( .A(n_874), .Y(n_881) );
BUFx4f_ASAP7_75t_L g915 ( .A(n_874), .Y(n_915) );
INVx1_ASAP7_75t_L g960 ( .A(n_874), .Y(n_960) );
OAI221xp5_ASAP7_75t_L g877 ( .A1(n_878), .A2(n_879), .B1(n_880), .B2(n_882), .C(n_883), .Y(n_877) );
INVx2_ASAP7_75t_SL g880 ( .A(n_881), .Y(n_880) );
INVx1_ASAP7_75t_L g950 ( .A(n_899), .Y(n_950) );
NAND3xp33_ASAP7_75t_L g900 ( .A(n_901), .B(n_937), .C(n_944), .Y(n_900) );
NOR2xp33_ASAP7_75t_L g901 ( .A(n_902), .B(n_924), .Y(n_901) );
OAI33xp33_ASAP7_75t_L g902 ( .A1(n_903), .A2(n_904), .A3(n_909), .B1(n_916), .B2(n_919), .B3(n_923), .Y(n_902) );
OAI22xp5_ASAP7_75t_L g904 ( .A1(n_905), .A2(n_906), .B1(n_907), .B2(n_908), .Y(n_904) );
OAI22xp5_ASAP7_75t_L g909 ( .A1(n_910), .A2(n_911), .B1(n_913), .B2(n_914), .Y(n_909) );
OAI22xp5_ASAP7_75t_L g916 ( .A1(n_911), .A2(n_914), .B1(n_917), .B2(n_918), .Y(n_916) );
INVx2_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
INVx2_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
OAI22xp33_ASAP7_75t_L g933 ( .A1(n_926), .A2(n_934), .B1(n_935), .B2(n_936), .Y(n_933) );
INVx2_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
INVx2_ASAP7_75t_L g951 ( .A(n_952), .Y(n_951) );
INVx1_ASAP7_75t_L g953 ( .A(n_954), .Y(n_953) );
NAND3xp33_ASAP7_75t_L g955 ( .A(n_956), .B(n_961), .C(n_964), .Y(n_955) );
INVx1_ASAP7_75t_L g958 ( .A(n_959), .Y(n_958) );
INVx1_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
NAND2xp5_ASAP7_75t_L g980 ( .A(n_981), .B(n_989), .Y(n_980) );
BUFx2_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
INVx1_ASAP7_75t_L g997 ( .A(n_998), .Y(n_997) );
INVx1_ASAP7_75t_L g998 ( .A(n_999), .Y(n_998) );
INVx1_ASAP7_75t_L g1001 ( .A(n_1002), .Y(n_1001) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1002), .Y(n_1262) );
OAI21xp5_ASAP7_75t_L g1004 ( .A1(n_1005), .A2(n_1013), .B(n_1214), .Y(n_1004) );
INVx1_ASAP7_75t_L g1005 ( .A(n_1006), .Y(n_1005) );
BUFx3_ASAP7_75t_L g1006 ( .A(n_1007), .Y(n_1006) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1007), .Y(n_1177) );
AND2x4_ASAP7_75t_L g1007 ( .A(n_1008), .B(n_1011), .Y(n_1007) );
AND2x2_ASAP7_75t_L g1064 ( .A(n_1008), .B(n_1011), .Y(n_1064) );
HB1xp67_ASAP7_75t_L g1315 ( .A(n_1008), .Y(n_1315) );
INVx1_ASAP7_75t_L g1008 ( .A(n_1009), .Y(n_1008) );
AND2x4_ASAP7_75t_L g1031 ( .A(n_1009), .B(n_1011), .Y(n_1031) );
INVx1_ASAP7_75t_L g1009 ( .A(n_1010), .Y(n_1009) );
NAND2xp5_ASAP7_75t_L g1023 ( .A(n_1010), .B(n_1024), .Y(n_1023) );
INVx1_ASAP7_75t_L g1024 ( .A(n_1012), .Y(n_1024) );
AND2x2_ASAP7_75t_L g1013 ( .A(n_1014), .B(n_1141), .Y(n_1013) );
NOR2xp33_ASAP7_75t_L g1014 ( .A(n_1015), .B(n_1123), .Y(n_1014) );
NAND3xp33_ASAP7_75t_L g1015 ( .A(n_1016), .B(n_1080), .C(n_1109), .Y(n_1015) );
O2A1O1Ixp33_ASAP7_75t_L g1016 ( .A1(n_1017), .A2(n_1047), .B(n_1052), .C(n_1066), .Y(n_1016) );
AND2x2_ASAP7_75t_L g1017 ( .A(n_1018), .B(n_1032), .Y(n_1017) );
AND2x2_ASAP7_75t_L g1068 ( .A(n_1018), .B(n_1069), .Y(n_1068) );
AND2x2_ASAP7_75t_L g1089 ( .A(n_1018), .B(n_1090), .Y(n_1089) );
NOR2xp33_ASAP7_75t_L g1107 ( .A(n_1018), .B(n_1053), .Y(n_1107) );
AND2x2_ASAP7_75t_L g1112 ( .A(n_1018), .B(n_1033), .Y(n_1112) );
AND2x2_ASAP7_75t_L g1122 ( .A(n_1018), .B(n_1108), .Y(n_1122) );
OAI332xp33_ASAP7_75t_L g1145 ( .A1(n_1018), .A2(n_1077), .A3(n_1096), .B1(n_1097), .B2(n_1146), .B3(n_1149), .C1(n_1150), .C2(n_1152), .Y(n_1145) );
OAI32xp33_ASAP7_75t_L g1207 ( .A1(n_1018), .A2(n_1138), .A3(n_1163), .B1(n_1193), .B2(n_1208), .Y(n_1207) );
INVx1_ASAP7_75t_L g1209 ( .A(n_1018), .Y(n_1209) );
INVx4_ASAP7_75t_L g1018 ( .A(n_1019), .Y(n_1018) );
NAND2xp5_ASAP7_75t_L g1049 ( .A(n_1019), .B(n_1050), .Y(n_1049) );
NAND2xp5_ASAP7_75t_L g1077 ( .A(n_1019), .B(n_1069), .Y(n_1077) );
INVx3_ASAP7_75t_L g1095 ( .A(n_1019), .Y(n_1095) );
AND2x2_ASAP7_75t_L g1103 ( .A(n_1019), .B(n_1097), .Y(n_1103) );
AND2x2_ASAP7_75t_L g1132 ( .A(n_1019), .B(n_1117), .Y(n_1132) );
OR2x2_ASAP7_75t_L g1161 ( .A(n_1019), .B(n_1069), .Y(n_1161) );
NOR2xp33_ASAP7_75t_L g1204 ( .A(n_1019), .B(n_1148), .Y(n_1204) );
NAND3xp33_ASAP7_75t_L g1211 ( .A(n_1019), .B(n_1194), .C(n_1205), .Y(n_1211) );
NOR3xp33_ASAP7_75t_L g1212 ( .A(n_1019), .B(n_1091), .C(n_1213), .Y(n_1212) );
AND2x4_ASAP7_75t_L g1019 ( .A(n_1020), .B(n_1030), .Y(n_1019) );
AND2x4_ASAP7_75t_L g1021 ( .A(n_1022), .B(n_1025), .Y(n_1021) );
INVx1_ASAP7_75t_L g1022 ( .A(n_1023), .Y(n_1022) );
OR2x2_ASAP7_75t_L g1042 ( .A(n_1023), .B(n_1026), .Y(n_1042) );
HB1xp67_ASAP7_75t_L g1314 ( .A(n_1024), .Y(n_1314) );
AND2x4_ASAP7_75t_L g1027 ( .A(n_1025), .B(n_1028), .Y(n_1027) );
INVx1_ASAP7_75t_L g1025 ( .A(n_1026), .Y(n_1025) );
OR2x2_ASAP7_75t_L g1043 ( .A(n_1026), .B(n_1029), .Y(n_1043) );
INVx1_ASAP7_75t_L g1028 ( .A(n_1029), .Y(n_1028) );
INVx2_ASAP7_75t_L g1056 ( .A(n_1031), .Y(n_1056) );
OAI21xp5_ASAP7_75t_L g1074 ( .A1(n_1032), .A2(n_1075), .B(n_1076), .Y(n_1074) );
INVx1_ASAP7_75t_L g1131 ( .A(n_1032), .Y(n_1131) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1032), .B(n_1094), .Y(n_1166) );
AOI221xp5_ASAP7_75t_L g1202 ( .A1(n_1032), .A2(n_1100), .B1(n_1196), .B2(n_1203), .C(n_1204), .Y(n_1202) );
AND2x2_ASAP7_75t_L g1032 ( .A(n_1033), .B(n_1037), .Y(n_1032) );
AND2x2_ASAP7_75t_L g1047 ( .A(n_1033), .B(n_1048), .Y(n_1047) );
NOR2x1_ASAP7_75t_L g1090 ( .A(n_1033), .B(n_1091), .Y(n_1090) );
NAND2xp5_ASAP7_75t_L g1105 ( .A(n_1033), .B(n_1091), .Y(n_1105) );
NAND2xp5_ASAP7_75t_L g1126 ( .A(n_1033), .B(n_1116), .Y(n_1126) );
AND2x2_ASAP7_75t_L g1151 ( .A(n_1033), .B(n_1086), .Y(n_1151) );
OR2x2_ASAP7_75t_L g1154 ( .A(n_1033), .B(n_1155), .Y(n_1154) );
INVx2_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
AND2x2_ASAP7_75t_L g1073 ( .A(n_1034), .B(n_1037), .Y(n_1073) );
AND2x2_ASAP7_75t_L g1075 ( .A(n_1034), .B(n_1050), .Y(n_1075) );
AND2x2_ASAP7_75t_L g1084 ( .A(n_1034), .B(n_1085), .Y(n_1084) );
BUFx3_ASAP7_75t_L g1097 ( .A(n_1034), .Y(n_1097) );
AND2x2_ASAP7_75t_L g1121 ( .A(n_1034), .B(n_1091), .Y(n_1121) );
AND2x2_ASAP7_75t_L g1130 ( .A(n_1034), .B(n_1116), .Y(n_1130) );
OR2x2_ASAP7_75t_L g1191 ( .A(n_1034), .B(n_1192), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1034 ( .A(n_1035), .B(n_1036), .Y(n_1034) );
AND2x2_ASAP7_75t_L g1102 ( .A(n_1037), .B(n_1103), .Y(n_1102) );
INVx1_ASAP7_75t_L g1148 ( .A(n_1037), .Y(n_1148) );
OAI21xp5_ASAP7_75t_L g1195 ( .A1(n_1037), .A2(n_1151), .B(n_1196), .Y(n_1195) );
AND2x2_ASAP7_75t_L g1037 ( .A(n_1038), .B(n_1044), .Y(n_1037) );
AND2x2_ASAP7_75t_L g1050 ( .A(n_1038), .B(n_1051), .Y(n_1050) );
INVx2_ASAP7_75t_L g1086 ( .A(n_1038), .Y(n_1086) );
OAI22xp33_ASAP7_75t_L g1057 ( .A1(n_1041), .A2(n_1058), .B1(n_1059), .B2(n_1060), .Y(n_1057) );
BUFx3_ASAP7_75t_L g1180 ( .A(n_1041), .Y(n_1180) );
BUFx6f_ASAP7_75t_L g1041 ( .A(n_1042), .Y(n_1041) );
HB1xp67_ASAP7_75t_L g1060 ( .A(n_1043), .Y(n_1060) );
INVx1_ASAP7_75t_L g1183 ( .A(n_1043), .Y(n_1183) );
INVx1_ASAP7_75t_L g1051 ( .A(n_1044), .Y(n_1051) );
AND2x2_ASAP7_75t_L g1085 ( .A(n_1044), .B(n_1086), .Y(n_1085) );
INVx1_ASAP7_75t_L g1091 ( .A(n_1044), .Y(n_1091) );
AOI221xp5_ASAP7_75t_L g1127 ( .A1(n_1047), .A2(n_1108), .B1(n_1128), .B2(n_1132), .C(n_1133), .Y(n_1127) );
INVx1_ASAP7_75t_L g1048 ( .A(n_1049), .Y(n_1048) );
INVx1_ASAP7_75t_L g1192 ( .A(n_1050), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1116 ( .A(n_1051), .B(n_1086), .Y(n_1116) );
NAND3xp33_ASAP7_75t_L g1101 ( .A(n_1052), .B(n_1099), .C(n_1102), .Y(n_1101) );
NAND2xp5_ASAP7_75t_L g1170 ( .A(n_1052), .B(n_1100), .Y(n_1170) );
AND2x4_ASAP7_75t_SL g1052 ( .A(n_1053), .B(n_1061), .Y(n_1052) );
AND2x2_ASAP7_75t_L g1082 ( .A(n_1053), .B(n_1062), .Y(n_1082) );
OR2x2_ASAP7_75t_L g1138 ( .A(n_1053), .B(n_1061), .Y(n_1138) );
INVx2_ASAP7_75t_SL g1053 ( .A(n_1054), .Y(n_1053) );
AND2x2_ASAP7_75t_L g1079 ( .A(n_1054), .B(n_1061), .Y(n_1079) );
OR2x2_ASAP7_75t_L g1098 ( .A(n_1054), .B(n_1099), .Y(n_1098) );
INVx2_ASAP7_75t_L g1135 ( .A(n_1054), .Y(n_1135) );
INVx2_ASAP7_75t_L g1055 ( .A(n_1056), .Y(n_1055) );
AND2x2_ASAP7_75t_L g1113 ( .A(n_1061), .B(n_1100), .Y(n_1113) );
AND2x2_ASAP7_75t_L g1194 ( .A(n_1061), .B(n_1069), .Y(n_1194) );
CKINVDCx6p67_ASAP7_75t_R g1061 ( .A(n_1062), .Y(n_1061) );
AND2x2_ASAP7_75t_L g1108 ( .A(n_1062), .B(n_1069), .Y(n_1108) );
AND2x2_ASAP7_75t_L g1117 ( .A(n_1062), .B(n_1118), .Y(n_1117) );
CKINVDCx5p33_ASAP7_75t_R g1152 ( .A(n_1062), .Y(n_1152) );
OR2x6_ASAP7_75t_L g1062 ( .A(n_1063), .B(n_1065), .Y(n_1062) );
O2A1O1Ixp33_ASAP7_75t_L g1066 ( .A1(n_1067), .A2(n_1072), .B(n_1074), .C(n_1078), .Y(n_1066) );
INVx1_ASAP7_75t_L g1067 ( .A(n_1068), .Y(n_1067) );
AND2x2_ASAP7_75t_L g1157 ( .A(n_1068), .B(n_1116), .Y(n_1157) );
INVx1_ASAP7_75t_L g1083 ( .A(n_1069), .Y(n_1083) );
CKINVDCx5p33_ASAP7_75t_R g1100 ( .A(n_1069), .Y(n_1100) );
INVx1_ASAP7_75t_SL g1118 ( .A(n_1069), .Y(n_1118) );
AND2x2_ASAP7_75t_L g1069 ( .A(n_1070), .B(n_1071), .Y(n_1069) );
AOI21xp33_ASAP7_75t_SL g1104 ( .A1(n_1072), .A2(n_1105), .B(n_1106), .Y(n_1104) );
NOR2xp33_ASAP7_75t_L g1189 ( .A(n_1072), .B(n_1100), .Y(n_1189) );
INVx1_ASAP7_75t_L g1072 ( .A(n_1073), .Y(n_1072) );
AOI21xp5_ASAP7_75t_L g1167 ( .A1(n_1073), .A2(n_1168), .B(n_1169), .Y(n_1167) );
NAND2xp5_ASAP7_75t_L g1188 ( .A(n_1073), .B(n_1144), .Y(n_1188) );
AND2x2_ASAP7_75t_L g1133 ( .A(n_1075), .B(n_1134), .Y(n_1133) );
INVx1_ASAP7_75t_L g1076 ( .A(n_1077), .Y(n_1076) );
INVx1_ASAP7_75t_L g1078 ( .A(n_1079), .Y(n_1078) );
NAND2xp5_ASAP7_75t_L g1124 ( .A(n_1079), .B(n_1118), .Y(n_1124) );
NAND2xp5_ASAP7_75t_L g1156 ( .A(n_1079), .B(n_1157), .Y(n_1156) );
NAND2xp5_ASAP7_75t_L g1187 ( .A(n_1079), .B(n_1095), .Y(n_1187) );
AOI211xp5_ASAP7_75t_SL g1080 ( .A1(n_1081), .A2(n_1084), .B(n_1087), .C(n_1104), .Y(n_1080) );
AND2x2_ASAP7_75t_L g1081 ( .A(n_1082), .B(n_1083), .Y(n_1081) );
INVx2_ASAP7_75t_L g1092 ( .A(n_1082), .Y(n_1092) );
NAND3xp33_ASAP7_75t_L g1208 ( .A(n_1083), .B(n_1203), .C(n_1209), .Y(n_1208) );
NAND2xp5_ASAP7_75t_L g1111 ( .A(n_1085), .B(n_1112), .Y(n_1111) );
NAND2xp5_ASAP7_75t_L g1155 ( .A(n_1085), .B(n_1095), .Y(n_1155) );
INVx1_ASAP7_75t_L g1172 ( .A(n_1085), .Y(n_1172) );
INVx2_ASAP7_75t_L g1203 ( .A(n_1086), .Y(n_1203) );
OAI221xp5_ASAP7_75t_L g1087 ( .A1(n_1088), .A2(n_1092), .B1(n_1093), .B2(n_1098), .C(n_1101), .Y(n_1087) );
INVx1_ASAP7_75t_L g1088 ( .A(n_1089), .Y(n_1088) );
OR2x2_ASAP7_75t_L g1096 ( .A(n_1091), .B(n_1097), .Y(n_1096) );
AOI222xp33_ASAP7_75t_L g1206 ( .A1(n_1091), .A2(n_1113), .B1(n_1175), .B2(n_1207), .C1(n_1210), .C2(n_1212), .Y(n_1206) );
OR2x2_ASAP7_75t_L g1093 ( .A(n_1094), .B(n_1096), .Y(n_1093) );
NAND2xp5_ASAP7_75t_L g1162 ( .A(n_1094), .B(n_1113), .Y(n_1162) );
INVx2_ASAP7_75t_L g1094 ( .A(n_1095), .Y(n_1094) );
OR2x2_ASAP7_75t_L g1125 ( .A(n_1095), .B(n_1126), .Y(n_1125) );
NAND2xp5_ASAP7_75t_L g1140 ( .A(n_1095), .B(n_1130), .Y(n_1140) );
NAND2xp5_ASAP7_75t_L g1200 ( .A(n_1095), .B(n_1151), .Y(n_1200) );
OR2x2_ASAP7_75t_L g1171 ( .A(n_1097), .B(n_1172), .Y(n_1171) );
INVx1_ASAP7_75t_L g1168 ( .A(n_1098), .Y(n_1168) );
INVx3_ASAP7_75t_L g1099 ( .A(n_1100), .Y(n_1099) );
NOR2xp33_ASAP7_75t_L g1198 ( .A(n_1100), .B(n_1140), .Y(n_1198) );
NAND2xp5_ASAP7_75t_L g1106 ( .A(n_1107), .B(n_1108), .Y(n_1106) );
AND2x2_ASAP7_75t_L g1134 ( .A(n_1108), .B(n_1135), .Y(n_1134) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1108), .Y(n_1149) );
AOI221xp5_ASAP7_75t_L g1109 ( .A1(n_1110), .A2(n_1113), .B1(n_1114), .B2(n_1117), .C(n_1119), .Y(n_1109) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1111), .Y(n_1110) );
NAND2xp5_ASAP7_75t_L g1115 ( .A(n_1112), .B(n_1116), .Y(n_1115) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1115), .Y(n_1114) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1116), .Y(n_1147) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1117), .Y(n_1201) );
INVxp67_ASAP7_75t_SL g1119 ( .A(n_1120), .Y(n_1119) );
NAND2xp5_ASAP7_75t_L g1120 ( .A(n_1121), .B(n_1122), .Y(n_1120) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1121), .Y(n_1163) );
OAI211xp5_ASAP7_75t_L g1123 ( .A1(n_1124), .A2(n_1125), .B(n_1127), .C(n_1136), .Y(n_1123) );
OAI221xp5_ASAP7_75t_L g1186 ( .A1(n_1124), .A2(n_1150), .B1(n_1171), .B2(n_1187), .C(n_1188), .Y(n_1186) );
NAND2xp5_ASAP7_75t_L g1128 ( .A(n_1129), .B(n_1131), .Y(n_1128) );
OAI221xp5_ASAP7_75t_L g1153 ( .A1(n_1129), .A2(n_1138), .B1(n_1152), .B2(n_1154), .C(n_1156), .Y(n_1153) );
INVx1_ASAP7_75t_L g1129 ( .A(n_1130), .Y(n_1129) );
INVx2_ASAP7_75t_L g1144 ( .A(n_1135), .Y(n_1144) );
NOR2xp33_ASAP7_75t_L g1160 ( .A(n_1135), .B(n_1161), .Y(n_1160) );
INVx2_ASAP7_75t_L g1165 ( .A(n_1135), .Y(n_1165) );
OAI31xp33_ASAP7_75t_L g1190 ( .A1(n_1135), .A2(n_1191), .A3(n_1193), .B(n_1195), .Y(n_1190) );
AND2x2_ASAP7_75t_L g1205 ( .A(n_1135), .B(n_1175), .Y(n_1205) );
NAND2xp5_ASAP7_75t_L g1136 ( .A(n_1137), .B(n_1139), .Y(n_1136) );
INVx1_ASAP7_75t_L g1137 ( .A(n_1138), .Y(n_1137) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1140), .Y(n_1139) );
AOI21xp5_ASAP7_75t_L g1141 ( .A1(n_1142), .A2(n_1173), .B(n_1184), .Y(n_1141) );
NAND3xp33_ASAP7_75t_L g1142 ( .A(n_1143), .B(n_1164), .C(n_1167), .Y(n_1142) );
AOI211xp5_ASAP7_75t_L g1143 ( .A1(n_1144), .A2(n_1145), .B(n_1153), .C(n_1158), .Y(n_1143) );
NAND2xp5_ASAP7_75t_L g1146 ( .A(n_1147), .B(n_1148), .Y(n_1146) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
OAI221xp5_ASAP7_75t_SL g1199 ( .A1(n_1152), .A2(n_1172), .B1(n_1200), .B2(n_1201), .C(n_1202), .Y(n_1199) );
AOI21xp33_ASAP7_75t_SL g1158 ( .A1(n_1159), .A2(n_1162), .B(n_1163), .Y(n_1158) );
INVx1_ASAP7_75t_L g1159 ( .A(n_1160), .Y(n_1159) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1161), .Y(n_1196) );
NAND2xp5_ASAP7_75t_L g1164 ( .A(n_1165), .B(n_1166), .Y(n_1164) );
NOR2xp33_ASAP7_75t_L g1169 ( .A(n_1170), .B(n_1171), .Y(n_1169) );
INVx2_ASAP7_75t_L g1173 ( .A(n_1174), .Y(n_1173) );
OAI31xp33_ASAP7_75t_L g1185 ( .A1(n_1174), .A2(n_1186), .A3(n_1189), .B(n_1190), .Y(n_1185) );
BUFx3_ASAP7_75t_L g1174 ( .A(n_1175), .Y(n_1174) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1175), .Y(n_1213) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1177), .Y(n_1176) );
OAI22xp33_ASAP7_75t_L g1178 ( .A1(n_1179), .A2(n_1180), .B1(n_1181), .B2(n_1182), .Y(n_1178) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1183), .Y(n_1182) );
NAND3xp33_ASAP7_75t_L g1184 ( .A(n_1185), .B(n_1197), .C(n_1206), .Y(n_1184) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1194), .Y(n_1193) );
OAI21xp33_ASAP7_75t_L g1197 ( .A1(n_1198), .A2(n_1199), .B(n_1205), .Y(n_1197) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1211), .Y(n_1210) );
INVx1_ASAP7_75t_L g1269 ( .A(n_1217), .Y(n_1269) );
AOI211x1_ASAP7_75t_L g1217 ( .A1(n_1218), .A2(n_1229), .B(n_1231), .C(n_1259), .Y(n_1217) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1230), .Y(n_1229) );
NAND2xp5_ASAP7_75t_L g1231 ( .A(n_1232), .B(n_1244), .Y(n_1231) );
INVx1_ASAP7_75t_L g1239 ( .A(n_1240), .Y(n_1239) );
INVx2_ASAP7_75t_SL g1242 ( .A(n_1243), .Y(n_1242) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1248), .Y(n_1247) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1254), .Y(n_1253) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1258), .Y(n_1257) );
BUFx2_ASAP7_75t_L g1270 ( .A(n_1271), .Y(n_1270) );
INVx1_ASAP7_75t_L g1273 ( .A(n_1274), .Y(n_1273) );
HB1xp67_ASAP7_75t_L g1274 ( .A(n_1275), .Y(n_1274) );
NAND3xp33_ASAP7_75t_L g1287 ( .A(n_1288), .B(n_1290), .C(n_1292), .Y(n_1287) );
NAND4xp25_ASAP7_75t_L g1295 ( .A(n_1296), .B(n_1299), .C(n_1302), .D(n_1306), .Y(n_1295) );
A2O1A1Ixp33_ASAP7_75t_L g1312 ( .A1(n_1311), .A2(n_1313), .B(n_1315), .C(n_1316), .Y(n_1312) );
INVx1_ASAP7_75t_L g1313 ( .A(n_1314), .Y(n_1313) );
endmodule