module real_aes_6315_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_119;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_449;
wire n_754;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_741;
wire n_283;
wire n_314;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g237 ( .A1(n_0), .A2(n_238), .B(n_239), .C(n_243), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_1), .B(n_179), .Y(n_244) );
INVx1_ASAP7_75t_L g107 ( .A(n_2), .Y(n_107) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_3), .B(n_151), .Y(n_227) );
A2O1A1Ixp33_ASAP7_75t_L g503 ( .A1(n_4), .A2(n_137), .B(n_142), .C(n_504), .Y(n_503) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_5), .A2(n_132), .B(n_542), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_6), .A2(n_132), .B(n_170), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_7), .B(n_179), .Y(n_548) );
AO21x2_ASAP7_75t_L g182 ( .A1(n_8), .A2(n_167), .B(n_183), .Y(n_182) );
AND2x6_ASAP7_75t_L g137 ( .A(n_9), .B(n_138), .Y(n_137) );
A2O1A1Ixp33_ASAP7_75t_L g252 ( .A1(n_10), .A2(n_137), .B(n_142), .C(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g486 ( .A(n_11), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_12), .B(n_113), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_12), .B(n_42), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_13), .A2(n_104), .B1(n_114), .B2(n_761), .Y(n_103) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_14), .B(n_242), .Y(n_506) );
INVx1_ASAP7_75t_L g161 ( .A(n_15), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_16), .B(n_151), .Y(n_189) );
A2O1A1Ixp33_ASAP7_75t_L g493 ( .A1(n_17), .A2(n_152), .B(n_494), .C(n_496), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_18), .B(n_179), .Y(n_497) );
AOI222xp33_ASAP7_75t_L g467 ( .A1(n_19), .A2(n_468), .B1(n_745), .B2(n_751), .C1(n_754), .C2(n_755), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_20), .B(n_216), .Y(n_585) );
A2O1A1Ixp33_ASAP7_75t_L g211 ( .A1(n_21), .A2(n_142), .B(n_193), .C(n_212), .Y(n_211) );
A2O1A1Ixp33_ASAP7_75t_L g515 ( .A1(n_22), .A2(n_191), .B(n_241), .C(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_23), .B(n_242), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_24), .B(n_242), .Y(n_526) );
CKINVDCx16_ASAP7_75t_R g533 ( .A(n_25), .Y(n_533) );
INVx1_ASAP7_75t_L g525 ( .A(n_26), .Y(n_525) );
A2O1A1Ixp33_ASAP7_75t_L g185 ( .A1(n_27), .A2(n_142), .B(n_186), .C(n_193), .Y(n_185) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_28), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_29), .Y(n_502) );
INVx1_ASAP7_75t_L g582 ( .A(n_30), .Y(n_582) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_31), .A2(n_132), .B(n_235), .Y(n_234) );
INVx2_ASAP7_75t_L g135 ( .A(n_32), .Y(n_135) );
A2O1A1Ixp33_ASAP7_75t_L g200 ( .A1(n_33), .A2(n_140), .B(n_155), .C(n_201), .Y(n_200) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_34), .Y(n_509) );
A2O1A1Ixp33_ASAP7_75t_L g544 ( .A1(n_35), .A2(n_241), .B(n_545), .C(n_547), .Y(n_544) );
INVxp67_ASAP7_75t_L g583 ( .A(n_36), .Y(n_583) );
OAI22xp5_ASAP7_75t_SL g122 ( .A1(n_37), .A2(n_47), .B1(n_123), .B2(n_124), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_37), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_38), .B(n_188), .Y(n_187) );
A2O1A1Ixp33_ASAP7_75t_L g523 ( .A1(n_39), .A2(n_142), .B(n_193), .C(n_524), .Y(n_523) );
CKINVDCx14_ASAP7_75t_R g543 ( .A(n_40), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g748 ( .A1(n_41), .A2(n_46), .B1(n_749), .B2(n_750), .Y(n_748) );
INVx1_ASAP7_75t_L g750 ( .A(n_41), .Y(n_750) );
INVx1_ASAP7_75t_L g113 ( .A(n_42), .Y(n_113) );
A2O1A1Ixp33_ASAP7_75t_L g483 ( .A1(n_43), .A2(n_243), .B(n_484), .C(n_485), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_44), .B(n_210), .Y(n_209) );
CKINVDCx20_ASAP7_75t_R g257 ( .A(n_45), .Y(n_257) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_46), .Y(n_749) );
INVx1_ASAP7_75t_L g124 ( .A(n_47), .Y(n_124) );
OAI321xp33_ASAP7_75t_L g120 ( .A1(n_48), .A2(n_121), .A3(n_455), .B1(n_461), .B2(n_462), .C(n_464), .Y(n_120) );
INVx1_ASAP7_75t_L g461 ( .A(n_48), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_49), .B(n_151), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_50), .B(n_132), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g528 ( .A(n_51), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g579 ( .A(n_52), .Y(n_579) );
A2O1A1Ixp33_ASAP7_75t_L g139 ( .A1(n_53), .A2(n_140), .B(n_145), .C(n_155), .Y(n_139) );
INVx1_ASAP7_75t_L g240 ( .A(n_54), .Y(n_240) );
INVx1_ASAP7_75t_L g146 ( .A(n_55), .Y(n_146) );
INVx1_ASAP7_75t_L g514 ( .A(n_56), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_57), .B(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_58), .B(n_132), .Y(n_131) );
CKINVDCx20_ASAP7_75t_R g219 ( .A(n_59), .Y(n_219) );
CKINVDCx14_ASAP7_75t_R g482 ( .A(n_60), .Y(n_482) );
INVx1_ASAP7_75t_L g138 ( .A(n_61), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_62), .B(n_132), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_63), .B(n_179), .Y(n_178) );
A2O1A1Ixp33_ASAP7_75t_L g172 ( .A1(n_64), .A2(n_173), .B(n_175), .C(n_177), .Y(n_172) );
INVx1_ASAP7_75t_L g160 ( .A(n_65), .Y(n_160) );
INVx1_ASAP7_75t_SL g546 ( .A(n_66), .Y(n_546) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_67), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_68), .B(n_151), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_69), .B(n_179), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_70), .B(n_152), .Y(n_254) );
INVx1_ASAP7_75t_L g536 ( .A(n_71), .Y(n_536) );
CKINVDCx16_ASAP7_75t_R g236 ( .A(n_72), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_73), .B(n_148), .Y(n_213) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_74), .A2(n_142), .B(n_155), .C(n_225), .Y(n_224) );
CKINVDCx16_ASAP7_75t_R g171 ( .A(n_75), .Y(n_171) );
INVx1_ASAP7_75t_L g111 ( .A(n_76), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_77), .A2(n_132), .B(n_481), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_78), .Y(n_539) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_79), .A2(n_132), .B(n_491), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_80), .A2(n_210), .B(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g492 ( .A(n_81), .Y(n_492) );
CKINVDCx16_ASAP7_75t_R g522 ( .A(n_82), .Y(n_522) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_83), .B(n_147), .Y(n_214) );
AOI22xp5_ASAP7_75t_L g745 ( .A1(n_84), .A2(n_746), .B1(n_747), .B2(n_748), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_84), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g205 ( .A(n_85), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_86), .A2(n_132), .B(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g495 ( .A(n_87), .Y(n_495) );
INVx2_ASAP7_75t_L g158 ( .A(n_88), .Y(n_158) );
INVx1_ASAP7_75t_L g505 ( .A(n_89), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g232 ( .A(n_90), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_91), .B(n_242), .Y(n_255) );
INVx2_ASAP7_75t_L g108 ( .A(n_92), .Y(n_108) );
OR2x2_ASAP7_75t_L g457 ( .A(n_92), .B(n_458), .Y(n_457) );
OR2x2_ASAP7_75t_L g744 ( .A(n_92), .B(n_459), .Y(n_744) );
A2O1A1Ixp33_ASAP7_75t_L g534 ( .A1(n_93), .A2(n_142), .B(n_155), .C(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_94), .B(n_132), .Y(n_199) );
INVx1_ASAP7_75t_L g202 ( .A(n_95), .Y(n_202) );
INVxp67_ASAP7_75t_L g176 ( .A(n_96), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_97), .B(n_167), .Y(n_487) );
INVx2_ASAP7_75t_L g517 ( .A(n_98), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_99), .B(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g226 ( .A(n_100), .Y(n_226) );
INVx1_ASAP7_75t_L g250 ( .A(n_101), .Y(n_250) );
AND2x2_ASAP7_75t_L g162 ( .A(n_102), .B(n_157), .Y(n_162) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g762 ( .A(n_105), .Y(n_762) );
OR2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_112), .Y(n_105) );
NAND3xp33_ASAP7_75t_SL g106 ( .A(n_107), .B(n_108), .C(n_109), .Y(n_106) );
AND2x2_ASAP7_75t_L g459 ( .A(n_107), .B(n_460), .Y(n_459) );
OR2x2_ASAP7_75t_L g473 ( .A(n_108), .B(n_459), .Y(n_473) );
NOR2x2_ASAP7_75t_L g753 ( .A(n_108), .B(n_458), .Y(n_753) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
OA21x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_120), .B(n_466), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
BUFx3_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_SL g760 ( .A(n_118), .Y(n_760) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_121), .B(n_463), .Y(n_462) );
XOR2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_125), .Y(n_121) );
AOI22xp5_ASAP7_75t_L g469 ( .A1(n_125), .A2(n_470), .B1(n_474), .B2(n_741), .Y(n_469) );
INVx4_ASAP7_75t_L g758 ( .A(n_125), .Y(n_758) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
OR5x1_ASAP7_75t_L g126 ( .A(n_127), .B(n_328), .C(n_406), .D(n_430), .E(n_447), .Y(n_126) );
OAI211xp5_ASAP7_75t_SL g127 ( .A1(n_128), .A2(n_194), .B(n_245), .C(n_305), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_129), .B(n_163), .Y(n_128) );
AND2x2_ASAP7_75t_L g259 ( .A(n_129), .B(n_165), .Y(n_259) );
INVx5_ASAP7_75t_SL g287 ( .A(n_129), .Y(n_287) );
AND2x2_ASAP7_75t_L g323 ( .A(n_129), .B(n_308), .Y(n_323) );
OR2x2_ASAP7_75t_L g362 ( .A(n_129), .B(n_164), .Y(n_362) );
OR2x2_ASAP7_75t_L g393 ( .A(n_129), .B(n_284), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_129), .B(n_297), .Y(n_429) );
AND2x2_ASAP7_75t_L g441 ( .A(n_129), .B(n_284), .Y(n_441) );
OR2x6_ASAP7_75t_L g129 ( .A(n_130), .B(n_162), .Y(n_129) );
AOI21xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_139), .B(n_157), .Y(n_130) );
BUFx2_ASAP7_75t_L g210 ( .A(n_132), .Y(n_210) );
AND2x4_ASAP7_75t_L g132 ( .A(n_133), .B(n_137), .Y(n_132) );
NAND2x1p5_ASAP7_75t_L g251 ( .A(n_133), .B(n_137), .Y(n_251) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_136), .Y(n_133) );
INVx1_ASAP7_75t_L g177 ( .A(n_134), .Y(n_177) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g143 ( .A(n_135), .Y(n_143) );
INVx1_ASAP7_75t_L g192 ( .A(n_135), .Y(n_192) );
INVx1_ASAP7_75t_L g144 ( .A(n_136), .Y(n_144) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_136), .Y(n_149) );
INVx3_ASAP7_75t_L g152 ( .A(n_136), .Y(n_152) );
INVx1_ASAP7_75t_L g188 ( .A(n_136), .Y(n_188) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_136), .Y(n_242) );
INVx4_ASAP7_75t_SL g156 ( .A(n_137), .Y(n_156) );
BUFx3_ASAP7_75t_L g193 ( .A(n_137), .Y(n_193) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
O2A1O1Ixp33_ASAP7_75t_L g170 ( .A1(n_141), .A2(n_156), .B(n_171), .C(n_172), .Y(n_170) );
O2A1O1Ixp33_ASAP7_75t_SL g235 ( .A1(n_141), .A2(n_156), .B(n_236), .C(n_237), .Y(n_235) );
O2A1O1Ixp33_ASAP7_75t_SL g481 ( .A1(n_141), .A2(n_156), .B(n_482), .C(n_483), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_SL g491 ( .A1(n_141), .A2(n_156), .B(n_492), .C(n_493), .Y(n_491) );
O2A1O1Ixp33_ASAP7_75t_SL g513 ( .A1(n_141), .A2(n_156), .B(n_514), .C(n_515), .Y(n_513) );
O2A1O1Ixp33_ASAP7_75t_L g542 ( .A1(n_141), .A2(n_156), .B(n_543), .C(n_544), .Y(n_542) );
O2A1O1Ixp33_ASAP7_75t_SL g578 ( .A1(n_141), .A2(n_156), .B(n_579), .C(n_580), .Y(n_578) );
INVx5_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x6_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
BUFx3_ASAP7_75t_L g154 ( .A(n_143), .Y(n_154) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_143), .Y(n_229) );
O2A1O1Ixp33_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_147), .B(n_150), .C(n_153), .Y(n_145) );
O2A1O1Ixp33_ASAP7_75t_L g201 ( .A1(n_147), .A2(n_153), .B(n_202), .C(n_203), .Y(n_201) );
O2A1O1Ixp5_ASAP7_75t_L g504 ( .A1(n_147), .A2(n_505), .B(n_506), .C(n_507), .Y(n_504) );
O2A1O1Ixp33_ASAP7_75t_L g535 ( .A1(n_147), .A2(n_507), .B(n_536), .C(n_537), .Y(n_535) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx4_ASAP7_75t_L g174 ( .A(n_149), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_151), .B(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g238 ( .A(n_151), .Y(n_238) );
O2A1O1Ixp33_ASAP7_75t_L g524 ( .A1(n_151), .A2(n_215), .B(n_525), .C(n_526), .Y(n_524) );
OAI22xp33_ASAP7_75t_L g581 ( .A1(n_151), .A2(n_174), .B1(n_582), .B2(n_583), .Y(n_581) );
INVx5_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_152), .B(n_486), .Y(n_485) );
HB1xp67_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g243 ( .A(n_154), .Y(n_243) );
INVx1_ASAP7_75t_L g496 ( .A(n_154), .Y(n_496) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_157), .A2(n_199), .B(n_200), .Y(n_198) );
INVx2_ASAP7_75t_L g217 ( .A(n_157), .Y(n_217) );
INVx1_ASAP7_75t_L g220 ( .A(n_157), .Y(n_220) );
OA21x2_ASAP7_75t_L g479 ( .A1(n_157), .A2(n_480), .B(n_487), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_L g521 ( .A1(n_157), .A2(n_251), .B(n_522), .C(n_523), .Y(n_521) );
AND2x2_ASAP7_75t_SL g157 ( .A(n_158), .B(n_159), .Y(n_157) );
AND2x2_ASAP7_75t_L g168 ( .A(n_158), .B(n_159), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_160), .B(n_161), .Y(n_159) );
AND2x2_ASAP7_75t_L g440 ( .A(n_163), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_SL g163 ( .A(n_164), .Y(n_163) );
OR2x2_ASAP7_75t_L g303 ( .A(n_164), .B(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g164 ( .A(n_165), .B(n_181), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_165), .B(n_284), .Y(n_283) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_165), .Y(n_296) );
INVx3_ASAP7_75t_L g311 ( .A(n_165), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_165), .B(n_181), .Y(n_335) );
OR2x2_ASAP7_75t_L g344 ( .A(n_165), .B(n_287), .Y(n_344) );
AND2x2_ASAP7_75t_L g348 ( .A(n_165), .B(n_308), .Y(n_348) );
AND2x2_ASAP7_75t_L g354 ( .A(n_165), .B(n_355), .Y(n_354) );
INVxp67_ASAP7_75t_L g391 ( .A(n_165), .Y(n_391) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_165), .B(n_248), .Y(n_405) );
OA21x2_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_169), .B(n_178), .Y(n_165) );
OA21x2_ASAP7_75t_L g489 ( .A1(n_166), .A2(n_490), .B(n_497), .Y(n_489) );
OA21x2_ASAP7_75t_L g511 ( .A1(n_166), .A2(n_512), .B(n_518), .Y(n_511) );
OA21x2_ASAP7_75t_L g540 ( .A1(n_166), .A2(n_541), .B(n_548), .Y(n_540) );
HB1xp67_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx4_ASAP7_75t_L g180 ( .A(n_167), .Y(n_180) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_167), .A2(n_184), .B(n_185), .Y(n_183) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g258 ( .A(n_168), .Y(n_258) );
O2A1O1Ixp33_ASAP7_75t_L g225 ( .A1(n_173), .A2(n_226), .B(n_227), .C(n_228), .Y(n_225) );
INVx1_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_174), .B(n_495), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_174), .B(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g215 ( .A(n_177), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g580 ( .A(n_177), .B(n_581), .Y(n_580) );
OA21x2_ASAP7_75t_L g233 ( .A1(n_179), .A2(n_234), .B(n_244), .Y(n_233) );
INVx3_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g204 ( .A(n_180), .B(n_205), .Y(n_204) );
AO21x2_ASAP7_75t_L g222 ( .A1(n_180), .A2(n_223), .B(n_231), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_180), .B(n_232), .Y(n_231) );
AO21x2_ASAP7_75t_L g248 ( .A1(n_180), .A2(n_249), .B(n_256), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_180), .B(n_509), .Y(n_508) );
NOR2xp33_ASAP7_75t_L g527 ( .A(n_180), .B(n_528), .Y(n_527) );
AO21x2_ASAP7_75t_L g531 ( .A1(n_180), .A2(n_532), .B(n_538), .Y(n_531) );
OR2x2_ASAP7_75t_L g297 ( .A(n_181), .B(n_248), .Y(n_297) );
AND2x2_ASAP7_75t_L g308 ( .A(n_181), .B(n_284), .Y(n_308) );
AND2x2_ASAP7_75t_L g320 ( .A(n_181), .B(n_311), .Y(n_320) );
NAND2xp5_ASAP7_75t_SL g343 ( .A(n_181), .B(n_248), .Y(n_343) );
INVx1_ASAP7_75t_SL g355 ( .A(n_181), .Y(n_355) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AND2x2_ASAP7_75t_L g247 ( .A(n_182), .B(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_182), .B(n_287), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_189), .B(n_190), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_190), .A2(n_254), .B(n_255), .Y(n_253) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx3_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
INVx1_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AND2x2_ASAP7_75t_L g195 ( .A(n_196), .B(n_206), .Y(n_195) );
AND2x2_ASAP7_75t_L g268 ( .A(n_196), .B(n_269), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_196), .B(n_221), .Y(n_272) );
AND2x2_ASAP7_75t_L g275 ( .A(n_196), .B(n_276), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_196), .B(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g300 ( .A(n_196), .B(n_291), .Y(n_300) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_196), .Y(n_319) );
AND2x2_ASAP7_75t_L g340 ( .A(n_196), .B(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g350 ( .A(n_196), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g396 ( .A(n_196), .B(n_279), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_196), .B(n_302), .Y(n_423) );
INVx5_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
BUFx2_ASAP7_75t_L g293 ( .A(n_197), .Y(n_293) );
AND2x2_ASAP7_75t_L g359 ( .A(n_197), .B(n_291), .Y(n_359) );
AND2x2_ASAP7_75t_L g443 ( .A(n_197), .B(n_311), .Y(n_443) );
OR2x6_ASAP7_75t_L g197 ( .A(n_198), .B(n_204), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_206), .B(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g432 ( .A(n_206), .Y(n_432) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_221), .Y(n_206) );
AND2x2_ASAP7_75t_L g262 ( .A(n_207), .B(n_263), .Y(n_262) );
AND2x4_ASAP7_75t_L g271 ( .A(n_207), .B(n_269), .Y(n_271) );
INVx5_ASAP7_75t_L g279 ( .A(n_207), .Y(n_279) );
AND2x2_ASAP7_75t_L g302 ( .A(n_207), .B(n_233), .Y(n_302) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_207), .Y(n_339) );
OR2x6_ASAP7_75t_L g207 ( .A(n_208), .B(n_218), .Y(n_207) );
AOI21xp5_ASAP7_75t_SL g208 ( .A1(n_209), .A2(n_211), .B(n_216), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_214), .B(n_215), .Y(n_212) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_217), .B(n_539), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_219), .B(n_220), .Y(n_218) );
AO21x2_ASAP7_75t_L g500 ( .A1(n_220), .A2(n_501), .B(n_508), .Y(n_500) );
INVx1_ASAP7_75t_L g380 ( .A(n_221), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_221), .B(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g413 ( .A(n_221), .B(n_279), .Y(n_413) );
A2O1A1Ixp33_ASAP7_75t_L g442 ( .A1(n_221), .A2(n_336), .B(n_443), .C(n_444), .Y(n_442) );
AND2x2_ASAP7_75t_L g221 ( .A(n_222), .B(n_233), .Y(n_221) );
BUFx2_ASAP7_75t_L g263 ( .A(n_222), .Y(n_263) );
INVx2_ASAP7_75t_L g267 ( .A(n_222), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_224), .B(n_230), .Y(n_223) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx3_ASAP7_75t_L g547 ( .A(n_229), .Y(n_547) );
INVx2_ASAP7_75t_L g269 ( .A(n_233), .Y(n_269) );
AND2x2_ASAP7_75t_L g276 ( .A(n_233), .B(n_267), .Y(n_276) );
AND2x2_ASAP7_75t_L g367 ( .A(n_233), .B(n_279), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g239 ( .A(n_240), .B(n_241), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_241), .B(n_546), .Y(n_545) );
INVx4_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx2_ASAP7_75t_L g484 ( .A(n_242), .Y(n_484) );
INVx2_ASAP7_75t_L g507 ( .A(n_243), .Y(n_507) );
AOI211x1_ASAP7_75t_SL g245 ( .A1(n_246), .A2(n_260), .B(n_273), .C(n_298), .Y(n_245) );
INVx1_ASAP7_75t_L g364 ( .A(n_246), .Y(n_364) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_259), .Y(n_246) );
INVx5_ASAP7_75t_SL g284 ( .A(n_248), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_248), .B(n_354), .Y(n_353) );
AOI311xp33_ASAP7_75t_L g372 ( .A1(n_248), .A2(n_373), .A3(n_375), .B(n_376), .C(n_382), .Y(n_372) );
A2O1A1Ixp33_ASAP7_75t_L g407 ( .A1(n_248), .A2(n_320), .B(n_408), .C(n_411), .Y(n_407) );
OAI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_251), .B(n_252), .Y(n_249) );
OAI21xp5_ASAP7_75t_L g501 ( .A1(n_251), .A2(n_502), .B(n_503), .Y(n_501) );
OAI21xp5_ASAP7_75t_L g532 ( .A1(n_251), .A2(n_533), .B(n_534), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
INVx2_ASAP7_75t_L g575 ( .A(n_258), .Y(n_575) );
INVxp67_ASAP7_75t_L g327 ( .A(n_259), .Y(n_327) );
NAND4xp25_ASAP7_75t_SL g260 ( .A(n_261), .B(n_264), .C(n_270), .D(n_272), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_261), .B(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g318 ( .A(n_262), .B(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_265), .B(n_268), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_265), .B(n_271), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_265), .B(n_278), .Y(n_398) );
BUFx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_266), .B(n_279), .Y(n_416) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g291 ( .A(n_267), .Y(n_291) );
INVxp67_ASAP7_75t_L g326 ( .A(n_268), .Y(n_326) );
AND2x4_ASAP7_75t_L g278 ( .A(n_269), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g352 ( .A(n_269), .B(n_291), .Y(n_352) );
INVx1_ASAP7_75t_L g379 ( .A(n_269), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_269), .B(n_366), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_270), .B(n_340), .Y(n_360) );
INVx1_ASAP7_75t_SL g270 ( .A(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_271), .B(n_293), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_271), .B(n_340), .Y(n_439) );
INVx1_ASAP7_75t_L g450 ( .A(n_272), .Y(n_450) );
A2O1A1Ixp33_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_277), .B(n_280), .C(n_288), .Y(n_273) );
INVx1_ASAP7_75t_SL g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g292 ( .A(n_276), .B(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g330 ( .A(n_276), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g312 ( .A(n_277), .Y(n_312) );
AND2x2_ASAP7_75t_L g289 ( .A(n_278), .B(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_278), .B(n_340), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_278), .B(n_359), .Y(n_383) );
OR2x2_ASAP7_75t_L g299 ( .A(n_279), .B(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g331 ( .A(n_279), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_279), .B(n_291), .Y(n_346) );
AND2x2_ASAP7_75t_L g403 ( .A(n_279), .B(n_359), .Y(n_403) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_279), .Y(n_410) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AOI221xp5_ASAP7_75t_L g414 ( .A1(n_281), .A2(n_293), .B1(n_415), .B2(n_417), .C(n_420), .Y(n_414) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_285), .Y(n_281) );
INVx1_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g304 ( .A(n_284), .B(n_287), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_284), .B(n_354), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_284), .B(n_311), .Y(n_419) );
INVx1_ASAP7_75t_SL g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g404 ( .A(n_286), .B(n_405), .Y(n_404) );
OR2x2_ASAP7_75t_L g418 ( .A(n_286), .B(n_419), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_287), .B(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g315 ( .A(n_287), .B(n_308), .Y(n_315) );
AND2x2_ASAP7_75t_L g385 ( .A(n_287), .B(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_287), .B(n_334), .Y(n_431) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_287), .B(n_435), .Y(n_434) );
OAI21xp5_ASAP7_75t_SL g288 ( .A1(n_289), .A2(n_292), .B(n_294), .Y(n_288) );
INVx2_ASAP7_75t_L g321 ( .A(n_289), .Y(n_321) );
HB1xp67_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g341 ( .A(n_291), .Y(n_341) );
OR2x2_ASAP7_75t_L g345 ( .A(n_293), .B(n_346), .Y(n_345) );
OR2x2_ASAP7_75t_L g448 ( .A(n_293), .B(n_416), .Y(n_448) );
INVx1_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
AOI21xp33_ASAP7_75t_SL g298 ( .A1(n_299), .A2(n_301), .B(n_303), .Y(n_298) );
INVx1_ASAP7_75t_L g452 ( .A(n_299), .Y(n_452) );
INVx2_ASAP7_75t_SL g366 ( .A(n_300), .Y(n_366) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
A2O1A1Ixp33_ASAP7_75t_L g447 ( .A1(n_303), .A2(n_384), .B(n_448), .C(n_449), .Y(n_447) );
OAI322xp33_ASAP7_75t_SL g316 ( .A1(n_304), .A2(n_317), .A3(n_320), .B1(n_321), .B2(n_322), .C1(n_324), .C2(n_327), .Y(n_316) );
INVx2_ASAP7_75t_L g336 ( .A(n_304), .Y(n_336) );
AOI221xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_312), .B1(n_313), .B2(n_315), .C(n_316), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
OAI22xp33_ASAP7_75t_SL g382 ( .A1(n_307), .A2(n_383), .B1(n_384), .B2(n_387), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_308), .B(n_311), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_308), .B(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
OR2x2_ASAP7_75t_L g381 ( .A(n_310), .B(n_343), .Y(n_381) );
INVx1_ASAP7_75t_L g371 ( .A(n_311), .Y(n_371) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g424 ( .A1(n_315), .A2(n_425), .B(n_427), .Y(n_424) );
AOI21xp33_ASAP7_75t_L g349 ( .A1(n_317), .A2(n_350), .B(n_353), .Y(n_349) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NOR2xp67_ASAP7_75t_SL g378 ( .A(n_319), .B(n_379), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_319), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_SL g435 ( .A(n_320), .Y(n_435) );
INVx1_ASAP7_75t_SL g322 ( .A(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND4xp25_ASAP7_75t_L g328 ( .A(n_329), .B(n_356), .C(n_372), .D(n_388), .Y(n_328) );
AOI211xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_332), .B(n_337), .C(n_349), .Y(n_329) );
INVx1_ASAP7_75t_L g421 ( .A(n_330), .Y(n_421) );
AND2x2_ASAP7_75t_L g369 ( .A(n_331), .B(n_352), .Y(n_369) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_334), .B(n_336), .Y(n_333) );
INVx1_ASAP7_75t_SL g334 ( .A(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_336), .B(n_371), .Y(n_370) );
OAI22xp33_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_342), .B1(n_345), .B2(n_347), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_339), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g387 ( .A(n_340), .Y(n_387) );
O2A1O1Ixp33_ASAP7_75t_L g401 ( .A1(n_340), .A2(n_379), .B(n_402), .C(n_404), .Y(n_401) );
OR2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx1_ASAP7_75t_L g386 ( .A(n_343), .Y(n_386) );
INVx1_ASAP7_75t_L g446 ( .A(n_344), .Y(n_446) );
NAND2xp33_ASAP7_75t_SL g436 ( .A(n_345), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_SL g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g375 ( .A(n_354), .Y(n_375) );
O2A1O1Ixp33_ASAP7_75t_L g356 ( .A1(n_357), .A2(n_360), .B(n_361), .C(n_363), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
OAI22xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_365), .B1(n_368), .B2(n_370), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_366), .B(n_367), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_366), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_371), .B(n_392), .Y(n_454) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AOI21xp33_ASAP7_75t_SL g376 ( .A1(n_377), .A2(n_380), .B(n_381), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
AOI221xp5_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_394), .B1(n_397), .B2(n_399), .C(n_401), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .Y(n_390) );
INVx1_ASAP7_75t_SL g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVxp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_404), .A2(n_421), .B1(n_422), .B2(n_423), .Y(n_420) );
NAND3xp33_ASAP7_75t_SL g406 ( .A(n_407), .B(n_414), .C(n_424), .Y(n_406) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_SL g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
CKINVDCx16_ASAP7_75t_R g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVxp67_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
OAI211xp5_ASAP7_75t_L g430 ( .A1(n_431), .A2(n_432), .B(n_433), .C(n_442), .Y(n_430) );
INVx1_ASAP7_75t_L g451 ( .A(n_431), .Y(n_451) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_436), .B1(n_438), .B2(n_440), .Y(n_433) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_451), .B1(n_452), .B2(n_453), .Y(n_449) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx2_ASAP7_75t_L g463 ( .A(n_457), .Y(n_463) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g465 ( .A(n_463), .Y(n_465) );
NAND3xp33_ASAP7_75t_L g466 ( .A(n_464), .B(n_467), .C(n_759), .Y(n_466) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AOI22x1_ASAP7_75t_SL g756 ( .A1(n_470), .A2(n_741), .B1(n_757), .B2(n_758), .Y(n_756) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g757 ( .A(n_474), .Y(n_757) );
OR2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_671), .Y(n_474) );
NAND5xp2_ASAP7_75t_L g475 ( .A(n_476), .B(n_586), .C(n_618), .D(n_635), .E(n_658), .Y(n_475) );
AOI221xp5_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_519), .B1(n_549), .B2(n_553), .C(n_557), .Y(n_476) );
INVx1_ASAP7_75t_L g698 ( .A(n_477), .Y(n_698) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_498), .Y(n_477) );
AND3x2_ASAP7_75t_L g673 ( .A(n_478), .B(n_500), .C(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_488), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_479), .B(n_555), .Y(n_554) );
BUFx3_ASAP7_75t_L g564 ( .A(n_479), .Y(n_564) );
AND2x2_ASAP7_75t_L g568 ( .A(n_479), .B(n_510), .Y(n_568) );
INVx2_ASAP7_75t_L g595 ( .A(n_479), .Y(n_595) );
OR2x2_ASAP7_75t_L g606 ( .A(n_479), .B(n_511), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g625 ( .A(n_479), .B(n_499), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_479), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g685 ( .A(n_479), .B(n_511), .Y(n_685) );
HB1xp67_ASAP7_75t_L g567 ( .A(n_488), .Y(n_567) );
AND2x2_ASAP7_75t_L g626 ( .A(n_488), .B(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_488), .B(n_499), .Y(n_645) );
INVx1_ASAP7_75t_SL g488 ( .A(n_489), .Y(n_488) );
OR2x2_ASAP7_75t_L g556 ( .A(n_489), .B(n_499), .Y(n_556) );
HB1xp67_ASAP7_75t_L g563 ( .A(n_489), .Y(n_563) );
AND2x2_ASAP7_75t_L g612 ( .A(n_489), .B(n_511), .Y(n_612) );
NAND3xp33_ASAP7_75t_L g637 ( .A(n_489), .B(n_498), .C(n_595), .Y(n_637) );
AND2x2_ASAP7_75t_L g702 ( .A(n_489), .B(n_500), .Y(n_702) );
AND2x2_ASAP7_75t_L g736 ( .A(n_489), .B(n_499), .Y(n_736) );
INVxp67_ASAP7_75t_L g565 ( .A(n_498), .Y(n_565) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_510), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_499), .B(n_595), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_499), .B(n_626), .Y(n_634) );
AND2x2_ASAP7_75t_L g684 ( .A(n_499), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g712 ( .A(n_499), .Y(n_712) );
INVx4_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g619 ( .A(n_500), .B(n_612), .Y(n_619) );
BUFx3_ASAP7_75t_L g651 ( .A(n_500), .Y(n_651) );
INVx2_ASAP7_75t_L g627 ( .A(n_510), .Y(n_627) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_511), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_519), .A2(n_687), .B1(n_689), .B2(n_690), .Y(n_686) );
AND2x2_ASAP7_75t_L g519 ( .A(n_520), .B(n_529), .Y(n_519) );
AND2x2_ASAP7_75t_L g549 ( .A(n_520), .B(n_550), .Y(n_549) );
INVx3_ASAP7_75t_SL g560 ( .A(n_520), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_520), .B(n_590), .Y(n_622) );
OR2x2_ASAP7_75t_L g641 ( .A(n_520), .B(n_530), .Y(n_641) );
AND2x2_ASAP7_75t_L g646 ( .A(n_520), .B(n_598), .Y(n_646) );
AND2x2_ASAP7_75t_L g649 ( .A(n_520), .B(n_591), .Y(n_649) );
AND2x2_ASAP7_75t_L g661 ( .A(n_520), .B(n_540), .Y(n_661) );
AND2x2_ASAP7_75t_L g677 ( .A(n_520), .B(n_531), .Y(n_677) );
AND2x4_ASAP7_75t_L g680 ( .A(n_520), .B(n_551), .Y(n_680) );
OR2x2_ASAP7_75t_L g697 ( .A(n_520), .B(n_633), .Y(n_697) );
OR2x2_ASAP7_75t_L g728 ( .A(n_520), .B(n_573), .Y(n_728) );
NAND2xp5_ASAP7_75t_SL g730 ( .A(n_520), .B(n_656), .Y(n_730) );
OR2x6_ASAP7_75t_L g520 ( .A(n_521), .B(n_527), .Y(n_520) );
AND2x2_ASAP7_75t_L g604 ( .A(n_529), .B(n_571), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_529), .B(n_591), .Y(n_723) );
AND2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_540), .Y(n_529) );
AND2x2_ASAP7_75t_L g559 ( .A(n_530), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g590 ( .A(n_530), .B(n_591), .Y(n_590) );
AND2x2_ASAP7_75t_L g598 ( .A(n_530), .B(n_573), .Y(n_598) );
AND2x2_ASAP7_75t_L g616 ( .A(n_530), .B(n_551), .Y(n_616) );
OR2x2_ASAP7_75t_L g633 ( .A(n_530), .B(n_591), .Y(n_633) );
INVx2_ASAP7_75t_SL g530 ( .A(n_531), .Y(n_530) );
BUFx2_ASAP7_75t_L g552 ( .A(n_531), .Y(n_552) );
AND2x2_ASAP7_75t_L g656 ( .A(n_531), .B(n_540), .Y(n_656) );
INVx2_ASAP7_75t_L g551 ( .A(n_540), .Y(n_551) );
INVx1_ASAP7_75t_L g668 ( .A(n_540), .Y(n_668) );
AND2x2_ASAP7_75t_L g718 ( .A(n_540), .B(n_560), .Y(n_718) );
AND2x2_ASAP7_75t_L g570 ( .A(n_550), .B(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g602 ( .A(n_550), .B(n_560), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_550), .B(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
AND2x2_ASAP7_75t_L g589 ( .A(n_551), .B(n_560), .Y(n_589) );
OR2x2_ASAP7_75t_L g705 ( .A(n_552), .B(n_679), .Y(n_705) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_555), .B(n_685), .Y(n_691) );
INVx2_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
OAI32xp33_ASAP7_75t_L g647 ( .A1(n_556), .A2(n_648), .A3(n_650), .B1(n_652), .B2(n_653), .Y(n_647) );
OR2x2_ASAP7_75t_L g664 ( .A(n_556), .B(n_606), .Y(n_664) );
OAI21xp33_ASAP7_75t_SL g689 ( .A1(n_556), .A2(n_566), .B(n_594), .Y(n_689) );
OAI22xp33_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_561), .B1(n_566), .B2(n_569), .Y(n_557) );
INVxp33_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_559), .B(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_560), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g615 ( .A(n_560), .B(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g715 ( .A(n_560), .B(n_656), .Y(n_715) );
OR2x2_ASAP7_75t_L g739 ( .A(n_560), .B(n_633), .Y(n_739) );
AOI21xp33_ASAP7_75t_L g722 ( .A1(n_561), .A2(n_621), .B(n_723), .Y(n_722) );
OR2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_565), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
INVx1_ASAP7_75t_L g599 ( .A(n_563), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_563), .B(n_568), .Y(n_617) );
AND2x2_ASAP7_75t_L g639 ( .A(n_564), .B(n_612), .Y(n_639) );
INVx1_ASAP7_75t_L g652 ( .A(n_564), .Y(n_652) );
OR2x2_ASAP7_75t_L g657 ( .A(n_564), .B(n_591), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_567), .B(n_606), .Y(n_605) );
OAI22xp33_ASAP7_75t_L g587 ( .A1(n_568), .A2(n_588), .B1(n_593), .B2(n_597), .Y(n_587) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_571), .A2(n_630), .B1(n_637), .B2(n_638), .Y(n_636) );
AND2x2_ASAP7_75t_L g714 ( .A(n_571), .B(n_715), .Y(n_714) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_573), .B(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g733 ( .A(n_573), .B(n_616), .Y(n_733) );
AO21x2_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_576), .B(n_584), .Y(n_573) );
INVx1_ASAP7_75t_L g592 ( .A(n_574), .Y(n_592) );
INVx1_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
OA21x2_ASAP7_75t_L g591 ( .A1(n_577), .A2(n_585), .B(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AOI221xp5_ASAP7_75t_L g586 ( .A1(n_587), .A2(n_599), .B1(n_600), .B2(n_605), .C(n_607), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_589), .B(n_591), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_589), .B(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g608 ( .A(n_590), .Y(n_608) );
O2A1O1Ixp33_ASAP7_75t_L g695 ( .A1(n_590), .A2(n_696), .B(n_697), .C(n_698), .Y(n_695) );
AND2x2_ASAP7_75t_L g700 ( .A(n_590), .B(n_680), .Y(n_700) );
O2A1O1Ixp33_ASAP7_75t_SL g738 ( .A1(n_590), .A2(n_679), .B(n_739), .C(n_740), .Y(n_738) );
BUFx3_ASAP7_75t_L g630 ( .A(n_591), .Y(n_630) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_594), .B(n_651), .Y(n_694) );
AOI211xp5_ASAP7_75t_L g713 ( .A1(n_594), .A2(n_714), .B(n_716), .C(n_722), .Y(n_713) );
AND2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_596), .Y(n_594) );
INVxp67_ASAP7_75t_L g674 ( .A(n_596), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_598), .B(n_718), .Y(n_717) );
NAND2xp5_ASAP7_75t_SL g600 ( .A(n_601), .B(n_603), .Y(n_600) );
INVx1_ASAP7_75t_SL g601 ( .A(n_602), .Y(n_601) );
AOI211xp5_ASAP7_75t_L g618 ( .A1(n_602), .A2(n_619), .B(n_620), .C(n_628), .Y(n_618) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g703 ( .A(n_606), .Y(n_703) );
OR2x2_ASAP7_75t_L g720 ( .A(n_606), .B(n_650), .Y(n_720) );
OAI22xp5_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_609), .B1(n_614), .B2(n_617), .Y(n_607) );
OAI22xp33_ASAP7_75t_L g620 ( .A1(n_609), .A2(n_621), .B1(n_622), .B2(n_623), .Y(n_620) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_611), .B(n_613), .Y(n_610) );
OR2x2_ASAP7_75t_L g707 ( .A(n_611), .B(n_651), .Y(n_707) );
INVx1_ASAP7_75t_SL g611 ( .A(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g662 ( .A(n_612), .B(n_652), .Y(n_662) );
INVx1_ASAP7_75t_L g670 ( .A(n_613), .Y(n_670) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_616), .B(n_630), .Y(n_678) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
NAND2xp5_ASAP7_75t_SL g669 ( .A(n_626), .B(n_670), .Y(n_669) );
INVx2_ASAP7_75t_L g735 ( .A(n_627), .Y(n_735) );
AOI21xp33_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_631), .B(n_634), .Y(n_628) );
INVx1_ASAP7_75t_L g665 ( .A(n_629), .Y(n_665) );
NAND2xp5_ASAP7_75t_SL g640 ( .A(n_630), .B(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_630), .B(n_661), .Y(n_660) );
NAND2x1p5_ASAP7_75t_L g681 ( .A(n_630), .B(n_656), .Y(n_681) );
NAND2xp5_ASAP7_75t_SL g688 ( .A(n_630), .B(n_677), .Y(n_688) );
OAI211xp5_ASAP7_75t_L g692 ( .A1(n_630), .A2(n_640), .B(n_680), .C(n_693), .Y(n_692) );
INVx1_ASAP7_75t_SL g632 ( .A(n_633), .Y(n_632) );
AOI221xp5_ASAP7_75t_SL g635 ( .A1(n_636), .A2(n_640), .B1(n_642), .B2(n_646), .C(n_647), .Y(n_635) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVxp67_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_644), .B(n_652), .Y(n_726) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
O2A1O1Ixp33_ASAP7_75t_L g737 ( .A1(n_646), .A2(n_661), .B(n_663), .C(n_738), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_649), .B(n_656), .Y(n_721) );
NAND2xp5_ASAP7_75t_SL g740 ( .A(n_650), .B(n_703), .Y(n_740) );
CKINVDCx16_ASAP7_75t_R g650 ( .A(n_651), .Y(n_650) );
INVxp33_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NOR2xp33_ASAP7_75t_L g654 ( .A(n_655), .B(n_657), .Y(n_654) );
AOI21xp33_ASAP7_75t_SL g666 ( .A1(n_655), .A2(n_667), .B(n_669), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g727 ( .A(n_655), .B(n_728), .Y(n_727) );
INVx2_ASAP7_75t_SL g655 ( .A(n_656), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_656), .B(n_710), .Y(n_709) );
AOI221xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_662), .B1(n_663), .B2(n_665), .C(n_666), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_662), .B(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g696 ( .A(n_668), .Y(n_696) );
NAND5xp2_ASAP7_75t_L g671 ( .A(n_672), .B(n_699), .C(n_713), .D(n_724), .E(n_737), .Y(n_671) );
AOI211xp5_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_675), .B(n_682), .C(n_695), .Y(n_672) );
INVx2_ASAP7_75t_SL g719 ( .A(n_673), .Y(n_719) );
NAND4xp25_ASAP7_75t_SL g675 ( .A(n_676), .B(n_678), .C(n_679), .D(n_681), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx3_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
OAI211xp5_ASAP7_75t_SL g682 ( .A1(n_681), .A2(n_683), .B(n_686), .C(n_692), .Y(n_682) );
CKINVDCx20_ASAP7_75t_R g683 ( .A(n_684), .Y(n_683) );
AOI221xp5_ASAP7_75t_L g724 ( .A1(n_684), .A2(n_725), .B1(n_727), .B2(n_729), .C(n_731), .Y(n_724) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AOI221xp5_ASAP7_75t_SL g699 ( .A1(n_700), .A2(n_701), .B1(n_704), .B2(n_706), .C(n_708), .Y(n_699) );
AND2x2_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
OAI22xp5_ASAP7_75t_L g731 ( .A1(n_707), .A2(n_730), .B1(n_732), .B2(n_734), .Y(n_731) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_SL g710 ( .A(n_711), .Y(n_710) );
OAI22xp5_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_719), .B1(n_720), .B2(n_721), .Y(n_716) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_SL g732 ( .A(n_733), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_735), .B(n_736), .Y(n_734) );
INVx1_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
INVx2_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_745), .Y(n_754) );
CKINVDCx16_ASAP7_75t_R g747 ( .A(n_748), .Y(n_747) );
INVx2_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_SL g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
endmodule