module real_aes_12740_n_78 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_77, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_78);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_78;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_673;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_528;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_236;
wire n_278;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_87;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_288;
wire n_147;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_662;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_653;
wire n_365;
wire n_290;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_633;
wire n_679;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
OA21x2_ASAP7_75t_L g109 ( .A1(n_0), .A2(n_41), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g185 ( .A(n_0), .Y(n_185) );
INVxp67_ASAP7_75t_SL g498 ( .A(n_1), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_1), .A2(n_54), .B1(n_643), .B2(n_644), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_2), .B(n_220), .Y(n_219) );
NAND2xp33_ASAP7_75t_L g241 ( .A(n_3), .B(n_242), .Y(n_241) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_4), .A2(n_29), .B1(n_517), .B2(n_535), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_4), .A2(n_10), .B1(n_630), .B2(n_633), .Y(n_629) );
BUFx3_ASAP7_75t_L g495 ( .A(n_5), .Y(n_495) );
INVx3_ASAP7_75t_L g566 ( .A(n_6), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_7), .B(n_163), .Y(n_162) );
XNOR2xp5_ASAP7_75t_L g482 ( .A(n_8), .B(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g491 ( .A(n_9), .Y(n_491) );
INVx1_ASAP7_75t_L g540 ( .A(n_9), .Y(n_540) );
AOI221xp5_ASAP7_75t_SL g505 ( .A1(n_10), .A2(n_70), .B1(n_506), .B2(n_508), .C(n_511), .Y(n_505) );
CKINVDCx5p33_ASAP7_75t_R g200 ( .A(n_11), .Y(n_200) );
INVx1_ASAP7_75t_L g96 ( .A(n_12), .Y(n_96) );
BUFx3_ASAP7_75t_L g116 ( .A(n_12), .Y(n_116) );
A2O1A1Ixp33_ASAP7_75t_L g176 ( .A1(n_13), .A2(n_128), .B(n_177), .C(n_180), .Y(n_176) );
INVx1_ASAP7_75t_L g553 ( .A(n_14), .Y(n_553) );
BUFx10_ASAP7_75t_L g691 ( .A(n_15), .Y(n_691) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_16), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_17), .B(n_118), .Y(n_168) );
AOI22xp5_ASAP7_75t_L g672 ( .A1(n_17), .A2(n_673), .B1(n_674), .B2(n_679), .Y(n_672) );
INVx1_ASAP7_75t_L g679 ( .A(n_17), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_18), .B(n_234), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_19), .B(n_155), .Y(n_267) );
A2O1A1Ixp33_ASAP7_75t_L g189 ( .A1(n_20), .A2(n_190), .B(n_191), .C(n_193), .Y(n_189) );
AND2x2_ASAP7_75t_L g144 ( .A(n_21), .B(n_108), .Y(n_144) );
AOI221xp5_ASAP7_75t_L g525 ( .A1(n_22), .A2(n_50), .B1(n_526), .B2(n_528), .C(n_532), .Y(n_525) );
INVxp33_ASAP7_75t_SL g591 ( .A(n_22), .Y(n_591) );
AND2x2_ASAP7_75t_L g577 ( .A(n_23), .B(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g603 ( .A(n_23), .B(n_33), .Y(n_603) );
INVxp33_ASAP7_75t_L g621 ( .A(n_23), .Y(n_621) );
INVx1_ASAP7_75t_L g638 ( .A(n_23), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_24), .B(n_136), .Y(n_169) );
AOI22xp33_ASAP7_75t_L g209 ( .A1(n_25), .A2(n_59), .B1(n_161), .B2(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g86 ( .A(n_26), .Y(n_86) );
INVx2_ASAP7_75t_L g574 ( .A(n_27), .Y(n_574) );
INVx1_ASAP7_75t_L g223 ( .A(n_28), .Y(n_223) );
INVx1_ASAP7_75t_L g624 ( .A(n_29), .Y(n_624) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_30), .B(n_161), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_31), .B(n_136), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_32), .B(n_179), .Y(n_266) );
INVx2_ASAP7_75t_L g578 ( .A(n_33), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_33), .B(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_34), .B(n_136), .Y(n_135) );
NAND2xp5_ASAP7_75t_SL g153 ( .A(n_35), .B(n_94), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_36), .Y(n_178) );
AND2x4_ASAP7_75t_L g85 ( .A(n_37), .B(n_86), .Y(n_85) );
HB1xp67_ASAP7_75t_L g656 ( .A(n_37), .Y(n_656) );
INVx1_ASAP7_75t_L g492 ( .A(n_38), .Y(n_492) );
INVx1_ASAP7_75t_L g524 ( .A(n_38), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g207 ( .A1(n_39), .A2(n_66), .B1(n_161), .B2(n_163), .Y(n_207) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_40), .A2(n_72), .B1(n_517), .B2(n_521), .Y(n_516) );
INVxp33_ASAP7_75t_L g579 ( .A(n_40), .Y(n_579) );
INVx1_ASAP7_75t_L g184 ( .A(n_41), .Y(n_184) );
INVx1_ASAP7_75t_L g110 ( .A(n_42), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g678 ( .A(n_43), .Y(n_678) );
OAI22xp5_ASAP7_75t_L g661 ( .A1(n_44), .A2(n_662), .B1(n_663), .B2(n_664), .Y(n_661) );
INVx1_ASAP7_75t_L g663 ( .A(n_44), .Y(n_663) );
INVx1_ASAP7_75t_L g548 ( .A(n_45), .Y(n_548) );
OAI22xp5_ASAP7_75t_L g536 ( .A1(n_46), .A2(n_74), .B1(n_537), .B2(n_543), .Y(n_536) );
INVx1_ASAP7_75t_L g605 ( .A(n_46), .Y(n_605) );
AND2x2_ASAP7_75t_L g274 ( .A(n_47), .B(n_137), .Y(n_274) );
BUFx2_ASAP7_75t_L g676 ( .A(n_48), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_49), .B(n_155), .Y(n_154) );
BUFx2_ASAP7_75t_L g696 ( .A(n_49), .Y(n_696) );
INVxp33_ASAP7_75t_SL g586 ( .A(n_50), .Y(n_586) );
NAND2x1_ASAP7_75t_L g127 ( .A(n_51), .B(n_128), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_52), .B(n_240), .Y(n_239) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_52), .Y(n_667) );
CKINVDCx5p33_ASAP7_75t_R g669 ( .A(n_53), .Y(n_669) );
INVxp33_ASAP7_75t_SL g556 ( .A(n_54), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g166 ( .A(n_55), .B(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_56), .B(n_125), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g113 ( .A(n_57), .B(n_114), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_58), .B(n_196), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g273 ( .A(n_60), .B(n_179), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_61), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_62), .B(n_118), .Y(n_117) );
NAND2xp33_ASAP7_75t_SL g218 ( .A(n_63), .B(n_119), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_64), .B(n_150), .Y(n_215) );
INVx1_ASAP7_75t_L g560 ( .A(n_65), .Y(n_560) );
OAI21xp5_ASAP7_75t_L g596 ( .A1(n_65), .A2(n_597), .B(n_604), .Y(n_596) );
INVx1_ASAP7_75t_L g90 ( .A(n_67), .Y(n_90) );
INVx1_ASAP7_75t_L g132 ( .A(n_67), .Y(n_132) );
BUFx3_ASAP7_75t_L g151 ( .A(n_67), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_68), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_69), .B(n_272), .Y(n_271) );
INVxp67_ASAP7_75t_L g584 ( .A(n_70), .Y(n_584) );
INVx2_ASAP7_75t_L g575 ( .A(n_71), .Y(n_575) );
INVxp67_ASAP7_75t_SL g589 ( .A(n_71), .Y(n_589) );
AND2x2_ASAP7_75t_L g594 ( .A(n_71), .B(n_574), .Y(n_594) );
INVx1_ASAP7_75t_L g628 ( .A(n_72), .Y(n_628) );
NAND2xp33_ASAP7_75t_L g235 ( .A(n_73), .B(n_236), .Y(n_235) );
INVx1_ASAP7_75t_L g641 ( .A(n_74), .Y(n_641) );
INVx2_ASAP7_75t_L g497 ( .A(n_75), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g149 ( .A(n_76), .B(n_150), .Y(n_149) );
HB1xp67_ASAP7_75t_L g662 ( .A(n_77), .Y(n_662) );
AOI21xp5_ASAP7_75t_L g78 ( .A1(n_79), .A2(n_97), .B(n_481), .Y(n_78) );
CKINVDCx6p67_ASAP7_75t_R g79 ( .A(n_80), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_81), .Y(n_80) );
AND2x2_ASAP7_75t_L g81 ( .A(n_82), .B(n_87), .Y(n_81) );
BUFx2_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
NAND3xp33_ASAP7_75t_L g202 ( .A(n_83), .B(n_203), .C(n_205), .Y(n_202) );
NAND3xp33_ASAP7_75t_L g208 ( .A(n_83), .B(n_131), .C(n_205), .Y(n_208) );
INVx1_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
INVx2_ASAP7_75t_L g134 ( .A(n_85), .Y(n_134) );
BUFx6f_ASAP7_75t_SL g142 ( .A(n_85), .Y(n_142) );
INVx1_ASAP7_75t_L g264 ( .A(n_85), .Y(n_264) );
HB1xp67_ASAP7_75t_L g654 ( .A(n_86), .Y(n_654) );
INVxp67_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
AO21x2_ASAP7_75t_L g709 ( .A1(n_88), .A2(n_653), .B(n_710), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g88 ( .A(n_89), .B(n_91), .Y(n_88) );
BUFx3_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx1_ASAP7_75t_L g121 ( .A(n_90), .Y(n_121) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_94), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
INVx2_ASAP7_75t_L g119 ( .A(n_95), .Y(n_119) );
INVx2_ASAP7_75t_L g150 ( .A(n_95), .Y(n_150) );
INVx1_ASAP7_75t_L g236 ( .A(n_95), .Y(n_236) );
BUFx6f_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
INVx2_ASAP7_75t_L g130 ( .A(n_96), .Y(n_130) );
INVx1_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
AND2x4_ASAP7_75t_L g98 ( .A(n_99), .B(n_389), .Y(n_98) );
NOR3xp33_ASAP7_75t_L g99 ( .A(n_100), .B(n_321), .C(n_357), .Y(n_99) );
NAND2xp5_ASAP7_75t_L g100 ( .A(n_101), .B(n_288), .Y(n_100) );
AOI221xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_170), .B1(n_244), .B2(n_255), .C(n_258), .Y(n_101) );
INVx1_ASAP7_75t_L g316 ( .A(n_102), .Y(n_316) );
AND2x2_ASAP7_75t_L g102 ( .A(n_103), .B(n_139), .Y(n_102) );
AND2x2_ASAP7_75t_L g422 ( .A(n_103), .B(n_360), .Y(n_422) );
HB1xp67_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_104), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g367 ( .A(n_104), .B(n_310), .Y(n_367) );
AND2x2_ASAP7_75t_L g404 ( .A(n_104), .B(n_293), .Y(n_404) );
INVx1_ASAP7_75t_L g426 ( .A(n_104), .Y(n_426) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g285 ( .A(n_105), .Y(n_285) );
INVx1_ASAP7_75t_L g292 ( .A(n_105), .Y(n_292) );
OAI21x1_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_111), .B(n_135), .Y(n_105) );
OAI21xp5_ASAP7_75t_L g157 ( .A1(n_106), .A2(n_158), .B(n_169), .Y(n_157) );
OAI21x1_ASAP7_75t_L g294 ( .A1(n_106), .A2(n_158), .B(n_169), .Y(n_294) );
BUFx6f_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
BUFx6f_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVxp67_ASAP7_75t_SL g143 ( .A(n_108), .Y(n_143) );
NOR2xp67_ASAP7_75t_SL g263 ( .A(n_108), .B(n_264), .Y(n_263) );
BUFx6f_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g138 ( .A(n_109), .Y(n_138) );
INVxp33_ASAP7_75t_L g224 ( .A(n_109), .Y(n_224) );
BUFx2_ASAP7_75t_L g227 ( .A(n_109), .Y(n_227) );
INVx1_ASAP7_75t_L g186 ( .A(n_110), .Y(n_186) );
OAI21xp5_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_122), .B(n_133), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_117), .B(n_120), .Y(n_112) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g161 ( .A(n_115), .Y(n_161) );
INVx2_ASAP7_75t_L g242 ( .A(n_115), .Y(n_242) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_116), .Y(n_126) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_116), .Y(n_156) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_120), .A2(n_153), .B(n_154), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_120), .A2(n_166), .B(n_168), .Y(n_165) );
AO21x1_ASAP7_75t_L g214 ( .A1(n_120), .A2(n_215), .B(n_216), .Y(n_214) );
BUFx10_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
O2A1O1Ixp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_124), .B(n_127), .C(n_131), .Y(n_122) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx2_ASAP7_75t_L g210 ( .A(n_126), .Y(n_210) );
INVx2_ASAP7_75t_L g234 ( .A(n_126), .Y(n_234) );
INVx2_ASAP7_75t_L g272 ( .A(n_126), .Y(n_272) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx2_ASAP7_75t_L g148 ( .A(n_129), .Y(n_148) );
INVx2_ASAP7_75t_L g167 ( .A(n_129), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_129), .B(n_192), .Y(n_191) );
INVx3_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_130), .Y(n_179) );
INVx2_ASAP7_75t_L g268 ( .A(n_131), .Y(n_268) );
BUFx3_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g181 ( .A(n_132), .Y(n_181) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx2_ASAP7_75t_SL g187 ( .A(n_134), .Y(n_187) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
NAND2x1_ASAP7_75t_L g473 ( .A(n_139), .B(n_382), .Y(n_473) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_157), .Y(n_139) );
HB1xp67_ASAP7_75t_L g257 ( .A(n_140), .Y(n_257) );
BUFx2_ASAP7_75t_L g281 ( .A(n_140), .Y(n_281) );
INVx2_ASAP7_75t_L g297 ( .A(n_140), .Y(n_297) );
AND2x2_ASAP7_75t_L g341 ( .A(n_140), .B(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g361 ( .A(n_140), .Y(n_361) );
INVx2_ASAP7_75t_L g371 ( .A(n_140), .Y(n_371) );
INVx1_ASAP7_75t_L g419 ( .A(n_140), .Y(n_419) );
AND2x2_ASAP7_75t_L g436 ( .A(n_140), .B(n_296), .Y(n_436) );
OR2x6_ASAP7_75t_L g140 ( .A(n_141), .B(n_145), .Y(n_140) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_143), .B(n_144), .Y(n_141) );
OAI21x1_ASAP7_75t_L g158 ( .A1(n_142), .A2(n_159), .B(n_165), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_142), .A2(n_222), .B(n_226), .Y(n_225) );
OAI21x1_ASAP7_75t_L g231 ( .A1(n_142), .A2(n_232), .B(n_238), .Y(n_231) );
AOI211x1_ASAP7_75t_L g145 ( .A1(n_144), .A2(n_146), .B(n_151), .C(n_152), .Y(n_145) );
OAI21xp5_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_148), .B(n_149), .Y(n_146) );
INVx2_ASAP7_75t_L g164 ( .A(n_151), .Y(n_164) );
INVx2_ASAP7_75t_L g194 ( .A(n_151), .Y(n_194) );
INVx1_ASAP7_75t_L g237 ( .A(n_151), .Y(n_237) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g163 ( .A(n_156), .Y(n_163) );
INVx2_ASAP7_75t_L g220 ( .A(n_156), .Y(n_220) );
INVx2_ASAP7_75t_L g240 ( .A(n_156), .Y(n_240) );
INVx1_ASAP7_75t_L g283 ( .A(n_157), .Y(n_283) );
AND2x2_ASAP7_75t_L g340 ( .A(n_157), .B(n_296), .Y(n_340) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_162), .B(n_164), .Y(n_159) );
AO21x1_ASAP7_75t_L g217 ( .A1(n_164), .A2(n_218), .B(n_219), .Y(n_217) );
INVx1_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
OAI221xp5_ASAP7_75t_L g301 ( .A1(n_171), .A2(n_295), .B1(n_302), .B2(n_305), .C(n_308), .Y(n_301) );
OR2x2_ASAP7_75t_L g171 ( .A(n_172), .B(n_211), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
AND2x2_ASAP7_75t_L g313 ( .A(n_173), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g173 ( .A(n_174), .B(n_197), .Y(n_173) );
INVx2_ASAP7_75t_L g278 ( .A(n_174), .Y(n_278) );
OR2x2_ASAP7_75t_L g307 ( .A(n_174), .B(n_213), .Y(n_307) );
AND2x2_ASAP7_75t_L g398 ( .A(n_174), .B(n_198), .Y(n_398) );
AND2x2_ASAP7_75t_L g415 ( .A(n_174), .B(n_213), .Y(n_415) );
NAND2x1p5_ASAP7_75t_L g174 ( .A(n_175), .B(n_188), .Y(n_174) );
NAND2x1p5_ASAP7_75t_L g248 ( .A(n_175), .B(n_188), .Y(n_248) );
OR2x2_ASAP7_75t_L g175 ( .A(n_176), .B(n_182), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_178), .B(n_179), .Y(n_177) );
INVx1_ASAP7_75t_L g190 ( .A(n_179), .Y(n_190) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx2_ASAP7_75t_L g204 ( .A(n_181), .Y(n_204) );
OA21x2_ASAP7_75t_L g188 ( .A1(n_182), .A2(n_189), .B(n_195), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_183), .B(n_187), .Y(n_182) );
INVx2_ASAP7_75t_L g196 ( .A(n_183), .Y(n_196) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_183), .B(n_200), .Y(n_199) );
AO21x2_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_185), .B(n_186), .Y(n_183) );
AOI21x1_ASAP7_75t_L g206 ( .A1(n_184), .A2(n_185), .B(n_186), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_193), .A2(n_239), .B(n_241), .Y(n_238) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx1_ASAP7_75t_L g324 ( .A(n_197), .Y(n_324) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx1_ASAP7_75t_L g252 ( .A(n_198), .Y(n_252) );
AND2x2_ASAP7_75t_L g300 ( .A(n_198), .B(n_279), .Y(n_300) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_198), .Y(n_337) );
AND2x2_ASAP7_75t_L g344 ( .A(n_198), .B(n_229), .Y(n_344) );
INVx1_ASAP7_75t_L g388 ( .A(n_198), .Y(n_388) );
INVxp67_ASAP7_75t_L g480 ( .A(n_198), .Y(n_480) );
OR2x2_ASAP7_75t_L g198 ( .A(n_199), .B(n_201), .Y(n_198) );
OAI22xp5_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_207), .B1(n_208), .B2(n_209), .Y(n_201) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
OR2x2_ASAP7_75t_L g416 ( .A(n_211), .B(n_246), .Y(n_416) );
OR2x2_ASAP7_75t_L g466 ( .A(n_211), .B(n_336), .Y(n_466) );
INVx3_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g287 ( .A(n_212), .B(n_246), .Y(n_287) );
AND2x2_ASAP7_75t_L g387 ( .A(n_212), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g397 ( .A(n_212), .B(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_228), .Y(n_212) );
INVx2_ASAP7_75t_L g251 ( .A(n_213), .Y(n_251) );
AND2x2_ASAP7_75t_L g314 ( .A(n_213), .B(n_229), .Y(n_314) );
AND2x2_ASAP7_75t_L g325 ( .A(n_213), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g356 ( .A(n_213), .Y(n_356) );
AO31x2_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_217), .A3(n_221), .B(n_225), .Y(n_213) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_223), .B(n_224), .Y(n_222) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
BUFx3_ASAP7_75t_L g230 ( .A(n_227), .Y(n_230) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx1_ASAP7_75t_L g254 ( .A(n_229), .Y(n_254) );
INVx1_ASAP7_75t_L g279 ( .A(n_229), .Y(n_279) );
AND2x2_ASAP7_75t_L g365 ( .A(n_229), .B(n_252), .Y(n_365) );
AND2x2_ASAP7_75t_L g380 ( .A(n_229), .B(n_278), .Y(n_380) );
OAI21x1_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_243), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_235), .B(n_237), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_237), .A2(n_271), .B(n_273), .Y(n_270) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
NAND2x1p5_ASAP7_75t_L g245 ( .A(n_246), .B(n_249), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_247), .Y(n_353) );
AND2x2_ASAP7_75t_L g364 ( .A(n_247), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g299 ( .A(n_248), .B(n_251), .Y(n_299) );
INVx1_ASAP7_75t_L g326 ( .A(n_248), .Y(n_326) );
BUFx2_ASAP7_75t_L g338 ( .A(n_248), .Y(n_338) );
AND2x2_ASAP7_75t_L g346 ( .A(n_248), .B(n_297), .Y(n_346) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_248), .Y(n_429) );
AOI22xp5_ASAP7_75t_L g446 ( .A1(n_249), .A2(n_328), .B1(n_387), .B2(n_447), .Y(n_446) );
AND2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_253), .Y(n_249) );
AND2x2_ASAP7_75t_L g276 ( .A(n_250), .B(n_277), .Y(n_276) );
AND2x4_ASAP7_75t_L g379 ( .A(n_250), .B(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
INVx1_ASAP7_75t_L g376 ( .A(n_251), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_253), .B(n_306), .Y(n_305) );
INVx2_ASAP7_75t_L g396 ( .A(n_253), .Y(n_396) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_253), .B(n_414), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_253), .B(n_307), .Y(n_439) );
BUFx3_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_254), .B(n_356), .Y(n_355) );
INVxp67_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
OAI22xp5_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_275), .B1(n_280), .B2(n_286), .Y(n_258) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g304 ( .A(n_260), .Y(n_304) );
OR2x2_ASAP7_75t_L g373 ( .A(n_260), .B(n_349), .Y(n_373) );
INVx2_ASAP7_75t_L g296 ( .A(n_261), .Y(n_296) );
OR2x2_ASAP7_75t_L g312 ( .A(n_261), .B(n_294), .Y(n_312) );
AND2x2_ASAP7_75t_L g320 ( .A(n_261), .B(n_293), .Y(n_320) );
AND2x4_ASAP7_75t_L g360 ( .A(n_261), .B(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g383 ( .A(n_261), .Y(n_383) );
AND2x4_ASAP7_75t_L g261 ( .A(n_262), .B(n_269), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_263), .B(n_265), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_263), .A2(n_270), .B(n_274), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_267), .B(n_268), .Y(n_265) );
AOI21xp33_ASAP7_75t_SL g315 ( .A1(n_275), .A2(n_316), .B(n_317), .Y(n_315) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_281), .B(n_282), .Y(n_280) );
INVx1_ASAP7_75t_L g318 ( .A(n_281), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_281), .B(n_311), .Y(n_333) );
INVx1_ASAP7_75t_L g438 ( .A(n_281), .Y(n_438) );
INVx2_ASAP7_75t_L g462 ( .A(n_282), .Y(n_462) );
AND2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
INVx1_ASAP7_75t_L g303 ( .A(n_283), .Y(n_303) );
INVx2_ASAP7_75t_L g330 ( .A(n_284), .Y(n_330) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx2_ASAP7_75t_L g342 ( .A(n_285), .Y(n_342) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AOI211xp5_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_298), .B(n_301), .C(n_315), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_295), .Y(n_290) );
INVx2_ASAP7_75t_L g384 ( .A(n_291), .Y(n_384) );
INVx1_ASAP7_75t_L g433 ( .A(n_291), .Y(n_433) );
INVx2_ASAP7_75t_SL g478 ( .A(n_291), .Y(n_478) );
OR2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
INVx1_ASAP7_75t_L g310 ( .A(n_293), .Y(n_310) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g394 ( .A(n_295), .Y(n_394) );
OR2x2_ASAP7_75t_L g451 ( .A(n_295), .B(n_330), .Y(n_451) );
NAND2xp33_ASAP7_75t_L g477 ( .A(n_295), .B(n_478), .Y(n_477) );
OR2x2_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
AND2x4_ASAP7_75t_SL g370 ( .A(n_296), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g309 ( .A(n_297), .B(n_310), .Y(n_309) );
BUFx3_ASAP7_75t_L g349 ( .A(n_297), .Y(n_349) );
AND2x4_ASAP7_75t_SL g298 ( .A(n_299), .B(n_300), .Y(n_298) );
AND2x2_ASAP7_75t_L g409 ( .A(n_299), .B(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g463 ( .A(n_299), .B(n_344), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_299), .B(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_303), .B(n_360), .Y(n_448) );
INVx1_ASAP7_75t_L g458 ( .A(n_303), .Y(n_458) );
INVx1_ASAP7_75t_L g395 ( .A(n_306), .Y(n_395) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_L g400 ( .A(n_307), .B(n_401), .Y(n_400) );
OAI21xp33_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_311), .B(n_313), .Y(n_308) );
AND2x4_ASAP7_75t_L g328 ( .A(n_311), .B(n_329), .Y(n_328) );
AOI322xp5_ASAP7_75t_L g391 ( .A1(n_311), .A2(n_392), .A3(n_395), .B1(n_396), .B2(n_397), .C1(n_399), .C2(n_402), .Y(n_391) );
NAND3xp33_ASAP7_75t_L g407 ( .A(n_311), .B(n_329), .C(n_408), .Y(n_407) );
INVx4_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
OAI33xp33_ASAP7_75t_L g335 ( .A1(n_312), .A2(n_336), .A3(n_338), .B1(n_339), .B2(n_343), .B3(n_345), .Y(n_335) );
NOR2x1_ASAP7_75t_L g431 ( .A(n_312), .B(n_418), .Y(n_431) );
OR2x2_ASAP7_75t_L g445 ( .A(n_312), .B(n_426), .Y(n_445) );
AND2x2_ASAP7_75t_L g452 ( .A(n_314), .B(n_398), .Y(n_452) );
OR2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
OR2x2_ASAP7_75t_L g456 ( .A(n_319), .B(n_330), .Y(n_456) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g348 ( .A(n_320), .B(n_349), .Y(n_348) );
OAI211xp5_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_327), .B(n_331), .C(n_347), .Y(n_321) );
INVx1_ASAP7_75t_L g334 ( .A(n_322), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_323), .B(n_325), .Y(n_322) );
OR2x2_ASAP7_75t_L g413 ( .A(n_323), .B(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_325), .B(n_344), .Y(n_454) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_330), .B(n_340), .Y(n_351) );
AND2x2_ASAP7_75t_L g378 ( .A(n_330), .B(n_370), .Y(n_378) );
OR2x2_ASAP7_75t_L g475 ( .A(n_330), .B(n_476), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_334), .B(n_335), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
NAND4xp25_ASAP7_75t_L g468 ( .A(n_333), .B(n_469), .C(n_472), .D(n_473), .Y(n_468) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_L g424 ( .A(n_338), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
AND2x2_ASAP7_75t_L g425 ( .A(n_340), .B(n_426), .Y(n_425) );
AND2x2_ASAP7_75t_L g437 ( .A(n_340), .B(n_438), .Y(n_437) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_342), .Y(n_362) );
OR2x2_ASAP7_75t_L g418 ( .A(n_342), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx2_ASAP7_75t_L g401 ( .A(n_344), .Y(n_401) );
AND2x2_ASAP7_75t_L g423 ( .A(n_344), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
OAI21xp33_ASAP7_75t_SL g347 ( .A1(n_348), .A2(n_350), .B(n_352), .Y(n_347) );
INVx2_ASAP7_75t_L g408 ( .A(n_349), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_349), .B(n_433), .Y(n_432) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_349), .Y(n_443) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OAI32xp33_ASAP7_75t_L g464 ( .A1(n_351), .A2(n_401), .A3(n_415), .B1(n_465), .B2(n_466), .Y(n_464) );
NOR2x1p5_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
BUFx3_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OAI211xp5_ASAP7_75t_SL g357 ( .A1(n_358), .A2(n_363), .B(n_366), .C(n_377), .Y(n_357) );
NAND3xp33_ASAP7_75t_SL g461 ( .A(n_358), .B(n_373), .C(n_462), .Y(n_461) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_362), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_360), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_365), .B(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_365), .B(n_429), .Y(n_428) );
A2O1A1Ixp33_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_368), .B(n_372), .C(n_374), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_367), .B(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g476 ( .A(n_370), .Y(n_476) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AOI22xp33_ASAP7_75t_SL g377 ( .A1(n_378), .A2(n_379), .B1(n_381), .B2(n_385), .Y(n_377) );
INVx2_ASAP7_75t_L g459 ( .A(n_379), .Y(n_459) );
AND2x4_ASAP7_75t_SL g381 ( .A(n_382), .B(n_384), .Y(n_381) );
OR2x2_ASAP7_75t_L g417 ( .A(n_382), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g470 ( .A(n_382), .Y(n_470) );
INVx4_ASAP7_75t_R g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g472 ( .A(n_384), .Y(n_472) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx2_ASAP7_75t_L g410 ( .A(n_388), .Y(n_410) );
NOR2x1_ASAP7_75t_L g389 ( .A(n_390), .B(n_440), .Y(n_389) );
NAND3xp33_ASAP7_75t_L g390 ( .A(n_391), .B(n_405), .C(n_411), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
O2A1O1Ixp33_ASAP7_75t_L g457 ( .A1(n_394), .A2(n_456), .B(n_458), .C(n_459), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_399), .A2(n_468), .B(n_474), .Y(n_467) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_SL g405 ( .A(n_406), .B(n_409), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_412), .B(n_427), .Y(n_411) );
A2O1A1Ixp33_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_416), .B(n_417), .C(n_420), .Y(n_412) );
OAI221xp5_ASAP7_75t_L g427 ( .A1(n_413), .A2(n_428), .B1(n_430), .B2(n_432), .C(n_434), .Y(n_427) );
OA21x2_ASAP7_75t_L g441 ( .A1(n_414), .A2(n_442), .B(n_446), .Y(n_441) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AOI22xp5_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_422), .B1(n_423), .B2(n_425), .Y(n_420) );
AND2x2_ASAP7_75t_L g435 ( .A(n_426), .B(n_436), .Y(n_435) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_426), .Y(n_471) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OAI21xp33_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_437), .B(n_439), .Y(n_434) );
INVx1_ASAP7_75t_L g465 ( .A(n_435), .Y(n_465) );
NAND4xp75_ASAP7_75t_L g440 ( .A(n_441), .B(n_449), .C(n_460), .D(n_467), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_443), .B(n_444), .Y(n_442) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
AOI221xp5_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_452), .B1(n_453), .B2(n_455), .C(n_457), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_463), .B(n_464), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
AOI21xp33_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_477), .B(n_479), .Y(n_474) );
OAI221xp5_ASAP7_75t_L g481 ( .A1(n_482), .A2(n_483), .B1(n_648), .B2(n_657), .C(n_703), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g703 ( .A1(n_483), .A2(n_696), .B1(n_704), .B2(n_707), .Y(n_703) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_562), .B(n_567), .Y(n_484) );
NAND4xp25_ASAP7_75t_L g485 ( .A(n_486), .B(n_504), .C(n_547), .D(n_555), .Y(n_485) );
AOI21xp33_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_498), .B(n_499), .Y(n_486) );
AND2x4_ASAP7_75t_L g487 ( .A(n_488), .B(n_493), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx3_ASAP7_75t_L g507 ( .A(n_489), .Y(n_507) );
INVx1_ASAP7_75t_SL g535 ( .A(n_489), .Y(n_535) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
BUFx6f_ASAP7_75t_L g550 ( .A(n_490), .Y(n_550) );
AND2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
INVx2_ASAP7_75t_L g502 ( .A(n_491), .Y(n_502) );
AND2x2_ASAP7_75t_L g520 ( .A(n_491), .B(n_503), .Y(n_520) );
INVx2_ASAP7_75t_L g503 ( .A(n_492), .Y(n_503) );
AND2x4_ASAP7_75t_L g499 ( .A(n_493), .B(n_500), .Y(n_499) );
NAND2x1p5_ASAP7_75t_L g543 ( .A(n_493), .B(n_544), .Y(n_543) );
BUFx3_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx1_ASAP7_75t_L g542 ( .A(n_494), .Y(n_542) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_496), .Y(n_494) );
AND2x4_ASAP7_75t_L g514 ( .A(n_495), .B(n_515), .Y(n_514) );
OR2x2_ASAP7_75t_L g533 ( .A(n_495), .B(n_496), .Y(n_533) );
OR2x6_ASAP7_75t_L g552 ( .A(n_495), .B(n_497), .Y(n_552) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
BUFx2_ASAP7_75t_L g515 ( .A(n_497), .Y(n_515) );
AND2x4_ASAP7_75t_L g554 ( .A(n_500), .B(n_551), .Y(n_554) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx2_ASAP7_75t_L g510 ( .A(n_501), .Y(n_510) );
BUFx6f_ASAP7_75t_L g531 ( .A(n_501), .Y(n_531) );
AND2x4_ASAP7_75t_L g501 ( .A(n_502), .B(n_503), .Y(n_501) );
AND2x4_ASAP7_75t_L g523 ( .A(n_502), .B(n_524), .Y(n_523) );
AOI221xp5_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_516), .B1(n_525), .B2(n_534), .C(n_536), .Y(n_504) );
BUFx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
BUFx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx4_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
BUFx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx3_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx3_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
BUFx6f_ASAP7_75t_L g559 ( .A(n_520), .Y(n_559) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
CKINVDCx5p33_ASAP7_75t_R g527 ( .A(n_522), .Y(n_527) );
AND2x2_ASAP7_75t_L g561 ( .A(n_522), .B(n_551), .Y(n_561) );
BUFx12f_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g546 ( .A(n_524), .Y(n_546) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
NAND3xp33_ASAP7_75t_L g689 ( .A(n_532), .B(n_539), .C(n_690), .Y(n_689) );
BUFx6f_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx2_ASAP7_75t_SL g695 ( .A(n_537), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_537), .B(n_689), .Y(n_702) );
INVx2_ASAP7_75t_SL g537 ( .A(n_538), .Y(n_537) );
AND2x4_ASAP7_75t_L g538 ( .A(n_539), .B(n_541), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g547 ( .A1(n_548), .A2(n_549), .B1(n_553), .B2(n_554), .Y(n_547) );
OAI221xp5_ASAP7_75t_L g639 ( .A1(n_548), .A2(n_623), .B1(n_640), .B2(n_641), .C(n_642), .Y(n_639) );
AND2x4_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
AND2x4_ASAP7_75t_L g558 ( .A(n_551), .B(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_553), .A2(n_605), .B1(n_606), .B2(n_610), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_557), .B1(n_560), .B2(n_561), .Y(n_555) );
BUFx3_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
CKINVDCx5p33_ASAP7_75t_R g562 ( .A(n_563), .Y(n_562) );
BUFx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
OR2x6_ASAP7_75t_L g636 ( .A(n_565), .B(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x4_ASAP7_75t_L g576 ( .A(n_566), .B(n_577), .Y(n_576) );
NAND2x1p5_ASAP7_75t_L g602 ( .A(n_566), .B(n_603), .Y(n_602) );
AND2x4_ASAP7_75t_SL g609 ( .A(n_566), .B(n_603), .Y(n_609) );
AND3x1_ASAP7_75t_L g618 ( .A(n_566), .B(n_619), .C(n_621), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_595), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_569), .B(n_585), .Y(n_568) );
AOI22xp33_ASAP7_75t_SL g569 ( .A1(n_570), .A2(n_579), .B1(n_580), .B2(n_584), .Y(n_569) );
AND2x4_ASAP7_75t_L g570 ( .A(n_571), .B(n_576), .Y(n_570) );
BUFx6f_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx5_ASAP7_75t_L g634 ( .A(n_572), .Y(n_634) );
AND2x4_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .Y(n_572) );
INVx1_ASAP7_75t_L g590 ( .A(n_573), .Y(n_590) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx2_ASAP7_75t_L g582 ( .A(n_574), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_574), .B(n_575), .Y(n_601) );
INVx2_ASAP7_75t_L g583 ( .A(n_575), .Y(n_583) );
AND2x2_ASAP7_75t_L g580 ( .A(n_576), .B(n_581), .Y(n_580) );
AND2x6_ASAP7_75t_L g587 ( .A(n_576), .B(n_588), .Y(n_587) );
AND2x4_ASAP7_75t_L g592 ( .A(n_576), .B(n_593), .Y(n_592) );
INVx2_ASAP7_75t_L g620 ( .A(n_578), .Y(n_620) );
AND2x2_ASAP7_75t_L g647 ( .A(n_581), .B(n_609), .Y(n_647) );
AND2x4_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
BUFx3_ASAP7_75t_L g608 ( .A(n_582), .Y(n_608) );
NAND2x1p5_ASAP7_75t_L g627 ( .A(n_582), .B(n_583), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_587), .B1(n_591), .B2(n_592), .Y(n_585) );
AND2x4_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
INVx1_ASAP7_75t_L g613 ( .A(n_589), .Y(n_613) );
BUFx3_ASAP7_75t_L g643 ( .A(n_593), .Y(n_643) );
BUFx6f_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
BUFx4f_ASAP7_75t_L g632 ( .A(n_594), .Y(n_632) );
NOR3xp33_ASAP7_75t_L g595 ( .A(n_596), .B(n_614), .C(n_645), .Y(n_595) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
OR2x4_ASAP7_75t_L g599 ( .A(n_600), .B(n_602), .Y(n_599) );
BUFx6f_ASAP7_75t_L g623 ( .A(n_600), .Y(n_623) );
BUFx6f_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NAND2x1p5_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
AND2x4_ASAP7_75t_L g610 ( .A(n_609), .B(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
OAI22xp5_ASAP7_75t_SL g614 ( .A1(n_615), .A2(n_622), .B1(n_635), .B2(n_639), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx3_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OAI221xp5_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_624), .B1(n_625), .B2(n_628), .C(n_629), .Y(n_622) );
BUFx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
BUFx3_ASAP7_75t_L g640 ( .A(n_626), .Y(n_640) );
BUFx6f_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx4_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx3_ASAP7_75t_L g644 ( .A(n_634), .Y(n_644) );
BUFx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
CKINVDCx20_ASAP7_75t_R g648 ( .A(n_649), .Y(n_648) );
CKINVDCx20_ASAP7_75t_R g649 ( .A(n_650), .Y(n_649) );
BUFx6f_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_655), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
BUFx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g687 ( .A(n_654), .Y(n_687) );
AND2x2_ASAP7_75t_L g710 ( .A(n_655), .B(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_656), .B(n_687), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_681), .B1(n_696), .B2(n_697), .Y(n_657) );
OAI22xp5_ASAP7_75t_L g704 ( .A1(n_658), .A2(n_696), .B1(n_705), .B2(n_706), .Y(n_704) );
AOI22xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_671), .B1(n_672), .B2(n_680), .Y(n_658) );
INVx1_ASAP7_75t_L g680 ( .A(n_659), .Y(n_680) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_661), .B1(n_665), .B2(n_670), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g664 ( .A(n_662), .Y(n_664) );
INVx1_ASAP7_75t_L g670 ( .A(n_665), .Y(n_670) );
OAI22xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_667), .B1(n_668), .B2(n_669), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OAI22xp5_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_676), .B1(n_677), .B2(n_678), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
BUFx3_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx5_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx3_ASAP7_75t_L g705 ( .A(n_684), .Y(n_705) );
AND2x6_ASAP7_75t_L g684 ( .A(n_685), .B(n_692), .Y(n_684) );
NOR2xp33_ASAP7_75t_L g685 ( .A(n_686), .B(n_688), .Y(n_685) );
INVxp67_ASAP7_75t_L g701 ( .A(n_686), .Y(n_701) );
INVx1_ASAP7_75t_L g711 ( .A(n_687), .Y(n_711) );
INVxp67_ASAP7_75t_SL g688 ( .A(n_689), .Y(n_688) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
CKINVDCx11_ASAP7_75t_R g694 ( .A(n_691), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_693), .B(n_695), .Y(n_692) );
CKINVDCx5p33_ASAP7_75t_R g693 ( .A(n_694), .Y(n_693) );
INVx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
BUFx6f_ASAP7_75t_SL g698 ( .A(n_699), .Y(n_698) );
BUFx6f_ASAP7_75t_L g706 ( .A(n_699), .Y(n_706) );
INVx4_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
CKINVDCx20_ASAP7_75t_R g707 ( .A(n_708), .Y(n_707) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_709), .Y(n_708) );
endmodule