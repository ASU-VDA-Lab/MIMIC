module fake_netlist_6_143_n_779 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_127, n_125, n_77, n_106, n_92, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_779);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_779;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_144;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_142;
wire n_724;
wire n_143;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_698;
wire n_617;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_141;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_147;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_153;
wire n_720;
wire n_525;
wire n_758;
wire n_611;
wire n_156;
wire n_491;
wire n_145;
wire n_656;
wire n_772;
wire n_666;
wire n_371;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_260;
wire n_265;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_719;
wire n_594;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_152;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_767;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_550;
wire n_487;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_146;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_193;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_151;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_515;
wire n_434;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_778;
wire n_332;
wire n_336;
wire n_410;
wire n_398;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g141 ( 
.A(n_99),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_11),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_27),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_52),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_106),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_90),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_14),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_86),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_93),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_94),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_4),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_124),
.Y(n_153)
);

BUFx10_ASAP7_75t_L g154 ( 
.A(n_55),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_136),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_19),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_77),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_96),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_107),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_45),
.Y(n_160)
);

BUFx8_ASAP7_75t_SL g161 ( 
.A(n_134),
.Y(n_161)
);

NOR2xp67_ASAP7_75t_L g162 ( 
.A(n_50),
.B(n_139),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_47),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_54),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_12),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_114),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_138),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_126),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_48),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

INVx2_ASAP7_75t_SL g171 ( 
.A(n_30),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_64),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_131),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_84),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_105),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_91),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_111),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_82),
.Y(n_178)
);

BUFx10_ASAP7_75t_L g179 ( 
.A(n_85),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_62),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_10),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_25),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_137),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_87),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_122),
.Y(n_185)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_5),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_0),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_42),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_0),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_1),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_135),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_59),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_46),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_123),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_125),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_24),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_154),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_1),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_165),
.Y(n_199)
);

AND2x4_ASAP7_75t_L g200 ( 
.A(n_151),
.B(n_20),
.Y(n_200)
);

OAI22x1_ASAP7_75t_L g201 ( 
.A1(n_186),
.A2(n_187),
.B1(n_152),
.B2(n_142),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_175),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_147),
.B(n_2),
.Y(n_203)
);

BUFx8_ASAP7_75t_L g204 ( 
.A(n_175),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_147),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_175),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_154),
.B(n_2),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_141),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_154),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_175),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_151),
.B(n_3),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_163),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_163),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_156),
.Y(n_214)
);

BUFx8_ASAP7_75t_L g215 ( 
.A(n_170),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_181),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_170),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_146),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_176),
.B(n_3),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_189),
.Y(n_220)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_179),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_176),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_148),
.Y(n_223)
);

AND2x4_ASAP7_75t_L g224 ( 
.A(n_149),
.B(n_21),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_190),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_143),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_155),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_161),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_161),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_179),
.Y(n_230)
);

OAI21x1_ASAP7_75t_L g231 ( 
.A1(n_159),
.A2(n_9),
.B(n_10),
.Y(n_231)
);

OA21x2_ASAP7_75t_L g232 ( 
.A1(n_164),
.A2(n_11),
.B(n_12),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_166),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_143),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_179),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_167),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_168),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_150),
.B(n_13),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_172),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_202),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_213),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_213),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_229),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_213),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_229),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_202),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_213),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_234),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_234),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_202),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_199),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_216),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_216),
.Y(n_253)
);

BUFx10_ASAP7_75t_L g254 ( 
.A(n_214),
.Y(n_254)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_202),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_227),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_228),
.Y(n_257)
);

INVx6_ASAP7_75t_L g258 ( 
.A(n_204),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_197),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_197),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_209),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_209),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_235),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_235),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_199),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_220),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_230),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_230),
.B(n_144),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_205),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_227),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_230),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_R g272 ( 
.A(n_204),
.B(n_145),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_R g273 ( 
.A(n_204),
.B(n_169),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_212),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_221),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_221),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_221),
.Y(n_277)
);

BUFx10_ASAP7_75t_L g278 ( 
.A(n_208),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_201),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_219),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_212),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_212),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_R g283 ( 
.A(n_221),
.B(n_153),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_221),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_215),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_206),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_225),
.A2(n_169),
.B1(n_195),
.B2(n_194),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_215),
.Y(n_288)
);

INVxp33_ASAP7_75t_L g289 ( 
.A(n_273),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_267),
.B(n_238),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_255),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_241),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_268),
.B(n_224),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_255),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_246),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_271),
.B(n_238),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_250),
.Y(n_297)
);

INVx2_ASAP7_75t_SL g298 ( 
.A(n_254),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_242),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_244),
.Y(n_300)
);

AND2x4_ASAP7_75t_L g301 ( 
.A(n_256),
.B(n_224),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_259),
.B(n_224),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_275),
.B(n_215),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_260),
.B(n_207),
.Y(n_304)
);

NOR3xp33_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_207),
.C(n_198),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_240),
.Y(n_306)
);

OR2x2_ASAP7_75t_SL g307 ( 
.A(n_280),
.B(n_232),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_240),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_247),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_261),
.B(n_239),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_262),
.B(n_201),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_276),
.B(n_200),
.Y(n_312)
);

NAND2xp33_ASAP7_75t_L g313 ( 
.A(n_277),
.B(n_203),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_286),
.Y(n_314)
);

BUFx5_ASAP7_75t_L g315 ( 
.A(n_274),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_263),
.B(n_200),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_278),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_240),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_264),
.B(n_239),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g320 ( 
.A(n_278),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_266),
.B(n_237),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_240),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_284),
.B(n_211),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_270),
.B(n_218),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_288),
.B(n_200),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_281),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_282),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_254),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_283),
.B(n_212),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_283),
.B(n_212),
.Y(n_330)
);

NOR3xp33_ASAP7_75t_L g331 ( 
.A(n_279),
.B(n_222),
.C(n_203),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_258),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_258),
.B(n_218),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_258),
.B(n_218),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_252),
.Y(n_335)
);

NAND3xp33_ASAP7_75t_L g336 ( 
.A(n_253),
.B(n_226),
.C(n_233),
.Y(n_336)
);

AO221x1_ASAP7_75t_L g337 ( 
.A1(n_257),
.A2(n_173),
.B1(n_178),
.B2(n_174),
.C(n_183),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_272),
.B(n_218),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_285),
.B(n_223),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_272),
.B(n_157),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_269),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_243),
.B(n_223),
.Y(n_342)
);

NAND2xp33_ASAP7_75t_L g343 ( 
.A(n_245),
.B(n_158),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_248),
.B(n_223),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_249),
.B(n_223),
.Y(n_345)
);

AND2x4_ASAP7_75t_L g346 ( 
.A(n_251),
.B(n_217),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_265),
.B(n_160),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_268),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_268),
.B(n_233),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_268),
.B(n_233),
.Y(n_350)
);

NAND2x1p5_ASAP7_75t_L g351 ( 
.A(n_268),
.B(n_232),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_268),
.B(n_233),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_268),
.B(n_236),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_241),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_290),
.B(n_217),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_314),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_295),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_348),
.B(n_236),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_306),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_305),
.A2(n_232),
.B1(n_231),
.B2(n_162),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_297),
.Y(n_361)
);

OR2x6_ASAP7_75t_L g362 ( 
.A(n_298),
.B(n_231),
.Y(n_362)
);

AND2x4_ASAP7_75t_L g363 ( 
.A(n_301),
.B(n_185),
.Y(n_363)
);

INVx8_ASAP7_75t_L g364 ( 
.A(n_346),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_291),
.Y(n_365)
);

NAND2x1p5_ASAP7_75t_L g366 ( 
.A(n_320),
.B(n_188),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_301),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_290),
.B(n_236),
.Y(n_368)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_318),
.Y(n_369)
);

HB1xp67_ASAP7_75t_L g370 ( 
.A(n_346),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_348),
.B(n_236),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_296),
.B(n_177),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_293),
.B(n_236),
.Y(n_373)
);

OR2x2_ASAP7_75t_L g374 ( 
.A(n_321),
.B(n_341),
.Y(n_374)
);

NAND3xp33_ASAP7_75t_SL g375 ( 
.A(n_305),
.B(n_192),
.C(n_182),
.Y(n_375)
);

NAND3xp33_ASAP7_75t_SL g376 ( 
.A(n_331),
.B(n_196),
.C(n_193),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_310),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_336),
.A2(n_191),
.B1(n_184),
.B2(n_180),
.Y(n_378)
);

NAND2x1p5_ASAP7_75t_L g379 ( 
.A(n_335),
.B(n_206),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_306),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_296),
.B(n_210),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_292),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_300),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_349),
.B(n_210),
.Y(n_384)
);

HB1xp67_ASAP7_75t_L g385 ( 
.A(n_321),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_294),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_350),
.B(n_22),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_319),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_354),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_352),
.B(n_23),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_326),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_299),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_309),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_353),
.B(n_26),
.Y(n_394)
);

AOI22xp33_ASAP7_75t_L g395 ( 
.A1(n_331),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_395)
);

BUFx4f_ASAP7_75t_L g396 ( 
.A(n_328),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g397 ( 
.A(n_344),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_319),
.B(n_15),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_304),
.B(n_16),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_327),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_306),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_308),
.Y(n_402)
);

AOI22xp33_ASAP7_75t_L g403 ( 
.A1(n_351),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_322),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_344),
.B(n_17),
.Y(n_405)
);

OR2x4_ASAP7_75t_L g406 ( 
.A(n_345),
.B(n_18),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_308),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_351),
.B(n_28),
.Y(n_408)
);

INVxp67_ASAP7_75t_SL g409 ( 
.A(n_308),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_323),
.B(n_29),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_337),
.A2(n_19),
.B1(n_31),
.B2(n_32),
.Y(n_411)
);

BUFx4f_ASAP7_75t_L g412 ( 
.A(n_332),
.Y(n_412)
);

INVx2_ASAP7_75t_SL g413 ( 
.A(n_316),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_323),
.B(n_33),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_312),
.B(n_34),
.Y(n_415)
);

OR2x6_ASAP7_75t_L g416 ( 
.A(n_317),
.B(n_35),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_345),
.B(n_36),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_R g418 ( 
.A(n_343),
.B(n_37),
.Y(n_418)
);

BUFx8_ASAP7_75t_L g419 ( 
.A(n_289),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_342),
.B(n_38),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_324),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_324),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_342),
.B(n_39),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_370),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_395),
.A2(n_307),
.B1(n_317),
.B2(n_311),
.Y(n_425)
);

OAI21xp33_ASAP7_75t_L g426 ( 
.A1(n_399),
.A2(n_302),
.B(n_325),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_385),
.B(n_347),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_382),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_368),
.B(n_339),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_383),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_388),
.B(n_397),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_410),
.A2(n_414),
.B1(n_372),
.B2(n_421),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_408),
.A2(n_330),
.B(n_329),
.Y(n_433)
);

NOR2x1_ASAP7_75t_L g434 ( 
.A(n_374),
.B(n_338),
.Y(n_434)
);

INVx5_ASAP7_75t_L g435 ( 
.A(n_364),
.Y(n_435)
);

BUFx12f_ASAP7_75t_L g436 ( 
.A(n_419),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_356),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_389),
.Y(n_438)
);

NOR3xp33_ASAP7_75t_SL g439 ( 
.A(n_376),
.B(n_339),
.C(n_340),
.Y(n_439)
);

INVx4_ASAP7_75t_L g440 ( 
.A(n_359),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_422),
.A2(n_303),
.B1(n_333),
.B2(n_334),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_357),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_403),
.A2(n_313),
.B1(n_315),
.B2(n_43),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_361),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_413),
.B(n_315),
.Y(n_445)
);

O2A1O1Ixp33_ASAP7_75t_SL g446 ( 
.A1(n_390),
.A2(n_315),
.B(n_41),
.C(n_44),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_367),
.B(n_363),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_398),
.B(n_315),
.Y(n_448)
);

A2O1A1Ixp33_ASAP7_75t_L g449 ( 
.A1(n_375),
.A2(n_315),
.B(n_49),
.C(n_51),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_400),
.Y(n_450)
);

INVx4_ASAP7_75t_L g451 ( 
.A(n_359),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_377),
.B(n_315),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_355),
.B(n_40),
.Y(n_453)
);

AND2x2_ASAP7_75t_SL g454 ( 
.A(n_396),
.B(n_53),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_358),
.B(n_56),
.Y(n_455)
);

INVx5_ASAP7_75t_L g456 ( 
.A(n_364),
.Y(n_456)
);

O2A1O1Ixp5_ASAP7_75t_L g457 ( 
.A1(n_381),
.A2(n_57),
.B(n_58),
.C(n_60),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_373),
.A2(n_61),
.B(n_63),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_371),
.B(n_65),
.Y(n_459)
);

INVx4_ASAP7_75t_L g460 ( 
.A(n_359),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_384),
.B(n_66),
.Y(n_461)
);

OR2x6_ASAP7_75t_L g462 ( 
.A(n_364),
.B(n_67),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_363),
.B(n_68),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_360),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_408),
.A2(n_72),
.B(n_73),
.Y(n_465)
);

BUFx2_ASAP7_75t_L g466 ( 
.A(n_406),
.Y(n_466)
);

OR2x6_ASAP7_75t_L g467 ( 
.A(n_416),
.B(n_74),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_369),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_396),
.B(n_75),
.Y(n_469)
);

A2O1A1Ixp33_ASAP7_75t_L g470 ( 
.A1(n_417),
.A2(n_76),
.B(n_78),
.C(n_79),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_392),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_366),
.B(n_80),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_360),
.A2(n_81),
.B1(n_83),
.B2(n_88),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_416),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_369),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_401),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_420),
.A2(n_89),
.B1(n_92),
.B2(n_95),
.Y(n_477)
);

AO21x1_ASAP7_75t_L g478 ( 
.A1(n_423),
.A2(n_97),
.B(n_98),
.Y(n_478)
);

A2O1A1Ixp33_ASAP7_75t_SL g479 ( 
.A1(n_415),
.A2(n_100),
.B(n_101),
.C(n_102),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_416),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_402),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_405),
.A2(n_103),
.B1(n_104),
.B2(n_108),
.Y(n_482)
);

AND2x4_ASAP7_75t_L g483 ( 
.A(n_435),
.B(n_393),
.Y(n_483)
);

OAI21x1_ASAP7_75t_L g484 ( 
.A1(n_433),
.A2(n_390),
.B(n_394),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_427),
.B(n_379),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_436),
.Y(n_486)
);

OAI21x1_ASAP7_75t_L g487 ( 
.A1(n_455),
.A2(n_387),
.B(n_404),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_431),
.B(n_378),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_468),
.Y(n_489)
);

AO21x1_ASAP7_75t_L g490 ( 
.A1(n_432),
.A2(n_411),
.B(n_378),
.Y(n_490)
);

OAI21x1_ASAP7_75t_SL g491 ( 
.A1(n_478),
.A2(n_411),
.B(n_407),
.Y(n_491)
);

AO21x2_ASAP7_75t_L g492 ( 
.A1(n_459),
.A2(n_418),
.B(n_391),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_435),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_440),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_424),
.Y(n_495)
);

AOI21x1_ASAP7_75t_L g496 ( 
.A1(n_461),
.A2(n_386),
.B(n_365),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_435),
.B(n_409),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_456),
.Y(n_498)
);

NAND2x1p5_ASAP7_75t_L g499 ( 
.A(n_456),
.B(n_380),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_428),
.Y(n_500)
);

OAI21x1_ASAP7_75t_L g501 ( 
.A1(n_465),
.A2(n_362),
.B(n_380),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_430),
.Y(n_502)
);

INVxp67_ASAP7_75t_SL g503 ( 
.A(n_440),
.Y(n_503)
);

INVx6_ASAP7_75t_L g504 ( 
.A(n_456),
.Y(n_504)
);

INVx3_ASAP7_75t_SL g505 ( 
.A(n_467),
.Y(n_505)
);

OAI21x1_ASAP7_75t_L g506 ( 
.A1(n_457),
.A2(n_362),
.B(n_380),
.Y(n_506)
);

OAI21x1_ASAP7_75t_SL g507 ( 
.A1(n_473),
.A2(n_412),
.B(n_362),
.Y(n_507)
);

OR2x2_ASAP7_75t_L g508 ( 
.A(n_438),
.B(n_419),
.Y(n_508)
);

INVx1_ASAP7_75t_SL g509 ( 
.A(n_466),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_475),
.Y(n_510)
);

OR2x6_ASAP7_75t_L g511 ( 
.A(n_462),
.B(n_412),
.Y(n_511)
);

INVx4_ASAP7_75t_L g512 ( 
.A(n_451),
.Y(n_512)
);

INVx1_ASAP7_75t_SL g513 ( 
.A(n_474),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_451),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_437),
.Y(n_515)
);

BUFx2_ASAP7_75t_SL g516 ( 
.A(n_460),
.Y(n_516)
);

OAI21x1_ASAP7_75t_L g517 ( 
.A1(n_445),
.A2(n_109),
.B(n_110),
.Y(n_517)
);

AO21x2_ASAP7_75t_L g518 ( 
.A1(n_429),
.A2(n_112),
.B(n_113),
.Y(n_518)
);

OAI21x1_ASAP7_75t_L g519 ( 
.A1(n_464),
.A2(n_115),
.B(n_116),
.Y(n_519)
);

BUFx2_ASAP7_75t_SL g520 ( 
.A(n_460),
.Y(n_520)
);

NOR2x1_ASAP7_75t_R g521 ( 
.A(n_447),
.B(n_117),
.Y(n_521)
);

AND2x6_ASAP7_75t_L g522 ( 
.A(n_473),
.B(n_118),
.Y(n_522)
);

OR3x4_ASAP7_75t_SL g523 ( 
.A(n_425),
.B(n_119),
.C(n_120),
.Y(n_523)
);

INVx2_ASAP7_75t_SL g524 ( 
.A(n_480),
.Y(n_524)
);

INVx1_ASAP7_75t_SL g525 ( 
.A(n_442),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_450),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_462),
.Y(n_527)
);

OAI21x1_ASAP7_75t_L g528 ( 
.A1(n_463),
.A2(n_121),
.B(n_127),
.Y(n_528)
);

AOI21x1_ASAP7_75t_L g529 ( 
.A1(n_441),
.A2(n_128),
.B(n_129),
.Y(n_529)
);

BUFx12f_ASAP7_75t_L g530 ( 
.A(n_467),
.Y(n_530)
);

BUFx8_ASAP7_75t_SL g531 ( 
.A(n_486),
.Y(n_531)
);

AOI22xp33_ASAP7_75t_L g532 ( 
.A1(n_522),
.A2(n_425),
.B1(n_426),
.B2(n_443),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_500),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_502),
.Y(n_534)
);

AO21x1_ASAP7_75t_L g535 ( 
.A1(n_529),
.A2(n_448),
.B(n_477),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_515),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_488),
.B(n_434),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_515),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_526),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_489),
.Y(n_540)
);

AOI22xp33_ASAP7_75t_L g541 ( 
.A1(n_522),
.A2(n_426),
.B1(n_454),
.B2(n_447),
.Y(n_541)
);

AOI22xp33_ASAP7_75t_L g542 ( 
.A1(n_522),
.A2(n_467),
.B1(n_453),
.B2(n_444),
.Y(n_542)
);

AO21x1_ASAP7_75t_L g543 ( 
.A1(n_519),
.A2(n_448),
.B(n_482),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_485),
.B(n_469),
.Y(n_544)
);

OAI21x1_ASAP7_75t_L g545 ( 
.A1(n_501),
.A2(n_458),
.B(n_481),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_SL g546 ( 
.A1(n_522),
.A2(n_472),
.B1(n_462),
.B2(n_452),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_495),
.Y(n_547)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_495),
.Y(n_548)
);

BUFx4f_ASAP7_75t_SL g549 ( 
.A(n_486),
.Y(n_549)
);

HB1xp67_ASAP7_75t_SL g550 ( 
.A(n_527),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_489),
.Y(n_551)
);

OAI22xp33_ASAP7_75t_SL g552 ( 
.A1(n_523),
.A2(n_482),
.B1(n_471),
.B2(n_476),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_510),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_514),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_510),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_514),
.Y(n_556)
);

CKINVDCx11_ASAP7_75t_R g557 ( 
.A(n_509),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_496),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_514),
.Y(n_559)
);

OR2x6_ASAP7_75t_L g560 ( 
.A(n_511),
.B(n_507),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_501),
.Y(n_561)
);

AO21x2_ASAP7_75t_L g562 ( 
.A1(n_484),
.A2(n_449),
.B(n_479),
.Y(n_562)
);

BUFx2_ASAP7_75t_L g563 ( 
.A(n_503),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_L g564 ( 
.A1(n_522),
.A2(n_481),
.B1(n_476),
.B2(n_439),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_517),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_525),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_506),
.Y(n_567)
);

INVx2_ASAP7_75t_SL g568 ( 
.A(n_514),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_506),
.Y(n_569)
);

BUFx3_ASAP7_75t_L g570 ( 
.A(n_504),
.Y(n_570)
);

BUFx2_ASAP7_75t_L g571 ( 
.A(n_503),
.Y(n_571)
);

BUFx3_ASAP7_75t_L g572 ( 
.A(n_504),
.Y(n_572)
);

INVx4_ASAP7_75t_L g573 ( 
.A(n_554),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_537),
.B(n_488),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_536),
.Y(n_575)
);

CKINVDCx16_ASAP7_75t_R g576 ( 
.A(n_550),
.Y(n_576)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_544),
.B(n_566),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_547),
.Y(n_578)
);

NAND2xp33_ASAP7_75t_R g579 ( 
.A(n_544),
.B(n_508),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_533),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_548),
.B(n_513),
.Y(n_581)
);

HB1xp67_ASAP7_75t_L g582 ( 
.A(n_563),
.Y(n_582)
);

BUFx3_ASAP7_75t_L g583 ( 
.A(n_557),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_533),
.B(n_524),
.Y(n_584)
);

AND2x4_ASAP7_75t_L g585 ( 
.A(n_570),
.B(n_527),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_532),
.B(n_490),
.Y(n_586)
);

NAND2xp33_ASAP7_75t_R g587 ( 
.A(n_560),
.B(n_511),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_536),
.Y(n_588)
);

AND2x2_ASAP7_75t_L g589 ( 
.A(n_534),
.B(n_505),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_R g590 ( 
.A(n_549),
.B(n_504),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_570),
.B(n_572),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_SL g592 ( 
.A1(n_552),
.A2(n_530),
.B1(n_523),
.B2(n_511),
.Y(n_592)
);

NAND2x1_ASAP7_75t_L g593 ( 
.A(n_563),
.B(n_494),
.Y(n_593)
);

BUFx10_ASAP7_75t_L g594 ( 
.A(n_554),
.Y(n_594)
);

NAND2x1_ASAP7_75t_L g595 ( 
.A(n_571),
.B(n_494),
.Y(n_595)
);

AOI21xp33_ASAP7_75t_L g596 ( 
.A1(n_552),
.A2(n_491),
.B(n_519),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_534),
.B(n_505),
.Y(n_597)
);

A2O1A1Ixp33_ASAP7_75t_L g598 ( 
.A1(n_541),
.A2(n_484),
.B(n_470),
.C(n_483),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_539),
.B(n_492),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_539),
.B(n_483),
.Y(n_600)
);

INVxp67_ASAP7_75t_L g601 ( 
.A(n_570),
.Y(n_601)
);

OR2x6_ASAP7_75t_L g602 ( 
.A(n_560),
.B(n_530),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_546),
.A2(n_483),
.B1(n_518),
.B2(n_493),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_538),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_538),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_572),
.B(n_493),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_571),
.B(n_492),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_542),
.B(n_497),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_531),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_554),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_551),
.Y(n_611)
);

O2A1O1Ixp33_ASAP7_75t_L g612 ( 
.A1(n_543),
.A2(n_446),
.B(n_518),
.C(n_499),
.Y(n_612)
);

AOI21xp33_ASAP7_75t_L g613 ( 
.A1(n_543),
.A2(n_487),
.B(n_521),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_572),
.B(n_520),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_554),
.Y(n_615)
);

NAND2xp33_ASAP7_75t_SL g616 ( 
.A(n_554),
.B(n_498),
.Y(n_616)
);

AND2x4_ASAP7_75t_SL g617 ( 
.A(n_554),
.B(n_498),
.Y(n_617)
);

OR2x6_ASAP7_75t_L g618 ( 
.A(n_560),
.B(n_498),
.Y(n_618)
);

OR2x6_ASAP7_75t_L g619 ( 
.A(n_560),
.B(n_498),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_540),
.B(n_497),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_551),
.B(n_516),
.Y(n_621)
);

INVx5_ASAP7_75t_L g622 ( 
.A(n_618),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_599),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_599),
.Y(n_624)
);

HB1xp67_ASAP7_75t_L g625 ( 
.A(n_578),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_582),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_580),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_602),
.B(n_560),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_574),
.B(n_569),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_604),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_605),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_577),
.B(n_569),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_575),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_586),
.B(n_561),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_607),
.Y(n_635)
);

AND2x4_ASAP7_75t_L g636 ( 
.A(n_602),
.B(n_556),
.Y(n_636)
);

HB1xp67_ASAP7_75t_L g637 ( 
.A(n_600),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_607),
.B(n_561),
.Y(n_638)
);

AOI21xp5_ASAP7_75t_L g639 ( 
.A1(n_598),
.A2(n_535),
.B(n_564),
.Y(n_639)
);

BUFx2_ASAP7_75t_L g640 ( 
.A(n_618),
.Y(n_640)
);

OR2x2_ASAP7_75t_L g641 ( 
.A(n_602),
.B(n_567),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_588),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_611),
.B(n_567),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_610),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_610),
.B(n_555),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_592),
.B(n_555),
.Y(n_646)
);

AND2x4_ASAP7_75t_L g647 ( 
.A(n_618),
.B(n_556),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_584),
.B(n_553),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_581),
.B(n_553),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_608),
.A2(n_535),
.B1(n_540),
.B2(n_565),
.Y(n_650)
);

OR2x2_ASAP7_75t_L g651 ( 
.A(n_608),
.B(n_558),
.Y(n_651)
);

BUFx2_ASAP7_75t_L g652 ( 
.A(n_619),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_620),
.B(n_558),
.Y(n_653)
);

OR2x2_ASAP7_75t_L g654 ( 
.A(n_619),
.B(n_562),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_620),
.B(n_556),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_589),
.B(n_556),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_615),
.Y(n_657)
);

OR2x2_ASAP7_75t_L g658 ( 
.A(n_619),
.B(n_562),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_597),
.B(n_559),
.Y(n_659)
);

BUFx2_ASAP7_75t_L g660 ( 
.A(n_573),
.Y(n_660)
);

AND2x2_ASAP7_75t_L g661 ( 
.A(n_596),
.B(n_559),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_612),
.Y(n_662)
);

OR2x2_ASAP7_75t_L g663 ( 
.A(n_635),
.B(n_596),
.Y(n_663)
);

AND2x4_ASAP7_75t_L g664 ( 
.A(n_628),
.B(n_573),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_627),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_625),
.B(n_632),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_632),
.B(n_576),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_630),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_630),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_628),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_627),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_638),
.B(n_613),
.Y(n_672)
);

OR2x2_ASAP7_75t_L g673 ( 
.A(n_651),
.B(n_603),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_631),
.Y(n_674)
);

AOI22xp33_ASAP7_75t_L g675 ( 
.A1(n_639),
.A2(n_583),
.B1(n_613),
.B2(n_585),
.Y(n_675)
);

INVx5_ASAP7_75t_L g676 ( 
.A(n_622),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_638),
.B(n_562),
.Y(n_677)
);

OR2x2_ASAP7_75t_L g678 ( 
.A(n_651),
.B(n_635),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_631),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_626),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_623),
.Y(n_681)
);

INVx1_ASAP7_75t_SL g682 ( 
.A(n_656),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_643),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_662),
.A2(n_585),
.B1(n_591),
.B2(n_606),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_655),
.B(n_601),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_623),
.Y(n_686)
);

INVxp67_ASAP7_75t_L g687 ( 
.A(n_649),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_661),
.B(n_615),
.Y(n_688)
);

OR2x2_ASAP7_75t_L g689 ( 
.A(n_663),
.B(n_624),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_688),
.B(n_661),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_668),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_669),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_665),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_665),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_687),
.B(n_629),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_680),
.B(n_629),
.Y(n_696)
);

BUFx3_ASAP7_75t_L g697 ( 
.A(n_664),
.Y(n_697)
);

OAI21x1_ASAP7_75t_L g698 ( 
.A1(n_675),
.A2(n_662),
.B(n_545),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_688),
.B(n_654),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_667),
.B(n_659),
.Y(n_700)
);

HB1xp67_ASAP7_75t_L g701 ( 
.A(n_678),
.Y(n_701)
);

NOR2x1p5_ASAP7_75t_L g702 ( 
.A(n_670),
.B(n_609),
.Y(n_702)
);

CKINVDCx20_ASAP7_75t_R g703 ( 
.A(n_666),
.Y(n_703)
);

OR2x2_ASAP7_75t_L g704 ( 
.A(n_663),
.B(n_624),
.Y(n_704)
);

AND2x4_ASAP7_75t_L g705 ( 
.A(n_697),
.B(n_699),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_691),
.Y(n_706)
);

INVx1_ASAP7_75t_SL g707 ( 
.A(n_689),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_701),
.B(n_672),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_695),
.B(n_672),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_700),
.B(n_685),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_692),
.Y(n_711)
);

NAND2x1_ASAP7_75t_SL g712 ( 
.A(n_690),
.B(n_670),
.Y(n_712)
);

OAI22xp5_ASAP7_75t_L g713 ( 
.A1(n_703),
.A2(n_675),
.B1(n_684),
.B2(n_673),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_693),
.Y(n_714)
);

AOI21xp33_ASAP7_75t_L g715 ( 
.A1(n_713),
.A2(n_579),
.B(n_704),
.Y(n_715)
);

NAND3xp33_ASAP7_75t_L g716 ( 
.A(n_706),
.B(n_684),
.C(n_704),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_711),
.Y(n_717)
);

OAI21xp33_ASAP7_75t_L g718 ( 
.A1(n_709),
.A2(n_696),
.B(n_689),
.Y(n_718)
);

OR2x2_ASAP7_75t_L g719 ( 
.A(n_708),
.B(n_690),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_L g720 ( 
.A1(n_715),
.A2(n_628),
.B1(n_710),
.B2(n_703),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_718),
.B(n_705),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_717),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_719),
.Y(n_723)
);

OAI211xp5_ASAP7_75t_SL g724 ( 
.A1(n_716),
.A2(n_707),
.B(n_714),
.C(n_694),
.Y(n_724)
);

OAI222xp33_ASAP7_75t_L g725 ( 
.A1(n_719),
.A2(n_707),
.B1(n_705),
.B2(n_670),
.C1(n_682),
.C2(n_699),
.Y(n_725)
);

OAI211xp5_ASAP7_75t_L g726 ( 
.A1(n_720),
.A2(n_724),
.B(n_722),
.C(n_721),
.Y(n_726)
);

OAI322xp33_ASAP7_75t_L g727 ( 
.A1(n_723),
.A2(n_686),
.A3(n_681),
.B1(n_674),
.B2(n_671),
.C1(n_683),
.C2(n_654),
.Y(n_727)
);

AOI21xp5_ASAP7_75t_L g728 ( 
.A1(n_720),
.A2(n_698),
.B(n_646),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_725),
.B(n_712),
.Y(n_729)
);

AOI21xp5_ASAP7_75t_L g730 ( 
.A1(n_726),
.A2(n_728),
.B(n_729),
.Y(n_730)
);

A2O1A1Ixp33_ASAP7_75t_L g731 ( 
.A1(n_727),
.A2(n_702),
.B(n_698),
.C(n_697),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_730),
.Y(n_732)
);

OAI221xp5_ASAP7_75t_L g733 ( 
.A1(n_731),
.A2(n_587),
.B1(n_650),
.B2(n_652),
.C(n_640),
.Y(n_733)
);

AOI221x1_ASAP7_75t_L g734 ( 
.A1(n_730),
.A2(n_616),
.B1(n_621),
.B2(n_657),
.C(n_591),
.Y(n_734)
);

OAI211xp5_ASAP7_75t_L g735 ( 
.A1(n_732),
.A2(n_590),
.B(n_614),
.C(n_646),
.Y(n_735)
);

NOR2x1_ASAP7_75t_L g736 ( 
.A(n_733),
.B(n_734),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_732),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_732),
.Y(n_738)
);

AOI22xp5_ASAP7_75t_L g739 ( 
.A1(n_732),
.A2(n_664),
.B1(n_636),
.B2(n_656),
.Y(n_739)
);

NOR2x1_ASAP7_75t_L g740 ( 
.A(n_732),
.B(n_512),
.Y(n_740)
);

OAI211xp5_ASAP7_75t_L g741 ( 
.A1(n_736),
.A2(n_676),
.B(n_622),
.C(n_648),
.Y(n_741)
);

OAI22xp5_ASAP7_75t_L g742 ( 
.A1(n_739),
.A2(n_676),
.B1(n_622),
.B2(n_640),
.Y(n_742)
);

NOR3xp33_ASAP7_75t_L g743 ( 
.A(n_737),
.B(n_559),
.C(n_512),
.Y(n_743)
);

OAI221xp5_ASAP7_75t_L g744 ( 
.A1(n_735),
.A2(n_676),
.B1(n_652),
.B2(n_622),
.C(n_658),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_738),
.Y(n_745)
);

AOI221xp5_ASAP7_75t_L g746 ( 
.A1(n_740),
.A2(n_648),
.B1(n_636),
.B2(n_660),
.C(n_647),
.Y(n_746)
);

NAND3xp33_ASAP7_75t_L g747 ( 
.A(n_736),
.B(n_657),
.C(n_615),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_745),
.B(n_743),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_747),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_742),
.Y(n_750)
);

AOI222xp33_ASAP7_75t_L g751 ( 
.A1(n_741),
.A2(n_676),
.B1(n_636),
.B2(n_528),
.C1(n_622),
.C2(n_660),
.Y(n_751)
);

HB1xp67_ASAP7_75t_L g752 ( 
.A(n_744),
.Y(n_752)
);

INVx1_ASAP7_75t_SL g753 ( 
.A(n_746),
.Y(n_753)
);

INVxp67_ASAP7_75t_SL g754 ( 
.A(n_752),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_749),
.Y(n_755)
);

XNOR2xp5_ASAP7_75t_L g756 ( 
.A(n_753),
.B(n_664),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_748),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_750),
.A2(n_751),
.B1(n_676),
.B2(n_647),
.Y(n_758)
);

INVxp67_ASAP7_75t_L g759 ( 
.A(n_752),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_749),
.Y(n_760)
);

AO22x2_ASAP7_75t_L g761 ( 
.A1(n_753),
.A2(n_568),
.B1(n_559),
.B2(n_647),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_L g762 ( 
.A1(n_759),
.A2(n_754),
.B1(n_760),
.B2(n_755),
.Y(n_762)
);

AOI22xp5_ASAP7_75t_L g763 ( 
.A1(n_756),
.A2(n_757),
.B1(n_758),
.B2(n_761),
.Y(n_763)
);

OAI31xp33_ASAP7_75t_L g764 ( 
.A1(n_759),
.A2(n_617),
.A3(n_499),
.B(n_568),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_754),
.A2(n_655),
.B1(n_644),
.B2(n_677),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_761),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_754),
.A2(n_644),
.B1(n_677),
.B2(n_637),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_SL g768 ( 
.A1(n_754),
.A2(n_497),
.B1(n_645),
.B2(n_679),
.Y(n_768)
);

OAI31xp33_ASAP7_75t_L g769 ( 
.A1(n_759),
.A2(n_658),
.A3(n_641),
.B(n_565),
.Y(n_769)
);

OAI22xp5_ASAP7_75t_L g770 ( 
.A1(n_762),
.A2(n_641),
.B1(n_679),
.B2(n_683),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_SL g771 ( 
.A1(n_763),
.A2(n_595),
.B1(n_593),
.B2(n_642),
.Y(n_771)
);

OAI221xp5_ASAP7_75t_L g772 ( 
.A1(n_764),
.A2(n_642),
.B1(n_633),
.B2(n_653),
.C(n_645),
.Y(n_772)
);

AOI22x1_ASAP7_75t_L g773 ( 
.A1(n_766),
.A2(n_633),
.B1(n_130),
.B2(n_132),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_R g774 ( 
.A1(n_771),
.A2(n_768),
.B1(n_769),
.B2(n_765),
.Y(n_774)
);

INVxp67_ASAP7_75t_L g775 ( 
.A(n_773),
.Y(n_775)
);

NAND3xp33_ASAP7_75t_SL g776 ( 
.A(n_775),
.B(n_767),
.C(n_772),
.Y(n_776)
);

AOI22xp5_ASAP7_75t_SL g777 ( 
.A1(n_776),
.A2(n_770),
.B1(n_774),
.B2(n_594),
.Y(n_777)
);

OR2x6_ASAP7_75t_L g778 ( 
.A(n_777),
.B(n_528),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_778),
.A2(n_594),
.B1(n_653),
.B2(n_634),
.Y(n_779)
);


endmodule