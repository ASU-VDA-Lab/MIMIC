module fake_jpeg_20198_n_164 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_164);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx4f_ASAP7_75t_SL g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx24_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_34),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_8),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_38),
.Y(n_60)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_20),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx8_ASAP7_75t_L g64 ( 
.A(n_13),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVxp33_ASAP7_75t_L g69 ( 
.A(n_14),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_44),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_24),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_3),
.Y(n_72)
);

INVx8_ASAP7_75t_SL g73 ( 
.A(n_1),
.Y(n_73)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_16),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_46),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_15),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_19),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

BUFx16f_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_81),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_73),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_85),
.A2(n_61),
.B1(n_56),
.B2(n_53),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_86),
.A2(n_87),
.B1(n_64),
.B2(n_54),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_81),
.A2(n_69),
.B1(n_74),
.B2(n_75),
.Y(n_87)
);

O2A1O1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_80),
.A2(n_57),
.B(n_69),
.C(n_55),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_58),
.Y(n_103)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_96),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_75),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_97),
.B(n_108),
.Y(n_116)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_99),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g100 ( 
.A(n_88),
.B(n_71),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_58),
.C(n_54),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_95),
.B(n_60),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_101),
.B(n_105),
.Y(n_111)
);

OA22x2_ASAP7_75t_L g122 ( 
.A1(n_102),
.A2(n_49),
.B1(n_52),
.B2(n_72),
.Y(n_122)
);

NAND3xp33_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_47),
.C(n_51),
.Y(n_112)
);

OR2x2_ASAP7_75t_SL g104 ( 
.A(n_86),
.B(n_64),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_104),
.A2(n_107),
.B(n_59),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_77),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_94),
.A2(n_63),
.B(n_70),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_93),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_92),
.A2(n_52),
.B1(n_68),
.B2(n_66),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_109),
.A2(n_48),
.B1(n_62),
.B2(n_2),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_98),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_110),
.B(n_115),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_118),
.Y(n_139)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_109),
.Y(n_114)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_100),
.Y(n_117)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_119),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_106),
.Y(n_120)
);

BUFx24_ASAP7_75t_SL g127 ( 
.A(n_120),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_104),
.A2(n_92),
.B1(n_49),
.B2(n_65),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_121),
.A2(n_122),
.B1(n_3),
.B2(n_4),
.Y(n_133)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_123),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_0),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_124),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_125),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_126),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_116),
.A2(n_0),
.B(n_1),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_9),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_122),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_135),
.A2(n_140),
.B1(n_122),
.B2(n_113),
.Y(n_144)
);

AND2x4_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_5),
.Y(n_137)
);

OAI32xp33_ASAP7_75t_L g147 ( 
.A1(n_137),
.A2(n_112),
.A3(n_10),
.B1(n_11),
.B2(n_9),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_126),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_142),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_111),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_143),
.A2(n_144),
.B(n_145),
.Y(n_149)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_138),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_146),
.A2(n_147),
.B(n_148),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_149),
.A2(n_144),
.B1(n_137),
.B2(n_130),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_152),
.A2(n_150),
.B1(n_137),
.B2(n_147),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_153),
.A2(n_151),
.B(n_131),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_154),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_155),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_139),
.B1(n_127),
.B2(n_132),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_136),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_139),
.Y(n_159)
);

AOI321xp33_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_10),
.A3(n_12),
.B1(n_21),
.B2(n_25),
.C(n_26),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_27),
.B(n_28),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_161),
.A2(n_30),
.B(n_31),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_32),
.B(n_35),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_163),
.Y(n_164)
);


endmodule