module fake_jpeg_26463_n_59 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_59);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_59;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx12_ASAP7_75t_L g8 ( 
.A(n_7),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g9 ( 
.A(n_4),
.B(n_6),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_5),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_SL g14 ( 
.A(n_0),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

AOI21xp33_ASAP7_75t_SL g16 ( 
.A1(n_14),
.A2(n_1),
.B(n_2),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_16),
.B(n_17),
.Y(n_23)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_19),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_9),
.B(n_1),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_20),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_20),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_22),
.B(n_14),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_17),
.A2(n_15),
.B1(n_10),
.B2(n_12),
.Y(n_25)
);

OA22x2_ASAP7_75t_L g31 ( 
.A1(n_25),
.A2(n_15),
.B1(n_12),
.B2(n_8),
.Y(n_31)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_30),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_27),
.B(n_28),
.Y(n_35)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_13),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_31),
.A2(n_21),
.B(n_11),
.Y(n_36)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_34),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_31),
.B1(n_8),
.B2(n_18),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_11),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_28),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_41),
.Y(n_45)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_42),
.A2(n_31),
.B1(n_12),
.B2(n_6),
.Y(n_47)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_38),
.C(n_34),
.Y(n_44)
);

FAx1_ASAP7_75t_SL g46 ( 
.A(n_44),
.B(n_31),
.CI(n_13),
.CON(n_46),
.SN(n_46)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_39),
.C(n_2),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_47),
.A2(n_44),
.B1(n_40),
.B2(n_7),
.Y(n_49)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_51),
.C(n_45),
.Y(n_53)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_46),
.Y(n_51)
);

A2O1A1Ixp33_ASAP7_75t_SL g55 ( 
.A1(n_53),
.A2(n_50),
.B(n_48),
.C(n_3),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_52),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_55),
.Y(n_56)
);

INVxp33_ASAP7_75t_L g57 ( 
.A(n_56),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_48),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_3),
.Y(n_59)
);


endmodule