module fake_jpeg_24350_n_256 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_256);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_256;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_9),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_38),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_34),
.A2(n_28),
.B1(n_25),
.B2(n_27),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_49),
.B1(n_57),
.B2(n_36),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_26),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_18),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_34),
.A2(n_28),
.B1(n_22),
.B2(n_23),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_44),
.A2(n_52),
.B(n_29),
.C(n_37),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_26),
.Y(n_47)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_34),
.A2(n_25),
.B1(n_27),
.B2(n_22),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_22),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_23),
.Y(n_53)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_22),
.C(n_31),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_54),
.B(n_16),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_36),
.A2(n_25),
.B1(n_22),
.B2(n_18),
.Y(n_57)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_59),
.B(n_65),
.Y(n_91)
);

OAI22x1_ASAP7_75t_L g111 ( 
.A1(n_60),
.A2(n_29),
.B1(n_16),
.B2(n_3),
.Y(n_111)
);

OAI21xp33_ASAP7_75t_L g87 ( 
.A1(n_61),
.A2(n_83),
.B(n_26),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_43),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_62),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_44),
.A2(n_35),
.B1(n_25),
.B2(n_18),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_63),
.A2(n_56),
.B1(n_48),
.B2(n_23),
.Y(n_94)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_66),
.A2(n_85),
.B(n_36),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_68),
.Y(n_93)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx4_ASAP7_75t_SL g69 ( 
.A(n_51),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_70),
.Y(n_98)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_33),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_78),
.Y(n_100)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_52),
.A2(n_17),
.B1(n_32),
.B2(n_31),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_74),
.A2(n_30),
.B1(n_19),
.B2(n_21),
.Y(n_108)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_75),
.Y(n_101)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_16),
.Y(n_77)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_33),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_50),
.B(n_33),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_80),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_33),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_16),
.Y(n_81)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_55),
.B(n_39),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_55),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_41),
.B(n_17),
.Y(n_83)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_84),
.A2(n_48),
.B1(n_56),
.B2(n_86),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_87),
.B(n_108),
.Y(n_137)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_88),
.B(n_105),
.Y(n_120)
);

OAI21xp33_ASAP7_75t_L g92 ( 
.A1(n_78),
.A2(n_1),
.B(n_2),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_92),
.A2(n_102),
.B(n_110),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_94),
.A2(n_109),
.B1(n_111),
.B2(n_65),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_73),
.A2(n_63),
.B1(n_85),
.B2(n_60),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_95),
.A2(n_72),
.B1(n_64),
.B2(n_79),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_SL g102 ( 
.A1(n_67),
.A2(n_29),
.B(n_36),
.C(n_48),
.Y(n_102)
);

BUFx4f_ASAP7_75t_SL g103 ( 
.A(n_68),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_64),
.C(n_82),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_106),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_90),
.B(n_61),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_113),
.B(n_133),
.Y(n_142)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_114),
.B(n_119),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_71),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_116),
.B(n_134),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_117),
.A2(n_135),
.B1(n_112),
.B2(n_97),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_118),
.B(n_112),
.Y(n_150)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_96),
.A2(n_84),
.B1(n_75),
.B2(n_58),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_121),
.A2(n_123),
.B1(n_138),
.B2(n_30),
.Y(n_165)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_122),
.B(n_124),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_96),
.A2(n_58),
.B1(n_70),
.B2(n_86),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_103),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_126),
.Y(n_144)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_127),
.B(n_131),
.Y(n_158)
);

NAND2xp33_ASAP7_75t_SL g128 ( 
.A(n_111),
.B(n_83),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_128),
.A2(n_130),
.B(n_102),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_100),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_129),
.Y(n_147)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_88),
.B(n_76),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_102),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_139),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_107),
.A2(n_59),
.B1(n_39),
.B2(n_37),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_89),
.B(n_39),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_139),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_145),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_115),
.A2(n_110),
.B(n_89),
.Y(n_141)
);

NOR2x1_ASAP7_75t_R g183 ( 
.A(n_141),
.B(n_153),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_102),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_137),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_151),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_162),
.C(n_119),
.Y(n_169)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_120),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_115),
.A2(n_97),
.B(n_101),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_157),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_134),
.A2(n_136),
.B(n_116),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_155),
.A2(n_161),
.B1(n_164),
.B2(n_24),
.Y(n_178)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_138),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_159),
.B(n_160),
.Y(n_179)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_123),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_131),
.A2(n_105),
.B(n_99),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_118),
.B(n_117),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_132),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_165),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_127),
.A2(n_99),
.B1(n_37),
.B2(n_32),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_113),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_166),
.Y(n_174)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_161),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_172),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_169),
.B(n_175),
.C(n_142),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_144),
.Y(n_172)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_173),
.Y(n_197)
);

A2O1A1O1Ixp25_ASAP7_75t_L g175 ( 
.A1(n_141),
.A2(n_122),
.B(n_125),
.C(n_114),
.D(n_126),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_176),
.B(n_177),
.Y(n_194)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_158),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_178),
.A2(n_181),
.B1(n_187),
.B2(n_188),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_148),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_180),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_152),
.A2(n_24),
.B1(n_21),
.B2(n_19),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_147),
.B(n_1),
.Y(n_184)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_184),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_147),
.B(n_140),
.Y(n_185)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_185),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_2),
.Y(n_186)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_186),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_152),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_156),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_170),
.A2(n_160),
.B1(n_157),
.B2(n_159),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_190),
.A2(n_206),
.B1(n_173),
.B2(n_185),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_162),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_195),
.Y(n_217)
);

NOR3xp33_ASAP7_75t_SL g193 ( 
.A(n_174),
.B(n_166),
.C(n_153),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_198),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_150),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_145),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_199),
.C(n_202),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_171),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_164),
.Y(n_201)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_201),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_155),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_167),
.A2(n_156),
.B1(n_165),
.B2(n_146),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_206),
.A2(n_189),
.B(n_197),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_209),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_204),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_210),
.A2(n_214),
.B1(n_218),
.B2(n_207),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_211),
.B(n_212),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_190),
.A2(n_179),
.B1(n_192),
.B2(n_202),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_212),
.A2(n_215),
.B1(n_199),
.B2(n_195),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_184),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_213),
.B(n_216),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_200),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_192),
.A2(n_149),
.B1(n_177),
.B2(n_182),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_180),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_SL g218 ( 
.A1(n_196),
.A2(n_178),
.B(n_176),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_203),
.A2(n_151),
.B1(n_172),
.B2(n_175),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_219),
.A2(n_187),
.B1(n_188),
.B2(n_181),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_191),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_221),
.B(n_224),
.C(n_230),
.Y(n_235)
);

NAND4xp25_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_208),
.C(n_219),
.D(n_163),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_222),
.A2(n_6),
.B(n_8),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_225),
.B(n_227),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_228),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_209),
.B(n_205),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_211),
.B(n_217),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_4),
.C(n_6),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_224),
.C(n_229),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_228),
.A2(n_220),
.B(n_7),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_234),
.B(n_12),
.Y(n_244)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_236),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_237),
.B(n_221),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_8),
.C(n_9),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_238),
.B(n_11),
.Y(n_241)
);

NOR2xp67_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_10),
.Y(n_239)
);

XOR2x2_ASAP7_75t_L g242 ( 
.A(n_239),
.B(n_223),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_13),
.C(n_14),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_241),
.B(n_245),
.Y(n_248)
);

A2O1A1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_242),
.A2(n_233),
.B(n_239),
.C(n_232),
.Y(n_246)
);

AO21x1_ASAP7_75t_L g249 ( 
.A1(n_244),
.A2(n_13),
.B(n_14),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_12),
.Y(n_245)
);

NAND3xp33_ASAP7_75t_SL g252 ( 
.A(n_246),
.B(n_247),
.C(n_249),
.Y(n_252)
);

A2O1A1Ixp33_ASAP7_75t_L g250 ( 
.A1(n_248),
.A2(n_244),
.B(n_243),
.C(n_15),
.Y(n_250)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_250),
.Y(n_253)
);

AOI21x1_ASAP7_75t_L g251 ( 
.A1(n_246),
.A2(n_13),
.B(n_14),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_251),
.B(n_15),
.C(n_252),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_254),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_253),
.Y(n_256)
);


endmodule