module fake_jpeg_2457_n_55 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_55);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_55;

wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

AND2x2_ASAP7_75t_L g16 ( 
.A(n_2),
.B(n_12),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_19),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_20),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_19),
.A2(n_14),
.B1(n_13),
.B2(n_10),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g29 ( 
.A1(n_23),
.A2(n_16),
.B(n_20),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_20),
.Y(n_25)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_16),
.B(n_22),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_SL g32 ( 
.A1(n_28),
.A2(n_16),
.B(n_23),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_33),
.C(n_21),
.Y(n_40)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_35),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_34),
.A2(n_29),
.B1(n_24),
.B2(n_26),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_37),
.A2(n_24),
.B1(n_17),
.B2(n_21),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_27),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_SL g41 ( 
.A(n_38),
.B(n_39),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_SL g39 ( 
.A(n_31),
.B(n_27),
.Y(n_39)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_18),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_44),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_45),
.Y(n_49)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_38),
.A2(n_17),
.B1(n_18),
.B2(n_2),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_39),
.C(n_9),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_47),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_0),
.C(n_1),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_49),
.B(n_41),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_51),
.A2(n_52),
.B(n_1),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_48),
.B(n_0),
.Y(n_52)
);

AOI322xp5_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_51),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_3),
.C2(n_8),
.Y(n_54)
);

OAI321xp33_ASAP7_75t_L g55 ( 
.A1(n_54),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_50),
.C(n_52),
.Y(n_55)
);


endmodule