module fake_jpeg_1902_n_317 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx6_ASAP7_75t_SL g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_5),
.B(n_12),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_36),
.Y(n_47)
);

NAND2xp33_ASAP7_75t_SL g107 ( 
.A(n_47),
.B(n_78),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_18),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_48),
.B(n_63),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_49),
.Y(n_150)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_50),
.Y(n_109)
);

BUFx4f_ASAP7_75t_SL g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx4f_ASAP7_75t_SL g117 ( 
.A(n_51),
.Y(n_117)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g149 ( 
.A(n_52),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

BUFx4f_ASAP7_75t_SL g54 ( 
.A(n_20),
.Y(n_54)
);

INVx13_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_55),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_15),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_56),
.B(n_57),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_0),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_44),
.B(n_0),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_58),
.B(n_64),
.Y(n_135)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_60),
.Y(n_140)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_61),
.Y(n_124)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_62),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_18),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_3),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_18),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_65),
.B(n_68),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_66),
.Y(n_137)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_67),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_28),
.B(n_5),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_69),
.Y(n_141)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

BUFx12_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_72),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_73),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_28),
.B(n_25),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_74),
.B(n_83),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_22),
.Y(n_75)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_76),
.Y(n_136)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_17),
.Y(n_77)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_77),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_79),
.Y(n_138)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_80),
.Y(n_143)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_81),
.Y(n_148)
);

BUFx16f_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_82),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_17),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_84),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_19),
.B(n_6),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_85),
.B(n_87),
.Y(n_146)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_86),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_19),
.B(n_6),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_88),
.B(n_89),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_25),
.B(n_31),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_90),
.B(n_91),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_20),
.Y(n_91)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_92),
.B(n_93),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_31),
.B(n_7),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_94),
.B(n_33),
.C(n_43),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_37),
.B(n_7),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_95),
.A2(n_96),
.B1(n_98),
.B2(n_9),
.Y(n_126)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_30),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_97),
.A2(n_99),
.B1(n_82),
.B2(n_55),
.Y(n_119)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_32),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_33),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_100),
.B(n_59),
.Y(n_153)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_84),
.A2(n_37),
.B1(n_45),
.B2(n_42),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_101),
.A2(n_102),
.B1(n_149),
.B2(n_150),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_57),
.A2(n_20),
.B1(n_43),
.B2(n_42),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_105),
.A2(n_112),
.B1(n_128),
.B2(n_130),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_53),
.A2(n_45),
.B1(n_40),
.B2(n_35),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_66),
.A2(n_40),
.B1(n_35),
.B2(n_27),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_114),
.A2(n_140),
.B1(n_134),
.B2(n_100),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_119),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_68),
.A2(n_27),
.B1(n_10),
.B2(n_11),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_123),
.A2(n_127),
.B1(n_147),
.B2(n_114),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_107),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_99),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_58),
.A2(n_13),
.B1(n_56),
.B2(n_95),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_76),
.A2(n_13),
.B1(n_88),
.B2(n_89),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_47),
.A2(n_13),
.B1(n_74),
.B2(n_54),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_131),
.A2(n_139),
.B1(n_126),
.B2(n_117),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_91),
.A2(n_51),
.B1(n_59),
.B2(n_72),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_79),
.A2(n_24),
.B1(n_36),
.B2(n_46),
.Y(n_147)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_109),
.Y(n_151)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_151),
.Y(n_191)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_144),
.Y(n_152)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_152),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_153),
.B(n_162),
.Y(n_190)
);

INVx6_ASAP7_75t_SL g154 ( 
.A(n_103),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_154),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_155),
.A2(n_158),
.B1(n_164),
.B2(n_171),
.Y(n_195)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_133),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_156),
.Y(n_204)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_148),
.Y(n_157)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_157),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_160),
.B(n_161),
.Y(n_201)
);

NAND2xp33_ASAP7_75t_SL g161 ( 
.A(n_132),
.B(n_111),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_L g162 ( 
.A1(n_115),
.A2(n_125),
.B(n_116),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_120),
.B(n_146),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_163),
.B(n_170),
.Y(n_203)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_165),
.Y(n_200)
);

INVx13_ASAP7_75t_L g166 ( 
.A(n_117),
.Y(n_166)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_166),
.Y(n_196)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_110),
.Y(n_167)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_167),
.Y(n_199)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_124),
.Y(n_168)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_168),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_135),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_129),
.A2(n_124),
.B1(n_143),
.B2(n_104),
.Y(n_171)
);

NAND2x1_ASAP7_75t_SL g172 ( 
.A(n_117),
.B(n_107),
.Y(n_172)
);

O2A1O1Ixp33_ASAP7_75t_L g197 ( 
.A1(n_172),
.A2(n_179),
.B(n_169),
.C(n_186),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g173 ( 
.A(n_132),
.Y(n_173)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_173),
.Y(n_208)
);

OA22x2_ASAP7_75t_L g188 ( 
.A1(n_174),
.A2(n_186),
.B1(n_110),
.B2(n_138),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_175),
.B(n_176),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_121),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_113),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_178),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_136),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_106),
.B(n_108),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_179),
.B(n_182),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_122),
.A2(n_136),
.B1(n_137),
.B2(n_104),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_180),
.A2(n_183),
.B1(n_165),
.B2(n_171),
.Y(n_207)
);

AOI21xp33_ASAP7_75t_L g181 ( 
.A1(n_121),
.A2(n_118),
.B(n_111),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_181),
.B(n_172),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_108),
.B(n_106),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_137),
.A2(n_142),
.B1(n_141),
.B2(n_133),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_142),
.B(n_141),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_184),
.B(n_185),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_138),
.B(n_113),
.Y(n_185)
);

CKINVDCx6p67_ASAP7_75t_R g186 ( 
.A(n_118),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_188),
.Y(n_216)
);

AND2x6_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_122),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_189),
.B(n_160),
.Y(n_213)
);

OAI21xp33_ASAP7_75t_L g212 ( 
.A1(n_193),
.A2(n_197),
.B(n_164),
.Y(n_212)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_207),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_L g209 ( 
.A1(n_174),
.A2(n_155),
.B1(n_183),
.B2(n_169),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_209),
.A2(n_201),
.B1(n_207),
.B2(n_190),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_151),
.B(n_164),
.C(n_178),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_177),
.C(n_166),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_212),
.A2(n_230),
.B(n_192),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_213),
.B(n_215),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_195),
.A2(n_159),
.B1(n_180),
.B2(n_168),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_214),
.A2(n_224),
.B1(n_228),
.B2(n_229),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_175),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_196),
.Y(n_217)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_217),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_194),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_232),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_205),
.B(n_152),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_221),
.Y(n_243)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_191),
.Y(n_220)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_220),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_201),
.A2(n_157),
.B1(n_156),
.B2(n_161),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_186),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_222),
.B(n_225),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_201),
.A2(n_154),
.B1(n_186),
.B2(n_167),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_176),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_231),
.C(n_225),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_197),
.A2(n_173),
.B(n_193),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_227),
.A2(n_188),
.B(n_208),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_198),
.A2(n_209),
.B1(n_188),
.B2(n_211),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_210),
.A2(n_198),
.B(n_194),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_203),
.B(n_189),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_206),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_233),
.B(n_241),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_222),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_234),
.B(n_248),
.Y(n_265)
);

BUFx24_ASAP7_75t_SL g236 ( 
.A(n_231),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_236),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_219),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_245),
.C(n_226),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_240),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_215),
.B(n_188),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_199),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_220),
.Y(n_246)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_246),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_232),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_224),
.Y(n_249)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_249),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_250),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_218),
.B(n_187),
.Y(n_251)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_251),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_262),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_250),
.Y(n_255)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_255),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_239),
.A2(n_223),
.B1(n_228),
.B2(n_213),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_259),
.A2(n_263),
.B1(n_239),
.B2(n_249),
.Y(n_271)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_242),
.Y(n_260)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_260),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_244),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_264),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_237),
.A2(n_223),
.B1(n_229),
.B2(n_216),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_237),
.A2(n_223),
.B(n_214),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_265),
.B(n_248),
.Y(n_270)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_270),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_271),
.A2(n_264),
.B(n_259),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_262),
.B(n_233),
.C(n_238),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_272),
.B(n_275),
.C(n_276),
.Y(n_281)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_253),
.Y(n_273)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_273),
.Y(n_286)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_265),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_251),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_245),
.C(n_247),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_266),
.B(n_243),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_277),
.B(n_278),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_255),
.B(n_243),
.C(n_234),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_276),
.B(n_257),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_283),
.Y(n_291)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_282),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_268),
.B(n_258),
.Y(n_283)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_284),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_278),
.B(n_242),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_277),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_275),
.C(n_272),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_290),
.Y(n_299)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_287),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_292),
.B(n_279),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_267),
.C(n_266),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_293),
.B(n_279),
.C(n_267),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g301 ( 
.A(n_295),
.B(n_296),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_294),
.A2(n_282),
.B(n_271),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g302 ( 
.A1(n_297),
.A2(n_254),
.B(n_263),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_286),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_298),
.B(n_300),
.Y(n_304)
);

BUFx10_ASAP7_75t_L g300 ( 
.A(n_289),
.Y(n_300)
);

NOR2xp67_ASAP7_75t_SL g309 ( 
.A(n_302),
.B(n_241),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_288),
.C(n_293),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_303),
.B(n_305),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_256),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_304),
.B(n_269),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_307),
.B(n_309),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_200),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_308),
.B(n_235),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_310),
.Y(n_313)
);

AOI322xp5_ASAP7_75t_L g311 ( 
.A1(n_306),
.A2(n_300),
.A3(n_254),
.B1(n_246),
.B2(n_240),
.C1(n_235),
.C2(n_221),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_311),
.B(n_217),
.C(n_204),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_217),
.C(n_312),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_315),
.B(n_204),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_313),
.Y(n_317)
);


endmodule