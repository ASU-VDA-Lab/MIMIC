module real_aes_12987_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_673;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_363;
wire n_182;
wire n_449;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_87;
wire n_171;
wire n_658;
wire n_676;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_193;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_541;
wire n_166;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_84;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
OA21x2_ASAP7_75t_L g109 ( .A1(n_0), .A2(n_42), .B(n_110), .Y(n_109) );
INVx1_ASAP7_75t_L g204 ( .A(n_0), .Y(n_204) );
INVx1_ASAP7_75t_L g564 ( .A(n_1), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_2), .A2(n_21), .B1(n_496), .B2(n_502), .Y(n_495) );
INVxp67_ASAP7_75t_SL g596 ( .A(n_2), .Y(n_596) );
AND2x2_ASAP7_75t_L g165 ( .A(n_3), .B(n_155), .Y(n_165) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_4), .A2(n_73), .B1(n_529), .B2(n_538), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_4), .A2(n_36), .B1(n_598), .B2(n_601), .Y(n_597) );
AOI22xp5_ASAP7_75t_L g672 ( .A1(n_5), .A2(n_43), .B1(n_673), .B2(n_674), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_5), .Y(n_673) );
AOI221xp5_ASAP7_75t_L g197 ( .A1(n_6), .A2(n_70), .B1(n_95), .B2(n_186), .C(n_198), .Y(n_197) );
BUFx3_ASAP7_75t_L g521 ( .A(n_7), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_8), .B(n_140), .Y(n_159) );
INVx3_ASAP7_75t_L g573 ( .A(n_9), .Y(n_573) );
INVx2_ASAP7_75t_L g501 ( .A(n_10), .Y(n_501) );
INVx1_ASAP7_75t_L g548 ( .A(n_10), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_11), .B(n_114), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_12), .B(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g93 ( .A(n_13), .Y(n_93) );
BUFx3_ASAP7_75t_L g116 ( .A(n_13), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_14), .B(n_126), .Y(n_172) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_14), .Y(n_698) );
INVx1_ASAP7_75t_L g530 ( .A(n_15), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_15), .A2(n_75), .B1(n_616), .B2(n_618), .Y(n_615) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_16), .Y(n_245) );
BUFx10_ASAP7_75t_L g687 ( .A(n_17), .Y(n_687) );
INVx1_ASAP7_75t_L g535 ( .A(n_18), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_19), .B(n_185), .Y(n_184) );
INVx1_ASAP7_75t_L g666 ( .A(n_19), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_20), .B(n_132), .Y(n_242) );
OAI21xp33_ASAP7_75t_L g286 ( .A1(n_20), .A2(n_55), .B(n_287), .Y(n_286) );
INVxp33_ASAP7_75t_SL g628 ( .A(n_21), .Y(n_628) );
O2A1O1Ixp5_ASAP7_75t_L g199 ( .A1(n_22), .A2(n_91), .B(n_157), .C(n_200), .Y(n_199) );
OAI221xp5_ASAP7_75t_L g555 ( .A1(n_23), .A2(n_48), .B1(n_556), .B2(n_560), .C(n_562), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_23), .B(n_644), .Y(n_643) );
INVxp33_ASAP7_75t_L g581 ( .A(n_24), .Y(n_581) );
INVx1_ASAP7_75t_L g608 ( .A(n_24), .Y(n_608) );
HB1xp67_ASAP7_75t_L g648 ( .A(n_24), .Y(n_648) );
INVx1_ASAP7_75t_L g87 ( .A(n_25), .Y(n_87) );
INVx2_ASAP7_75t_L g588 ( .A(n_26), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_27), .B(n_119), .Y(n_248) );
INVx1_ASAP7_75t_L g675 ( .A(n_28), .Y(n_675) );
INVx1_ASAP7_75t_L g667 ( .A(n_29), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_30), .B(n_183), .Y(n_182) );
INVx2_ASAP7_75t_L g580 ( .A(n_31), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_31), .B(n_608), .Y(n_607) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_31), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_32), .B(n_126), .Y(n_125) );
AND2x4_ASAP7_75t_L g86 ( .A(n_33), .B(n_87), .Y(n_86) );
HB1xp67_ASAP7_75t_L g660 ( .A(n_33), .Y(n_660) );
NAND2x1_ASAP7_75t_L g154 ( .A(n_34), .B(n_155), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g251 ( .A(n_35), .Y(n_251) );
AOI221xp5_ASAP7_75t_L g507 ( .A1(n_36), .A2(n_52), .B1(n_508), .B2(n_511), .C(n_517), .Y(n_507) );
INVx1_ASAP7_75t_L g149 ( .A(n_37), .Y(n_149) );
INVx1_ASAP7_75t_L g500 ( .A(n_38), .Y(n_500) );
INVx1_ASAP7_75t_L g505 ( .A(n_38), .Y(n_505) );
CKINVDCx5p33_ASAP7_75t_R g221 ( .A(n_39), .Y(n_221) );
AND2x2_ASAP7_75t_L g164 ( .A(n_40), .B(n_124), .Y(n_164) );
INVx1_ASAP7_75t_L g711 ( .A(n_40), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_41), .B(n_118), .Y(n_267) );
INVx1_ASAP7_75t_L g203 ( .A(n_42), .Y(n_203) );
INVx1_ASAP7_75t_L g674 ( .A(n_43), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_44), .B(n_140), .Y(n_232) );
INVx1_ASAP7_75t_L g110 ( .A(n_45), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_46), .B(n_124), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_47), .B(n_132), .Y(n_276) );
INVx1_ASAP7_75t_L g612 ( .A(n_48), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_49), .B(n_153), .Y(n_152) );
NAND2xp5_ASAP7_75t_SL g117 ( .A(n_50), .B(n_118), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_51), .B(n_225), .Y(n_224) );
INVxp67_ASAP7_75t_SL g634 ( .A(n_52), .Y(n_634) );
INVx1_ASAP7_75t_L g566 ( .A(n_53), .Y(n_566) );
AND2x2_ASAP7_75t_L g169 ( .A(n_54), .B(n_140), .Y(n_169) );
CKINVDCx5p33_ASAP7_75t_R g207 ( .A(n_55), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_56), .B(n_91), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_57), .B(n_114), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_58), .B(n_118), .Y(n_222) );
CKINVDCx5p33_ASAP7_75t_R g201 ( .A(n_59), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_60), .B(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_61), .B(n_132), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_62), .B(n_133), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g123 ( .A(n_63), .B(n_124), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g253 ( .A(n_64), .Y(n_253) );
AOI22xp5_ASAP7_75t_L g488 ( .A1(n_65), .A2(n_489), .B1(n_490), .B2(n_650), .Y(n_488) );
CKINVDCx5p33_ASAP7_75t_R g489 ( .A(n_65), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_66), .B(n_185), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_67), .B(n_269), .Y(n_268) );
INVx1_ASAP7_75t_L g96 ( .A(n_68), .Y(n_96) );
BUFx3_ASAP7_75t_L g129 ( .A(n_68), .Y(n_129) );
INVx1_ASAP7_75t_L g158 ( .A(n_68), .Y(n_158) );
INVx2_ASAP7_75t_L g587 ( .A(n_69), .Y(n_587) );
AND2x2_ASAP7_75t_L g600 ( .A(n_69), .B(n_588), .Y(n_600) );
INVxp67_ASAP7_75t_SL g640 ( .A(n_69), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_71), .B(n_228), .Y(n_227) );
INVx2_ASAP7_75t_L g523 ( .A(n_72), .Y(n_523) );
INVxp67_ASAP7_75t_SL g589 ( .A(n_73), .Y(n_589) );
AOI21xp33_ASAP7_75t_L g540 ( .A1(n_74), .A2(n_541), .B(n_543), .Y(n_540) );
OAI21xp5_ASAP7_75t_SL g621 ( .A1(n_74), .A2(n_622), .B(n_625), .Y(n_621) );
INVx1_ASAP7_75t_L g549 ( .A(n_75), .Y(n_549) );
INVx1_ASAP7_75t_L g545 ( .A(n_76), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_97), .B(n_487), .Y(n_77) );
CKINVDCx6p67_ASAP7_75t_R g78 ( .A(n_79), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g79 ( .A(n_80), .Y(n_79) );
BUFx2_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
NOR2x1_ASAP7_75t_L g81 ( .A(n_82), .B(n_88), .Y(n_81) );
INVx1_ASAP7_75t_SL g82 ( .A(n_83), .Y(n_82) );
BUFx2_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_86), .Y(n_85) );
BUFx6f_ASAP7_75t_SL g130 ( .A(n_86), .Y(n_130) );
INVx3_ASAP7_75t_L g177 ( .A(n_86), .Y(n_177) );
INVx2_ASAP7_75t_L g231 ( .A(n_86), .Y(n_231) );
INVx1_ASAP7_75t_L g256 ( .A(n_86), .Y(n_256) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_87), .Y(n_658) );
AO21x2_ASAP7_75t_L g714 ( .A1(n_88), .A2(n_657), .B(n_715), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g88 ( .A(n_89), .B(n_94), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx2_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx2_ASAP7_75t_L g124 ( .A(n_92), .Y(n_124) );
INVx1_ASAP7_75t_L g150 ( .A(n_92), .Y(n_150) );
INVx2_ASAP7_75t_L g229 ( .A(n_92), .Y(n_229) );
BUFx6f_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx2_ASAP7_75t_L g187 ( .A(n_93), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_94), .B(n_220), .Y(n_219) );
INVx2_ASAP7_75t_SL g94 ( .A(n_95), .Y(n_94) );
OAI22xp5_ASAP7_75t_L g216 ( .A1(n_95), .A2(n_217), .B1(n_219), .B2(n_222), .Y(n_216) );
INVx1_ASAP7_75t_L g254 ( .A(n_95), .Y(n_254) );
BUFx3_ASAP7_75t_L g95 ( .A(n_96), .Y(n_95) );
INVx1_ASAP7_75t_L g121 ( .A(n_96), .Y(n_121) );
INVx2_ASAP7_75t_SL g97 ( .A(n_98), .Y(n_97) );
AND2x2_ASAP7_75t_L g98 ( .A(n_99), .B(n_416), .Y(n_98) );
NOR3xp33_ASAP7_75t_L g99 ( .A(n_100), .B(n_363), .C(n_393), .Y(n_99) );
NAND4xp25_ASAP7_75t_L g100 ( .A(n_101), .B(n_291), .C(n_330), .D(n_343), .Y(n_100) );
AOI332xp33_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_193), .A3(n_209), .B1(n_233), .B2(n_238), .B3(n_259), .C1(n_277), .C2(n_281), .Y(n_101) );
AND2x2_ASAP7_75t_L g102 ( .A(n_103), .B(n_160), .Y(n_102) );
AND2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_135), .Y(n_103) );
INVx2_ASAP7_75t_L g234 ( .A(n_104), .Y(n_234) );
AND2x2_ASAP7_75t_L g348 ( .A(n_104), .B(n_136), .Y(n_348) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
BUFx3_ASAP7_75t_L g303 ( .A(n_105), .Y(n_303) );
OAI21x1_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_111), .B(n_131), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
BUFx3_ASAP7_75t_L g287 ( .A(n_108), .Y(n_287) );
BUFx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g134 ( .A(n_109), .Y(n_134) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_109), .Y(n_140) );
INVx1_ASAP7_75t_L g205 ( .A(n_110), .Y(n_205) );
OAI21xp5_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_122), .B(n_130), .Y(n_111) );
AOI21xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_117), .B(n_120), .Y(n_112) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_115), .B(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g218 ( .A(n_115), .Y(n_218) );
INVx2_ASAP7_75t_L g226 ( .A(n_115), .Y(n_226) );
INVx2_ASAP7_75t_L g252 ( .A(n_115), .Y(n_252) );
BUFx6f_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g119 ( .A(n_116), .Y(n_119) );
BUFx6f_ASAP7_75t_L g127 ( .A(n_116), .Y(n_127) );
INVx2_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g153 ( .A(n_119), .Y(n_153) );
INVx1_ASAP7_75t_L g183 ( .A(n_119), .Y(n_183) );
INVx2_ASAP7_75t_L g247 ( .A(n_119), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_120), .A2(n_182), .B(n_184), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g223 ( .A1(n_120), .A2(n_224), .B(n_227), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_120), .A2(n_272), .B(n_274), .Y(n_271) );
BUFx10_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
AOI21xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_125), .B(n_128), .Y(n_122) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx3_ASAP7_75t_L g146 ( .A(n_127), .Y(n_146) );
INVx3_ASAP7_75t_L g155 ( .A(n_127), .Y(n_155) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx2_ASAP7_75t_L g144 ( .A(n_129), .Y(n_144) );
NOR2xp33_ASAP7_75t_L g148 ( .A(n_129), .B(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g249 ( .A(n_129), .Y(n_249) );
OAI21x1_ASAP7_75t_L g141 ( .A1(n_130), .A2(n_142), .B(n_151), .Y(n_141) );
INVx1_ASAP7_75t_L g192 ( .A(n_130), .Y(n_192) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_133), .B(n_192), .Y(n_191) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g354 ( .A(n_135), .B(n_303), .Y(n_354) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g237 ( .A(n_136), .Y(n_237) );
AND2x4_ASAP7_75t_SL g278 ( .A(n_136), .B(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_136), .B(n_162), .Y(n_306) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_136), .Y(n_324) );
AND2x2_ASAP7_75t_L g350 ( .A(n_136), .B(n_303), .Y(n_350) );
INVx1_ASAP7_75t_L g397 ( .A(n_136), .Y(n_397) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
OAI21x1_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_141), .B(n_159), .Y(n_137) );
INVx1_ASAP7_75t_SL g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVxp33_ASAP7_75t_L g175 ( .A(n_140), .Y(n_175) );
INVx1_ASAP7_75t_L g208 ( .A(n_140), .Y(n_208) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_140), .Y(n_214) );
OAI21xp5_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_145), .B(n_147), .Y(n_142) );
INVx1_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_148), .B(n_150), .Y(n_147) );
AOI21x1_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_154), .B(n_156), .Y(n_151) );
INVx1_ASAP7_75t_L g269 ( .A(n_153), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_156), .A2(n_189), .B(n_190), .Y(n_188) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g270 ( .A(n_157), .Y(n_270) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
BUFx3_ASAP7_75t_L g167 ( .A(n_158), .Y(n_167) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g320 ( .A(n_161), .Y(n_320) );
INVx1_ASAP7_75t_L g451 ( .A(n_161), .Y(n_451) );
OR2x2_ASAP7_75t_L g161 ( .A(n_162), .B(n_178), .Y(n_161) );
INVx2_ASAP7_75t_L g279 ( .A(n_162), .Y(n_279) );
AND2x2_ASAP7_75t_L g325 ( .A(n_162), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g380 ( .A(n_162), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_162), .B(n_397), .Y(n_428) );
AO21x2_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_168), .B(n_174), .Y(n_162) );
OAI21xp5_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_165), .B(n_166), .Y(n_163) );
INVx1_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
INVx2_ASAP7_75t_L g173 ( .A(n_167), .Y(n_173) );
NOR2xp67_ASAP7_75t_L g168 ( .A(n_169), .B(n_170), .Y(n_168) );
AOI21xp33_ASAP7_75t_L g174 ( .A1(n_169), .A2(n_175), .B(n_176), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B(n_173), .Y(n_170) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NOR3xp33_ASAP7_75t_L g196 ( .A(n_177), .B(n_197), .C(n_199), .Y(n_196) );
INVx1_ASAP7_75t_L g236 ( .A(n_178), .Y(n_236) );
AND2x2_ASAP7_75t_L g301 ( .A(n_178), .B(n_302), .Y(n_301) );
INVx3_ASAP7_75t_L g326 ( .A(n_178), .Y(n_326) );
INVx1_ASAP7_75t_L g347 ( .A(n_178), .Y(n_347) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_178), .Y(n_351) );
AND2x2_ASAP7_75t_L g361 ( .A(n_178), .B(n_279), .Y(n_361) );
AND2x4_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
OAI21xp5_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_188), .B(n_191), .Y(n_180) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx3_ASAP7_75t_L g198 ( .A(n_187), .Y(n_198) );
INVx1_ASAP7_75t_L g403 ( .A(n_193), .Y(n_403) );
HB1xp67_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
AND2x4_ASAP7_75t_L g261 ( .A(n_194), .B(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g412 ( .A(n_194), .B(n_386), .Y(n_412) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AND2x2_ASAP7_75t_L g297 ( .A(n_195), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g336 ( .A(n_195), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g369 ( .A(n_195), .B(n_263), .Y(n_369) );
INVx1_ASAP7_75t_L g459 ( .A(n_195), .Y(n_459) );
AO21x2_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_202), .B(n_206), .Y(n_195) );
NAND2xp33_ASAP7_75t_L g288 ( .A(n_196), .B(n_289), .Y(n_288) );
INVx2_ASAP7_75t_L g273 ( .A(n_198), .Y(n_273) );
AO21x2_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_204), .B(n_205), .Y(n_202) );
AOI21x1_ASAP7_75t_L g257 ( .A1(n_203), .A2(n_204), .B(n_205), .Y(n_257) );
NOR2xp33_ASAP7_75t_R g206 ( .A(n_207), .B(n_208), .Y(n_206) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
HB1xp67_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_211), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g335 ( .A(n_211), .Y(n_335) );
INVx2_ASAP7_75t_L g357 ( .A(n_211), .Y(n_357) );
OR2x2_ASAP7_75t_L g431 ( .A(n_211), .B(n_285), .Y(n_431) );
AND2x2_ASAP7_75t_L g470 ( .A(n_211), .B(n_261), .Y(n_470) );
BUFx3_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g310 ( .A(n_212), .Y(n_310) );
OAI21x1_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_215), .B(n_232), .Y(n_212) );
OAI21x1_ASAP7_75t_L g258 ( .A1(n_213), .A2(n_215), .B(n_232), .Y(n_258) );
OAI21x1_ASAP7_75t_L g264 ( .A1(n_213), .A2(n_265), .B(n_276), .Y(n_264) );
OAI21xp5_ASAP7_75t_L g298 ( .A1(n_213), .A2(n_265), .B(n_276), .Y(n_298) );
BUFx6f_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
OAI21x1_ASAP7_75t_L g215 ( .A1(n_216), .A2(n_223), .B(n_230), .Y(n_215) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
OAI221xp5_ASAP7_75t_L g250 ( .A1(n_229), .A2(n_251), .B1(n_252), .B2(n_253), .C(n_254), .Y(n_250) );
INVx2_ASAP7_75t_SL g230 ( .A(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g275 ( .A(n_231), .Y(n_275) );
NOR2x1_ASAP7_75t_L g233 ( .A(n_234), .B(n_235), .Y(n_233) );
INVx1_ASAP7_75t_L g280 ( .A(n_234), .Y(n_280) );
AND2x2_ASAP7_75t_L g402 ( .A(n_234), .B(n_387), .Y(n_402) );
AND2x2_ASAP7_75t_L g407 ( .A(n_234), .B(n_278), .Y(n_407) );
AND2x2_ASAP7_75t_L g482 ( .A(n_234), .B(n_325), .Y(n_482) );
OR2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_237), .Y(n_235) );
INVx2_ASAP7_75t_L g374 ( .A(n_236), .Y(n_374) );
INVx1_ASAP7_75t_L g433 ( .A(n_237), .Y(n_433) );
AND2x2_ASAP7_75t_L g448 ( .A(n_237), .B(n_449), .Y(n_448) );
OAI211xp5_ASAP7_75t_SL g466 ( .A1(n_238), .A2(n_467), .B(n_469), .C(n_471), .Y(n_466) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
AND2x4_ASAP7_75t_SL g352 ( .A(n_239), .B(n_261), .Y(n_352) );
AND2x2_ASAP7_75t_L g392 ( .A(n_239), .B(n_297), .Y(n_392) );
AND2x2_ASAP7_75t_L g404 ( .A(n_239), .B(n_369), .Y(n_404) );
AND2x2_ASAP7_75t_L g411 ( .A(n_239), .B(n_412), .Y(n_411) );
AND2x4_ASAP7_75t_L g239 ( .A(n_240), .B(n_258), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx2_ASAP7_75t_L g296 ( .A(n_241), .Y(n_296) );
AND2x2_ASAP7_75t_L g309 ( .A(n_241), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g338 ( .A(n_241), .Y(n_338) );
AND2x2_ASAP7_75t_L g441 ( .A(n_241), .B(n_258), .Y(n_441) );
AND2x4_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
NAND3xp33_ASAP7_75t_L g285 ( .A(n_243), .B(n_286), .C(n_288), .Y(n_285) );
NAND3xp33_ASAP7_75t_L g243 ( .A(n_244), .B(n_250), .C(n_255), .Y(n_243) );
A2O1A1Ixp33_ASAP7_75t_L g244 ( .A1(n_245), .A2(n_246), .B(n_248), .C(n_249), .Y(n_244) );
INVx2_ASAP7_75t_SL g246 ( .A(n_247), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
INVx2_ASAP7_75t_L g290 ( .A(n_257), .Y(n_290) );
INVx1_ASAP7_75t_L g388 ( .A(n_258), .Y(n_388) );
A2O1A1Ixp33_ASAP7_75t_L g406 ( .A1(n_259), .A2(n_387), .B(n_407), .C(n_408), .Y(n_406) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g311 ( .A(n_262), .Y(n_311) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVxp67_ASAP7_75t_L g283 ( .A(n_264), .Y(n_283) );
OAI21x1_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_271), .B(n_275), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_268), .B(n_270), .Y(n_266) );
AND2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_280), .Y(n_277) );
INVx2_ASAP7_75t_L g445 ( .A(n_278), .Y(n_445) );
AND2x2_ASAP7_75t_L g465 ( .A(n_278), .B(n_351), .Y(n_465) );
BUFx2_ASAP7_75t_L g414 ( .A(n_279), .Y(n_414) );
OR2x2_ASAP7_75t_L g427 ( .A(n_280), .B(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g475 ( .A(n_281), .Y(n_475) );
AND2x2_ASAP7_75t_L g281 ( .A(n_282), .B(n_284), .Y(n_281) );
INVx1_ASAP7_75t_L g333 ( .A(n_282), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_282), .B(n_334), .Y(n_362) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g328 ( .A(n_283), .B(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g329 ( .A(n_285), .Y(n_329) );
OR2x2_ASAP7_75t_L g356 ( .A(n_285), .B(n_357), .Y(n_356) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AOI221xp5_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_299), .B1(n_307), .B2(n_312), .C(n_314), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_297), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x4_ASAP7_75t_L g387 ( .A(n_296), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g398 ( .A(n_297), .B(n_335), .Y(n_398) );
AND2x2_ASAP7_75t_L g434 ( .A(n_297), .B(n_387), .Y(n_434) );
AND2x2_ASAP7_75t_L g481 ( .A(n_297), .B(n_441), .Y(n_481) );
INVx1_ASAP7_75t_L g386 ( .A(n_298), .Y(n_386) );
NOR2xp67_ASAP7_75t_SL g299 ( .A(n_300), .B(n_304), .Y(n_299) );
NAND4xp25_ASAP7_75t_L g425 ( .A(n_300), .B(n_379), .C(n_426), .D(n_427), .Y(n_425) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g312 ( .A(n_301), .B(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_301), .B(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g318 ( .A(n_302), .Y(n_318) );
INVx1_ASAP7_75t_L g360 ( .A(n_302), .Y(n_360) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_302), .Y(n_415) );
AND2x2_ASAP7_75t_L g424 ( .A(n_302), .B(n_313), .Y(n_424) );
INVx3_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g449 ( .A(n_303), .B(n_380), .Y(n_449) );
INVx1_ASAP7_75t_L g372 ( .A(n_304), .Y(n_372) );
BUFx3_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g390 ( .A(n_305), .B(n_347), .Y(n_390) );
AND2x4_ASAP7_75t_L g405 ( .A(n_305), .B(n_374), .Y(n_405) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g313 ( .A(n_306), .Y(n_313) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_311), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_309), .B(n_369), .Y(n_376) );
INVx1_ASAP7_75t_L g473 ( .A(n_309), .Y(n_473) );
BUFx3_ASAP7_75t_L g367 ( .A(n_310), .Y(n_367) );
NAND2xp5_ASAP7_75t_SL g479 ( .A(n_311), .B(n_402), .Y(n_479) );
O2A1O1Ixp33_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_319), .B(n_321), .C(n_327), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OAI21xp33_ASAP7_75t_L g474 ( .A1(n_317), .A2(n_475), .B(n_476), .Y(n_474) );
INVx1_ASAP7_75t_L g342 ( .A(n_318), .Y(n_342) );
INVxp67_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g353 ( .A(n_320), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g395 ( .A(n_320), .B(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g399 ( .A(n_320), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NAND2x1_ASAP7_75t_L g340 ( .A(n_322), .B(n_341), .Y(n_340) );
AND2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_325), .Y(n_322) );
INVxp67_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_324), .Y(n_382) );
INVx1_ASAP7_75t_L g364 ( .A(n_325), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_325), .B(n_342), .Y(n_439) );
OR2x2_ASAP7_75t_L g379 ( .A(n_326), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g454 ( .A(n_326), .Y(n_454) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OAI21xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_336), .B(n_339), .Y(n_330) );
INVxp33_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AOI22xp5_ASAP7_75t_L g394 ( .A1(n_336), .A2(n_395), .B1(n_398), .B2(n_399), .Y(n_394) );
AND2x2_ASAP7_75t_L g368 ( .A(n_337), .B(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g422 ( .A(n_337), .Y(n_422) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AOI222xp33_ASAP7_75t_L g343 ( .A1(n_344), .A2(n_352), .B1(n_353), .B2(n_355), .C1(n_358), .C2(n_362), .Y(n_343) );
NAND2xp33_ASAP7_75t_L g344 ( .A(n_345), .B(n_349), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
AND2x2_ASAP7_75t_L g391 ( .A(n_347), .B(n_350), .Y(n_391) );
AND2x2_ASAP7_75t_L g462 ( .A(n_347), .B(n_433), .Y(n_462) );
INVx1_ASAP7_75t_L g426 ( .A(n_348), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_350), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_354), .B(n_378), .Y(n_409) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AOI22xp5_ASAP7_75t_L g480 ( .A1(n_358), .A2(n_392), .B1(n_481), .B2(n_482), .Y(n_480) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
INVx1_ASAP7_75t_L g400 ( .A(n_360), .Y(n_400) );
OAI211xp5_ASAP7_75t_L g363 ( .A1(n_364), .A2(n_365), .B(n_370), .C(n_389), .Y(n_363) );
NAND2x1p5_ASAP7_75t_L g365 ( .A(n_366), .B(n_368), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_368), .A2(n_407), .B1(n_411), .B2(n_413), .Y(n_410) );
INVx1_ASAP7_75t_L g468 ( .A(n_369), .Y(n_468) );
AOI22xp5_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_375), .B1(n_377), .B2(n_383), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
AND2x2_ASAP7_75t_L g423 ( .A(n_373), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OR2x2_ASAP7_75t_L g486 ( .A(n_374), .B(n_445), .Y(n_486) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x4_ASAP7_75t_L g377 ( .A(n_378), .B(n_381), .Y(n_377) );
AOI32xp33_ASAP7_75t_L g401 ( .A1(n_378), .A2(n_402), .A3(n_403), .B1(n_404), .B2(n_405), .Y(n_401) );
INVx3_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_SL g384 ( .A(n_385), .B(n_387), .Y(n_384) );
INVx2_ASAP7_75t_L g421 ( .A(n_385), .Y(n_421) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_387), .B(n_403), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_387), .B(n_421), .Y(n_476) );
OAI21xp33_ASAP7_75t_L g389 ( .A1(n_390), .A2(n_391), .B(n_392), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_390), .A2(n_465), .B1(n_466), .B2(n_474), .Y(n_464) );
NAND4xp25_ASAP7_75t_SL g393 ( .A(n_394), .B(n_401), .C(n_406), .D(n_410), .Y(n_393) );
HB1xp67_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_403), .B(n_472), .Y(n_471) );
INVx2_ASAP7_75t_SL g452 ( .A(n_404), .Y(n_452) );
OAI21xp5_ASAP7_75t_SL g453 ( .A1(n_404), .A2(n_454), .B(n_455), .Y(n_453) );
INVxp67_ASAP7_75t_SL g408 ( .A(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_417), .B(n_463), .Y(n_416) );
NAND3xp33_ASAP7_75t_L g417 ( .A(n_418), .B(n_435), .C(n_453), .Y(n_417) );
AOI222xp33_ASAP7_75t_L g418 ( .A1(n_419), .A2(n_423), .B1(n_425), .B2(n_429), .C1(n_432), .C2(n_434), .Y(n_418) );
INVxp67_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
OR2x2_ASAP7_75t_L g430 ( .A(n_421), .B(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g440 ( .A(n_421), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g484 ( .A(n_431), .Y(n_484) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
AOI221xp5_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_438), .B1(n_440), .B2(n_442), .C(n_446), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
AND2x2_ASAP7_75t_L g457 ( .A(n_441), .B(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_450), .B(n_452), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
O2A1O1Ixp33_ASAP7_75t_L g455 ( .A1(n_454), .A2(n_456), .B(n_460), .C(n_462), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_454), .B(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
NAND4xp25_ASAP7_75t_L g463 ( .A(n_464), .B(n_477), .C(n_480), .D(n_483), .Y(n_463) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVxp67_ASAP7_75t_SL g478 ( .A(n_479), .Y(n_478) );
OAI21xp33_ASAP7_75t_SL g483 ( .A1(n_481), .A2(n_484), .B(n_485), .Y(n_483) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
OAI221xp5_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_651), .B1(n_661), .B2(n_705), .C(n_706), .Y(n_487) );
INVx1_ASAP7_75t_L g650 ( .A(n_490), .Y(n_650) );
INVxp33_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_492), .B(n_620), .Y(n_491) );
O2A1O1Ixp33_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_555), .B(n_567), .C(n_574), .Y(n_492) );
NAND4xp25_ASAP7_75t_L g493 ( .A(n_494), .B(n_524), .C(n_534), .D(n_544), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_495), .B(n_507), .Y(n_494) );
BUFx12f_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x4_ASAP7_75t_L g563 ( .A(n_497), .B(n_561), .Y(n_563) );
BUFx6f_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx3_ASAP7_75t_L g539 ( .A(n_498), .Y(n_539) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_501), .Y(n_498) );
AND2x4_ASAP7_75t_L g516 ( .A(n_499), .B(n_506), .Y(n_516) );
INVx1_ASAP7_75t_L g552 ( .A(n_499), .Y(n_552) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AND2x2_ASAP7_75t_L g510 ( .A(n_500), .B(n_501), .Y(n_510) );
INVx2_ASAP7_75t_L g506 ( .A(n_501), .Y(n_506) );
NAND2x1_ASAP7_75t_L g560 ( .A(n_502), .B(n_561), .Y(n_560) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx4_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
BUFx12f_ASAP7_75t_L g542 ( .A(n_504), .Y(n_542) );
AND2x4_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
AND2x4_ASAP7_75t_L g558 ( .A(n_505), .B(n_548), .Y(n_558) );
INVx3_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx5_ASAP7_75t_L g529 ( .A(n_509), .Y(n_529) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx3_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx5_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g536 ( .A(n_515), .Y(n_536) );
AND2x4_ASAP7_75t_L g565 ( .A(n_515), .B(n_561), .Y(n_565) );
BUFx6f_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
BUFx6f_ASAP7_75t_L g533 ( .A(n_516), .Y(n_533) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AND2x4_ASAP7_75t_L g520 ( .A(n_521), .B(n_522), .Y(n_520) );
AND2x2_ASAP7_75t_L g527 ( .A(n_521), .B(n_528), .Y(n_527) );
OR2x2_ASAP7_75t_L g543 ( .A(n_521), .B(n_528), .Y(n_543) );
OR2x6_ASAP7_75t_L g559 ( .A(n_521), .B(n_523), .Y(n_559) );
BUFx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g528 ( .A(n_523), .Y(n_528) );
AOI21xp33_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_530), .B(n_531), .Y(n_524) );
AND2x4_ASAP7_75t_L g525 ( .A(n_526), .B(n_529), .Y(n_525) );
AND2x2_ASAP7_75t_SL g531 ( .A(n_526), .B(n_532), .Y(n_531) );
AND2x4_ASAP7_75t_L g546 ( .A(n_526), .B(n_547), .Y(n_546) );
BUFx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g554 ( .A(n_527), .Y(n_554) );
BUFx6f_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
OAI211xp5_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_536), .B(n_537), .C(n_540), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_535), .A2(n_626), .B1(n_628), .B2(n_629), .Y(n_625) );
INVx5_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
BUFx6f_ASAP7_75t_L g688 ( .A(n_543), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_546), .B1(n_549), .B2(n_550), .Y(n_544) );
AOI222xp33_ASAP7_75t_L g633 ( .A1(n_545), .A2(n_566), .B1(n_634), .B2(n_635), .C1(n_636), .C2(n_638), .Y(n_633) );
NAND3xp33_ASAP7_75t_L g685 ( .A(n_547), .B(n_686), .C(n_688), .Y(n_685) );
AND2x4_ASAP7_75t_L g694 ( .A(n_547), .B(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
AND2x4_ASAP7_75t_L g550 ( .A(n_551), .B(n_553), .Y(n_550) );
INVx3_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g695 ( .A(n_554), .Y(n_695) );
OR2x2_ASAP7_75t_L g556 ( .A(n_557), .B(n_559), .Y(n_556) );
INVx8_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx2_ASAP7_75t_L g561 ( .A(n_559), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_564), .B1(n_565), .B2(n_566), .Y(n_562) );
OAI221xp5_ASAP7_75t_L g610 ( .A1(n_564), .A2(n_611), .B1(n_612), .B2(n_613), .C(n_615), .Y(n_610) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVxp67_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx2_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
BUFx3_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g649 ( .A(n_572), .Y(n_649) );
INVx2_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND3x1_ASAP7_75t_L g577 ( .A(n_573), .B(n_578), .C(n_581), .Y(n_577) );
INVx2_ASAP7_75t_L g609 ( .A(n_573), .Y(n_609) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_582), .B1(n_606), .B2(n_610), .Y(n_574) );
BUFx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
INVx3_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g627 ( .A(n_579), .Y(n_627) );
AND2x4_ASAP7_75t_L g636 ( .A(n_579), .B(n_637), .Y(n_636) );
AND2x4_ASAP7_75t_SL g638 ( .A(n_579), .B(n_639), .Y(n_638) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OAI221xp5_ASAP7_75t_SL g582 ( .A1(n_583), .A2(n_589), .B1(n_590), .B2(n_596), .C(n_597), .Y(n_582) );
HB1xp67_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
BUFx6f_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
BUFx3_ASAP7_75t_L g611 ( .A(n_585), .Y(n_611) );
OR2x2_ASAP7_75t_SL g622 ( .A(n_585), .B(n_623), .Y(n_622) );
OR2x6_ASAP7_75t_L g644 ( .A(n_585), .B(n_627), .Y(n_644) );
BUFx6f_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_587), .B(n_588), .Y(n_586) );
INVx2_ASAP7_75t_L g594 ( .A(n_587), .Y(n_594) );
AND2x4_ASAP7_75t_L g604 ( .A(n_587), .B(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g595 ( .A(n_588), .Y(n_595) );
INVx2_ASAP7_75t_L g605 ( .A(n_588), .Y(n_605) );
INVx3_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx1_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
BUFx12f_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
NAND2x1p5_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
AND2x4_ASAP7_75t_L g619 ( .A(n_594), .B(n_595), .Y(n_619) );
BUFx3_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
BUFx6f_ASAP7_75t_L g614 ( .A(n_599), .Y(n_614) );
AND2x2_ASAP7_75t_L g626 ( .A(n_599), .B(n_627), .Y(n_626) );
BUFx6f_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
BUFx6f_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx4_ASAP7_75t_L g631 ( .A(n_603), .Y(n_631) );
INVx5_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
BUFx6f_ASAP7_75t_L g617 ( .A(n_604), .Y(n_617) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_605), .Y(n_637) );
OR2x6_ASAP7_75t_L g606 ( .A(n_607), .B(n_609), .Y(n_606) );
CKINVDCx5p33_ASAP7_75t_R g613 ( .A(n_614), .Y(n_613) );
BUFx6f_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
BUFx2_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
BUFx2_ASAP7_75t_L g635 ( .A(n_619), .Y(n_635) );
AND2x4_ASAP7_75t_L g642 ( .A(n_619), .B(n_623), .Y(n_642) );
OAI31xp33_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_632), .A3(n_643), .B(n_645), .Y(n_620) );
INVx3_ASAP7_75t_R g630 ( .A(n_623), .Y(n_630) );
BUFx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
AND2x4_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_633), .B(n_641), .Y(n_632) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
CKINVDCx8_ASAP7_75t_R g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
INVx1_ASAP7_75t_L g705 ( .A(n_650), .Y(n_705) );
CKINVDCx16_ASAP7_75t_R g651 ( .A(n_652), .Y(n_651) );
CKINVDCx16_ASAP7_75t_R g652 ( .A(n_653), .Y(n_652) );
HB1xp67_ASAP7_75t_SL g653 ( .A(n_654), .Y(n_653) );
BUFx6f_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_656), .B(n_659), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
BUFx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g683 ( .A(n_658), .Y(n_683) );
AND2x2_ASAP7_75t_L g715 ( .A(n_659), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_660), .B(n_683), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_677), .B1(n_696), .B2(n_699), .Y(n_661) );
OAI22xp5_ASAP7_75t_L g707 ( .A1(n_662), .A2(n_696), .B1(n_708), .B2(n_709), .Y(n_707) );
AOI22xp5_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_664), .B1(n_669), .B2(n_670), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_666), .B1(n_667), .B2(n_668), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g668 ( .A(n_667), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_672), .B1(n_675), .B2(n_676), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g676 ( .A(n_675), .Y(n_676) );
INVx3_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
BUFx3_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx5_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx5_ASAP7_75t_L g708 ( .A(n_680), .Y(n_708) );
AND2x6_ASAP7_75t_L g680 ( .A(n_681), .B(n_689), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_682), .B(n_684), .Y(n_681) );
INVxp67_ASAP7_75t_L g703 ( .A(n_682), .Y(n_703) );
INVx1_ASAP7_75t_L g716 ( .A(n_683), .Y(n_716) );
INVxp67_ASAP7_75t_SL g684 ( .A(n_685), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_685), .B(n_693), .Y(n_704) );
INVx2_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
CKINVDCx11_ASAP7_75t_R g691 ( .A(n_687), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_690), .B(n_692), .Y(n_689) );
CKINVDCx5p33_ASAP7_75t_R g690 ( .A(n_691), .Y(n_690) );
INVx2_ASAP7_75t_SL g692 ( .A(n_693), .Y(n_692) );
INVx2_ASAP7_75t_SL g693 ( .A(n_694), .Y(n_693) );
CKINVDCx5p33_ASAP7_75t_R g696 ( .A(n_697), .Y(n_696) );
INVx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx2_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
BUFx4f_ASAP7_75t_SL g700 ( .A(n_701), .Y(n_700) );
BUFx6f_ASAP7_75t_L g709 ( .A(n_701), .Y(n_709) );
INVx4_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g702 ( .A(n_703), .B(n_704), .Y(n_702) );
AOI22xp5_ASAP7_75t_L g706 ( .A1(n_705), .A2(n_707), .B1(n_710), .B2(n_712), .Y(n_706) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g712 ( .A(n_713), .Y(n_712) );
CKINVDCx20_ASAP7_75t_R g713 ( .A(n_714), .Y(n_713) );
endmodule