module fake_jpeg_22769_n_79 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_79);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_79;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx2_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_7),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_3),
.B(n_2),
.Y(n_14)
);

BUFx12_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_15),
.B(n_0),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_19),
.B(n_21),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_20),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_12),
.B(n_1),
.Y(n_21)
);

BUFx4f_ASAP7_75t_SL g22 ( 
.A(n_13),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_23),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_24),
.B(n_25),
.Y(n_31)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_21),
.B(n_18),
.Y(n_26)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_11),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_30),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_14),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_11),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_18),
.Y(n_39)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_35),
.Y(n_44)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_39),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_30),
.A2(n_9),
.B1(n_25),
.B2(n_17),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_43),
.B1(n_36),
.B2(n_40),
.Y(n_48)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_33),
.A2(n_9),
.B1(n_22),
.B2(n_25),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_32),
.A2(n_22),
.B1(n_24),
.B2(n_23),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_12),
.B1(n_10),
.B2(n_16),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_45),
.A2(n_49),
.B(n_51),
.Y(n_53)
);

NOR2xp67_ASAP7_75t_R g46 ( 
.A(n_40),
.B(n_24),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_46),
.B(n_1),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_48),
.B(n_49),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_24),
.B(n_23),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_42),
.A2(n_23),
.B(n_16),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_47),
.B(n_37),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_52),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_50),
.A2(n_35),
.B1(n_43),
.B2(n_34),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_55),
.B(n_57),
.Y(n_61)
);

INVxp33_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_59),
.Y(n_60)
);

OAI21xp33_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_10),
.B(n_4),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_51),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_64),
.Y(n_69)
);

NAND3xp33_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_52),
.C(n_8),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_65),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_53),
.C(n_20),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_15),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_68),
.B(n_61),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_70),
.A2(n_72),
.B(n_69),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_71),
.A2(n_69),
.B(n_15),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_67),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_73),
.A2(n_4),
.B(n_5),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_71),
.C(n_70),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_75),
.B(n_76),
.C(n_6),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_6),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_5),
.Y(n_79)
);


endmodule