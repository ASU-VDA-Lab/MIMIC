module fake_jpeg_22378_n_318 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_318);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_16),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

INVx11_ASAP7_75t_SL g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx10_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_0),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_37),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_44),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_41),
.Y(n_63)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_34),
.B1(n_20),
.B2(n_26),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_46),
.A2(n_55),
.B1(n_31),
.B2(n_22),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_34),
.B1(n_19),
.B2(n_20),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_51),
.A2(n_54),
.B1(n_72),
.B2(n_25),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_37),
.B(n_32),
.Y(n_52)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_37),
.B(n_21),
.Y(n_53)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_34),
.B1(n_20),
.B2(n_19),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_34),
.B1(n_26),
.B2(n_19),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_56),
.B(n_60),
.Y(n_74)
);

BUFx4f_ASAP7_75t_SL g58 ( 
.A(n_42),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_58),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_32),
.Y(n_59)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_22),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_22),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_64),
.Y(n_75)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_32),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_65),
.B(n_68),
.Y(n_77)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_44),
.Y(n_69)
);

AOI21xp33_ASAP7_75t_L g93 ( 
.A1(n_69),
.A2(n_44),
.B(n_18),
.Y(n_93)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_42),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_43),
.A2(n_33),
.B1(n_25),
.B2(n_31),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g82 ( 
.A1(n_71),
.A2(n_25),
.B(n_42),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_43),
.A2(n_33),
.B1(n_35),
.B2(n_27),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_73),
.B(n_86),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_76),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_61),
.A2(n_33),
.B1(n_35),
.B2(n_27),
.Y(n_78)
);

A2O1A1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_78),
.A2(n_93),
.B(n_29),
.C(n_21),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_57),
.A2(n_31),
.B1(n_30),
.B2(n_35),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_79),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_80),
.B(n_83),
.Y(n_132)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_82),
.A2(n_23),
.B(n_24),
.Y(n_135)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_L g84 ( 
.A1(n_47),
.A2(n_43),
.B1(n_42),
.B2(n_45),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_84),
.A2(n_88),
.B1(n_96),
.B2(n_63),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_47),
.B(n_45),
.C(n_41),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_87),
.B(n_89),
.Y(n_134)
);

AO22x1_ASAP7_75t_L g88 ( 
.A1(n_54),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_50),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_92),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_49),
.B(n_29),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_101),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_97),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_57),
.A2(n_27),
.B1(n_30),
.B2(n_23),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_98),
.A2(n_24),
.B1(n_21),
.B2(n_28),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_72),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_100),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_63),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_49),
.B(n_29),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_32),
.Y(n_103)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

INVx5_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_105),
.Y(n_128)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_51),
.B(n_45),
.C(n_41),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_107),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_53),
.B(n_29),
.Y(n_107)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_48),
.B(n_32),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_109),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_73),
.B(n_48),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_110),
.B(n_125),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_99),
.A2(n_66),
.B1(n_67),
.B2(n_63),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_112),
.A2(n_104),
.B1(n_108),
.B2(n_105),
.Y(n_142)
);

AND2x6_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_11),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_115),
.B(n_85),
.C(n_44),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_116),
.A2(n_120),
.B1(n_129),
.B2(n_100),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_74),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_117),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_96),
.A2(n_66),
.B1(n_18),
.B2(n_30),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_124),
.A2(n_130),
.B(n_129),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_29),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_106),
.A2(n_18),
.B1(n_23),
.B2(n_24),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_101),
.B(n_95),
.Y(n_130)
);

AO21x1_ASAP7_75t_L g166 ( 
.A1(n_135),
.A2(n_28),
.B(n_76),
.Y(n_166)
);

NAND2xp33_ASAP7_75t_SL g139 ( 
.A(n_136),
.B(n_88),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_78),
.B(n_95),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_138),
.B(n_84),
.Y(n_144)
);

AO21x1_ASAP7_75t_L g171 ( 
.A1(n_139),
.A2(n_166),
.B(n_168),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_118),
.A2(n_88),
.B1(n_107),
.B2(n_82),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_140),
.A2(n_167),
.B1(n_62),
.B2(n_45),
.Y(n_199)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_114),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_141),
.B(n_151),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_142),
.A2(n_145),
.B1(n_164),
.B2(n_133),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_144),
.A2(n_159),
.B(n_169),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_122),
.A2(n_102),
.B1(n_91),
.B2(n_77),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_134),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_146),
.B(n_148),
.Y(n_193)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_128),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_102),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_149),
.B(n_165),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_150),
.B(n_154),
.Y(n_197)
);

BUFx24_ASAP7_75t_SL g152 ( 
.A(n_130),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_153),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_117),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_155),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_110),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_156),
.Y(n_200)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_131),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_161),
.Y(n_185)
);

OAI21xp33_ASAP7_75t_L g158 ( 
.A1(n_138),
.A2(n_91),
.B(n_11),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_158),
.A2(n_135),
.B(n_133),
.Y(n_174)
);

INVx5_ASAP7_75t_SL g160 ( 
.A(n_114),
.Y(n_160)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_160),
.Y(n_180)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_114),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_162),
.B(n_163),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_116),
.A2(n_89),
.B1(n_75),
.B2(n_87),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_126),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_123),
.A2(n_80),
.B1(n_83),
.B2(n_81),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_119),
.Y(n_168)
);

NOR2xp67_ASAP7_75t_SL g169 ( 
.A(n_124),
.B(n_40),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_112),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_170),
.B(n_92),
.Y(n_198)
);

AO21x1_ASAP7_75t_L g207 ( 
.A1(n_174),
.A2(n_175),
.B(n_191),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_169),
.A2(n_122),
.B(n_113),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_145),
.B(n_127),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_176),
.B(n_182),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_159),
.A2(n_113),
.B(n_127),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_178),
.A2(n_181),
.B1(n_186),
.B2(n_188),
.Y(n_225)
);

OAI32xp33_ASAP7_75t_L g179 ( 
.A1(n_147),
.A2(n_120),
.A3(n_127),
.B1(n_125),
.B2(n_115),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_194),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_147),
.B(n_121),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_161),
.A2(n_121),
.B(n_111),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_140),
.B(n_136),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_187),
.B(n_192),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_150),
.A2(n_111),
.B(n_137),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_170),
.A2(n_137),
.B1(n_131),
.B2(n_28),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_189),
.A2(n_190),
.B1(n_199),
.B2(n_141),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_163),
.A2(n_62),
.B1(n_60),
.B2(n_45),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_156),
.A2(n_32),
.B(n_1),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_151),
.B(n_40),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_164),
.B(n_40),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_160),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_195),
.B(n_196),
.Y(n_205)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_142),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_198),
.B(n_148),
.Y(n_208)
);

AO21x1_ASAP7_75t_L g201 ( 
.A1(n_166),
.A2(n_41),
.B(n_40),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_201),
.B(n_154),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_173),
.B(n_143),
.Y(n_203)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_203),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_202),
.A2(n_183),
.B1(n_196),
.B2(n_199),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_206),
.A2(n_212),
.B1(n_201),
.B2(n_171),
.Y(n_235)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_208),
.Y(n_242)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_185),
.Y(n_209)
);

OAI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_209),
.A2(n_211),
.B1(n_213),
.B2(n_216),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_177),
.B(n_157),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_210),
.Y(n_246)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_198),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_193),
.Y(n_213)
);

INVx13_ASAP7_75t_L g214 ( 
.A(n_180),
.Y(n_214)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_214),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_215),
.A2(n_217),
.B1(n_218),
.B2(n_228),
.Y(n_244)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_197),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_180),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_186),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_190),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_220),
.A2(n_221),
.B1(n_223),
.B2(n_227),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_188),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_189),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_146),
.Y(n_224)
);

AND2x2_ASAP7_75t_SL g238 ( 
.A(n_224),
.B(n_226),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_167),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_195),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_181),
.B(n_162),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_221),
.A2(n_179),
.B1(n_172),
.B2(n_187),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_229),
.A2(n_38),
.B1(n_1),
.B2(n_2),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_175),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_230),
.B(n_233),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_178),
.C(n_176),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_231),
.B(n_232),
.C(n_236),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_225),
.C(n_172),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_204),
.B(n_182),
.Y(n_233)
);

OA21x2_ASAP7_75t_SL g234 ( 
.A1(n_207),
.A2(n_171),
.B(n_174),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_234),
.B(n_207),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_235),
.B(n_16),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_192),
.C(n_191),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_194),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_248),
.C(n_249),
.Y(n_254)
);

NAND2x1_ASAP7_75t_SL g241 ( 
.A(n_205),
.B(n_153),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_241),
.A2(n_0),
.B(n_1),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_220),
.A2(n_184),
.B1(n_126),
.B2(n_10),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_243),
.A2(n_213),
.B1(n_216),
.B2(n_223),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_211),
.B(n_41),
.C(n_40),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_219),
.B(n_41),
.C(n_40),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_215),
.B(n_41),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_250),
.B(n_208),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_252),
.B(n_258),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_253),
.B(n_264),
.Y(n_278)
);

AO221x1_ASAP7_75t_L g255 ( 
.A1(n_241),
.A2(n_217),
.B1(n_214),
.B2(n_227),
.C(n_209),
.Y(n_255)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_255),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_224),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_257),
.Y(n_275)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_240),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_245),
.Y(n_258)
);

OR2x2_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_267),
.Y(n_277)
);

XOR2x1_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_226),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_261),
.A2(n_262),
.B(n_263),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_8),
.Y(n_262)
);

BUFx12_ASAP7_75t_L g263 ( 
.A(n_247),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_246),
.A2(n_8),
.B1(n_15),
.B2(n_3),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_265),
.A2(n_229),
.B1(n_248),
.B2(n_4),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_265),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_268),
.A2(n_242),
.B1(n_232),
.B2(n_236),
.Y(n_269)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_269),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_268),
.A2(n_238),
.B(n_244),
.Y(n_270)
);

AO21x1_ASAP7_75t_L g293 ( 
.A1(n_270),
.A2(n_3),
.B(n_5),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_271),
.B(n_259),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_239),
.C(n_249),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_273),
.C(n_281),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_254),
.B(n_231),
.C(n_233),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_261),
.A2(n_250),
.B1(n_230),
.B2(n_0),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_279),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_0),
.C(n_3),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_282),
.B(n_253),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_260),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_285),
.C(n_292),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_284),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_251),
.C(n_266),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_291),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_263),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_290),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_263),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_275),
.B(n_251),
.Y(n_291)
);

AO21x1_ASAP7_75t_L g303 ( 
.A1(n_293),
.A2(n_6),
.B(n_7),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_5),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_294),
.B(n_293),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_296),
.B(n_297),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_286),
.A2(n_269),
.B1(n_279),
.B2(n_274),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_298),
.B(n_12),
.Y(n_308)
);

OAI321xp33_ASAP7_75t_L g300 ( 
.A1(n_286),
.A2(n_282),
.A3(n_271),
.B1(n_270),
.B2(n_280),
.C(n_278),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_300),
.A2(n_302),
.B1(n_10),
.B2(n_12),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_289),
.A2(n_278),
.B1(n_281),
.B2(n_9),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_303),
.B(n_7),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_299),
.A2(n_292),
.B1(n_283),
.B2(n_12),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_305),
.A2(n_302),
.B1(n_303),
.B2(n_301),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_306),
.B(n_309),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_307),
.A2(n_308),
.B(n_13),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_295),
.B(n_13),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_310),
.A2(n_298),
.B(n_14),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_311),
.A2(n_312),
.B(n_304),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_305),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_314),
.A2(n_315),
.B(n_313),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_13),
.B(n_15),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_16),
.Y(n_318)
);


endmodule