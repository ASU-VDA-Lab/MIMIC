module fake_jpeg_22962_n_321 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_321);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_321;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_38),
.Y(n_54)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_34),
.Y(n_57)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_0),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_23),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_41),
.B(n_22),
.Y(n_45)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_25),
.B(n_9),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_44),
.B(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_45),
.B(n_51),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_20),
.B1(n_17),
.B2(n_26),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_20),
.B1(n_17),
.B2(n_26),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_47),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_40),
.A2(n_22),
.B1(n_24),
.B2(n_26),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_53),
.Y(n_70)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_20),
.B1(n_24),
.B2(n_33),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g74 ( 
.A1(n_50),
.A2(n_30),
.B(n_31),
.C(n_35),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_24),
.B1(n_33),
.B2(n_27),
.Y(n_53)
);

CKINVDCx6p67_ASAP7_75t_R g55 ( 
.A(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_41),
.A2(n_27),
.B1(n_33),
.B2(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_58),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_57),
.B(n_61),
.Y(n_71)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_23),
.B1(n_33),
.B2(n_27),
.Y(n_60)
);

AO22x1_ASAP7_75t_L g77 ( 
.A1(n_60),
.A2(n_31),
.B1(n_30),
.B2(n_35),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_33),
.C(n_27),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_44),
.A2(n_27),
.B1(n_21),
.B2(n_29),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_67),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_36),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_65),
.Y(n_81)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g67 ( 
.A(n_36),
.B(n_32),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_31),
.Y(n_80)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_72),
.Y(n_99)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_74),
.A2(n_77),
.B1(n_47),
.B2(n_46),
.Y(n_97)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_78),
.B(n_79),
.Y(n_111)
);

INVx6_ASAP7_75t_SL g79 ( 
.A(n_49),
.Y(n_79)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_82),
.B(n_84),
.Y(n_114)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

AND2x6_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_14),
.Y(n_85)
);

AND2x6_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_55),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_87),
.Y(n_109)
);

NAND3xp33_ASAP7_75t_L g90 ( 
.A(n_55),
.B(n_14),
.C(n_16),
.Y(n_90)
);

OR2x2_ASAP7_75t_SL g122 ( 
.A(n_90),
.B(n_16),
.Y(n_122)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_95),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_55),
.B(n_19),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_92),
.B(n_67),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_63),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_93),
.Y(n_112)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_96),
.A2(n_85),
.B1(n_92),
.B2(n_72),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_97),
.A2(n_107),
.B1(n_115),
.B2(n_77),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_87),
.Y(n_100)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_100),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_61),
.C(n_45),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_101),
.B(n_43),
.Y(n_152)
);

MAJx3_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_61),
.C(n_56),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_102),
.A2(n_113),
.B(n_75),
.Y(n_137)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_87),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g151 ( 
.A(n_103),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_57),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_105),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_66),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_106),
.B(n_118),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_76),
.A2(n_53),
.B1(n_60),
.B2(n_50),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_110),
.Y(n_128)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_75),
.B(n_64),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_94),
.A2(n_54),
.B1(n_65),
.B2(n_68),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_121),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_86),
.B(n_51),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_67),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_119),
.B(n_86),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_19),
.Y(n_120)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_120),
.Y(n_124)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_74),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_28),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_81),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_123),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_102),
.A2(n_94),
.B1(n_83),
.B2(n_91),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_125),
.A2(n_134),
.B1(n_143),
.B2(n_144),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_114),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_126),
.B(n_133),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_102),
.A2(n_77),
.B1(n_88),
.B2(n_70),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_127),
.A2(n_141),
.B(n_145),
.Y(n_161)
);

AND2x2_ASAP7_75t_SL g129 ( 
.A(n_102),
.B(n_91),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_129),
.A2(n_101),
.B(n_119),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_114),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_123),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_135),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_136),
.B(n_142),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_152),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_97),
.A2(n_117),
.B(n_121),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_138),
.A2(n_149),
.B(n_139),
.Y(n_163)
);

OA21x2_ASAP7_75t_L g141 ( 
.A1(n_115),
.A2(n_81),
.B(n_48),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_99),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_113),
.A2(n_69),
.B1(n_92),
.B2(n_82),
.Y(n_144)
);

OA21x2_ASAP7_75t_L g145 ( 
.A1(n_107),
.A2(n_63),
.B(n_79),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_99),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_148),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_98),
.B(n_108),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_104),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_111),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_117),
.A2(n_78),
.B(n_43),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_150),
.Y(n_182)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_111),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_146),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_156),
.A2(n_136),
.B(n_131),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_159),
.B(n_174),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_152),
.B(n_129),
.C(n_137),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_160),
.B(n_170),
.C(n_184),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_105),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_162),
.B(n_178),
.Y(n_202)
);

AOI221xp5_ASAP7_75t_L g205 ( 
.A1(n_163),
.A2(n_127),
.B1(n_142),
.B2(n_153),
.C(n_132),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_140),
.Y(n_164)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_164),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_130),
.B(n_98),
.Y(n_165)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_128),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_167),
.B(n_172),
.Y(n_188)
);

OA21x2_ASAP7_75t_L g168 ( 
.A1(n_145),
.A2(n_96),
.B(n_106),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_168),
.A2(n_177),
.B(n_141),
.Y(n_200)
);

INVxp67_ASAP7_75t_SL g169 ( 
.A(n_140),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_169),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_129),
.B(n_96),
.C(n_118),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_130),
.B(n_120),
.Y(n_171)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_171),
.Y(n_195)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_128),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_139),
.Y(n_173)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_173),
.Y(n_204)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_147),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_149),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_175),
.Y(n_206)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_176),
.Y(n_211)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_144),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_138),
.B(n_122),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_145),
.A2(n_84),
.B1(n_73),
.B2(n_110),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_179),
.A2(n_180),
.B1(n_181),
.B2(n_126),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_145),
.A2(n_112),
.B1(n_109),
.B2(n_62),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_143),
.A2(n_62),
.B1(n_112),
.B2(n_109),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_129),
.B(n_103),
.C(n_100),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_184),
.B(n_135),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_185),
.A2(n_196),
.B(n_207),
.Y(n_227)
);

BUFx5_ASAP7_75t_L g187 ( 
.A(n_164),
.Y(n_187)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_187),
.Y(n_212)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_189),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_160),
.B(n_134),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_190),
.B(n_199),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_157),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_192),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_194),
.A2(n_197),
.B1(n_177),
.B2(n_174),
.Y(n_220)
);

BUFx12f_ASAP7_75t_SL g196 ( 
.A(n_168),
.Y(n_196)
);

AO22x1_ASAP7_75t_L g197 ( 
.A1(n_161),
.A2(n_141),
.B1(n_127),
.B2(n_132),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_200),
.A2(n_158),
.B1(n_179),
.B2(n_167),
.Y(n_230)
);

NOR2x1_ASAP7_75t_R g201 ( 
.A(n_156),
.B(n_141),
.Y(n_201)
);

XOR2x1_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_163),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_155),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_203),
.Y(n_229)
);

XNOR2x1_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_178),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_161),
.A2(n_131),
.B(n_150),
.Y(n_207)
);

BUFx12_ASAP7_75t_L g209 ( 
.A(n_168),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_210),
.Y(n_217)
);

INVx13_ASAP7_75t_L g210 ( 
.A(n_181),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_170),
.C(n_165),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_214),
.C(n_216),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_202),
.B(n_154),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_202),
.C(n_193),
.Y(n_216)
);

XNOR2x2_ASAP7_75t_SL g251 ( 
.A(n_218),
.B(n_219),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_220),
.A2(n_221),
.B1(n_233),
.B2(n_204),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_196),
.A2(n_197),
.B1(n_210),
.B2(n_194),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_190),
.C(n_199),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_223),
.B(n_225),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_189),
.B(n_124),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_224),
.B(n_235),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_158),
.C(n_159),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_154),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_226),
.B(n_234),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_230),
.A2(n_211),
.B1(n_191),
.B2(n_186),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_187),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_231),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_201),
.B(n_162),
.Y(n_232)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_232),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_206),
.A2(n_195),
.B1(n_200),
.B2(n_209),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_185),
.B(n_171),
.C(n_183),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_188),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_198),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_172),
.Y(n_239)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_239),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_227),
.A2(n_207),
.B(n_209),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_240),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_217),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_243),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_212),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_140),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_244),
.B(n_250),
.Y(n_260)
);

NOR3xp33_ASAP7_75t_SL g245 ( 
.A(n_218),
.B(n_185),
.C(n_198),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_255),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_246),
.A2(n_234),
.B1(n_213),
.B2(n_216),
.Y(n_262)
);

A2O1A1O1Ixp25_ASAP7_75t_L g247 ( 
.A1(n_219),
.A2(n_232),
.B(n_226),
.C(n_215),
.D(n_223),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_10),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_248),
.A2(n_249),
.B1(n_253),
.B2(n_220),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_236),
.A2(n_211),
.B1(n_151),
.B2(n_182),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_229),
.B(n_124),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_225),
.A2(n_151),
.B1(n_109),
.B2(n_116),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_233),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_221),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_257),
.A2(n_28),
.B1(n_32),
.B2(n_30),
.Y(n_269)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_259),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_262),
.Y(n_281)
);

A2O1A1Ixp33_ASAP7_75t_L g263 ( 
.A1(n_257),
.A2(n_215),
.B(n_214),
.C(n_222),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_263),
.A2(n_256),
.B(n_248),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_151),
.C(n_62),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_265),
.C(n_268),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_93),
.C(n_52),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_237),
.B(n_93),
.C(n_29),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_249),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_238),
.B(n_21),
.C(n_31),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_270),
.B(n_252),
.C(n_240),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_10),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_271),
.B(n_245),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_272),
.B(n_251),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_251),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_273),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_267),
.A2(n_242),
.B(n_254),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_274),
.A2(n_282),
.B(n_275),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_276),
.B(n_277),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_278),
.A2(n_283),
.B(n_284),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_286),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_239),
.C(n_247),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_282),
.B(n_287),
.C(n_270),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_264),
.A2(n_256),
.B(n_243),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_260),
.B(n_15),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_1),
.C(n_2),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_278),
.B(n_268),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_289),
.B(n_298),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_258),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_290),
.B(n_294),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_292),
.C(n_297),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_279),
.A2(n_261),
.B1(n_263),
.B2(n_272),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_269),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_283),
.A2(n_15),
.B(n_14),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_296),
.A2(n_12),
.B(n_11),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_285),
.A2(n_13),
.B(n_12),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_275),
.B(n_13),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_299),
.B(n_281),
.Y(n_302)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_301),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_303),
.C(n_305),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_12),
.C(n_11),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_11),
.C(n_2),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_293),
.A2(n_292),
.B(n_288),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_7),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_1),
.C(n_4),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_307),
.B(n_4),
.Y(n_312)
);

AOI322xp5_ASAP7_75t_L g310 ( 
.A1(n_308),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_294),
.C2(n_304),
.Y(n_310)
);

AOI322xp5_ASAP7_75t_L g318 ( 
.A1(n_310),
.A2(n_312),
.A3(n_313),
.B1(n_309),
.B2(n_6),
.C1(n_7),
.C2(n_5),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_300),
.Y(n_311)
);

A2O1A1Ixp33_ASAP7_75t_L g317 ( 
.A1(n_311),
.A2(n_315),
.B(n_5),
.C(n_6),
.Y(n_317)
);

A2O1A1Ixp33_ASAP7_75t_L g313 ( 
.A1(n_302),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_315),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_316),
.B(n_317),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_314),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_318),
.Y(n_321)
);


endmodule