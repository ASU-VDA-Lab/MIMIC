module fake_jpeg_17917_n_251 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_251);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_251;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_6),
.B(n_12),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_1),
.B(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_7),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_38),
.B(n_40),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_26),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_7),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_42),
.Y(n_51)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_24),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_58),
.Y(n_82)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_20),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_56),
.Y(n_73)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_37),
.A2(n_26),
.B1(n_18),
.B2(n_28),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_57),
.A2(n_18),
.B1(n_32),
.B2(n_26),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_24),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_60),
.B(n_62),
.Y(n_76)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_40),
.A2(n_17),
.B1(n_29),
.B2(n_21),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_64),
.A2(n_21),
.B1(n_29),
.B2(n_17),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_20),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_29),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_36),
.B(n_25),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_16),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_67),
.B(n_78),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_72),
.A2(n_19),
.B1(n_44),
.B2(n_60),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_46),
.A2(n_31),
.B1(n_23),
.B2(n_25),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_74),
.A2(n_86),
.B1(n_87),
.B2(n_91),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_31),
.C(n_23),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_75),
.B(n_59),
.C(n_52),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_84),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_47),
.B(n_24),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

OR2x2_ASAP7_75t_SL g83 ( 
.A(n_51),
.B(n_27),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_83),
.A2(n_88),
.B(n_82),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_66),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_45),
.A2(n_25),
.B1(n_16),
.B2(n_27),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_49),
.A2(n_63),
.B1(n_54),
.B2(n_53),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_88),
.B(n_90),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_51),
.A2(n_28),
.B1(n_18),
.B2(n_21),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_15),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_54),
.A2(n_31),
.B1(n_23),
.B2(n_17),
.Y(n_91)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_78),
.A2(n_61),
.B(n_50),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_94),
.A2(n_117),
.B(n_69),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_96),
.A2(n_98),
.B(n_102),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_82),
.A2(n_27),
.B(n_19),
.C(n_16),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_103),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_89),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_75),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_84),
.A2(n_50),
.B1(n_62),
.B2(n_56),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_101),
.A2(n_107),
.B1(n_91),
.B2(n_70),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_73),
.A2(n_0),
.B(n_1),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_43),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_19),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_105),
.Y(n_118)
);

INVx4_ASAP7_75t_SL g109 ( 
.A(n_76),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_73),
.B(n_31),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_44),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_0),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_111),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_121),
.Y(n_140)
);

AO21x2_ASAP7_75t_L g120 ( 
.A1(n_109),
.A2(n_87),
.B(n_74),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_120),
.A2(n_136),
.B1(n_93),
.B2(n_99),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_110),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_122),
.B(n_128),
.Y(n_149)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_124),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_127),
.A2(n_100),
.B(n_98),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_69),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_129),
.Y(n_145)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_92),
.Y(n_130)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_112),
.Y(n_147)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_92),
.Y(n_133)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_133),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_134),
.A2(n_94),
.B(n_102),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_106),
.B(n_86),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_135),
.B(n_94),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_98),
.A2(n_100),
.B1(n_99),
.B2(n_115),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

OAI32xp33_ASAP7_75t_L g139 ( 
.A1(n_131),
.A2(n_95),
.A3(n_104),
.B1(n_106),
.B2(n_96),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_139),
.B(n_134),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_141),
.A2(n_147),
.B(n_158),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_93),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_142),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_118),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_143),
.B(n_151),
.Y(n_174)
);

A2O1A1Ixp33_ASAP7_75t_L g144 ( 
.A1(n_131),
.A2(n_117),
.B(n_103),
.C(n_95),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_144),
.B(n_160),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_125),
.C(n_127),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_148),
.A2(n_153),
.B1(n_155),
.B2(n_132),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_120),
.A2(n_112),
.B1(n_109),
.B2(n_107),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_118),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_156),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_120),
.A2(n_117),
.B1(n_85),
.B2(n_71),
.Y(n_155)
);

BUFx24_ASAP7_75t_SL g156 ( 
.A(n_133),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_120),
.A2(n_97),
.B1(n_85),
.B2(n_71),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_123),
.Y(n_159)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_159),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_122),
.B(n_116),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_136),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_165),
.B(n_167),
.C(n_152),
.Y(n_190)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_138),
.Y(n_168)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_168),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_119),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_169),
.B(n_173),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_148),
.A2(n_127),
.B(n_137),
.Y(n_170)
);

BUFx12_ASAP7_75t_L g171 ( 
.A(n_138),
.Y(n_171)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_171),
.Y(n_186)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_145),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_175),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_129),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_176),
.B(n_177),
.Y(n_184)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_159),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_140),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_179),
.A2(n_147),
.B1(n_157),
.B2(n_153),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_180),
.A2(n_181),
.B1(n_188),
.B2(n_195),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_179),
.A2(n_147),
.B1(n_157),
.B2(n_150),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_151),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_187),
.C(n_189),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_163),
.Y(n_187)
);

AO22x2_ASAP7_75t_L g188 ( 
.A1(n_170),
.A2(n_158),
.B1(n_155),
.B2(n_143),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_144),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_190),
.B(n_191),
.C(n_193),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_152),
.C(n_150),
.Y(n_191)
);

AO21x1_ASAP7_75t_L g192 ( 
.A1(n_164),
.A2(n_154),
.B(n_126),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_192),
.B(n_172),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_174),
.B(n_123),
.C(n_108),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_164),
.A2(n_124),
.B1(n_114),
.B2(n_11),
.Y(n_195)
);

INVx13_ASAP7_75t_L g196 ( 
.A(n_186),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_198),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_176),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_185),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_201),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_182),
.B(n_169),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_194),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_202),
.B(n_203),
.Y(n_218)
);

FAx1_ASAP7_75t_SL g203 ( 
.A(n_189),
.B(n_161),
.CI(n_178),
.CON(n_203),
.SN(n_203)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_183),
.B(n_162),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_204),
.B(n_207),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_188),
.A2(n_177),
.B1(n_175),
.B2(n_173),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_205),
.A2(n_108),
.B1(n_80),
.B2(n_79),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_190),
.B(n_172),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_208),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_192),
.B(n_168),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_209),
.B(n_188),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_191),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_211),
.C(n_213),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_199),
.B(n_187),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_207),
.B(n_188),
.C(n_171),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_219),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_108),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_217),
.C(n_203),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_10),
.Y(n_217)
);

A2O1A1Ixp33_ASAP7_75t_SL g224 ( 
.A1(n_220),
.A2(n_196),
.B(n_198),
.C(n_206),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_221),
.A2(n_205),
.B(n_201),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_0),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_224),
.A2(n_212),
.B1(n_211),
.B2(n_2),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_218),
.Y(n_226)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_226),
.Y(n_232)
);

AOI31xp33_ASAP7_75t_L g227 ( 
.A1(n_213),
.A2(n_203),
.A3(n_206),
.B(n_11),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_227),
.B(n_13),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_6),
.C(n_14),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_80),
.C(n_79),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_229),
.B(n_230),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_210),
.B(n_6),
.Y(n_230)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_231),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_233),
.B(n_236),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_225),
.B(n_212),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_235),
.B(n_238),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_5),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_232),
.A2(n_223),
.B1(n_224),
.B2(n_8),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_239),
.B(n_236),
.C(n_237),
.Y(n_244)
);

OAI21xp33_ASAP7_75t_L g243 ( 
.A1(n_242),
.A2(n_234),
.B(n_238),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_243),
.A2(n_245),
.B(n_246),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_244),
.A2(n_5),
.B(n_15),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_240),
.B(n_242),
.Y(n_245)
);

OAI211xp5_ASAP7_75t_L g246 ( 
.A1(n_241),
.A2(n_5),
.B(n_13),
.C(n_11),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_248),
.B(n_0),
.C(n_1),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_249),
.A2(n_247),
.B1(n_2),
.B2(n_3),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_3),
.Y(n_251)
);


endmodule