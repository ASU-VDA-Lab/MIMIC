module fake_jpeg_5462_n_281 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_281);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_281;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx6_ASAP7_75t_SL g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_29),
.B(n_7),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_32),
.B(n_38),
.Y(n_58)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_37),
.Y(n_52)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx13_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_15),
.B(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_19),
.Y(n_39)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_41),
.Y(n_44)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_43),
.B(n_48),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_40),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_45),
.B(n_22),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_41),
.Y(n_48)
);

AOI21xp33_ASAP7_75t_L g49 ( 
.A1(n_32),
.A2(n_22),
.B(n_25),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_56),
.Y(n_83)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_55),
.Y(n_66)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx5_ASAP7_75t_SL g69 ( 
.A(n_53),
.Y(n_69)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_28),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_40),
.A2(n_26),
.B1(n_31),
.B2(n_20),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_59),
.A2(n_63),
.B1(n_65),
.B2(n_22),
.Y(n_78)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_42),
.A2(n_26),
.B1(n_31),
.B2(n_20),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_34),
.A2(n_16),
.B1(n_30),
.B2(n_15),
.Y(n_65)
);

AO22x1_ASAP7_75t_L g67 ( 
.A1(n_45),
.A2(n_34),
.B1(n_35),
.B2(n_22),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_67),
.A2(n_48),
.B(n_60),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVxp67_ASAP7_75t_SL g91 ( 
.A(n_68),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_56),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_71),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_56),
.A2(n_51),
.B1(n_39),
.B2(n_55),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_72),
.A2(n_86),
.B1(n_54),
.B2(n_48),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_36),
.C(n_30),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_24),
.B(n_43),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_53),
.A2(n_16),
.B1(n_36),
.B2(n_21),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_75),
.B(n_76),
.Y(n_87)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_58),
.A2(n_27),
.B1(n_21),
.B2(n_18),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_77),
.A2(n_79),
.B1(n_67),
.B2(n_71),
.Y(n_95)
);

O2A1O1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_78),
.A2(n_25),
.B(n_24),
.C(n_47),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_50),
.A2(n_27),
.B1(n_21),
.B2(n_18),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_84),
.B(n_60),
.Y(n_88)
);

O2A1O1Ixp33_ASAP7_75t_SL g85 ( 
.A1(n_46),
.A2(n_27),
.B(n_36),
.C(n_25),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_85),
.A2(n_47),
.B1(n_44),
.B2(n_61),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_50),
.A2(n_36),
.B1(n_25),
.B2(n_24),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_88),
.B(n_96),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_89),
.A2(n_101),
.B(n_105),
.Y(n_131)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_92),
.Y(n_115)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_93),
.A2(n_85),
.B(n_76),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_94),
.Y(n_114)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_67),
.A2(n_62),
.B1(n_64),
.B2(n_61),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_98),
.Y(n_117)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_60),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_99),
.B(n_103),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_69),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_100),
.Y(n_130)
);

AND2x2_ASAP7_75t_SL g101 ( 
.A(n_83),
.B(n_61),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_102),
.A2(n_79),
.B(n_85),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_47),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_77),
.Y(n_119)
);

AND2x2_ASAP7_75t_SL g105 ( 
.A(n_83),
.B(n_57),
.Y(n_105)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

BUFx12_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_120),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_111),
.A2(n_113),
.B1(n_105),
.B2(n_89),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_87),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_112),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_101),
.A2(n_83),
.B(n_84),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_116),
.A2(n_105),
.B1(n_108),
.B2(n_95),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_119),
.B(n_94),
.Y(n_139)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_87),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_122),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_90),
.B(n_68),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_128),
.Y(n_147)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_125),
.Y(n_156)
);

BUFx12_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_126),
.B(n_129),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_92),
.B(n_82),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_106),
.B(n_86),
.Y(n_129)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_132),
.A2(n_75),
.B1(n_120),
.B2(n_130),
.Y(n_141)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_128),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_134),
.Y(n_163)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_109),
.A2(n_105),
.B1(n_104),
.B2(n_101),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_135),
.A2(n_127),
.B(n_102),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_131),
.C(n_113),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_136),
.B(n_143),
.C(n_155),
.Y(n_177)
);

AND2x6_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_101),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_137),
.B(n_138),
.Y(n_165)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_115),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_151),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_141),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_105),
.C(n_88),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_145),
.B(n_148),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_115),
.B(n_106),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_154),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_109),
.A2(n_107),
.B1(n_102),
.B2(n_108),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_150),
.A2(n_114),
.B1(n_116),
.B2(n_126),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_123),
.Y(n_151)
);

INVx13_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_152),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_112),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_99),
.C(n_93),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_144),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_157),
.B(n_167),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_158),
.A2(n_166),
.B1(n_171),
.B2(n_175),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_147),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_159),
.B(n_169),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_137),
.B(n_125),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g188 ( 
.A(n_160),
.B(n_142),
.Y(n_188)
);

NAND3xp33_ASAP7_75t_L g162 ( 
.A(n_142),
.B(n_122),
.C(n_125),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_162),
.B(n_152),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_156),
.A2(n_111),
.B(n_129),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_147),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_168),
.B(n_173),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_146),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_145),
.A2(n_114),
.B1(n_121),
.B2(n_119),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_139),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_174),
.B(n_143),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_150),
.A2(n_121),
.B1(n_127),
.B2(n_96),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_135),
.A2(n_148),
.B1(n_155),
.B2(n_136),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_179),
.A2(n_174),
.B1(n_160),
.B2(n_165),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_130),
.Y(n_180)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_180),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_181),
.B(n_70),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_177),
.B(n_133),
.C(n_153),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_183),
.C(n_185),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_177),
.B(n_154),
.C(n_153),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_188),
.B(n_197),
.Y(n_207)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_172),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_195),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_164),
.A2(n_140),
.B1(n_138),
.B2(n_134),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_190),
.A2(n_192),
.B1(n_198),
.B2(n_0),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_179),
.B(n_110),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_202),
.C(n_44),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_164),
.A2(n_173),
.B1(n_161),
.B2(n_167),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_163),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_199),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_110),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_161),
.A2(n_132),
.B1(n_110),
.B2(n_100),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_157),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_176),
.B(n_98),
.Y(n_200)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_200),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_171),
.A2(n_80),
.B1(n_81),
.B2(n_100),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_201),
.A2(n_168),
.B1(n_180),
.B2(n_170),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_178),
.B(n_57),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_170),
.Y(n_203)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_203),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_204),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_185),
.A2(n_166),
.B(n_158),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_205),
.A2(n_211),
.B(n_215),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_175),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_197),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_193),
.B(n_176),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_183),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_212),
.B(n_213),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_187),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_182),
.B(n_98),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_214),
.B(n_220),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_44),
.C(n_70),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_216),
.B(n_217),
.C(n_192),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_202),
.B(n_44),
.C(n_70),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_218),
.B(n_1),
.Y(n_235)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_194),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_221),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_210),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_223),
.B(n_234),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_208),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_230),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_231),
.C(n_235),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_206),
.B(n_186),
.Y(n_229)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_229),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_184),
.C(n_181),
.Y(n_231)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_232),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_216),
.B(n_13),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_1),
.C(n_2),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_236),
.B(n_205),
.C(n_218),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_219),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_237),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_222),
.A2(n_217),
.B(n_204),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_241),
.C(n_235),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_207),
.C(n_203),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_6),
.C(n_7),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_228),
.A2(n_207),
.B(n_5),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_249),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_3),
.Y(n_247)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_247),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_233),
.A2(n_5),
.B(n_6),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_224),
.B(n_5),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_250),
.B(n_225),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_243),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_255),
.C(n_257),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_248),
.Y(n_254)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_254),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_236),
.C(n_223),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_237),
.Y(n_256)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_256),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_240),
.B(n_230),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_259),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_6),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_261),
.B(n_263),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_244),
.Y(n_263)
);

AO21x1_ASAP7_75t_L g266 ( 
.A1(n_259),
.A2(n_241),
.B(n_238),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_267),
.Y(n_272)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_7),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_264),
.A2(n_253),
.B1(n_260),
.B2(n_10),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_270),
.B(n_273),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_268),
.B(n_8),
.Y(n_271)
);

AOI21xp33_ASAP7_75t_L g275 ( 
.A1(n_271),
.A2(n_267),
.B(n_266),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_262),
.A2(n_8),
.B1(n_9),
.B2(n_12),
.Y(n_273)
);

AO21x1_ASAP7_75t_L g278 ( 
.A1(n_275),
.A2(n_9),
.B(n_12),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_269),
.B(n_265),
.Y(n_276)
);

OAI21x1_ASAP7_75t_L g277 ( 
.A1(n_276),
.A2(n_272),
.B(n_270),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_277),
.A2(n_278),
.B1(n_274),
.B2(n_9),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_279),
.B(n_13),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_280),
.Y(n_281)
);


endmodule