module fake_jpeg_29329_n_314 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_314);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_314;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_2),
.B(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_32),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_43),
.Y(n_90)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_32),
.Y(n_44)
);

BUFx4f_ASAP7_75t_SL g78 ( 
.A(n_44),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_30),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_46),
.B(n_54),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_19),
.B(n_0),
.Y(n_47)
);

OR2x2_ASAP7_75t_SL g70 ( 
.A(n_47),
.B(n_61),
.Y(n_70)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_25),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_56),
.B(n_57),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_19),
.B(n_18),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_30),
.B(n_0),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_58),
.B(n_69),
.Y(n_102)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_30),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_42),
.Y(n_98)
);

HAxp5_ASAP7_75t_SL g61 ( 
.A(n_38),
.B(n_1),
.CON(n_61),
.SN(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

BUFx24_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

CKINVDCx9p33_ASAP7_75t_R g103 ( 
.A(n_64),
.Y(n_103)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_67),
.Y(n_72)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_68),
.B(n_20),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_30),
.B(n_2),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_53),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_71),
.B(n_88),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_47),
.A2(n_34),
.B1(n_33),
.B2(n_23),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_74),
.A2(n_75),
.B1(n_80),
.B2(n_83),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_61),
.A2(n_31),
.B1(n_40),
.B2(n_35),
.Y(n_75)
);

CKINVDCx5p33_ASAP7_75t_R g79 ( 
.A(n_64),
.Y(n_79)
);

INVx2_ASAP7_75t_R g121 ( 
.A(n_79),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_67),
.A2(n_31),
.B1(n_40),
.B2(n_23),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_47),
.A2(n_33),
.B1(n_35),
.B2(n_23),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_50),
.A2(n_33),
.B1(n_22),
.B2(n_35),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_85),
.B(n_89),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_58),
.A2(n_22),
.B1(n_34),
.B2(n_42),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_86),
.A2(n_92),
.B1(n_99),
.B2(n_108),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_87),
.B(n_26),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_68),
.B(n_28),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_65),
.A2(n_22),
.B1(n_34),
.B2(n_39),
.Y(n_89)
);

CKINVDCx12_ASAP7_75t_R g91 ( 
.A(n_64),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_91),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_55),
.A2(n_40),
.B1(n_42),
.B2(n_39),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_100),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_69),
.A2(n_20),
.B1(n_36),
.B2(n_21),
.Y(n_99)
);

NAND3xp33_ASAP7_75t_L g100 ( 
.A(n_51),
.B(n_21),
.C(n_36),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_49),
.B(n_28),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_101),
.B(n_109),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_66),
.A2(n_42),
.B1(n_27),
.B2(n_37),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_56),
.B(n_27),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_45),
.A2(n_37),
.B1(n_26),
.B2(n_42),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_85),
.Y(n_114)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_73),
.Y(n_111)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_111),
.Y(n_151)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_73),
.Y(n_112)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_112),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_93),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_113),
.B(n_116),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_114),
.B(n_143),
.Y(n_170)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_115),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_103),
.Y(n_116)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_77),
.Y(n_118)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_118),
.Y(n_166)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_119),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_120),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_30),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_123),
.B(n_129),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_130),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_106),
.Y(n_125)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_125),
.Y(n_160)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_127),
.Y(n_169)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_128),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_102),
.B(n_63),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_103),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_104),
.Y(n_131)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_131),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_84),
.Y(n_134)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_134),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_86),
.B(n_62),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_135),
.B(n_137),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_95),
.B(n_18),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_136),
.B(n_138),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_83),
.B(n_43),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_70),
.B(n_56),
.Y(n_138)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_70),
.A2(n_44),
.B(n_43),
.C(n_16),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_139),
.A2(n_90),
.B(n_78),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_79),
.B(n_29),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_138),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_59),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_141),
.B(n_142),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_72),
.B(n_3),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_89),
.B(n_107),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_76),
.Y(n_144)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_144),
.Y(n_165)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_105),
.Y(n_146)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

OAI32xp33_ASAP7_75t_L g148 ( 
.A1(n_129),
.A2(n_72),
.A3(n_107),
.B1(n_96),
.B2(n_77),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_148),
.B(n_141),
.Y(n_183)
);

NAND2x1_ASAP7_75t_SL g149 ( 
.A(n_121),
.B(n_78),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_149),
.A2(n_131),
.B(n_143),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g155 ( 
.A1(n_132),
.A2(n_81),
.B1(n_76),
.B2(n_52),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_155),
.A2(n_176),
.B1(n_168),
.B2(n_96),
.Y(n_200)
);

AOI21xp33_ASAP7_75t_L g158 ( 
.A1(n_122),
.A2(n_78),
.B(n_4),
.Y(n_158)
);

OAI21xp33_ASAP7_75t_L g207 ( 
.A1(n_158),
.A2(n_178),
.B(n_147),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_123),
.B(n_105),
.C(n_82),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_159),
.B(n_97),
.C(n_82),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_171),
.B(n_139),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_121),
.Y(n_174)
);

INVx13_ASAP7_75t_L g203 ( 
.A(n_174),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_90),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_175),
.B(n_179),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_133),
.A2(n_81),
.B1(n_97),
.B2(n_90),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_118),
.Y(n_177)
);

BUFx24_ASAP7_75t_L g191 ( 
.A(n_177),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_126),
.B(n_96),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_161),
.B(n_126),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_190),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_163),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_182),
.B(n_185),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_183),
.A2(n_198),
.B1(n_200),
.B2(n_206),
.Y(n_218)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_156),
.Y(n_184)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_184),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_150),
.B(n_157),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_186),
.A2(n_192),
.B(n_196),
.Y(n_221)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_156),
.Y(n_187)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_187),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_149),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_188),
.B(n_189),
.Y(n_226)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_167),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_167),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_149),
.A2(n_134),
.B1(n_119),
.B2(n_131),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_161),
.B(n_135),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_193),
.B(n_154),
.C(n_153),
.Y(n_224)
);

AND2x6_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_145),
.Y(n_194)
);

A2O1A1O1Ixp25_ASAP7_75t_L g228 ( 
.A1(n_194),
.A2(n_48),
.B(n_177),
.C(n_169),
.D(n_7),
.Y(n_228)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_152),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_205),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_117),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_197),
.B(n_199),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_164),
.A2(n_114),
.B1(n_133),
.B2(n_137),
.Y(n_198)
);

INVx8_ASAP7_75t_L g199 ( 
.A(n_162),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_170),
.A2(n_133),
.B1(n_143),
.B2(n_115),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_201),
.A2(n_176),
.B1(n_170),
.B2(n_171),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_173),
.B(n_112),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_202),
.B(n_204),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g204 ( 
.A(n_173),
.B(n_159),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_175),
.B(n_164),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_170),
.A2(n_128),
.B1(n_144),
.B2(n_111),
.Y(n_206)
);

NAND3xp33_ASAP7_75t_L g214 ( 
.A(n_207),
.B(n_147),
.C(n_152),
.Y(n_214)
);

XNOR2x1_ASAP7_75t_L g209 ( 
.A(n_208),
.B(n_148),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_209),
.B(n_224),
.C(n_190),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_213),
.Y(n_234)
);

OAI21xp33_ASAP7_75t_L g240 ( 
.A1(n_214),
.A2(n_228),
.B(n_203),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_191),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_220),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_180),
.A2(n_168),
.B(n_151),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_217),
.A2(n_227),
.B(n_196),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_181),
.A2(n_165),
.B1(n_125),
.B2(n_120),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_219),
.A2(n_231),
.B1(n_191),
.B2(n_199),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_172),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_180),
.A2(n_153),
.B(n_169),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_200),
.A2(n_160),
.B1(n_162),
.B2(n_166),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_230),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_166),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_201),
.A2(n_160),
.B1(n_127),
.B2(n_84),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_29),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_232),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_3),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_233),
.B(n_5),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_235),
.B(n_242),
.Y(n_261)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_222),
.Y(n_236)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_236),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_221),
.A2(n_208),
.B(n_194),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_238),
.B(n_248),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_221),
.A2(n_206),
.B(n_184),
.Y(n_239)
);

O2A1O1Ixp33_ASAP7_75t_L g265 ( 
.A1(n_239),
.A2(n_241),
.B(n_253),
.C(n_216),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_240),
.A2(n_245),
.B1(n_215),
.B2(n_229),
.Y(n_257)
);

OAI21xp33_ASAP7_75t_L g241 ( 
.A1(n_226),
.A2(n_204),
.B(n_195),
.Y(n_241)
);

AO21x1_ASAP7_75t_L g244 ( 
.A1(n_212),
.A2(n_189),
.B(n_187),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_244),
.B(n_217),
.Y(n_254)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_222),
.Y(n_246)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_246),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_211),
.B(n_191),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_225),
.Y(n_249)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_249),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_250),
.B(n_248),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_210),
.B(n_224),
.C(n_209),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_252),
.C(n_233),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_210),
.B(n_29),
.C(n_7),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_212),
.A2(n_6),
.B(n_7),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_256),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_257),
.B(n_265),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_267),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_223),
.C(n_230),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_263),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_234),
.A2(n_213),
.B1(n_219),
.B2(n_218),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_262),
.A2(n_266),
.B1(n_245),
.B2(n_243),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_223),
.C(n_227),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_239),
.A2(n_218),
.B1(n_231),
.B2(n_225),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_242),
.B(n_228),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_237),
.B(n_8),
.Y(n_269)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_269),
.Y(n_274)
);

OAI21xp33_ASAP7_75t_L g271 ( 
.A1(n_254),
.A2(n_235),
.B(n_243),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_261),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_272),
.A2(n_246),
.B1(n_267),
.B2(n_261),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_265),
.A2(n_253),
.B(n_237),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_273),
.A2(n_276),
.B(n_262),
.Y(n_283)
);

OAI322xp33_ASAP7_75t_L g275 ( 
.A1(n_258),
.A2(n_247),
.A3(n_252),
.B1(n_238),
.B2(n_250),
.C1(n_244),
.C2(n_236),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_275),
.B(n_252),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_266),
.A2(n_244),
.B(n_247),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g278 ( 
.A(n_255),
.Y(n_278)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_278),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_249),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_281),
.Y(n_290)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_268),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_283),
.B(n_286),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_282),
.B(n_260),
.C(n_263),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_285),
.B(n_288),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_289),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_277),
.B(n_259),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_276),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_292),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_9),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_270),
.C(n_279),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_293),
.B(n_295),
.Y(n_304)
);

AOI322xp5_ASAP7_75t_L g295 ( 
.A1(n_283),
.A2(n_271),
.A3(n_273),
.B1(n_280),
.B2(n_278),
.C1(n_270),
.C2(n_14),
.Y(n_295)
);

AOI21xp33_ASAP7_75t_L g296 ( 
.A1(n_290),
.A2(n_278),
.B(n_10),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_296),
.A2(n_9),
.B(n_11),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_301),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_299),
.B(n_284),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_287),
.C(n_286),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_302),
.A2(n_11),
.B(n_12),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_298),
.B(n_9),
.Y(n_303)
);

AOI21x1_ASAP7_75t_L g309 ( 
.A1(n_303),
.A2(n_11),
.B(n_14),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_297),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_305),
.A2(n_295),
.B1(n_12),
.B2(n_13),
.Y(n_307)
);

AO21x1_ASAP7_75t_L g312 ( 
.A1(n_307),
.A2(n_308),
.B(n_309),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_306),
.A2(n_304),
.B(n_305),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_310),
.A2(n_311),
.B(n_29),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_307),
.A2(n_15),
.B(n_29),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_312),
.Y(n_314)
);


endmodule