module real_jpeg_24366_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_1),
.A2(n_26),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_1),
.A2(n_32),
.B1(n_37),
.B2(n_39),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_2),
.A2(n_36),
.B1(n_37),
.B2(n_39),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_2),
.A2(n_36),
.B1(n_60),
.B2(n_65),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_2),
.A2(n_26),
.B1(n_31),
.B2(n_36),
.Y(n_152)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g64 ( 
.A(n_5),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_6),
.A2(n_53),
.B1(n_56),
.B2(n_57),
.Y(n_52)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_6),
.A2(n_57),
.B1(n_60),
.B2(n_65),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_6),
.A2(n_37),
.B1(n_39),
.B2(n_57),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g206 ( 
.A1(n_6),
.A2(n_26),
.B1(n_31),
.B2(n_57),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_7),
.A2(n_37),
.B1(n_39),
.B2(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_7),
.A2(n_26),
.B1(n_31),
.B2(n_46),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_7),
.A2(n_46),
.B1(n_60),
.B2(n_65),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_8),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_9),
.A2(n_60),
.B1(n_65),
.B2(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_9),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_9),
.A2(n_37),
.B1(n_39),
.B2(n_84),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_9),
.A2(n_69),
.B1(n_74),
.B2(n_84),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_9),
.A2(n_26),
.B1(n_31),
.B2(n_84),
.Y(n_173)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_11),
.A2(n_56),
.B1(n_69),
.B2(n_71),
.Y(n_68)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_11),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_11),
.A2(n_60),
.B1(n_65),
.B2(n_71),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_11),
.A2(n_37),
.B1(n_39),
.B2(n_71),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_11),
.A2(n_26),
.B1(n_31),
.B2(n_71),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_13),
.A2(n_54),
.B1(n_55),
.B2(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_13),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_13),
.A2(n_60),
.B1(n_65),
.B2(n_144),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_13),
.A2(n_37),
.B1(n_39),
.B2(n_144),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_13),
.A2(n_26),
.B1(n_31),
.B2(n_144),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_14),
.A2(n_55),
.B1(n_74),
.B2(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_14),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_14),
.A2(n_60),
.B1(n_65),
.B2(n_107),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_14),
.A2(n_37),
.B1(n_39),
.B2(n_107),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_14),
.A2(n_26),
.B1(n_31),
.B2(n_107),
.Y(n_255)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_15),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_15),
.B(n_59),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_15),
.B(n_37),
.C(n_80),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_15),
.A2(n_60),
.B1(n_65),
.B2(n_168),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_15),
.B(n_122),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_15),
.A2(n_37),
.B1(n_39),
.B2(n_168),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_15),
.B(n_26),
.C(n_42),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_15),
.A2(n_25),
.B(n_256),
.Y(n_286)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_16),
.Y(n_97)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_16),
.Y(n_175)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_16),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_134),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_132),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_111),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_21),
.B(n_111),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_75),
.C(n_91),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_22),
.A2(n_75),
.B1(n_76),
.B2(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_22),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_48),
.Y(n_22)
);

AOI21xp33_ASAP7_75t_L g112 ( 
.A1(n_23),
.A2(n_24),
.B(n_50),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_33),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_24),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_24),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_24),
.A2(n_33),
.B1(n_34),
.B2(n_49),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_28),
.B(n_30),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_25),
.A2(n_30),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_25),
.A2(n_28),
.B1(n_96),
.B2(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_25),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_25),
.A2(n_173),
.B1(n_175),
.B2(n_206),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_25),
.B(n_226),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_25),
.A2(n_255),
.B(n_256),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

OA22x2_ASAP7_75t_L g44 ( 
.A1(n_26),
.A2(n_31),
.B1(n_42),
.B2(n_43),
.Y(n_44)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_31),
.B(n_283),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_40),
.B1(n_45),
.B2(n_47),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_35),
.A2(n_40),
.B1(n_47),
.B2(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_SL g39 ( 
.A(n_37),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_39),
.B1(n_42),
.B2(n_43),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_37),
.A2(n_39),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_37),
.B(n_265),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_40),
.A2(n_47),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_40),
.B(n_195),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_40),
.A2(n_47),
.B1(n_228),
.B2(n_230),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_44),
.Y(n_40)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_44),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_44),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_44),
.A2(n_87),
.B1(n_101),
.B2(n_154),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_44),
.A2(n_154),
.B(n_194),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_44),
.A2(n_194),
.B(n_229),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_44),
.B(n_168),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_45),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_47),
.B(n_195),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_58),
.B(n_66),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_52),
.A2(n_58),
.B1(n_108),
.B2(n_130),
.Y(n_129)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_55),
.Y(n_56)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_55),
.A2(n_63),
.B1(n_64),
.B2(n_74),
.Y(n_73)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

HAxp5_ASAP7_75t_SL g167 ( 
.A(n_56),
.B(n_168),
.CON(n_167),
.SN(n_167)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_58),
.B(n_68),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_58),
.A2(n_66),
.B(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_59),
.A2(n_72),
.B1(n_106),
.B2(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_59)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_60),
.A2(n_65),
.B1(n_80),
.B2(n_81),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_60),
.A2(n_64),
.B(n_167),
.C(n_169),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_60),
.B(n_221),
.Y(n_220)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND3xp33_ASAP7_75t_SL g169 ( 
.A(n_63),
.B(n_65),
.C(n_74),
.Y(n_169)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_72),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_72),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_72),
.A2(n_110),
.B(n_167),
.Y(n_196)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_86),
.B(n_90),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_86),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_78),
.A2(n_79),
.B1(n_83),
.B2(n_85),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_78),
.A2(n_79),
.B1(n_83),
.B2(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_78),
.A2(n_161),
.B(n_163),
.Y(n_160)
);

OAI21xp33_ASAP7_75t_L g232 ( 
.A1(n_78),
.A2(n_163),
.B(n_233),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_82),
.Y(n_78)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_79),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_79),
.A2(n_103),
.B(n_147),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_79),
.A2(n_147),
.B(n_202),
.Y(n_201)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_85),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_87),
.A2(n_243),
.B(n_244),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_87),
.A2(n_244),
.B(n_263),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_89),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_90),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_91),
.A2(n_92),
.B1(n_313),
.B2(n_315),
.Y(n_312)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_102),
.C(n_104),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_93),
.A2(n_94),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_98),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_95),
.A2(n_98),
.B1(n_99),
.B2(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_95),
.Y(n_156)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_97),
.Y(n_271)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_102),
.B(n_104),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_108),
.B(n_109),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_113),
.Y(n_111)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_129),
.B2(n_131),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_125),
.B1(n_126),
.B2(n_128),
.Y(n_118)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_119),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_121),
.A2(n_122),
.B1(n_162),
.B2(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_122),
.B(n_148),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_129),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_311),
.B(n_317),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_183),
.B(n_310),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_176),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_137),
.B(n_176),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_155),
.C(n_157),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_138),
.A2(n_139),
.B1(n_155),
.B2(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_149),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_145),
.B2(n_146),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_142),
.B(n_145),
.C(n_149),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_143),
.Y(n_159)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_153),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_150),
.B(n_153),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_152),
.A2(n_171),
.B1(n_172),
.B2(n_174),
.Y(n_170)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_155),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_157),
.B(n_307),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.C(n_164),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_158),
.B(n_160),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_164),
.B(n_209),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_170),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_165),
.A2(n_166),
.B1(n_170),
.B2(n_199),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_168),
.B(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_170),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_171),
.A2(n_269),
.B1(n_271),
.B2(n_272),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx3_ASAP7_75t_SL g174 ( 
.A(n_175),
.Y(n_174)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_175),
.Y(n_224)
);

INVx5_ASAP7_75t_L g285 ( 
.A(n_175),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_182),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_178),
.B(n_179),
.C(n_182),
.Y(n_316)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

O2A1O1Ixp33_ASAP7_75t_SL g183 ( 
.A1(n_184),
.A2(n_213),
.B(n_304),
.C(n_309),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_207),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_207),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_197),
.C(n_200),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_186),
.A2(n_187),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_196),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_192),
.B2(n_193),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_190),
.B(n_192),
.C(n_196),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_191),
.Y(n_202)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_197),
.A2(n_198),
.B1(n_200),
.B2(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_200),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_203),
.C(n_205),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_201),
.B(n_237),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_203),
.A2(n_204),
.B1(n_205),
.B2(n_238),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_205),
.Y(n_238)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_206),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_208),
.B(n_211),
.C(n_212),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_216),
.A2(n_297),
.B(n_303),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_245),
.B(n_296),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_234),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_218),
.B(n_234),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_227),
.C(n_231),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_219),
.B(n_292),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_222),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_222),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B(n_225),
.Y(n_222)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_225),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_226),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_227),
.A2(n_231),
.B1(n_232),
.B2(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_227),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_230),
.Y(n_243)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_239),
.B2(n_240),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_235),
.B(n_241),
.C(n_242),
.Y(n_302)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_290),
.B(n_295),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_266),
.B(n_289),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_260),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_248),
.B(n_260),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_254),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_252),
.B2(n_253),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_250),
.B(n_253),
.C(n_254),
.Y(n_294)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_255),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_259),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g279 ( 
.A(n_258),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_264),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_261),
.A2(n_262),
.B1(n_264),
.B2(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_264),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_275),
.B(n_288),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_273),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_268),
.B(n_273),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_270),
.A2(n_279),
.B(n_280),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_276),
.A2(n_281),
.B(n_287),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_278),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_286),
.Y(n_281)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_291),
.B(n_294),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_291),
.B(n_294),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_302),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_298),
.B(n_302),
.Y(n_303)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_306),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_312),
.B(n_316),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_316),
.Y(n_317)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_313),
.Y(n_315)
);


endmodule