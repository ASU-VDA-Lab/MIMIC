module fake_jpeg_25310_n_93 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_93);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_93;

wire n_10;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx5_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g17 ( 
.A(n_13),
.B(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_17),
.B(n_19),
.Y(n_29)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_22),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g27 ( 
.A(n_21),
.Y(n_27)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

AO22x1_ASAP7_75t_L g25 ( 
.A1(n_17),
.A2(n_13),
.B1(n_12),
.B2(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

NAND3xp33_ASAP7_75t_SL g26 ( 
.A(n_19),
.B(n_16),
.C(n_14),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_19),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_17),
.A2(n_16),
.B1(n_14),
.B2(n_10),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_28),
.A2(n_22),
.B1(n_18),
.B2(n_16),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_31),
.B(n_25),
.Y(n_44)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_35),
.Y(n_38)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_21),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_29),
.B(n_20),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_29),
.B(n_17),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_37),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_41),
.B(n_27),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_30),
.A2(n_25),
.B(n_28),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g49 ( 
.A1(n_43),
.A2(n_44),
.B(n_30),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_23),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_27),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_47),
.B(n_52),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_50),
.Y(n_55)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_14),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_51),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_15),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_9),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_12),
.Y(n_57)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_41),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_22),
.C(n_21),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_21),
.C(n_18),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_61),
.Y(n_69)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_66),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_64),
.B(n_65),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_61),
.A2(n_10),
.B1(n_15),
.B2(n_12),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_55),
.Y(n_66)
);

OAI322xp33_ASAP7_75t_L g67 ( 
.A1(n_56),
.A2(n_10),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_0),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_60),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_70),
.B(n_72),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_69),
.Y(n_71)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_SL g80 ( 
.A(n_75),
.B(n_54),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_63),
.C(n_62),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_78),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_69),
.C(n_56),
.Y(n_78)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_76),
.A2(n_68),
.B1(n_70),
.B2(n_4),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_79),
.A2(n_68),
.B(n_3),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_1),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_85),
.B(n_87),
.C(n_84),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_1),
.C(n_4),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_88),
.A2(n_89),
.B(n_5),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_86),
.A2(n_81),
.B1(n_6),
.B2(n_7),
.Y(n_89)
);

AOI21x1_ASAP7_75t_L g91 ( 
.A1(n_90),
.A2(n_6),
.B(n_7),
.Y(n_91)
);

AO21x1_ASAP7_75t_L g92 ( 
.A1(n_91),
.A2(n_7),
.B(n_8),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_8),
.Y(n_93)
);


endmodule