module fake_jpeg_9038_n_73 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_73);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_73;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_69;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_28;
wire n_38;
wire n_44;
wire n_36;
wire n_62;
wire n_31;
wire n_56;
wire n_67;
wire n_37;
wire n_29;
wire n_50;
wire n_43;
wire n_32;
wire n_70;
wire n_66;

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_18),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_1),
.B(n_26),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_33),
.A2(n_1),
.B1(n_27),
.B2(n_3),
.Y(n_35)
);

CKINVDCx6p67_ASAP7_75t_R g42 ( 
.A(n_35),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_2),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_15),
.Y(n_55)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_9),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_28),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_40),
.B(n_41),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_8),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_34),
.C(n_31),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_45),
.A2(n_16),
.B(n_17),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_46),
.A2(n_53),
.B(n_54),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_10),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_11),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_12),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_50),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_13),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_14),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_51),
.B(n_52),
.Y(n_59)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_SL g62 ( 
.A(n_55),
.B(n_19),
.Y(n_62)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_57),
.Y(n_65)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_62),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_42),
.A2(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_64),
.A2(n_42),
.B1(n_63),
.B2(n_44),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_58),
.C(n_65),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_61),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_68),
.B(n_59),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_69),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_70),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_71),
.A2(n_60),
.B(n_59),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_64),
.Y(n_73)
);


endmodule