module fake_netlist_1_6535_n_38 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_38);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_38;
wire n_20;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
INVx1_ASAP7_75t_L g11 ( .A(n_2), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_1), .Y(n_12) );
CKINVDCx16_ASAP7_75t_R g13 ( .A(n_8), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_8), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_10), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_1), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_3), .Y(n_17) );
AOI21xp5_ASAP7_75t_L g18 ( .A1(n_12), .A2(n_0), .B(n_2), .Y(n_18) );
CKINVDCx8_ASAP7_75t_R g19 ( .A(n_13), .Y(n_19) );
O2A1O1Ixp5_ASAP7_75t_L g20 ( .A1(n_12), .A2(n_0), .B(n_3), .C(n_4), .Y(n_20) );
NAND2xp5_ASAP7_75t_L g21 ( .A(n_13), .B(n_4), .Y(n_21) );
A2O1A1Ixp33_ASAP7_75t_L g22 ( .A1(n_12), .A2(n_5), .B(n_6), .C(n_7), .Y(n_22) );
NOR2x1_ASAP7_75t_L g23 ( .A(n_21), .B(n_11), .Y(n_23) );
NOR2xp33_ASAP7_75t_R g24 ( .A(n_19), .B(n_17), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_18), .B(n_17), .Y(n_25) );
AOI22xp33_ASAP7_75t_L g26 ( .A1(n_20), .A2(n_11), .B1(n_14), .B2(n_15), .Y(n_26) );
NAND2xp5_ASAP7_75t_L g27 ( .A(n_23), .B(n_14), .Y(n_27) );
OR2x2_ASAP7_75t_L g28 ( .A(n_25), .B(n_16), .Y(n_28) );
NAND2xp5_ASAP7_75t_L g29 ( .A(n_23), .B(n_22), .Y(n_29) );
AND2x2_ASAP7_75t_L g30 ( .A(n_28), .B(n_24), .Y(n_30) );
AOI22xp5_ASAP7_75t_L g31 ( .A1(n_29), .A2(n_26), .B1(n_22), .B2(n_7), .Y(n_31) );
NAND2xp33_ASAP7_75t_SL g32 ( .A(n_30), .B(n_27), .Y(n_32) );
AND2x2_ASAP7_75t_L g33 ( .A(n_31), .B(n_5), .Y(n_33) );
CKINVDCx5p33_ASAP7_75t_R g34 ( .A(n_32), .Y(n_34) );
INVx2_ASAP7_75t_L g35 ( .A(n_33), .Y(n_35) );
INVx2_ASAP7_75t_L g36 ( .A(n_35), .Y(n_36) );
CKINVDCx20_ASAP7_75t_R g37 ( .A(n_34), .Y(n_37) );
AOI22xp5_ASAP7_75t_SL g38 ( .A1(n_36), .A2(n_6), .B1(n_9), .B2(n_37), .Y(n_38) );
endmodule