module fake_netlist_1_7641_n_39 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_39);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_39;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_8), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_3), .Y(n_12) );
NOR2xp33_ASAP7_75t_R g13 ( .A(n_9), .B(n_10), .Y(n_13) );
BUFx3_ASAP7_75t_L g14 ( .A(n_6), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_5), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_0), .Y(n_16) );
BUFx6f_ASAP7_75t_L g17 ( .A(n_3), .Y(n_17) );
AND2x2_ASAP7_75t_L g18 ( .A(n_14), .B(n_0), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_14), .Y(n_19) );
O2A1O1Ixp33_ASAP7_75t_L g20 ( .A1(n_15), .A2(n_1), .B(n_2), .C(n_4), .Y(n_20) );
NOR2xp33_ASAP7_75t_SL g21 ( .A(n_11), .B(n_7), .Y(n_21) );
INVx5_ASAP7_75t_L g22 ( .A(n_17), .Y(n_22) );
INVxp67_ASAP7_75t_L g23 ( .A(n_18), .Y(n_23) );
AOI22xp33_ASAP7_75t_L g24 ( .A1(n_18), .A2(n_15), .B1(n_14), .B2(n_17), .Y(n_24) );
AND2x2_ASAP7_75t_L g25 ( .A(n_19), .B(n_16), .Y(n_25) );
OAI21xp5_ASAP7_75t_SL g26 ( .A1(n_20), .A2(n_17), .B(n_12), .Y(n_26) );
INVx2_ASAP7_75t_L g27 ( .A(n_25), .Y(n_27) );
NAND2xp5_ASAP7_75t_L g28 ( .A(n_23), .B(n_19), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_25), .Y(n_29) );
HB1xp67_ASAP7_75t_L g30 ( .A(n_27), .Y(n_30) );
OAI221xp5_ASAP7_75t_L g31 ( .A1(n_29), .A2(n_26), .B1(n_24), .B2(n_21), .C(n_17), .Y(n_31) );
OAI211xp5_ASAP7_75t_L g32 ( .A1(n_31), .A2(n_27), .B(n_28), .C(n_13), .Y(n_32) );
AOI222xp33_ASAP7_75t_L g33 ( .A1(n_30), .A2(n_17), .B1(n_22), .B2(n_4), .C1(n_5), .C2(n_6), .Y(n_33) );
INVx2_ASAP7_75t_L g34 ( .A(n_33), .Y(n_34) );
CKINVDCx5p33_ASAP7_75t_R g35 ( .A(n_32), .Y(n_35) );
CKINVDCx5p33_ASAP7_75t_R g36 ( .A(n_33), .Y(n_36) );
AOI22xp5_ASAP7_75t_L g37 ( .A1(n_36), .A2(n_22), .B1(n_1), .B2(n_2), .Y(n_37) );
OAI22x1_ASAP7_75t_L g38 ( .A1(n_34), .A2(n_22), .B1(n_36), .B2(n_35), .Y(n_38) );
AOI22xp5_ASAP7_75t_L g39 ( .A1(n_38), .A2(n_22), .B1(n_34), .B2(n_37), .Y(n_39) );
endmodule