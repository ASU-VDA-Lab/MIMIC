module real_aes_16435_n_267 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_267);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_267;
wire n_476;
wire n_887;
wire n_599;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1284;
wire n_1250;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_1380;
wire n_488;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_564;
wire n_638;
wire n_1361;
wire n_510;
wire n_1358;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_856;
wire n_594;
wire n_1146;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_1378;
wire n_524;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1143;
wire n_929;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1156;
wire n_988;
wire n_921;
wire n_1396;
wire n_1176;
wire n_640;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_578;
wire n_372;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_1049;
wire n_466;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_269;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_1390;
wire n_272;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp5_ASAP7_75t_L g1167 ( .A1(n_0), .A2(n_206), .B1(n_1140), .B2(n_1155), .Y(n_1167) );
AOI22xp33_ASAP7_75t_SL g940 ( .A1(n_1), .A2(n_83), .B1(n_477), .B2(n_680), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_1), .A2(n_247), .B1(n_415), .B2(n_418), .Y(n_948) );
INVx1_ASAP7_75t_L g557 ( .A(n_2), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g577 ( .A1(n_2), .A2(n_110), .B1(n_418), .B2(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g944 ( .A(n_3), .Y(n_944) );
OAI211xp5_ASAP7_75t_L g647 ( .A1(n_4), .A2(n_648), .B(n_651), .C(n_662), .Y(n_647) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_4), .B(n_300), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g1105 ( .A1(n_5), .A2(n_128), .B1(n_1031), .B2(n_1033), .Y(n_1105) );
AOI22xp33_ASAP7_75t_SL g1119 ( .A1(n_5), .A2(n_135), .B1(n_415), .B2(n_417), .Y(n_1119) );
AOI22xp33_ASAP7_75t_L g1163 ( .A1(n_6), .A2(n_57), .B1(n_1140), .B2(n_1155), .Y(n_1163) );
AOI22xp33_ASAP7_75t_SL g470 ( .A1(n_7), .A2(n_157), .B1(n_351), .B2(n_471), .Y(n_470) );
INVxp67_ASAP7_75t_SL g521 ( .A(n_7), .Y(n_521) );
INVx1_ASAP7_75t_L g1025 ( .A(n_8), .Y(n_1025) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_9), .A2(n_84), .B1(n_680), .B2(n_877), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g896 ( .A1(n_9), .A2(n_58), .B1(n_897), .B2(n_898), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g1070 ( .A1(n_10), .A2(n_219), .B1(n_418), .B2(n_1071), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g1088 ( .A1(n_10), .A2(n_252), .B1(n_340), .B2(n_874), .Y(n_1088) );
INVx1_ASAP7_75t_L g730 ( .A(n_11), .Y(n_730) );
AO22x1_ASAP7_75t_L g769 ( .A1(n_11), .A2(n_155), .B1(n_403), .B2(n_658), .Y(n_769) );
INVx1_ASAP7_75t_L g281 ( .A(n_12), .Y(n_281) );
AND2x2_ASAP7_75t_L g332 ( .A(n_12), .B(n_229), .Y(n_332) );
AND2x2_ASAP7_75t_L g393 ( .A(n_12), .B(n_394), .Y(n_393) );
NOR2xp33_ASAP7_75t_L g767 ( .A(n_12), .B(n_291), .Y(n_767) );
INVx1_ASAP7_75t_L g742 ( .A(n_13), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_13), .A2(n_108), .B1(n_408), .B2(n_654), .Y(n_768) );
AOI221xp5_ASAP7_75t_L g938 ( .A1(n_14), .A2(n_159), .B1(n_632), .B2(n_935), .C(n_939), .Y(n_938) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_14), .A2(n_68), .B1(n_418), .B2(n_826), .Y(n_950) );
AOI22xp33_ASAP7_75t_SL g1104 ( .A1(n_15), .A2(n_167), .B1(n_457), .B2(n_471), .Y(n_1104) );
AOI221xp5_ASAP7_75t_L g1117 ( .A1(n_15), .A2(n_20), .B1(n_412), .B2(n_430), .C(n_1118), .Y(n_1117) );
INVx1_ASAP7_75t_L g1356 ( .A(n_16), .Y(n_1356) );
OAI221xp5_ASAP7_75t_L g1369 ( .A1(n_16), .A2(n_165), .B1(n_612), .B2(n_1048), .C(n_1370), .Y(n_1369) );
INVx2_ASAP7_75t_L g1143 ( .A(n_17), .Y(n_1143) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_17), .B(n_114), .Y(n_1145) );
AND2x2_ASAP7_75t_L g1151 ( .A(n_17), .B(n_1149), .Y(n_1151) );
CKINVDCx5p33_ASAP7_75t_R g932 ( .A(n_18), .Y(n_932) );
OAI22xp5_ASAP7_75t_L g1082 ( .A1(n_19), .A2(n_101), .B1(n_300), .B2(n_544), .Y(n_1082) );
AOI22xp33_ASAP7_75t_SL g1109 ( .A1(n_20), .A2(n_35), .B1(n_353), .B2(n_844), .Y(n_1109) );
INVx1_ASAP7_75t_L g1102 ( .A(n_21), .Y(n_1102) );
OAI22xp33_ASAP7_75t_L g1110 ( .A1(n_22), .A2(n_212), .B1(n_481), .B2(n_487), .Y(n_1110) );
INVx1_ASAP7_75t_L g1122 ( .A(n_22), .Y(n_1122) );
AOI22xp5_ASAP7_75t_L g1180 ( .A1(n_23), .A2(n_34), .B1(n_1147), .B2(n_1150), .Y(n_1180) );
XNOR2xp5_ASAP7_75t_L g597 ( .A(n_24), .B(n_598), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g1032 ( .A1(n_25), .A2(n_51), .B1(n_366), .B2(n_1033), .Y(n_1032) );
AOI22xp33_ASAP7_75t_L g1045 ( .A1(n_25), .A2(n_265), .B1(n_593), .B2(n_897), .Y(n_1045) );
INVx1_ASAP7_75t_L g583 ( .A(n_26), .Y(n_583) );
AOI22xp33_ASAP7_75t_SL g558 ( .A1(n_27), .A2(n_82), .B1(n_351), .B2(n_559), .Y(n_558) );
AOI221xp5_ASAP7_75t_L g576 ( .A1(n_27), .A2(n_262), .B1(n_411), .B2(n_412), .C(n_500), .Y(n_576) );
AOI22xp5_ASAP7_75t_L g1166 ( .A1(n_28), .A2(n_152), .B1(n_1147), .B2(n_1150), .Y(n_1166) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_29), .A2(n_163), .B1(n_355), .B2(n_360), .Y(n_354) );
AOI221xp5_ASAP7_75t_L g425 ( .A1(n_29), .A2(n_227), .B1(n_426), .B2(n_430), .C(n_434), .Y(n_425) );
INVx1_ASAP7_75t_L g582 ( .A(n_30), .Y(n_582) );
OAI211xp5_ASAP7_75t_L g663 ( .A1(n_31), .A2(n_664), .B(n_665), .C(n_666), .Y(n_663) );
INVx1_ASAP7_75t_L g706 ( .A(n_31), .Y(n_706) );
INVx1_ASAP7_75t_L g1023 ( .A(n_32), .Y(n_1023) );
OAI221xp5_ASAP7_75t_L g1047 ( .A1(n_32), .A2(n_149), .B1(n_509), .B2(n_1048), .C(n_1049), .Y(n_1047) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_33), .A2(n_262), .B1(n_351), .B2(n_559), .Y(n_568) );
AOI22xp33_ASAP7_75t_SL g592 ( .A1(n_33), .A2(n_82), .B1(n_424), .B2(n_593), .Y(n_592) );
A2O1A1Ixp33_ASAP7_75t_L g1123 ( .A1(n_35), .A2(n_914), .B(n_1124), .C(n_1130), .Y(n_1123) );
AOI22xp33_ASAP7_75t_SL g1029 ( .A1(n_36), .A2(n_265), .B1(n_1030), .B2(n_1031), .Y(n_1029) );
AOI221xp5_ASAP7_75t_L g1056 ( .A1(n_36), .A2(n_51), .B1(n_654), .B2(n_656), .C(n_1057), .Y(n_1056) );
AOI22xp33_ASAP7_75t_SL g1363 ( .A1(n_37), .A2(n_98), .B1(n_374), .B2(n_844), .Y(n_1363) );
AOI221xp5_ASAP7_75t_L g1380 ( .A1(n_37), .A2(n_174), .B1(n_412), .B2(n_426), .C(n_530), .Y(n_1380) );
NAND2xp5_ASAP7_75t_SL g827 ( .A(n_38), .B(n_407), .Y(n_827) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_38), .A2(n_168), .B1(n_374), .B2(n_851), .Y(n_850) );
XNOR2xp5_ASAP7_75t_L g1061 ( .A(n_39), .B(n_1062), .Y(n_1061) );
AOI22xp33_ASAP7_75t_L g1139 ( .A1(n_39), .A2(n_103), .B1(n_1140), .B2(n_1144), .Y(n_1139) );
INVx1_ASAP7_75t_L g395 ( .A(n_40), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g831 ( .A1(n_41), .A2(n_168), .B1(n_403), .B2(n_580), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g843 ( .A1(n_41), .A2(n_245), .B1(n_374), .B2(n_844), .Y(n_843) );
AOI22xp5_ASAP7_75t_L g1175 ( .A1(n_42), .A2(n_100), .B1(n_1140), .B2(n_1176), .Y(n_1175) );
OAI22xp5_ASAP7_75t_L g1113 ( .A1(n_43), .A2(n_67), .B1(n_300), .B2(n_446), .Y(n_1113) );
OAI211xp5_ASAP7_75t_L g1115 ( .A1(n_43), .A2(n_495), .B(n_1116), .C(n_1120), .Y(n_1115) );
XOR2x2_ASAP7_75t_L g955 ( .A(n_44), .B(n_956), .Y(n_955) );
AOI22xp33_ASAP7_75t_L g1075 ( .A1(n_45), .A2(n_176), .B1(n_418), .B2(n_1076), .Y(n_1075) );
AOI22xp33_ASAP7_75t_SL g1090 ( .A1(n_45), .A2(n_129), .B1(n_357), .B2(n_477), .Y(n_1090) );
AOI21xp33_ASAP7_75t_L g618 ( .A1(n_46), .A2(n_411), .B(n_434), .Y(n_618) );
INVx1_ASAP7_75t_L g626 ( .A(n_46), .Y(n_626) );
XNOR2x2_ASAP7_75t_L g1096 ( .A(n_47), .B(n_1097), .Y(n_1096) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_48), .A2(n_227), .B1(n_355), .B2(n_366), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_48), .A2(n_163), .B1(n_415), .B2(n_417), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_49), .A2(n_73), .B1(n_580), .B2(n_607), .Y(n_652) );
AOI22xp33_ASAP7_75t_SL g678 ( .A1(n_49), .A2(n_259), .B1(n_351), .B2(n_559), .Y(n_678) );
AOI22xp33_ASAP7_75t_SL g881 ( .A1(n_50), .A2(n_140), .B1(n_882), .B2(n_883), .Y(n_881) );
INVxp67_ASAP7_75t_SL g912 ( .A(n_50), .Y(n_912) );
INVx1_ASAP7_75t_L g307 ( .A(n_52), .Y(n_307) );
INVx1_ASAP7_75t_L g324 ( .A(n_52), .Y(n_324) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_53), .A2(n_134), .B1(n_351), .B2(n_374), .Y(n_373) );
AOI221xp5_ASAP7_75t_L g406 ( .A1(n_53), .A2(n_80), .B1(n_407), .B2(n_410), .C(n_412), .Y(n_406) );
INVx1_ASAP7_75t_L g542 ( .A(n_54), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_55), .A2(n_204), .B1(n_415), .B2(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g627 ( .A(n_55), .Y(n_627) );
INVx1_ASAP7_75t_L g812 ( .A(n_56), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_58), .A2(n_146), .B1(n_476), .B2(n_680), .Y(n_878) );
AOI22xp5_ASAP7_75t_L g1189 ( .A1(n_59), .A2(n_142), .B1(n_1140), .B2(n_1176), .Y(n_1189) );
AOI22xp33_ASAP7_75t_L g1146 ( .A1(n_60), .A2(n_228), .B1(n_1147), .B2(n_1150), .Y(n_1146) );
AOI22xp33_ASAP7_75t_L g1106 ( .A1(n_61), .A2(n_135), .B1(n_1031), .B2(n_1107), .Y(n_1106) );
AOI221xp5_ASAP7_75t_L g1125 ( .A1(n_61), .A2(n_128), .B1(n_532), .B2(n_1126), .C(n_1127), .Y(n_1125) );
INVx1_ASAP7_75t_L g1026 ( .A(n_62), .Y(n_1026) );
INVx1_ASAP7_75t_L g274 ( .A(n_63), .Y(n_274) );
AOI221xp5_ASAP7_75t_L g602 ( .A1(n_64), .A2(n_236), .B1(n_412), .B2(n_603), .C(n_604), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_64), .A2(n_261), .B1(n_340), .B2(n_351), .Y(n_628) );
INVx2_ASAP7_75t_L g310 ( .A(n_65), .Y(n_310) );
INVx1_ASAP7_75t_L g801 ( .A(n_66), .Y(n_801) );
AOI221xp5_ASAP7_75t_L g934 ( .A1(n_68), .A2(n_78), .B1(n_353), .B2(n_935), .C(n_936), .Y(n_934) );
AOI221xp5_ASAP7_75t_L g961 ( .A1(n_69), .A2(n_125), .B1(n_501), .B2(n_962), .C(n_964), .Y(n_961) );
INVx1_ASAP7_75t_L g1004 ( .A(n_69), .Y(n_1004) );
INVx1_ASAP7_75t_L g887 ( .A(n_70), .Y(n_887) );
CKINVDCx5p33_ASAP7_75t_R g1018 ( .A(n_71), .Y(n_1018) );
INVx1_ASAP7_75t_L g928 ( .A(n_72), .Y(n_928) );
AOI22xp33_ASAP7_75t_SL g683 ( .A1(n_73), .A2(n_107), .B1(n_351), .B2(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g927 ( .A(n_74), .Y(n_927) );
AOI22xp33_ASAP7_75t_SL g479 ( .A1(n_75), .A2(n_77), .B1(n_351), .B2(n_353), .Y(n_479) );
AOI221xp5_ASAP7_75t_L g497 ( .A1(n_75), .A2(n_157), .B1(n_410), .B2(n_498), .C(n_501), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g971 ( .A1(n_76), .A2(n_137), .B1(n_415), .B2(n_967), .Y(n_971) );
INVx1_ASAP7_75t_L g991 ( .A(n_76), .Y(n_991) );
INVxp67_ASAP7_75t_SL g526 ( .A(n_77), .Y(n_526) );
AOI221xp5_ASAP7_75t_L g947 ( .A1(n_78), .A2(n_159), .B1(n_432), .B2(n_500), .C(n_661), .Y(n_947) );
AOI22xp33_ASAP7_75t_SL g472 ( .A1(n_79), .A2(n_193), .B1(n_473), .B2(n_476), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_79), .A2(n_141), .B1(n_415), .B2(n_417), .Y(n_502) );
AOI22xp33_ASAP7_75t_SL g350 ( .A1(n_80), .A2(n_221), .B1(n_351), .B2(n_353), .Y(n_350) );
INVx1_ASAP7_75t_L g853 ( .A(n_81), .Y(n_853) );
AOI221xp5_ASAP7_75t_L g951 ( .A1(n_83), .A2(n_87), .B1(n_432), .B2(n_591), .C(n_603), .Y(n_951) );
INVx1_ASAP7_75t_L g909 ( .A(n_84), .Y(n_909) );
OAI22xp5_ASAP7_75t_L g1019 ( .A1(n_85), .A2(n_214), .B1(n_446), .B2(n_492), .Y(n_1019) );
OAI211xp5_ASAP7_75t_L g1039 ( .A1(n_85), .A2(n_574), .B(n_1040), .C(n_1046), .Y(n_1039) );
OAI22xp33_ASAP7_75t_L g480 ( .A1(n_86), .A2(n_254), .B1(n_481), .B2(n_487), .Y(n_480) );
INVx1_ASAP7_75t_L g505 ( .A(n_86), .Y(n_505) );
AOI22xp33_ASAP7_75t_SL g937 ( .A1(n_87), .A2(n_247), .B1(n_477), .B2(n_680), .Y(n_937) );
AOI22xp33_ASAP7_75t_L g1362 ( .A1(n_88), .A2(n_184), .B1(n_366), .B2(n_737), .Y(n_1362) );
AOI22xp33_ASAP7_75t_L g1379 ( .A1(n_88), .A2(n_96), .B1(n_898), .B2(n_1071), .Y(n_1379) );
OAI222xp33_ASAP7_75t_L g753 ( .A1(n_89), .A2(n_211), .B1(n_754), .B2(n_756), .C1(n_758), .C2(n_760), .Y(n_753) );
INVx1_ASAP7_75t_L g773 ( .A(n_89), .Y(n_773) );
AOI22xp5_ASAP7_75t_L g1156 ( .A1(n_90), .A2(n_132), .B1(n_1147), .B2(n_1150), .Y(n_1156) );
INVx1_ASAP7_75t_L g867 ( .A(n_91), .Y(n_867) );
OAI222xp33_ASAP7_75t_L g901 ( .A1(n_91), .A2(n_131), .B1(n_512), .B2(n_902), .C1(n_903), .C2(n_910), .Y(n_901) );
OAI22xp5_ASAP7_75t_SL g820 ( .A1(n_92), .A2(n_112), .B1(n_821), .B2(n_822), .Y(n_820) );
OAI21xp33_ASAP7_75t_L g833 ( .A1(n_92), .A2(n_693), .B(n_834), .Y(n_833) );
INVx1_ASAP7_75t_L g973 ( .A(n_93), .Y(n_973) );
INVx1_ASAP7_75t_L g317 ( .A(n_94), .Y(n_317) );
AOI22xp33_ASAP7_75t_L g1172 ( .A1(n_95), .A2(n_116), .B1(n_1140), .B2(n_1155), .Y(n_1172) );
AOI22xp33_ASAP7_75t_L g1361 ( .A1(n_96), .A2(n_118), .B1(n_366), .B2(n_473), .Y(n_1361) );
INVx1_ASAP7_75t_L g1066 ( .A(n_97), .Y(n_1066) );
INVxp67_ASAP7_75t_SL g1372 ( .A(n_98), .Y(n_1372) );
CKINVDCx5p33_ASAP7_75t_R g735 ( .A(n_99), .Y(n_735) );
OAI211xp5_ASAP7_75t_L g1072 ( .A1(n_101), .A2(n_574), .B(n_1073), .C(n_1077), .Y(n_1072) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_102), .Y(n_276) );
AND2x2_ASAP7_75t_L g1141 ( .A(n_102), .B(n_274), .Y(n_1141) );
CKINVDCx5p33_ASAP7_75t_R g719 ( .A(n_104), .Y(n_719) );
CKINVDCx5p33_ASAP7_75t_R g931 ( .A(n_105), .Y(n_931) );
CKINVDCx5p33_ASAP7_75t_R g614 ( .A(n_106), .Y(n_614) );
AOI221xp5_ASAP7_75t_SL g659 ( .A1(n_107), .A2(n_259), .B1(n_408), .B2(n_660), .C(n_661), .Y(n_659) );
INVx1_ASAP7_75t_L g738 ( .A(n_108), .Y(n_738) );
CKINVDCx5p33_ASAP7_75t_R g564 ( .A(n_109), .Y(n_564) );
INVx1_ASAP7_75t_L g567 ( .A(n_110), .Y(n_567) );
OAI211xp5_ASAP7_75t_L g814 ( .A1(n_111), .A2(n_815), .B(n_816), .C(n_817), .Y(n_814) );
INVxp33_ASAP7_75t_SL g835 ( .A(n_111), .Y(n_835) );
INVxp67_ASAP7_75t_SL g857 ( .A(n_112), .Y(n_857) );
CKINVDCx5p33_ASAP7_75t_R g862 ( .A(n_113), .Y(n_862) );
AND2x2_ASAP7_75t_L g1142 ( .A(n_114), .B(n_1143), .Y(n_1142) );
INVx1_ASAP7_75t_L g1149 ( .A(n_114), .Y(n_1149) );
CKINVDCx5p33_ASAP7_75t_R g670 ( .A(n_115), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g1188 ( .A1(n_117), .A2(n_178), .B1(n_1147), .B2(n_1150), .Y(n_1188) );
AOI221xp5_ASAP7_75t_L g1373 ( .A1(n_118), .A2(n_184), .B1(n_591), .B2(n_1374), .C(n_1375), .Y(n_1373) );
OAI22xp33_ASAP7_75t_L g1364 ( .A1(n_119), .A2(n_180), .B1(n_487), .B2(n_1094), .Y(n_1364) );
INVx1_ASAP7_75t_L g1383 ( .A(n_119), .Y(n_1383) );
INVx1_ASAP7_75t_L g976 ( .A(n_120), .Y(n_976) );
INVx1_ASAP7_75t_L g552 ( .A(n_121), .Y(n_552) );
AOI21xp33_ASAP7_75t_L g590 ( .A1(n_121), .A2(n_411), .B(n_591), .Y(n_590) );
INVx2_ASAP7_75t_L g312 ( .A(n_122), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_122), .B(n_310), .Y(n_327) );
INVx1_ASAP7_75t_L g372 ( .A(n_122), .Y(n_372) );
AOI21xp33_ASAP7_75t_L g1069 ( .A1(n_123), .A2(n_531), .B(n_656), .Y(n_1069) );
AOI22xp33_ASAP7_75t_L g1089 ( .A1(n_123), .A2(n_176), .B1(n_477), .B2(n_695), .Y(n_1089) );
OAI22xp5_ASAP7_75t_L g673 ( .A1(n_124), .A2(n_148), .B1(n_664), .B2(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g690 ( .A(n_124), .Y(n_690) );
INVx1_ASAP7_75t_L g992 ( .A(n_125), .Y(n_992) );
INVx1_ASAP7_75t_L g748 ( .A(n_126), .Y(n_748) );
NAND2xp33_ASAP7_75t_SL g791 ( .A(n_126), .B(n_408), .Y(n_791) );
NOR2xp33_ASAP7_75t_L g1010 ( .A(n_127), .B(n_319), .Y(n_1010) );
INVxp67_ASAP7_75t_SL g1068 ( .A(n_129), .Y(n_1068) );
OAI22xp5_ASAP7_75t_L g543 ( .A1(n_130), .A2(n_231), .B1(n_492), .B2(n_544), .Y(n_543) );
OAI211xp5_ASAP7_75t_L g573 ( .A1(n_130), .A2(n_574), .B(n_575), .C(n_581), .Y(n_573) );
INVx1_ASAP7_75t_L g866 ( .A(n_131), .Y(n_866) );
INVx1_ASAP7_75t_L g1081 ( .A(n_133), .Y(n_1081) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_134), .A2(n_221), .B1(n_417), .B2(n_424), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g1173 ( .A1(n_136), .A2(n_240), .B1(n_1147), .B2(n_1150), .Y(n_1173) );
INVx1_ASAP7_75t_L g1000 ( .A(n_137), .Y(n_1000) );
AOI22xp5_ASAP7_75t_L g1154 ( .A1(n_138), .A2(n_139), .B1(n_1140), .B2(n_1155), .Y(n_1154) );
XOR2x2_ASAP7_75t_L g1350 ( .A(n_139), .B(n_1351), .Y(n_1350) );
AOI22xp33_ASAP7_75t_L g1388 ( .A1(n_139), .A2(n_1389), .B1(n_1392), .B2(n_1395), .Y(n_1388) );
AOI221xp5_ASAP7_75t_L g895 ( .A1(n_140), .A2(n_256), .B1(n_501), .B2(n_528), .C(n_530), .Y(n_895) );
AOI22xp33_ASAP7_75t_SL g478 ( .A1(n_141), .A2(n_239), .B1(n_473), .B2(n_476), .Y(n_478) );
AOI22xp33_ASAP7_75t_SL g1036 ( .A1(n_143), .A2(n_161), .B1(n_353), .B2(n_1037), .Y(n_1036) );
AOI221xp5_ASAP7_75t_L g1041 ( .A1(n_143), .A2(n_187), .B1(n_501), .B2(n_1042), .C(n_1043), .Y(n_1041) );
INVx1_ASAP7_75t_L g1079 ( .A(n_144), .Y(n_1079) );
OAI22xp33_ASAP7_75t_L g1093 ( .A1(n_144), .A2(n_188), .B1(n_693), .B2(n_1094), .Y(n_1093) );
INVx1_ASAP7_75t_L g610 ( .A(n_145), .Y(n_610) );
INVx1_ASAP7_75t_L g905 ( .A(n_146), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g1162 ( .A1(n_147), .A2(n_151), .B1(n_1147), .B2(n_1150), .Y(n_1162) );
INVx1_ASAP7_75t_L g704 ( .A(n_148), .Y(n_704) );
INVx1_ASAP7_75t_L g1022 ( .A(n_149), .Y(n_1022) );
CKINVDCx16_ASAP7_75t_R g755 ( .A(n_150), .Y(n_755) );
NAND5xp2_ASAP7_75t_L g645 ( .A(n_153), .B(n_646), .C(n_676), .D(n_691), .E(n_701), .Y(n_645) );
INVx1_ASAP7_75t_L g710 ( .A(n_153), .Y(n_710) );
AOI22xp33_ASAP7_75t_SL g619 ( .A1(n_154), .A2(n_261), .B1(n_403), .B2(n_424), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_154), .A2(n_236), .B1(n_351), .B2(n_632), .Y(n_631) );
AOI21xp5_ASAP7_75t_L g749 ( .A1(n_155), .A2(n_687), .B(n_750), .Y(n_749) );
OAI22xp5_ASAP7_75t_L g491 ( .A1(n_156), .A2(n_181), .B1(n_446), .B2(n_492), .Y(n_491) );
OAI211xp5_ASAP7_75t_SL g494 ( .A1(n_156), .A2(n_495), .B(n_496), .C(n_503), .Y(n_494) );
INVx1_ASAP7_75t_L g795 ( .A(n_158), .Y(n_795) );
INVx1_ASAP7_75t_L g609 ( .A(n_160), .Y(n_609) );
INVxp67_ASAP7_75t_SL g1055 ( .A(n_161), .Y(n_1055) );
BUFx3_ASAP7_75t_L g304 ( .A(n_162), .Y(n_304) );
AOI22xp5_ASAP7_75t_L g1177 ( .A1(n_164), .A2(n_166), .B1(n_1147), .B2(n_1150), .Y(n_1177) );
INVx1_ASAP7_75t_L g1355 ( .A(n_165), .Y(n_1355) );
NAND2xp5_ASAP7_75t_L g1128 ( .A(n_167), .B(n_1129), .Y(n_1128) );
AOI22xp5_ASAP7_75t_L g1181 ( .A1(n_169), .A2(n_230), .B1(n_1140), .B2(n_1155), .Y(n_1181) );
AOI221xp5_ASAP7_75t_L g1074 ( .A1(n_170), .A2(n_252), .B1(n_500), .B2(n_501), .C(n_962), .Y(n_1074) );
AOI22xp33_ASAP7_75t_L g1092 ( .A1(n_170), .A2(n_219), .B1(n_353), .B2(n_882), .Y(n_1092) );
INVx1_ASAP7_75t_L g981 ( .A(n_171), .Y(n_981) );
OAI21xp33_ASAP7_75t_L g885 ( .A1(n_172), .A2(n_446), .B(n_886), .Y(n_885) );
BUFx6f_ASAP7_75t_L g288 ( .A(n_173), .Y(n_288) );
AOI22xp33_ASAP7_75t_SL g1358 ( .A1(n_174), .A2(n_234), .B1(n_353), .B2(n_1359), .Y(n_1358) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_175), .A2(n_210), .B1(n_607), .B2(n_658), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_175), .A2(n_203), .B1(n_477), .B2(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g945 ( .A(n_177), .Y(n_945) );
CKINVDCx20_ASAP7_75t_R g376 ( .A(n_179), .Y(n_376) );
INVx1_ASAP7_75t_L g1382 ( .A(n_180), .Y(n_1382) );
AOI22xp33_ASAP7_75t_SL g1028 ( .A1(n_182), .A2(n_187), .B1(n_351), .B2(n_883), .Y(n_1028) );
INVx1_ASAP7_75t_L g1052 ( .A(n_182), .Y(n_1052) );
OAI21xp5_ASAP7_75t_SL g952 ( .A1(n_183), .A2(n_544), .B(n_953), .Y(n_952) );
INVx1_ASAP7_75t_L g888 ( .A(n_185), .Y(n_888) );
INVx1_ASAP7_75t_L g721 ( .A(n_186), .Y(n_721) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_186), .B(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g1078 ( .A(n_188), .Y(n_1078) );
XOR2xp5_ASAP7_75t_L g461 ( .A(n_189), .B(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g870 ( .A(n_190), .Y(n_870) );
XOR2xp5_ASAP7_75t_L g1393 ( .A(n_191), .B(n_1394), .Y(n_1393) );
OAI221xp5_ASAP7_75t_L g611 ( .A1(n_192), .A2(n_237), .B1(n_513), .B2(n_612), .C(n_613), .Y(n_611) );
OAI22xp33_ASAP7_75t_L g634 ( .A1(n_192), .A2(n_237), .B1(n_378), .B2(n_570), .Y(n_634) );
AOI221xp5_ASAP7_75t_L g527 ( .A1(n_193), .A2(n_239), .B1(n_528), .B2(n_530), .C(n_532), .Y(n_527) );
AOI21xp33_ASAP7_75t_L g830 ( .A1(n_194), .A2(n_411), .B(n_656), .Y(n_830) );
INVx1_ASAP7_75t_L g840 ( .A(n_194), .Y(n_840) );
INVx1_ASAP7_75t_L g700 ( .A(n_195), .Y(n_700) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_196), .Y(n_336) );
OAI211xp5_ASAP7_75t_L g959 ( .A1(n_197), .A2(n_902), .B(n_960), .C(n_968), .Y(n_959) );
INVx1_ASAP7_75t_L g1007 ( .A(n_197), .Y(n_1007) );
AOI221xp5_ASAP7_75t_L g972 ( .A1(n_198), .A2(n_249), .B1(n_500), .B2(n_532), .C(n_604), .Y(n_972) );
INVx1_ASAP7_75t_L g984 ( .A(n_198), .Y(n_984) );
INVx1_ASAP7_75t_L g978 ( .A(n_199), .Y(n_978) );
OAI332xp33_ASAP7_75t_SL g982 ( .A1(n_199), .A2(n_481), .A3(n_623), .B1(n_686), .B2(n_983), .B3(n_989), .C1(n_995), .C2(n_999), .Y(n_982) );
INVx1_ASAP7_75t_L g389 ( .A(n_200), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g1366 ( .A(n_201), .Y(n_1366) );
BUFx6f_ASAP7_75t_L g287 ( .A(n_202), .Y(n_287) );
AOI221xp5_ASAP7_75t_L g653 ( .A1(n_203), .A2(n_243), .B1(n_408), .B2(n_654), .C(n_656), .Y(n_653) );
INVx1_ASAP7_75t_L g630 ( .A(n_204), .Y(n_630) );
INVx1_ASAP7_75t_L g381 ( .A(n_205), .Y(n_381) );
XOR2x2_ASAP7_75t_L g807 ( .A(n_206), .B(n_808), .Y(n_807) );
AOI22xp33_ASAP7_75t_SL g825 ( .A1(n_207), .A2(n_250), .B1(n_403), .B2(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g842 ( .A(n_207), .Y(n_842) );
CKINVDCx5p33_ASAP7_75t_R g1112 ( .A(n_208), .Y(n_1112) );
CKINVDCx5p33_ASAP7_75t_R g490 ( .A(n_209), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_210), .A2(n_243), .B1(n_477), .B2(n_680), .Y(n_679) );
NOR2xp33_ASAP7_75t_R g780 ( .A(n_211), .B(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g1121 ( .A(n_212), .Y(n_1121) );
OAI22xp5_ASAP7_75t_L g1367 ( .A1(n_213), .A2(n_233), .B1(n_446), .B2(n_492), .Y(n_1367) );
INVx1_ASAP7_75t_L g715 ( .A(n_215), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_216), .A2(n_238), .B1(n_415), .B2(n_967), .Y(n_966) );
INVx1_ASAP7_75t_L g998 ( .A(n_216), .Y(n_998) );
INVx1_ASAP7_75t_L g466 ( .A(n_217), .Y(n_466) );
OAI221xp5_ASAP7_75t_SL g508 ( .A1(n_217), .A2(n_260), .B1(n_509), .B2(n_512), .C(n_517), .Y(n_508) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_218), .A2(n_263), .B1(n_492), .B2(n_544), .Y(n_637) );
INVx1_ASAP7_75t_L g1101 ( .A(n_220), .Y(n_1101) );
AOI22xp33_ASAP7_75t_SL g873 ( .A1(n_222), .A2(n_256), .B1(n_632), .B2(n_874), .Y(n_873) );
INVxp67_ASAP7_75t_SL g911 ( .A(n_222), .Y(n_911) );
INVx1_ASAP7_75t_L g636 ( .A(n_223), .Y(n_636) );
CKINVDCx5p33_ASAP7_75t_R g819 ( .A(n_224), .Y(n_819) );
INVx1_ASAP7_75t_L g975 ( .A(n_225), .Y(n_975) );
OAI211xp5_ASAP7_75t_L g1064 ( .A1(n_226), .A2(n_509), .B(n_1065), .C(n_1067), .Y(n_1064) );
INVx1_ASAP7_75t_L g1086 ( .A(n_226), .Y(n_1086) );
BUFx3_ASAP7_75t_L g291 ( .A(n_229), .Y(n_291) );
INVx1_ASAP7_75t_L g394 ( .A(n_229), .Y(n_394) );
XOR2x2_ASAP7_75t_L g1015 ( .A(n_232), .B(n_1016), .Y(n_1015) );
OAI211xp5_ASAP7_75t_L g1377 ( .A1(n_233), .A2(n_574), .B(n_1378), .C(n_1381), .Y(n_1377) );
INVxp67_ASAP7_75t_SL g1371 ( .A(n_234), .Y(n_1371) );
CKINVDCx5p33_ASAP7_75t_R g667 ( .A(n_235), .Y(n_667) );
INVx1_ASAP7_75t_L g986 ( .A(n_238), .Y(n_986) );
INVx1_ASAP7_75t_L g316 ( .A(n_241), .Y(n_316) );
INVx1_ASAP7_75t_L g330 ( .A(n_241), .Y(n_330) );
INVx2_ASAP7_75t_L g349 ( .A(n_241), .Y(n_349) );
XNOR2x1_ASAP7_75t_L g924 ( .A(n_242), .B(n_925), .Y(n_924) );
INVx1_ASAP7_75t_L g732 ( .A(n_244), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_244), .A2(n_266), .B1(n_607), .B2(n_658), .Y(n_790) );
NAND2xp5_ASAP7_75t_SL g824 ( .A(n_245), .B(n_411), .Y(n_824) );
INVx1_ASAP7_75t_L g460 ( .A(n_246), .Y(n_460) );
OAI21xp5_ASAP7_75t_L g445 ( .A1(n_248), .A2(n_446), .B(n_455), .Y(n_445) );
INVxp67_ASAP7_75t_SL g996 ( .A(n_249), .Y(n_996) );
INVxp67_ASAP7_75t_SL g849 ( .A(n_250), .Y(n_849) );
OAI22xp33_ASAP7_75t_SL g569 ( .A1(n_251), .A2(n_257), .B1(n_378), .B2(n_570), .Y(n_569) );
OAI221xp5_ASAP7_75t_L g584 ( .A1(n_251), .A2(n_257), .B1(n_509), .B2(n_513), .C(n_585), .Y(n_584) );
XNOR2xp5_ASAP7_75t_L g539 ( .A(n_253), .B(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g504 ( .A(n_254), .Y(n_504) );
INVx1_ASAP7_75t_L g915 ( .A(n_255), .Y(n_915) );
CKINVDCx5p33_ASAP7_75t_R g818 ( .A(n_258), .Y(n_818) );
INVx1_ASAP7_75t_L g468 ( .A(n_260), .Y(n_468) );
OAI211xp5_ASAP7_75t_L g600 ( .A1(n_263), .A2(n_574), .B(n_601), .C(n_608), .Y(n_600) );
INVx1_ASAP7_75t_L g829 ( .A(n_264), .Y(n_829) );
INVx1_ASAP7_75t_L g744 ( .A(n_266), .Y(n_744) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_292), .B(n_1133), .Y(n_267) );
BUFx4f_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx3_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g270 ( .A(n_271), .B(n_277), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g1387 ( .A(n_271), .B(n_280), .Y(n_1387) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
NOR2xp33_ASAP7_75t_L g1391 ( .A(n_273), .B(n_276), .Y(n_1391) );
INVx1_ASAP7_75t_L g1397 ( .A(n_273), .Y(n_1397) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g1399 ( .A(n_276), .B(n_1397), .Y(n_1399) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_282), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x4_ASAP7_75t_L g413 ( .A(n_281), .B(n_291), .Y(n_413) );
AND2x4_ASAP7_75t_L g435 ( .A(n_281), .B(n_290), .Y(n_435) );
AND2x4_ASAP7_75t_SL g1386 ( .A(n_282), .B(n_1387), .Y(n_1386) );
INVx3_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OR2x6_ASAP7_75t_L g283 ( .A(n_284), .B(n_289), .Y(n_283) );
INVxp67_ASAP7_75t_L g1129 ( .A(n_284), .Y(n_1129) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
BUFx4f_ASAP7_75t_L g520 ( .A(n_285), .Y(n_520) );
INVx3_ASAP7_75t_L g1051 ( .A(n_285), .Y(n_1051) );
INVx3_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
INVx2_ASAP7_75t_L g334 ( .A(n_287), .Y(n_334) );
AND2x2_ASAP7_75t_L g399 ( .A(n_287), .B(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g405 ( .A(n_287), .Y(n_405) );
AND2x2_ASAP7_75t_L g409 ( .A(n_287), .B(n_288), .Y(n_409) );
INVx1_ASAP7_75t_L g450 ( .A(n_287), .Y(n_450) );
NAND2x1_ASAP7_75t_L g589 ( .A(n_287), .B(n_288), .Y(n_589) );
INVx1_ASAP7_75t_L g335 ( .A(n_288), .Y(n_335) );
INVx2_ASAP7_75t_L g400 ( .A(n_288), .Y(n_400) );
AND2x2_ASAP7_75t_L g404 ( .A(n_288), .B(n_405), .Y(n_404) );
BUFx2_ASAP7_75t_L g440 ( .A(n_288), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_288), .B(n_405), .Y(n_525) );
OR2x2_ASAP7_75t_L g789 ( .A(n_288), .B(n_334), .Y(n_789) );
INVxp67_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OAI22xp33_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_919), .B1(n_1131), .B2(n_1132), .Y(n_292) );
INVx1_ASAP7_75t_L g1131 ( .A(n_293), .Y(n_1131) );
AO22x2_ASAP7_75t_L g293 ( .A1(n_294), .A2(n_640), .B1(n_641), .B2(n_918), .Y(n_293) );
INVx1_ASAP7_75t_L g918 ( .A(n_294), .Y(n_918) );
XNOR2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_537), .Y(n_294) );
XOR2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_461), .Y(n_295) );
XNOR2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_460), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_386), .Y(n_297) );
AOI221xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_317), .B1(n_318), .B2(n_336), .C(n_337), .Y(n_298) );
AOI221xp5_ASAP7_75t_L g926 ( .A1(n_299), .A2(n_318), .B1(n_927), .B2(n_928), .C(n_929), .Y(n_926) );
INVx3_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx5_ASAP7_75t_L g858 ( .A(n_300), .Y(n_858) );
OR2x6_ASAP7_75t_L g300 ( .A(n_301), .B(n_313), .Y(n_300) );
OR2x2_ASAP7_75t_L g492 ( .A(n_301), .B(n_313), .Y(n_492) );
NAND2x1p5_ASAP7_75t_L g301 ( .A(n_302), .B(n_308), .Y(n_301) );
INVx8_ASAP7_75t_L g352 ( .A(n_302), .Y(n_352) );
BUFx3_ASAP7_75t_L g750 ( .A(n_302), .Y(n_750) );
BUFx3_ASAP7_75t_L g844 ( .A(n_302), .Y(n_844) );
HB1xp67_ASAP7_75t_L g851 ( .A(n_302), .Y(n_851) );
AND2x4_ASAP7_75t_L g302 ( .A(n_303), .B(n_305), .Y(n_302) );
AND2x4_ASAP7_75t_L g358 ( .A(n_303), .B(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_304), .B(n_324), .Y(n_323) );
AND2x4_ASAP7_75t_L g341 ( .A(n_304), .B(n_342), .Y(n_341) );
BUFx6f_ASAP7_75t_L g363 ( .A(n_304), .Y(n_363) );
OR2x2_ASAP7_75t_L g484 ( .A(n_304), .B(n_306), .Y(n_484) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVxp67_ASAP7_75t_L g359 ( .A(n_307), .Y(n_359) );
AND2x4_ASAP7_75t_L g343 ( .A(n_308), .B(n_329), .Y(n_343) );
INVx1_ASAP7_75t_L g752 ( .A(n_308), .Y(n_752) );
AND2x6_ASAP7_75t_L g759 ( .A(n_308), .B(n_379), .Y(n_759) );
AND2x2_ASAP7_75t_L g761 ( .A(n_308), .B(n_385), .Y(n_761) );
AND2x4_ASAP7_75t_L g308 ( .A(n_309), .B(n_311), .Y(n_308) );
NAND3x1_ASAP7_75t_L g370 ( .A(n_309), .B(n_371), .C(n_372), .Y(n_370) );
NAND2x1p5_ASAP7_75t_L g687 ( .A(n_309), .B(n_372), .Y(n_687) );
INVx3_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
BUFx3_ASAP7_75t_L g347 ( .A(n_310), .Y(n_347) );
NAND2xp33_ASAP7_75t_SL g550 ( .A(n_310), .B(n_312), .Y(n_550) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND3x4_ASAP7_75t_L g346 ( .A(n_312), .B(n_347), .C(n_348), .Y(n_346) );
AND2x2_ASAP7_75t_L g739 ( .A(n_312), .B(n_347), .Y(n_739) );
INVxp67_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OR2x2_ASAP7_75t_L g447 ( .A(n_314), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g698 ( .A(n_314), .Y(n_698) );
OR2x2_ASAP7_75t_L g772 ( .A(n_314), .B(n_448), .Y(n_772) );
BUFx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx2_ASAP7_75t_L g326 ( .A(n_315), .Y(n_326) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AOI221xp5_ASAP7_75t_L g401 ( .A1(n_317), .A2(n_402), .B1(n_406), .B2(n_414), .C(n_419), .Y(n_401) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_318), .A2(n_490), .B(n_491), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_318), .A2(n_542), .B(n_543), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g635 ( .A1(n_318), .A2(n_636), .B(n_637), .Y(n_635) );
AOI211x1_ASAP7_75t_L g861 ( .A1(n_318), .A2(n_862), .B(n_863), .C(n_885), .Y(n_861) );
AOI21xp5_ASAP7_75t_L g1017 ( .A1(n_318), .A2(n_1018), .B(n_1019), .Y(n_1017) );
AOI21xp33_ASAP7_75t_L g1080 ( .A1(n_318), .A2(n_1081), .B(n_1082), .Y(n_1080) );
AOI21xp5_ASAP7_75t_L g1111 ( .A1(n_318), .A2(n_1112), .B(n_1113), .Y(n_1111) );
AOI21xp33_ASAP7_75t_SL g1365 ( .A1(n_318), .A2(n_1366), .B(n_1367), .Y(n_1365) );
INVx8_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x4_ASAP7_75t_L g319 ( .A(n_320), .B(n_328), .Y(n_319) );
INVx1_ASAP7_75t_L g705 ( .A(n_320), .Y(n_705) );
OR2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_325), .Y(n_320) );
BUFx3_ASAP7_75t_L g848 ( .A(n_321), .Y(n_848) );
INVx1_ASAP7_75t_L g988 ( .A(n_321), .Y(n_988) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
BUFx6f_ASAP7_75t_L g566 ( .A(n_322), .Y(n_566) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
BUFx2_ASAP7_75t_L g556 ( .A(n_323), .Y(n_556) );
INVx2_ASAP7_75t_L g342 ( .A(n_324), .Y(n_342) );
INVx1_ASAP7_75t_L g454 ( .A(n_324), .Y(n_454) );
OR2x2_ASAP7_75t_L g451 ( .A(n_325), .B(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g458 ( .A(n_325), .Y(n_458) );
INVx1_ASAP7_75t_L g486 ( .A(n_325), .Y(n_486) );
OR2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
OR2x2_ASAP7_75t_L g549 ( .A(n_326), .B(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_SL g785 ( .A(n_326), .B(n_413), .Y(n_785) );
INVx1_ASAP7_75t_L g726 ( .A(n_327), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_328), .B(n_803), .Y(n_802) );
OR2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_331), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g371 ( .A(n_330), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_330), .B(n_393), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
AND2x6_ASAP7_75t_L g419 ( .A(n_332), .B(n_408), .Y(n_419) );
AND2x2_ASAP7_75t_L g438 ( .A(n_332), .B(n_439), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_332), .B(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g516 ( .A(n_332), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_332), .B(n_349), .Y(n_777) );
AND2x2_ASAP7_75t_L g392 ( .A(n_333), .B(n_393), .Y(n_392) );
INVx3_ASAP7_75t_L g416 ( .A(n_333), .Y(n_416) );
BUFx6f_ASAP7_75t_L g580 ( .A(n_333), .Y(n_580) );
AND2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_334), .Y(n_669) );
NAND3xp33_ASAP7_75t_SL g337 ( .A(n_338), .B(n_344), .C(n_375), .Y(n_337) );
INVx2_ASAP7_75t_SL g488 ( .A(n_338), .Y(n_488) );
AND5x1_ASAP7_75t_L g808 ( .A(n_338), .B(n_809), .C(n_836), .D(n_852), .E(n_856), .Y(n_808) );
NAND3xp33_ASAP7_75t_SL g929 ( .A(n_338), .B(n_930), .C(n_933), .Y(n_929) );
NAND4xp75_ASAP7_75t_L g1016 ( .A(n_338), .B(n_1017), .C(n_1020), .D(n_1038), .Y(n_1016) );
INVx3_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_339), .Y(n_546) );
NOR3xp33_ASAP7_75t_L g621 ( .A(n_339), .B(n_622), .C(n_634), .Y(n_621) );
AOI221xp5_ASAP7_75t_L g688 ( .A1(n_339), .A2(n_571), .B1(n_667), .B2(n_689), .C(n_690), .Y(n_688) );
INVx3_ASAP7_75t_L g871 ( .A(n_339), .Y(n_871) );
AND2x4_ASAP7_75t_L g339 ( .A(n_340), .B(n_343), .Y(n_339) );
BUFx2_ASAP7_75t_L g471 ( .A(n_340), .Y(n_471) );
BUFx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
BUFx2_ASAP7_75t_L g353 ( .A(n_341), .Y(n_353) );
BUFx3_ASAP7_75t_L g374 ( .A(n_341), .Y(n_374) );
BUFx2_ASAP7_75t_L g559 ( .A(n_341), .Y(n_559) );
INVx2_ASAP7_75t_L g633 ( .A(n_341), .Y(n_633) );
INVx1_ASAP7_75t_L g364 ( .A(n_342), .Y(n_364) );
NAND2x1_ASAP7_75t_L g378 ( .A(n_343), .B(n_379), .Y(n_378) );
AND2x4_ASAP7_75t_L g382 ( .A(n_343), .B(n_383), .Y(n_382) );
AND2x2_ASAP7_75t_L g467 ( .A(n_343), .B(n_379), .Y(n_467) );
AND2x4_ASAP7_75t_SL g571 ( .A(n_343), .B(n_383), .Y(n_571) );
AND2x4_ASAP7_75t_SL g689 ( .A(n_343), .B(n_379), .Y(n_689) );
AOI33xp33_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_350), .A3(n_354), .B1(n_365), .B2(n_367), .B3(n_373), .Y(n_344) );
AOI33xp33_ASAP7_75t_L g469 ( .A1(n_345), .A2(n_367), .A3(n_470), .B1(n_472), .B2(n_478), .B3(n_479), .Y(n_469) );
AOI33xp33_ASAP7_75t_L g872 ( .A1(n_345), .A2(n_873), .A3(n_876), .B1(n_878), .B2(n_879), .B3(n_881), .Y(n_872) );
AOI33xp33_ASAP7_75t_L g1027 ( .A1(n_345), .A2(n_1028), .A3(n_1029), .B1(n_1032), .B2(n_1035), .B3(n_1036), .Y(n_1027) );
AOI33xp33_ASAP7_75t_L g1103 ( .A1(n_345), .A2(n_1104), .A3(n_1105), .B1(n_1106), .B2(n_1108), .B3(n_1109), .Y(n_1103) );
BUFx3_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AOI33xp33_ASAP7_75t_L g677 ( .A1(n_346), .A2(n_678), .A3(n_679), .B1(n_681), .B2(n_683), .B3(n_685), .Y(n_677) );
INVx1_ASAP7_75t_L g939 ( .A(n_346), .Y(n_939) );
AOI33xp33_ASAP7_75t_L g1087 ( .A1(n_346), .A2(n_1088), .A3(n_1089), .B1(n_1090), .B2(n_1091), .B3(n_1092), .Y(n_1087) );
AOI33xp33_ASAP7_75t_L g1357 ( .A1(n_346), .A2(n_1035), .A3(n_1358), .B1(n_1361), .B2(n_1362), .B3(n_1363), .Y(n_1357) );
INVx1_ASAP7_75t_L g536 ( .A(n_348), .Y(n_536) );
OAI31xp33_ASAP7_75t_L g722 ( .A1(n_348), .A2(n_723), .A3(n_727), .B(n_753), .Y(n_722) );
INVx2_ASAP7_75t_SL g1384 ( .A(n_348), .Y(n_1384) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
BUFx2_ASAP7_75t_L g444 ( .A(n_349), .Y(n_444) );
INVx8_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g457 ( .A(n_352), .Y(n_457) );
INVx3_ASAP7_75t_L g882 ( .A(n_352), .Y(n_882) );
INVx2_ASAP7_75t_L g935 ( .A(n_352), .Y(n_935) );
INVx1_ASAP7_75t_L g884 ( .A(n_353), .Y(n_884) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx2_ASAP7_75t_SL g356 ( .A(n_357), .Y(n_356) );
AND2x4_ASAP7_75t_L g459 ( .A(n_357), .B(n_458), .Y(n_459) );
INVx2_ASAP7_75t_SL g625 ( .A(n_357), .Y(n_625) );
INVx3_ASAP7_75t_L g985 ( .A(n_357), .Y(n_985) );
HB1xp67_ASAP7_75t_L g1030 ( .A(n_357), .Y(n_1030) );
BUFx8_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g475 ( .A(n_358), .Y(n_475) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_358), .Y(n_563) );
BUFx6f_ASAP7_75t_L g737 ( .A(n_358), .Y(n_737) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g877 ( .A(n_361), .Y(n_877) );
INVx5_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx3_ASAP7_75t_L g366 ( .A(n_362), .Y(n_366) );
BUFx12f_ASAP7_75t_L g477 ( .A(n_362), .Y(n_477) );
AND2x4_ASAP7_75t_L g804 ( .A(n_362), .B(n_726), .Y(n_804) );
BUFx3_ASAP7_75t_L g1031 ( .A(n_362), .Y(n_1031) );
AND2x4_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
INVx2_ASAP7_75t_L g380 ( .A(n_363), .Y(n_380) );
NAND2x1p5_ASAP7_75t_L g453 ( .A(n_363), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g385 ( .A(n_364), .Y(n_385) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
OAI22xp5_ASAP7_75t_SL g622 ( .A1(n_368), .A2(n_623), .B1(n_624), .B2(n_629), .Y(n_622) );
CKINVDCx5p33_ASAP7_75t_R g368 ( .A(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g560 ( .A(n_369), .Y(n_560) );
INVx2_ASAP7_75t_L g845 ( .A(n_369), .Y(n_845) );
INVx3_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx3_ASAP7_75t_L g880 ( .A(n_370), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_377), .B1(n_381), .B2(n_382), .Y(n_375) );
AOI222xp33_ASAP7_75t_L g420 ( .A1(n_376), .A2(n_381), .B1(n_421), .B2(n_423), .C1(n_425), .C2(n_436), .Y(n_420) );
AOI221x1_ASAP7_75t_L g836 ( .A1(n_377), .A2(n_382), .B1(n_812), .B2(n_818), .C(n_837), .Y(n_836) );
AOI22xp33_ASAP7_75t_L g1006 ( .A1(n_377), .A2(n_382), .B1(n_973), .B2(n_1007), .Y(n_1006) );
AOI22xp33_ASAP7_75t_L g1021 ( .A1(n_377), .A2(n_382), .B1(n_1022), .B2(n_1023), .Y(n_1021) );
AOI22xp33_ASAP7_75t_L g1354 ( .A1(n_377), .A2(n_382), .B1(n_1355), .B2(n_1356), .Y(n_1354) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx3_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_382), .A2(n_466), .B1(n_467), .B2(n_468), .Y(n_465) );
AO22x1_ASAP7_75t_L g865 ( .A1(n_382), .A2(n_467), .B1(n_866), .B2(n_867), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g1100 ( .A1(n_382), .A2(n_467), .B1(n_1101), .B2(n_1102), .Y(n_1100) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AOI21xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_441), .B(n_445), .Y(n_386) );
NAND3xp33_ASAP7_75t_L g387 ( .A(n_388), .B(n_401), .C(n_420), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_390), .B1(n_395), .B2(n_396), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_389), .A2(n_395), .B1(n_456), .B2(n_459), .Y(n_455) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_390), .A2(n_504), .B1(n_505), .B2(n_506), .Y(n_503) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_391), .A2(n_397), .B1(n_582), .B2(n_583), .Y(n_581) );
AOI22xp5_ASAP7_75t_L g943 ( .A1(n_391), .A2(n_397), .B1(n_944), .B2(n_945), .Y(n_943) );
NAND2xp5_ASAP7_75t_L g977 ( .A(n_391), .B(n_978), .Y(n_977) );
AOI22xp33_ASAP7_75t_L g1046 ( .A1(n_391), .A2(n_397), .B1(n_1025), .B2(n_1026), .Y(n_1046) );
AOI22xp33_ASAP7_75t_L g1077 ( .A1(n_391), .A2(n_396), .B1(n_1078), .B2(n_1079), .Y(n_1077) );
BUFx6f_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_392), .A2(n_397), .B1(n_609), .B2(n_610), .Y(n_608) );
AND2x4_ASAP7_75t_L g720 ( .A(n_392), .B(n_698), .Y(n_720) );
INVx1_ASAP7_75t_L g893 ( .A(n_392), .Y(n_893) );
AND2x4_ASAP7_75t_L g397 ( .A(n_393), .B(n_398), .Y(n_397) );
AND2x4_ASAP7_75t_L g402 ( .A(n_393), .B(n_403), .Y(n_402) );
AND2x4_ASAP7_75t_SL g422 ( .A(n_393), .B(n_408), .Y(n_422) );
AND2x2_ASAP7_75t_L g649 ( .A(n_393), .B(n_650), .Y(n_649) );
BUFx2_ASAP7_75t_L g672 ( .A(n_393), .Y(n_672) );
AND2x2_ASAP7_75t_L g699 ( .A(n_393), .B(n_398), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g1381 ( .A1(n_396), .A2(n_892), .B1(n_1382), .B2(n_1383), .Y(n_1381) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g507 ( .A(n_397), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_397), .A2(n_887), .B1(n_888), .B2(n_892), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g974 ( .A1(n_397), .A2(n_649), .B1(n_975), .B2(n_976), .Y(n_974) );
INVx2_ASAP7_75t_L g433 ( .A(n_398), .Y(n_433) );
BUFx6f_ASAP7_75t_L g531 ( .A(n_398), .Y(n_531) );
INVx1_ASAP7_75t_L g605 ( .A(n_398), .Y(n_605) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
BUFx3_ASAP7_75t_L g411 ( .A(n_399), .Y(n_411) );
INVx2_ASAP7_75t_L g655 ( .A(n_399), .Y(n_655) );
INVx3_ASAP7_75t_L g495 ( .A(n_402), .Y(n_495) );
INVx2_ASAP7_75t_SL g574 ( .A(n_402), .Y(n_574) );
NAND2xp5_ASAP7_75t_R g900 ( .A(n_402), .B(n_870), .Y(n_900) );
BUFx2_ASAP7_75t_L g967 ( .A(n_403), .Y(n_967) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
BUFx3_ASAP7_75t_L g418 ( .A(n_404), .Y(n_418) );
INVx2_ASAP7_75t_L g594 ( .A(n_404), .Y(n_594) );
BUFx3_ASAP7_75t_L g607 ( .A(n_404), .Y(n_607) );
BUFx3_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_408), .Y(n_500) );
BUFx3_ASAP7_75t_L g603 ( .A(n_408), .Y(n_603) );
INVx1_ASAP7_75t_L g965 ( .A(n_408), .Y(n_965) );
BUFx3_ASAP7_75t_L g1374 ( .A(n_408), .Y(n_1374) );
BUFx6f_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g429 ( .A(n_409), .Y(n_429) );
BUFx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g963 ( .A(n_411), .Y(n_963) );
INVx4_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_SL g501 ( .A(n_413), .Y(n_501) );
INVx4_ASAP7_75t_L g661 ( .A(n_413), .Y(n_661) );
NAND4xp25_ASAP7_75t_L g823 ( .A(n_413), .B(n_824), .C(n_825), .D(n_827), .Y(n_823) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_SL g424 ( .A(n_416), .Y(n_424) );
INVx2_ASAP7_75t_L g658 ( .A(n_416), .Y(n_658) );
INVx1_ASAP7_75t_L g826 ( .A(n_416), .Y(n_826) );
INVx2_ASAP7_75t_L g897 ( .A(n_416), .Y(n_897) );
INVx1_ASAP7_75t_L g1071 ( .A(n_416), .Y(n_1071) );
BUFx3_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_SL g899 ( .A(n_418), .Y(n_899) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_419), .A2(n_497), .B(n_502), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g575 ( .A1(n_419), .A2(n_576), .B(n_577), .Y(n_575) );
AOI21xp5_ASAP7_75t_L g601 ( .A1(n_419), .A2(n_602), .B(n_606), .Y(n_601) );
AOI21xp5_ASAP7_75t_L g894 ( .A1(n_419), .A2(n_895), .B(n_896), .Y(n_894) );
AOI221xp5_ASAP7_75t_L g946 ( .A1(n_419), .A2(n_649), .B1(n_927), .B2(n_947), .C(n_948), .Y(n_946) );
INVx1_ASAP7_75t_L g968 ( .A(n_419), .Y(n_968) );
AOI21xp5_ASAP7_75t_SL g1040 ( .A1(n_419), .A2(n_1041), .B(n_1045), .Y(n_1040) );
AOI21xp5_ASAP7_75t_L g1073 ( .A1(n_419), .A2(n_1074), .B(n_1075), .Y(n_1073) );
AOI21xp5_ASAP7_75t_L g1116 ( .A1(n_419), .A2(n_1117), .B(n_1119), .Y(n_1116) );
AOI21xp5_ASAP7_75t_L g1378 ( .A1(n_419), .A2(n_1379), .B(n_1380), .Y(n_1378) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_421), .B(n_812), .Y(n_811) );
AOI222xp33_ASAP7_75t_L g949 ( .A1(n_421), .A2(n_438), .B1(n_931), .B2(n_932), .C1(n_950), .C2(n_951), .Y(n_949) );
BUFx3_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g511 ( .A(n_422), .Y(n_511) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
BUFx2_ASAP7_75t_L g529 ( .A(n_429), .Y(n_529) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g1376 ( .A(n_433), .Y(n_1376) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g532 ( .A(n_435), .Y(n_532) );
INVx2_ASAP7_75t_L g591 ( .A(n_435), .Y(n_591) );
INVx3_ASAP7_75t_L g656 ( .A(n_435), .Y(n_656) );
OAI221xp5_ASAP7_75t_L g903 ( .A1(n_435), .A2(n_904), .B1(n_905), .B2(n_906), .C(n_909), .Y(n_903) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g970 ( .A1(n_438), .A2(n_971), .B1(n_972), .B2(n_973), .Y(n_970) );
NAND2xp5_ASAP7_75t_L g1065 ( .A(n_438), .B(n_1066), .Y(n_1065) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_439), .A2(n_667), .B1(n_668), .B2(n_670), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_439), .A2(n_668), .B1(n_818), .B2(n_819), .Y(n_817) );
BUFx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g515 ( .A(n_440), .Y(n_515) );
INVx1_ASAP7_75t_L g779 ( .A(n_440), .Y(n_779) );
OAI21xp5_ASAP7_75t_L g572 ( .A1(n_441), .A2(n_573), .B(n_584), .Y(n_572) );
OAI21xp5_ASAP7_75t_L g889 ( .A1(n_441), .A2(n_890), .B(n_901), .Y(n_889) );
AOI21xp5_ASAP7_75t_L g941 ( .A1(n_441), .A2(n_942), .B(n_952), .Y(n_941) );
OAI21xp5_ASAP7_75t_L g958 ( .A1(n_441), .A2(n_959), .B(n_969), .Y(n_958) );
OAI21xp5_ASAP7_75t_SL g1063 ( .A1(n_441), .A2(n_1064), .B(n_1072), .Y(n_1063) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
BUFx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_443), .B(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
OR2x6_ASAP7_75t_L g686 ( .A(n_444), .B(n_687), .Y(n_686) );
AND2x4_ASAP7_75t_L g766 ( .A(n_444), .B(n_767), .Y(n_766) );
OR2x2_ASAP7_75t_L g936 ( .A(n_444), .B(n_687), .Y(n_936) );
INVx2_ASAP7_75t_L g980 ( .A(n_446), .Y(n_980) );
AND2x4_ASAP7_75t_L g446 ( .A(n_447), .B(n_451), .Y(n_446) );
AND2x4_ASAP7_75t_L g544 ( .A(n_447), .B(n_451), .Y(n_544) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g702 ( .A(n_451), .Y(n_702) );
INVx3_ASAP7_75t_L g747 ( .A(n_452), .Y(n_747) );
INVx4_ASAP7_75t_L g994 ( .A(n_452), .Y(n_994) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx2_ASAP7_75t_L g734 ( .A(n_453), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_456), .A2(n_459), .B1(n_582), .B2(n_583), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g638 ( .A1(n_456), .A2(n_459), .B1(n_609), .B2(n_610), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g886 ( .A1(n_456), .A2(n_459), .B1(n_887), .B2(n_888), .Y(n_886) );
AND2x4_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
AND2x4_ASAP7_75t_L g703 ( .A(n_457), .B(n_458), .Y(n_703) );
AOI22xp5_ASAP7_75t_L g754 ( .A1(n_457), .A2(n_684), .B1(n_719), .B2(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g487 ( .A(n_459), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g1009 ( .A(n_459), .B(n_975), .Y(n_1009) );
AOI22xp33_ASAP7_75t_L g1024 ( .A1(n_459), .A2(n_703), .B1(n_1025), .B2(n_1026), .Y(n_1024) );
NAND3xp33_ASAP7_75t_L g462 ( .A(n_463), .B(n_489), .C(n_493), .Y(n_462) );
NOR3xp33_ASAP7_75t_L g463 ( .A(n_464), .B(n_480), .C(n_488), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_465), .B(n_469), .Y(n_464) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
BUFx2_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
OAI221xp5_ASAP7_75t_L g551 ( .A1(n_475), .A2(n_552), .B1(n_553), .B2(n_557), .C(n_558), .Y(n_551) );
INVx3_ASAP7_75t_L g695 ( .A(n_475), .Y(n_695) );
OR2x6_ASAP7_75t_SL g724 ( .A(n_475), .B(n_725), .Y(n_724) );
BUFx2_ASAP7_75t_L g1034 ( .A(n_475), .Y(n_1034) );
BUFx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g854 ( .A(n_481), .B(n_855), .Y(n_854) );
OR2x6_ASAP7_75t_L g481 ( .A(n_482), .B(n_485), .Y(n_481) );
OR2x2_ASAP7_75t_L g1094 ( .A(n_482), .B(n_485), .Y(n_1094) );
INVx2_ASAP7_75t_SL g482 ( .A(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
BUFx4f_ASAP7_75t_L g729 ( .A(n_484), .Y(n_729) );
BUFx3_ASAP7_75t_L g990 ( .A(n_484), .Y(n_990) );
BUFx3_ASAP7_75t_L g1001 ( .A(n_484), .Y(n_1001) );
INVxp67_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g694 ( .A(n_486), .B(n_695), .Y(n_694) );
NOR3xp33_ASAP7_75t_L g1352 ( .A(n_488), .B(n_1353), .C(n_1364), .Y(n_1352) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_492), .B(n_797), .Y(n_796) );
OAI21xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_508), .B(n_533), .Y(n_493) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
BUFx2_ASAP7_75t_L g1118 ( .A(n_500), .Y(n_1118) );
AOI22xp33_ASAP7_75t_L g1120 ( .A1(n_506), .A2(n_892), .B1(n_1121), .B2(n_1122), .Y(n_1120) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx2_ASAP7_75t_L g612 ( .A(n_510), .Y(n_612) );
INVx1_ASAP7_75t_L g902 ( .A(n_510), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g1130 ( .A1(n_510), .A2(n_514), .B1(n_1101), .B2(n_1102), .Y(n_1130) );
INVx4_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
BUFx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g1048 ( .A(n_514), .Y(n_1048) );
NOR2x1_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .Y(n_514) );
INVx1_ASAP7_75t_L g671 ( .A(n_516), .Y(n_671) );
OAI221xp5_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_521), .B1(n_522), .B2(n_526), .C(n_527), .Y(n_517) );
OAI22xp5_ASAP7_75t_L g910 ( .A1(n_518), .A2(n_911), .B1(n_912), .B2(n_913), .Y(n_910) );
OAI221xp5_ASAP7_75t_L g1370 ( .A1(n_518), .A2(n_913), .B1(n_1371), .B2(n_1372), .C(n_1373), .Y(n_1370) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx3_ASAP7_75t_L g664 ( .A(n_520), .Y(n_664) );
INVx4_ASAP7_75t_L g815 ( .A(n_520), .Y(n_815) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx4_ASAP7_75t_L g822 ( .A(n_523), .Y(n_822) );
BUFx6f_ASAP7_75t_L g914 ( .A(n_523), .Y(n_914) );
INVx2_ASAP7_75t_L g1054 ( .A(n_523), .Y(n_1054) );
INVx8_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g1126 ( .A(n_529), .Y(n_1126) );
BUFx3_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
OAI21xp5_ASAP7_75t_L g1114 ( .A1(n_533), .A2(n_1115), .B(n_1123), .Y(n_1114) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
HB1xp67_ASAP7_75t_L g832 ( .A(n_535), .Y(n_832) );
BUFx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
BUFx2_ASAP7_75t_L g620 ( .A(n_536), .Y(n_620) );
AOI21x1_ASAP7_75t_L g646 ( .A1(n_536), .A2(n_647), .B(n_675), .Y(n_646) );
HB1xp67_ASAP7_75t_L g1058 ( .A(n_536), .Y(n_1058) );
BUFx3_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
AO22x2_ASAP7_75t_L g538 ( .A1(n_539), .A2(n_596), .B1(n_597), .B2(n_639), .Y(n_538) );
INVx1_ASAP7_75t_L g639 ( .A(n_539), .Y(n_639) );
AND4x1_ASAP7_75t_L g540 ( .A(n_541), .B(n_545), .C(n_572), .D(n_595), .Y(n_540) );
NOR3xp33_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .C(n_569), .Y(n_545) );
NOR3xp33_ASAP7_75t_L g1083 ( .A(n_546), .B(n_1084), .C(n_1093), .Y(n_1083) );
NOR3xp33_ASAP7_75t_L g1098 ( .A(n_546), .B(n_1099), .C(n_1110), .Y(n_1098) );
OAI22xp5_ASAP7_75t_SL g547 ( .A1(n_548), .A2(n_551), .B1(n_560), .B2(n_561), .Y(n_547) );
BUFx4f_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
BUFx8_ASAP7_75t_L g623 ( .A(n_549), .Y(n_623) );
BUFx2_ASAP7_75t_L g838 ( .A(n_549), .Y(n_838) );
OAI221xp5_ASAP7_75t_L g624 ( .A1(n_553), .A2(n_625), .B1(n_626), .B2(n_627), .C(n_628), .Y(n_624) );
INVx3_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
BUFx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
OAI221xp5_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_564), .B1(n_565), .B2(n_567), .C(n_568), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
BUFx6f_ASAP7_75t_L g680 ( .A(n_563), .Y(n_680) );
BUFx6f_ASAP7_75t_L g682 ( .A(n_563), .Y(n_682) );
OAI211xp5_ASAP7_75t_L g585 ( .A1(n_564), .A2(n_586), .B(n_590), .C(n_592), .Y(n_585) );
OAI221xp5_ASAP7_75t_L g629 ( .A1(n_565), .A2(n_614), .B1(n_625), .B2(n_630), .C(n_631), .Y(n_629) );
CKINVDCx8_ASAP7_75t_R g565 ( .A(n_566), .Y(n_565) );
INVx3_ASAP7_75t_L g731 ( .A(n_566), .Y(n_731) );
INVx3_ASAP7_75t_L g743 ( .A(n_566), .Y(n_743) );
INVx3_ASAP7_75t_L g841 ( .A(n_566), .Y(n_841) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AOI22xp5_ASAP7_75t_L g930 ( .A1(n_571), .A2(n_689), .B1(n_931), .B2(n_932), .Y(n_930) );
AOI22xp33_ASAP7_75t_L g1085 ( .A1(n_571), .A2(n_689), .B1(n_1066), .B2(n_1086), .Y(n_1085) );
INVx2_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g1076 ( .A(n_579), .Y(n_1076) );
INVx3_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx2_ASAP7_75t_L g665 ( .A(n_587), .Y(n_665) );
INVx2_ASAP7_75t_L g816 ( .A(n_587), .Y(n_816) );
INVx4_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
BUFx4f_ASAP7_75t_L g674 ( .A(n_588), .Y(n_674) );
OR2x6_ASAP7_75t_L g792 ( .A(n_588), .B(n_793), .Y(n_792) );
BUFx4f_ASAP7_75t_L g904 ( .A(n_588), .Y(n_904) );
BUFx6f_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
BUFx3_ASAP7_75t_L g617 ( .A(n_589), .Y(n_617) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx3_ASAP7_75t_L g650 ( .A(n_594), .Y(n_650) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND4x1_ASAP7_75t_L g598 ( .A(n_599), .B(n_621), .C(n_635), .D(n_638), .Y(n_598) );
OAI21xp5_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_611), .B(n_620), .Y(n_599) );
INVx2_ASAP7_75t_SL g604 ( .A(n_605), .Y(n_604) );
OAI211xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_615), .B(n_618), .C(n_619), .Y(n_613) );
OAI211xp5_ASAP7_75t_L g828 ( .A1(n_615), .A2(n_829), .B(n_830), .C(n_831), .Y(n_828) );
INVx5_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx2_ASAP7_75t_SL g616 ( .A(n_617), .Y(n_616) );
OR2x2_ASAP7_75t_L g781 ( .A(n_617), .B(n_782), .Y(n_781) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g684 ( .A(n_633), .Y(n_684) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AO22x2_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_859), .B1(n_916), .B2(n_917), .Y(n_641) );
INVx1_ASAP7_75t_L g916 ( .A(n_642), .Y(n_916) );
XNOR2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_807), .Y(n_642) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_714), .B1(n_805), .B2(n_806), .Y(n_643) );
INVx1_ASAP7_75t_L g806 ( .A(n_644), .Y(n_806) );
NAND3xp33_ASAP7_75t_L g644 ( .A(n_645), .B(n_707), .C(n_711), .Y(n_644) );
INVx1_ASAP7_75t_L g708 ( .A(n_646), .Y(n_708) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AND2x4_ASAP7_75t_L g798 ( .A(n_650), .B(n_799), .Y(n_798) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_653), .B1(n_657), .B2(n_659), .Y(n_651) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx2_ASAP7_75t_L g660 ( .A(n_655), .Y(n_660) );
INVx2_ASAP7_75t_L g1044 ( .A(n_660), .Y(n_1044) );
HB1xp67_ASAP7_75t_L g1127 ( .A(n_660), .Y(n_1127) );
AOI22xp5_ASAP7_75t_L g662 ( .A1(n_663), .A2(n_671), .B1(n_672), .B2(n_673), .Y(n_662) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
AOI222xp33_ASAP7_75t_L g701 ( .A1(n_670), .A2(n_702), .B1(n_703), .B2(n_704), .C1(n_705), .C2(n_706), .Y(n_701) );
AOI22xp5_ASAP7_75t_L g813 ( .A1(n_671), .A2(n_672), .B1(n_814), .B2(n_820), .Y(n_813) );
OAI211xp5_ASAP7_75t_L g1067 ( .A1(n_674), .A2(n_1068), .B(n_1069), .C(n_1070), .Y(n_1067) );
INVx1_ASAP7_75t_L g709 ( .A(n_676), .Y(n_709) );
AND2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_688), .Y(n_676) );
INVx2_ASAP7_75t_L g997 ( .A(n_680), .Y(n_997) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_SL g1091 ( .A(n_686), .Y(n_1091) );
INVx1_ASAP7_75t_L g713 ( .A(n_691), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_692), .B(n_700), .Y(n_691) );
NAND2x1_ASAP7_75t_L g692 ( .A(n_693), .B(n_696), .Y(n_692) );
INVx2_ASAP7_75t_SL g693 ( .A(n_694), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g953 ( .A1(n_694), .A2(n_703), .B1(n_944), .B2(n_945), .Y(n_953) );
INVx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g718 ( .A1(n_697), .A2(n_719), .B1(n_720), .B2(n_721), .Y(n_718) );
AND2x4_ASAP7_75t_L g697 ( .A(n_698), .B(n_699), .Y(n_697) );
INVx1_ASAP7_75t_L g712 ( .A(n_701), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g834 ( .A1(n_702), .A2(n_705), .B1(n_819), .B2(n_835), .Y(n_834) );
OAI21xp5_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_709), .B(n_710), .Y(n_707) );
OAI21xp33_ASAP7_75t_L g711 ( .A1(n_710), .A2(n_712), .B(n_713), .Y(n_711) );
INVx1_ASAP7_75t_L g805 ( .A(n_714), .Y(n_805) );
XNOR2xp5_ASAP7_75t_L g714 ( .A(n_715), .B(n_716), .Y(n_714) );
NOR2x1_ASAP7_75t_L g716 ( .A(n_717), .B(n_762), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_718), .B(n_722), .Y(n_717) );
INVx3_ASAP7_75t_L g855 ( .A(n_720), .Y(n_855) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
HB1xp67_ASAP7_75t_L g757 ( .A(n_726), .Y(n_757) );
OAI221xp5_ASAP7_75t_L g727 ( .A1(n_728), .A2(n_733), .B1(n_740), .B2(n_745), .C(n_751), .Y(n_727) );
OAI22xp5_ASAP7_75t_L g728 ( .A1(n_729), .A2(n_730), .B1(n_731), .B2(n_732), .Y(n_728) );
OAI221xp5_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_735), .B1(n_736), .B2(n_738), .C(n_739), .Y(n_733) );
OR2x6_ASAP7_75t_L g751 ( .A(n_734), .B(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g1003 ( .A(n_734), .Y(n_1003) );
OAI211xp5_ASAP7_75t_L g786 ( .A1(n_735), .A2(n_787), .B(n_790), .C(n_791), .Y(n_786) );
INVx3_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
INVx2_ASAP7_75t_SL g741 ( .A(n_737), .Y(n_741) );
INVx5_ASAP7_75t_L g847 ( .A(n_737), .Y(n_847) );
OAI22xp5_ASAP7_75t_L g740 ( .A1(n_741), .A2(n_742), .B1(n_743), .B2(n_744), .Y(n_740) );
OAI221xp5_ASAP7_75t_L g839 ( .A1(n_741), .A2(n_840), .B1(n_841), .B2(n_842), .C(n_843), .Y(n_839) );
OAI21xp5_ASAP7_75t_SL g745 ( .A1(n_746), .A2(n_748), .B(n_749), .Y(n_745) );
INVx3_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
AOI22xp5_ASAP7_75t_L g770 ( .A1(n_755), .A2(n_771), .B1(n_773), .B2(n_774), .Y(n_770) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx4_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
NAND3xp33_ASAP7_75t_L g762 ( .A(n_763), .B(n_794), .C(n_800), .Y(n_762) );
NOR3xp33_ASAP7_75t_SL g763 ( .A(n_764), .B(n_780), .C(n_783), .Y(n_763) );
OAI21xp5_ASAP7_75t_SL g764 ( .A1(n_765), .A2(n_769), .B(n_770), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_766), .B(n_768), .Y(n_765) );
INVx1_ASAP7_75t_SL g771 ( .A(n_772), .Y(n_771) );
INVx2_ASAP7_75t_SL g774 ( .A(n_775), .Y(n_774) );
NAND2x2_ASAP7_75t_L g775 ( .A(n_776), .B(n_778), .Y(n_775) );
INVx1_ASAP7_75t_L g793 ( .A(n_776), .Y(n_793) );
INVx2_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx2_ASAP7_75t_SL g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g799 ( .A(n_782), .Y(n_799) );
OAI21xp5_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_786), .B(n_792), .Y(n_783) );
INVx2_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
INVx2_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
BUFx2_ASAP7_75t_L g821 ( .A(n_789), .Y(n_821) );
BUFx2_ASAP7_75t_L g908 ( .A(n_789), .Y(n_908) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_795), .B(n_796), .Y(n_794) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_801), .B(n_802), .Y(n_800) );
AOI21xp5_ASAP7_75t_L g809 ( .A1(n_810), .A2(n_832), .B(n_833), .Y(n_809) );
NAND4xp25_ASAP7_75t_L g810 ( .A(n_811), .B(n_813), .C(n_823), .D(n_828), .Y(n_810) );
OAI221xp5_ASAP7_75t_L g846 ( .A1(n_829), .A2(n_847), .B1(n_848), .B2(n_849), .C(n_850), .Y(n_846) );
OAI22xp5_ASAP7_75t_SL g837 ( .A1(n_838), .A2(n_839), .B1(n_845), .B2(n_846), .Y(n_837) );
INVx2_ASAP7_75t_SL g875 ( .A(n_844), .Y(n_875) );
BUFx3_ASAP7_75t_L g1037 ( .A(n_844), .Y(n_1037) );
INVx1_ASAP7_75t_L g1360 ( .A(n_844), .Y(n_1360) );
INVx8_ASAP7_75t_L g1107 ( .A(n_847), .Y(n_1107) );
OAI22xp5_ASAP7_75t_L g995 ( .A1(n_848), .A2(n_996), .B1(n_997), .B2(n_998), .Y(n_995) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_853), .B(n_854), .Y(n_852) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_857), .B(n_858), .Y(n_856) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_858), .B(n_870), .Y(n_869) );
NAND2xp5_ASAP7_75t_L g1008 ( .A(n_858), .B(n_976), .Y(n_1008) );
INVx2_ASAP7_75t_L g917 ( .A(n_859), .Y(n_917) );
XOR2x2_ASAP7_75t_L g859 ( .A(n_860), .B(n_915), .Y(n_859) );
NAND2xp5_ASAP7_75t_SL g860 ( .A(n_861), .B(n_889), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_864), .B(n_872), .Y(n_863) );
NOR2xp33_ASAP7_75t_L g864 ( .A(n_865), .B(n_868), .Y(n_864) );
NAND2xp5_ASAP7_75t_SL g868 ( .A(n_869), .B(n_871), .Y(n_868) );
NAND4xp25_ASAP7_75t_L g1005 ( .A(n_871), .B(n_1006), .C(n_1008), .D(n_1009), .Y(n_1005) );
INVx2_ASAP7_75t_L g874 ( .A(n_875), .Y(n_874) );
BUFx2_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
BUFx2_ASAP7_75t_L g1035 ( .A(n_880), .Y(n_1035) );
BUFx2_ASAP7_75t_L g1108 ( .A(n_880), .Y(n_1108) );
INVx1_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
NAND3xp33_ASAP7_75t_SL g890 ( .A(n_891), .B(n_894), .C(n_900), .Y(n_890) );
INVx2_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
INVx1_ASAP7_75t_SL g898 ( .A(n_899), .Y(n_898) );
INVx2_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
INVx4_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
INVx5_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
INVx1_ASAP7_75t_L g1132 ( .A(n_919), .Y(n_1132) );
XNOR2xp5_ASAP7_75t_L g919 ( .A(n_920), .B(n_1012), .Y(n_919) );
INVx1_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
INVx1_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
AOI22xp5_ASAP7_75t_L g922 ( .A1(n_923), .A2(n_954), .B1(n_955), .B2(n_1011), .Y(n_922) );
INVx1_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
HB1xp67_ASAP7_75t_L g1011 ( .A(n_924), .Y(n_1011) );
AND2x2_ASAP7_75t_L g925 ( .A(n_926), .B(n_941), .Y(n_925) );
AOI22xp5_ASAP7_75t_L g933 ( .A1(n_934), .A2(n_937), .B1(n_938), .B2(n_940), .Y(n_933) );
NAND3xp33_ASAP7_75t_L g942 ( .A(n_943), .B(n_946), .C(n_949), .Y(n_942) );
INVxp67_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
NOR3xp33_ASAP7_75t_L g956 ( .A(n_957), .B(n_1005), .C(n_1010), .Y(n_956) );
NAND2xp5_ASAP7_75t_L g957 ( .A(n_958), .B(n_979), .Y(n_957) );
NAND2xp5_ASAP7_75t_L g960 ( .A(n_961), .B(n_966), .Y(n_960) );
INVx1_ASAP7_75t_L g962 ( .A(n_963), .Y(n_962) );
INVx1_ASAP7_75t_L g964 ( .A(n_965), .Y(n_964) );
INVx1_ASAP7_75t_L g1042 ( .A(n_965), .Y(n_1042) );
INVx1_ASAP7_75t_L g1057 ( .A(n_965), .Y(n_1057) );
NAND3xp33_ASAP7_75t_L g969 ( .A(n_970), .B(n_974), .C(n_977), .Y(n_969) );
AOI21xp5_ASAP7_75t_L g979 ( .A1(n_980), .A2(n_981), .B(n_982), .Y(n_979) );
OAI22xp5_ASAP7_75t_L g983 ( .A1(n_984), .A2(n_985), .B1(n_986), .B2(n_987), .Y(n_983) );
INVx1_ASAP7_75t_L g987 ( .A(n_988), .Y(n_987) );
OAI22xp33_ASAP7_75t_L g989 ( .A1(n_990), .A2(n_991), .B1(n_992), .B2(n_993), .Y(n_989) );
INVx1_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
OAI22xp5_ASAP7_75t_L g999 ( .A1(n_1000), .A2(n_1001), .B1(n_1002), .B2(n_1004), .Y(n_999) );
INVx1_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
XNOR2xp5_ASAP7_75t_L g1012 ( .A(n_1013), .B(n_1095), .Y(n_1012) );
AOI22xp5_ASAP7_75t_L g1013 ( .A1(n_1014), .A2(n_1015), .B1(n_1059), .B2(n_1060), .Y(n_1013) );
INVx1_ASAP7_75t_L g1014 ( .A(n_1015), .Y(n_1014) );
AND3x1_ASAP7_75t_L g1020 ( .A(n_1021), .B(n_1024), .C(n_1027), .Y(n_1020) );
INVx2_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
OAI21xp5_ASAP7_75t_L g1038 ( .A1(n_1039), .A2(n_1047), .B(n_1058), .Y(n_1038) );
INVx2_ASAP7_75t_L g1043 ( .A(n_1044), .Y(n_1043) );
OAI221xp5_ASAP7_75t_L g1049 ( .A1(n_1050), .A2(n_1052), .B1(n_1053), .B2(n_1055), .C(n_1056), .Y(n_1049) );
BUFx6f_ASAP7_75t_L g1050 ( .A(n_1051), .Y(n_1050) );
BUFx6f_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
INVx1_ASAP7_75t_L g1059 ( .A(n_1060), .Y(n_1059) );
HB1xp67_ASAP7_75t_L g1060 ( .A(n_1061), .Y(n_1060) );
NAND3xp33_ASAP7_75t_L g1062 ( .A(n_1063), .B(n_1080), .C(n_1083), .Y(n_1062) );
NAND2xp5_ASAP7_75t_L g1084 ( .A(n_1085), .B(n_1087), .Y(n_1084) );
INVxp67_ASAP7_75t_SL g1095 ( .A(n_1096), .Y(n_1095) );
NAND3xp33_ASAP7_75t_L g1097 ( .A(n_1098), .B(n_1111), .C(n_1114), .Y(n_1097) );
NAND2xp5_ASAP7_75t_L g1099 ( .A(n_1100), .B(n_1103), .Y(n_1099) );
NAND2xp5_ASAP7_75t_L g1124 ( .A(n_1125), .B(n_1128), .Y(n_1124) );
OAI221xp5_ASAP7_75t_L g1133 ( .A1(n_1134), .A2(n_1347), .B1(n_1350), .B2(n_1385), .C(n_1388), .Y(n_1133) );
AND3x1_ASAP7_75t_L g1134 ( .A(n_1135), .B(n_1284), .C(n_1321), .Y(n_1134) );
AOI211xp5_ASAP7_75t_SL g1135 ( .A1(n_1136), .A2(n_1157), .B(n_1211), .C(n_1260), .Y(n_1135) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1137), .Y(n_1136) );
NAND2xp5_ASAP7_75t_L g1137 ( .A(n_1138), .B(n_1152), .Y(n_1137) );
INVx3_ASAP7_75t_L g1232 ( .A(n_1138), .Y(n_1232) );
A2O1A1Ixp33_ASAP7_75t_L g1250 ( .A1(n_1138), .A2(n_1251), .B(n_1252), .C(n_1253), .Y(n_1250) );
NAND2xp5_ASAP7_75t_L g1313 ( .A(n_1138), .B(n_1210), .Y(n_1313) );
AND2x2_ASAP7_75t_L g1138 ( .A(n_1139), .B(n_1146), .Y(n_1138) );
INVx2_ASAP7_75t_L g1349 ( .A(n_1140), .Y(n_1349) );
AND2x6_ASAP7_75t_L g1140 ( .A(n_1141), .B(n_1142), .Y(n_1140) );
AND2x2_ASAP7_75t_L g1144 ( .A(n_1141), .B(n_1145), .Y(n_1144) );
AND2x4_ASAP7_75t_L g1147 ( .A(n_1141), .B(n_1148), .Y(n_1147) );
AND2x6_ASAP7_75t_L g1150 ( .A(n_1141), .B(n_1151), .Y(n_1150) );
AND2x2_ASAP7_75t_L g1155 ( .A(n_1141), .B(n_1145), .Y(n_1155) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_1141), .B(n_1145), .Y(n_1176) );
OAI21xp5_ASAP7_75t_L g1396 ( .A1(n_1142), .A2(n_1397), .B(n_1398), .Y(n_1396) );
AND2x2_ASAP7_75t_L g1148 ( .A(n_1143), .B(n_1149), .Y(n_1148) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1152), .Y(n_1223) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1152), .Y(n_1247) );
AND2x2_ASAP7_75t_L g1252 ( .A(n_1152), .B(n_1192), .Y(n_1252) );
NAND2xp5_ASAP7_75t_L g1258 ( .A(n_1152), .B(n_1259), .Y(n_1258) );
AND2x2_ASAP7_75t_L g1292 ( .A(n_1152), .B(n_1174), .Y(n_1292) );
NAND3xp33_ASAP7_75t_L g1298 ( .A(n_1152), .B(n_1268), .C(n_1299), .Y(n_1298) );
INVx1_ASAP7_75t_L g1152 ( .A(n_1153), .Y(n_1152) );
AND2x2_ASAP7_75t_L g1219 ( .A(n_1153), .B(n_1210), .Y(n_1219) );
NAND2xp5_ASAP7_75t_L g1224 ( .A(n_1153), .B(n_1225), .Y(n_1224) );
INVx1_ASAP7_75t_L g1229 ( .A(n_1153), .Y(n_1229) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1153), .Y(n_1270) );
AND2x2_ASAP7_75t_L g1276 ( .A(n_1153), .B(n_1174), .Y(n_1276) );
NAND2xp5_ASAP7_75t_L g1153 ( .A(n_1154), .B(n_1156), .Y(n_1153) );
OAI211xp5_ASAP7_75t_SL g1157 ( .A1(n_1158), .A2(n_1168), .B(n_1182), .C(n_1199), .Y(n_1157) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1159), .Y(n_1158) );
AND2x2_ASAP7_75t_L g1159 ( .A(n_1160), .B(n_1164), .Y(n_1159) );
NOR2xp33_ASAP7_75t_L g1293 ( .A(n_1160), .B(n_1294), .Y(n_1293) );
INVx1_ASAP7_75t_L g1160 ( .A(n_1161), .Y(n_1160) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1161), .Y(n_1190) );
AND2x2_ASAP7_75t_L g1196 ( .A(n_1161), .B(n_1187), .Y(n_1196) );
INVx1_ASAP7_75t_L g1205 ( .A(n_1161), .Y(n_1205) );
OR2x2_ASAP7_75t_L g1226 ( .A(n_1161), .B(n_1186), .Y(n_1226) );
NAND2xp5_ASAP7_75t_L g1230 ( .A(n_1161), .B(n_1165), .Y(n_1230) );
NAND2xp5_ASAP7_75t_L g1237 ( .A(n_1161), .B(n_1164), .Y(n_1237) );
NAND2x1_ASAP7_75t_L g1161 ( .A(n_1162), .B(n_1163), .Y(n_1161) );
OR2x2_ASAP7_75t_L g1194 ( .A(n_1164), .B(n_1195), .Y(n_1194) );
OR2x2_ASAP7_75t_L g1203 ( .A(n_1164), .B(n_1204), .Y(n_1203) );
NAND2xp5_ASAP7_75t_L g1215 ( .A(n_1164), .B(n_1207), .Y(n_1215) );
AND2x2_ASAP7_75t_L g1256 ( .A(n_1164), .B(n_1196), .Y(n_1256) );
OR2x2_ASAP7_75t_L g1264 ( .A(n_1164), .B(n_1226), .Y(n_1264) );
AND2x2_ASAP7_75t_L g1283 ( .A(n_1164), .B(n_1244), .Y(n_1283) );
NAND2xp5_ASAP7_75t_L g1305 ( .A(n_1164), .B(n_1185), .Y(n_1305) );
INVx2_ASAP7_75t_L g1164 ( .A(n_1165), .Y(n_1164) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_1165), .B(n_1179), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1165), .B(n_1198), .Y(n_1197) );
AOI22xp5_ASAP7_75t_L g1199 ( .A1(n_1165), .A2(n_1200), .B1(n_1202), .B2(n_1206), .Y(n_1199) );
AND2x2_ASAP7_75t_L g1249 ( .A(n_1165), .B(n_1190), .Y(n_1249) );
NOR2xp33_ASAP7_75t_L g1266 ( .A(n_1165), .B(n_1267), .Y(n_1266) );
AND2x2_ASAP7_75t_L g1278 ( .A(n_1165), .B(n_1186), .Y(n_1278) );
OR2x2_ASAP7_75t_L g1312 ( .A(n_1165), .B(n_1226), .Y(n_1312) );
OR2x2_ASAP7_75t_L g1317 ( .A(n_1165), .B(n_1187), .Y(n_1317) );
NAND2xp5_ASAP7_75t_L g1337 ( .A(n_1165), .B(n_1187), .Y(n_1337) );
AND2x2_ASAP7_75t_L g1165 ( .A(n_1166), .B(n_1167), .Y(n_1165) );
OR2x2_ASAP7_75t_L g1168 ( .A(n_1169), .B(n_1178), .Y(n_1168) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1169), .Y(n_1259) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1169), .Y(n_1333) );
NAND2xp5_ASAP7_75t_L g1169 ( .A(n_1170), .B(n_1174), .Y(n_1169) );
INVx2_ASAP7_75t_L g1192 ( .A(n_1170), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1275 ( .A(n_1170), .B(n_1276), .Y(n_1275) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1171), .Y(n_1170) );
OR2x2_ASAP7_75t_L g1201 ( .A(n_1171), .B(n_1174), .Y(n_1201) );
INVx2_ASAP7_75t_SL g1209 ( .A(n_1171), .Y(n_1209) );
AND2x2_ASAP7_75t_L g1225 ( .A(n_1171), .B(n_1207), .Y(n_1225) );
NAND2xp5_ASAP7_75t_L g1274 ( .A(n_1171), .B(n_1210), .Y(n_1274) );
NAND2xp5_ASAP7_75t_L g1301 ( .A(n_1171), .B(n_1213), .Y(n_1301) );
AND2x2_ASAP7_75t_L g1171 ( .A(n_1172), .B(n_1173), .Y(n_1171) );
CKINVDCx5p33_ASAP7_75t_R g1210 ( .A(n_1174), .Y(n_1210) );
AOI221xp5_ASAP7_75t_L g1212 ( .A1(n_1174), .A2(n_1185), .B1(n_1213), .B2(n_1216), .C(n_1220), .Y(n_1212) );
AOI221xp5_ASAP7_75t_L g1233 ( .A1(n_1174), .A2(n_1187), .B1(n_1234), .B2(n_1238), .C(n_1241), .Y(n_1233) );
NAND2xp5_ASAP7_75t_L g1323 ( .A(n_1174), .B(n_1179), .Y(n_1323) );
NAND2xp5_ASAP7_75t_L g1340 ( .A(n_1174), .B(n_1341), .Y(n_1340) );
AND2x4_ASAP7_75t_L g1174 ( .A(n_1175), .B(n_1177), .Y(n_1174) );
AND2x2_ASAP7_75t_L g1198 ( .A(n_1178), .B(n_1185), .Y(n_1198) );
NAND2xp5_ASAP7_75t_L g1235 ( .A(n_1178), .B(n_1236), .Y(n_1235) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1178), .Y(n_1263) );
AND2x2_ASAP7_75t_L g1277 ( .A(n_1178), .B(n_1278), .Y(n_1277) );
OAI211xp5_ASAP7_75t_L g1286 ( .A1(n_1178), .A2(n_1287), .B(n_1289), .C(n_1291), .Y(n_1286) );
NAND2xp5_ASAP7_75t_L g1319 ( .A(n_1178), .B(n_1320), .Y(n_1319) );
OR2x2_ASAP7_75t_L g1339 ( .A(n_1178), .B(n_1237), .Y(n_1339) );
CKINVDCx5p33_ASAP7_75t_R g1178 ( .A(n_1179), .Y(n_1178) );
INVx3_ASAP7_75t_L g1207 ( .A(n_1179), .Y(n_1207) );
AND2x2_ASAP7_75t_L g1222 ( .A(n_1179), .B(n_1223), .Y(n_1222) );
NAND2xp5_ASAP7_75t_L g1343 ( .A(n_1179), .B(n_1218), .Y(n_1343) );
AND2x4_ASAP7_75t_SL g1179 ( .A(n_1180), .B(n_1181), .Y(n_1179) );
OAI22xp33_ASAP7_75t_L g1182 ( .A1(n_1183), .A2(n_1192), .B1(n_1193), .B2(n_1197), .Y(n_1182) );
NAND2xp5_ASAP7_75t_L g1183 ( .A(n_1184), .B(n_1192), .Y(n_1183) );
NAND2xp5_ASAP7_75t_L g1184 ( .A(n_1185), .B(n_1191), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1254 ( .A(n_1185), .B(n_1255), .Y(n_1254) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_1186), .B(n_1190), .Y(n_1185) );
OAI322xp33_ASAP7_75t_L g1220 ( .A1(n_1186), .A2(n_1192), .A3(n_1221), .B1(n_1224), .B2(n_1226), .C1(n_1227), .C2(n_1230), .Y(n_1220) );
INVx1_ASAP7_75t_L g1186 ( .A(n_1187), .Y(n_1186) );
OR2x2_ASAP7_75t_L g1204 ( .A(n_1187), .B(n_1205), .Y(n_1204) );
AND2x2_ASAP7_75t_L g1187 ( .A(n_1188), .B(n_1189), .Y(n_1187) );
AND2x2_ASAP7_75t_L g1243 ( .A(n_1191), .B(n_1244), .Y(n_1243) );
AND2x2_ASAP7_75t_L g1307 ( .A(n_1191), .B(n_1196), .Y(n_1307) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1192), .Y(n_1251) );
NAND2xp5_ASAP7_75t_L g1289 ( .A(n_1192), .B(n_1290), .Y(n_1289) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_1192), .B(n_1307), .Y(n_1306) );
NAND2xp5_ASAP7_75t_L g1329 ( .A(n_1192), .B(n_1202), .Y(n_1329) );
AND2x2_ASAP7_75t_L g1346 ( .A(n_1192), .B(n_1223), .Y(n_1346) );
O2A1O1Ixp33_ASAP7_75t_L g1330 ( .A1(n_1193), .A2(n_1331), .B(n_1333), .C(n_1334), .Y(n_1330) );
INVx1_ASAP7_75t_L g1193 ( .A(n_1194), .Y(n_1193) );
OR2x2_ASAP7_75t_L g1214 ( .A(n_1195), .B(n_1215), .Y(n_1214) );
OAI22xp5_ASAP7_75t_SL g1322 ( .A1(n_1195), .A2(n_1227), .B1(n_1323), .B2(n_1324), .Y(n_1322) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1196), .Y(n_1195) );
NAND2xp5_ASAP7_75t_L g1227 ( .A(n_1200), .B(n_1228), .Y(n_1227) );
AOI322xp5_ASAP7_75t_L g1248 ( .A1(n_1200), .A2(n_1222), .A3(n_1249), .B1(n_1250), .B2(n_1254), .C1(n_1256), .C2(n_1257), .Y(n_1248) );
INVx2_ASAP7_75t_L g1200 ( .A(n_1201), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1345 ( .A(n_1202), .B(n_1207), .Y(n_1345) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1203), .Y(n_1202) );
INVx1_ASAP7_75t_L g1244 ( .A(n_1204), .Y(n_1244) );
NOR2xp33_ASAP7_75t_L g1288 ( .A(n_1204), .B(n_1273), .Y(n_1288) );
NOR2xp33_ASAP7_75t_L g1206 ( .A(n_1207), .B(n_1208), .Y(n_1206) );
NAND2xp5_ASAP7_75t_L g1239 ( .A(n_1207), .B(n_1240), .Y(n_1239) );
CKINVDCx14_ASAP7_75t_R g1271 ( .A(n_1207), .Y(n_1271) );
NOR2xp33_ASAP7_75t_L g1295 ( .A(n_1207), .B(n_1218), .Y(n_1295) );
AND2x2_ASAP7_75t_L g1299 ( .A(n_1207), .B(n_1209), .Y(n_1299) );
INVx1_ASAP7_75t_L g1240 ( .A(n_1208), .Y(n_1240) );
OR2x2_ASAP7_75t_L g1208 ( .A(n_1209), .B(n_1210), .Y(n_1208) );
INVx2_ASAP7_75t_L g1218 ( .A(n_1209), .Y(n_1218) );
A2O1A1Ixp33_ASAP7_75t_L g1303 ( .A1(n_1209), .A2(n_1304), .B(n_1306), .C(n_1308), .Y(n_1303) );
A2O1A1Ixp33_ASAP7_75t_L g1335 ( .A1(n_1209), .A2(n_1276), .B(n_1336), .C(n_1338), .Y(n_1335) );
NAND2xp5_ASAP7_75t_L g1261 ( .A(n_1210), .B(n_1232), .Y(n_1261) );
AND2x2_ASAP7_75t_L g1269 ( .A(n_1210), .B(n_1270), .Y(n_1269) );
OAI221xp5_ASAP7_75t_SL g1211 ( .A1(n_1212), .A2(n_1231), .B1(n_1233), .B2(n_1245), .C(n_1248), .Y(n_1211) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1214), .Y(n_1213) );
INVx1_ASAP7_75t_L g1255 ( .A(n_1215), .Y(n_1255) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1217), .Y(n_1216) );
NAND2xp5_ASAP7_75t_L g1217 ( .A(n_1218), .B(n_1219), .Y(n_1217) );
NOR2xp33_ASAP7_75t_L g1325 ( .A(n_1218), .B(n_1326), .Y(n_1325) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1219), .Y(n_1253) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1222), .Y(n_1221) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1225), .Y(n_1281) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1226), .Y(n_1268) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1229), .Y(n_1228) );
CKINVDCx14_ASAP7_75t_R g1285 ( .A(n_1231), .Y(n_1285) );
OAI221xp5_ASAP7_75t_L g1309 ( .A1(n_1231), .A2(n_1310), .B1(n_1313), .B2(n_1314), .C(n_1315), .Y(n_1309) );
OAI31xp33_ASAP7_75t_SL g1321 ( .A1(n_1231), .A2(n_1322), .A3(n_1325), .B(n_1328), .Y(n_1321) );
CKINVDCx14_ASAP7_75t_R g1231 ( .A(n_1232), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1246 ( .A(n_1232), .B(n_1247), .Y(n_1246) );
AOI322xp5_ASAP7_75t_L g1265 ( .A1(n_1234), .A2(n_1266), .A3(n_1269), .B1(n_1271), .B2(n_1272), .C1(n_1275), .C2(n_1277), .Y(n_1265) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1235), .Y(n_1234) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1237), .Y(n_1236) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1239), .Y(n_1238) );
NAND2xp5_ASAP7_75t_L g1242 ( .A(n_1240), .B(n_1243), .Y(n_1242) );
NAND2xp5_ASAP7_75t_L g1314 ( .A(n_1240), .B(n_1311), .Y(n_1314) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1242), .Y(n_1241) );
NOR2xp33_ASAP7_75t_L g1267 ( .A(n_1244), .B(n_1268), .Y(n_1267) );
CKINVDCx14_ASAP7_75t_R g1245 ( .A(n_1246), .Y(n_1245) );
OR2x2_ASAP7_75t_L g1273 ( .A(n_1247), .B(n_1274), .Y(n_1273) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1249), .Y(n_1342) );
OAI211xp5_ASAP7_75t_SL g1328 ( .A1(n_1253), .A2(n_1329), .B(n_1330), .C(n_1344), .Y(n_1328) );
NAND2xp5_ASAP7_75t_L g1332 ( .A(n_1255), .B(n_1268), .Y(n_1332) );
NOR2xp33_ASAP7_75t_L g1324 ( .A(n_1256), .B(n_1296), .Y(n_1324) );
AND2x2_ASAP7_75t_L g1327 ( .A(n_1256), .B(n_1263), .Y(n_1327) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1258), .Y(n_1257) );
OAI211xp5_ASAP7_75t_SL g1260 ( .A1(n_1261), .A2(n_1262), .B(n_1265), .C(n_1279), .Y(n_1260) );
INVxp67_ASAP7_75t_SL g1308 ( .A(n_1261), .Y(n_1308) );
INVxp67_ASAP7_75t_L g1290 ( .A(n_1262), .Y(n_1290) );
OR2x2_ASAP7_75t_L g1262 ( .A(n_1263), .B(n_1264), .Y(n_1262) );
INVx2_ASAP7_75t_L g1296 ( .A(n_1264), .Y(n_1296) );
AOI221xp5_ASAP7_75t_SL g1291 ( .A1(n_1269), .A2(n_1292), .B1(n_1293), .B2(n_1296), .C(n_1297), .Y(n_1291) );
NAND2xp5_ASAP7_75t_L g1279 ( .A(n_1270), .B(n_1280), .Y(n_1279) );
NAND2xp5_ASAP7_75t_L g1310 ( .A(n_1271), .B(n_1311), .Y(n_1310) );
INVx1_ASAP7_75t_L g1272 ( .A(n_1273), .Y(n_1272) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1274), .Y(n_1320) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1276), .Y(n_1302) );
NOR2xp33_ASAP7_75t_L g1280 ( .A(n_1281), .B(n_1282), .Y(n_1280) );
INVx2_ASAP7_75t_L g1282 ( .A(n_1283), .Y(n_1282) );
AOI211xp5_ASAP7_75t_L g1284 ( .A1(n_1285), .A2(n_1286), .B(n_1300), .C(n_1309), .Y(n_1284) );
INVxp67_ASAP7_75t_L g1287 ( .A(n_1288), .Y(n_1287) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1295), .Y(n_1294) );
OAI21xp5_ASAP7_75t_L g1315 ( .A1(n_1296), .A2(n_1316), .B(n_1318), .Y(n_1315) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1298), .Y(n_1297) );
OAI21xp5_ASAP7_75t_L g1300 ( .A1(n_1301), .A2(n_1302), .B(n_1303), .Y(n_1300) );
OAI21xp33_ASAP7_75t_L g1344 ( .A1(n_1304), .A2(n_1345), .B(n_1346), .Y(n_1344) );
INVx1_ASAP7_75t_L g1304 ( .A(n_1305), .Y(n_1304) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1312), .Y(n_1311) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1317), .Y(n_1316) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1319), .Y(n_1318) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1327), .Y(n_1326) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1332), .Y(n_1331) );
NAND2xp5_ASAP7_75t_SL g1334 ( .A(n_1335), .B(n_1340), .Y(n_1334) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1337), .Y(n_1336) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1339), .Y(n_1338) );
NOR2xp33_ASAP7_75t_L g1341 ( .A(n_1342), .B(n_1343), .Y(n_1341) );
CKINVDCx20_ASAP7_75t_R g1347 ( .A(n_1348), .Y(n_1347) );
CKINVDCx20_ASAP7_75t_R g1348 ( .A(n_1349), .Y(n_1348) );
HB1xp67_ASAP7_75t_L g1394 ( .A(n_1351), .Y(n_1394) );
NAND3xp33_ASAP7_75t_L g1351 ( .A(n_1352), .B(n_1365), .C(n_1368), .Y(n_1351) );
NAND2xp5_ASAP7_75t_L g1353 ( .A(n_1354), .B(n_1357), .Y(n_1353) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1360), .Y(n_1359) );
OAI21xp5_ASAP7_75t_L g1368 ( .A1(n_1369), .A2(n_1377), .B(n_1384), .Y(n_1368) );
BUFx2_ASAP7_75t_L g1375 ( .A(n_1376), .Y(n_1375) );
CKINVDCx5p33_ASAP7_75t_R g1385 ( .A(n_1386), .Y(n_1385) );
HB1xp67_ASAP7_75t_SL g1389 ( .A(n_1390), .Y(n_1389) );
BUFx3_ASAP7_75t_L g1390 ( .A(n_1391), .Y(n_1390) );
INVxp33_ASAP7_75t_SL g1392 ( .A(n_1393), .Y(n_1392) );
HB1xp67_ASAP7_75t_L g1395 ( .A(n_1396), .Y(n_1395) );
INVx1_ASAP7_75t_L g1398 ( .A(n_1399), .Y(n_1398) );
endmodule