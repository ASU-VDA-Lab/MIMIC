module fake_jpeg_14917_n_355 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_355);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_355;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_12),
.B(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_43),
.Y(n_57)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_24),
.Y(n_44)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_16),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_45),
.B(n_46),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_22),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_51),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_1),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_53),
.Y(n_69)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_39),
.A2(n_32),
.B1(n_35),
.B2(n_18),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_54),
.A2(n_60),
.B1(n_31),
.B2(n_34),
.Y(n_101)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_37),
.B1(n_22),
.B2(n_36),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_46),
.B(n_18),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_63),
.B(n_17),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_36),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_30),
.Y(n_90)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_51),
.Y(n_70)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_50),
.A2(n_37),
.B1(n_38),
.B2(n_21),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_20),
.B1(n_23),
.B2(n_30),
.Y(n_88)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_76),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_24),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_77),
.B(n_79),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_69),
.A2(n_53),
.B(n_21),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_78),
.A2(n_65),
.B(n_57),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_29),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_29),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_81),
.B(n_87),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_19),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_82),
.B(n_85),
.Y(n_118)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_62),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_19),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_86),
.B(n_92),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_38),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_88),
.A2(n_111),
.B1(n_68),
.B2(n_66),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g89 ( 
.A(n_71),
.Y(n_89)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_90),
.B(n_103),
.Y(n_126)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

INVx3_ASAP7_75t_SL g138 ( 
.A(n_93),
.Y(n_138)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

NAND2xp33_ASAP7_75t_SL g95 ( 
.A(n_75),
.B(n_39),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_95),
.A2(n_75),
.B1(n_76),
.B2(n_67),
.Y(n_142)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_56),
.B(n_19),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_97),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_55),
.A2(n_31),
.B1(n_20),
.B2(n_23),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_98),
.A2(n_108),
.B1(n_68),
.B2(n_66),
.Y(n_115)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_100),
.Y(n_120)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_104),
.Y(n_134)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_71),
.Y(n_107)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_55),
.A2(n_34),
.B1(n_44),
.B2(n_13),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_54),
.A2(n_44),
.B1(n_28),
.B2(n_25),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_60),
.A2(n_44),
.B1(n_48),
.B2(n_49),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_114),
.A2(n_99),
.B1(n_80),
.B2(n_92),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_115),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_116),
.B(n_28),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_106),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_139),
.Y(n_152)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_77),
.B(n_57),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_129),
.B(n_141),
.C(n_17),
.Y(n_172)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_132),
.Y(n_163)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

INVx11_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_91),
.A2(n_75),
.B1(n_61),
.B2(n_67),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_106),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_79),
.B(n_43),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_142),
.A2(n_112),
.B(n_95),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_130),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_143),
.B(n_149),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_144),
.A2(n_167),
.B1(n_119),
.B2(n_120),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_141),
.B(n_78),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_145),
.B(n_146),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_129),
.B(n_81),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_147),
.A2(n_157),
.B(n_160),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_124),
.A2(n_90),
.B1(n_91),
.B2(n_101),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_148),
.A2(n_156),
.B1(n_159),
.B2(n_138),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_130),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_90),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_155),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_87),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_153),
.B(n_158),
.C(n_170),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_124),
.A2(n_109),
.B1(n_74),
.B2(n_80),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_154),
.A2(n_139),
.B1(n_127),
.B2(n_120),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_125),
.B(n_84),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_140),
.A2(n_112),
.B1(n_94),
.B2(n_83),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_140),
.A2(n_110),
.B(n_85),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_116),
.B(n_131),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_114),
.A2(n_83),
.B1(n_89),
.B2(n_110),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_142),
.A2(n_17),
.B(n_2),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_123),
.B(n_96),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_119),
.Y(n_182)
);

AO22x1_ASAP7_75t_L g165 ( 
.A1(n_138),
.A2(n_89),
.B1(n_48),
.B2(n_49),
.Y(n_165)
);

A2O1A1Ixp33_ASAP7_75t_SL g187 ( 
.A1(n_165),
.A2(n_136),
.B(n_134),
.C(n_121),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_113),
.A2(n_105),
.B1(n_61),
.B2(n_49),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_118),
.A2(n_43),
.B(n_47),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_168),
.A2(n_169),
.B(n_171),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_133),
.A2(n_137),
.B(n_118),
.Y(n_169)
);

MAJx2_ASAP7_75t_L g170 ( 
.A(n_126),
.B(n_47),
.C(n_17),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_172),
.B(n_123),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_126),
.B(n_17),
.C(n_93),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_26),
.C(n_35),
.Y(n_205)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_137),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_174),
.Y(n_188)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_152),
.Y(n_175)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_175),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_176),
.A2(n_183),
.B1(n_174),
.B2(n_166),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_178),
.B(n_186),
.C(n_205),
.Y(n_237)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_152),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_179),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_181),
.A2(n_185),
.B1(n_204),
.B2(n_207),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_182),
.B(n_195),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_160),
.A2(n_121),
.B1(n_117),
.B2(n_134),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_132),
.Y(n_186)
);

OA22x2_ASAP7_75t_L g211 ( 
.A1(n_187),
.A2(n_149),
.B1(n_157),
.B2(n_164),
.Y(n_211)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_150),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_189),
.Y(n_209)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_150),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_190),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_147),
.A2(n_136),
.B(n_117),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_191),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_163),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_193),
.B(n_194),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_163),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_161),
.B(n_128),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_169),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_196),
.B(n_197),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_146),
.B(n_122),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_153),
.B(n_122),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_202),
.Y(n_227)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_165),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_199),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_158),
.B(n_28),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_201),
.Y(n_212)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_165),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_155),
.B(n_156),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_203),
.A2(n_208),
.B(n_187),
.Y(n_213)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_143),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_144),
.A2(n_138),
.B1(n_35),
.B2(n_25),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_171),
.A2(n_26),
.B(n_25),
.Y(n_208)
);

OAI22x1_ASAP7_75t_L g239 ( 
.A1(n_211),
.A2(n_191),
.B1(n_183),
.B2(n_203),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_213),
.A2(n_228),
.B(n_200),
.Y(n_247)
);

OAI32xp33_ASAP7_75t_L g214 ( 
.A1(n_180),
.A2(n_151),
.A3(n_148),
.B1(n_170),
.B2(n_154),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_214),
.B(n_221),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_203),
.A2(n_162),
.B1(n_159),
.B2(n_173),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_215),
.A2(n_224),
.B1(n_234),
.B2(n_180),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_192),
.B(n_145),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_216),
.B(n_217),
.C(n_230),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_170),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_206),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_222),
.A2(n_202),
.B1(n_195),
.B2(n_190),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_176),
.A2(n_168),
.B1(n_166),
.B2(n_167),
.Y(n_224)
);

MAJx2_ASAP7_75t_L g225 ( 
.A(n_177),
.B(n_26),
.C(n_35),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_229),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_184),
.A2(n_1),
.B(n_2),
.Y(n_228)
);

AOI322xp5_ASAP7_75t_L g229 ( 
.A1(n_184),
.A2(n_16),
.A3(n_15),
.B1(n_14),
.B2(n_13),
.C1(n_6),
.C2(n_7),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_177),
.B(n_16),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_186),
.B(n_15),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_178),
.C(n_205),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_199),
.A2(n_14),
.B1(n_13),
.B2(n_4),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_182),
.B(n_2),
.Y(n_236)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_236),
.Y(n_243)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_188),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_2),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_239),
.A2(n_259),
.B1(n_218),
.B2(n_213),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_211),
.B(n_179),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_240),
.A2(n_219),
.B(n_215),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_231),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_241),
.B(n_264),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_221),
.B(n_175),
.Y(n_242)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_242),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_198),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_245),
.B(n_257),
.C(n_258),
.Y(n_271)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_220),
.Y(n_246)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_246),
.Y(n_267)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_247),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_223),
.A2(n_200),
.B(n_208),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_248),
.A2(n_256),
.B1(n_228),
.B2(n_211),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_232),
.Y(n_250)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_250),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_252),
.B(n_225),
.Y(n_282)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_220),
.Y(n_253)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_253),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_232),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_254),
.B(n_209),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_260),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_217),
.B(n_181),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_187),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_223),
.A2(n_189),
.B1(n_187),
.B2(n_4),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_237),
.B(n_3),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_261),
.B(n_263),
.C(n_236),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_227),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_262),
.B(n_210),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_214),
.B(n_3),
.Y(n_263)
);

INVx2_ASAP7_75t_SL g264 ( 
.A(n_238),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_257),
.B(n_230),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_269),
.B(n_272),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_245),
.B(n_233),
.Y(n_272)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_273),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_274),
.A2(n_280),
.B(n_247),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_249),
.A2(n_227),
.B1(n_219),
.B2(n_211),
.Y(n_275)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_275),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_251),
.B(n_235),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_282),
.C(n_251),
.Y(n_289)
);

NAND2x1_ASAP7_75t_L g278 ( 
.A(n_239),
.B(n_240),
.Y(n_278)
);

AND2x4_ASAP7_75t_L g288 ( 
.A(n_278),
.B(n_259),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_279),
.A2(n_258),
.B1(n_212),
.B2(n_252),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_241),
.A2(n_210),
.B1(n_209),
.B2(n_226),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_243),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_263),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_283),
.B(n_264),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_244),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_286),
.B(n_256),
.Y(n_291)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_287),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_288),
.B(n_289),
.Y(n_313)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_291),
.Y(n_316)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_292),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_303),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_295),
.B(n_297),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_271),
.B(n_261),
.C(n_244),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_296),
.B(n_301),
.C(n_302),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_268),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_265),
.A2(n_266),
.B1(n_270),
.B2(n_278),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_274),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_285),
.Y(n_308)
);

MAJx2_ASAP7_75t_L g300 ( 
.A(n_269),
.B(n_212),
.C(n_4),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_300),
.A2(n_275),
.B(n_6),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_271),
.B(n_272),
.C(n_276),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_3),
.C(n_5),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_277),
.B(n_5),
.Y(n_303)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_307),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_308),
.B(n_311),
.C(n_288),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_284),
.C(n_265),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_310),
.B(n_314),
.C(n_5),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_287),
.B(n_278),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_289),
.B(n_284),
.C(n_277),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_294),
.B(n_267),
.Y(n_315)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_315),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_288),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_296),
.B(n_273),
.C(n_6),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_319),
.B(n_288),
.C(n_299),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_318),
.B(n_302),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_321),
.B(n_322),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_304),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_323),
.B(n_324),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_313),
.B(n_304),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_325),
.B(n_327),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_316),
.B(n_290),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_326),
.B(n_330),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_319),
.A2(n_300),
.B1(n_6),
.B2(n_7),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_329),
.B(n_305),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_314),
.B(n_5),
.C(n_7),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_331),
.B(n_8),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_332),
.B(n_10),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_320),
.A2(n_312),
.B(n_311),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_333),
.B(n_336),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_331),
.B(n_310),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_337),
.B(n_339),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_328),
.B(n_309),
.Y(n_339)
);

AO21x1_ASAP7_75t_SL g341 ( 
.A1(n_335),
.A2(n_324),
.B(n_330),
.Y(n_341)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_341),
.Y(n_348)
);

O2A1O1Ixp33_ASAP7_75t_SL g343 ( 
.A1(n_338),
.A2(n_322),
.B(n_325),
.C(n_306),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_343),
.A2(n_345),
.B(n_334),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_340),
.B(n_306),
.C(n_308),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_346),
.A2(n_8),
.B1(n_9),
.B2(n_333),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_347),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_350),
.B(n_344),
.C(n_348),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_351),
.B(n_349),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_352),
.Y(n_353)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_353),
.A2(n_342),
.B(n_346),
.Y(n_354)
);

AOI31xp33_ASAP7_75t_L g355 ( 
.A1(n_354),
.A2(n_9),
.A3(n_347),
.B(n_353),
.Y(n_355)
);


endmodule