module fake_netlist_6_1386_n_1216 (n_52, n_1, n_91, n_326, n_256, n_209, n_367, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_350, n_78, n_84, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_65, n_230, n_141, n_383, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_111, n_314, n_378, n_377, n_35, n_183, n_79, n_375, n_338, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_39, n_344, n_73, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_213, n_294, n_302, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_155, n_109, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_381, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_352, n_9, n_107, n_6, n_14, n_89, n_374, n_366, n_103, n_272, n_185, n_348, n_69, n_376, n_293, n_31, n_334, n_53, n_370, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_83, n_363, n_323, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_102, n_204, n_261, n_312, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_61, n_237, n_244, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_345, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_277, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_317, n_149, n_90, n_347, n_24, n_54, n_328, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_135, n_165, n_351, n_259, n_177, n_364, n_295, n_385, n_190, n_262, n_187, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_1216);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_367;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_350;
input n_78;
input n_84;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_65;
input n_230;
input n_141;
input n_383;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_111;
input n_314;
input n_378;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_39;
input n_344;
input n_73;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_213;
input n_294;
input n_302;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_155;
input n_109;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_352;
input n_9;
input n_107;
input n_6;
input n_14;
input n_89;
input n_374;
input n_366;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_83;
input n_363;
input n_323;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_102;
input n_204;
input n_261;
input n_312;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_61;
input n_237;
input n_244;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_277;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_317;
input n_149;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_135;
input n_165;
input n_351;
input n_259;
input n_177;
input n_364;
input n_295;
input n_385;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_1216;

wire n_992;
wire n_591;
wire n_435;
wire n_1115;
wire n_793;
wire n_801;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_881;
wire n_1199;
wire n_875;
wire n_465;
wire n_680;
wire n_760;
wire n_741;
wire n_1008;
wire n_1027;
wire n_590;
wire n_625;
wire n_661;
wire n_1189;
wire n_1079;
wire n_1212;
wire n_828;
wire n_462;
wire n_1033;
wire n_607;
wire n_671;
wire n_726;
wire n_1052;
wire n_419;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_703;
wire n_578;
wire n_1003;
wire n_978;
wire n_1061;
wire n_595;
wire n_627;
wire n_1203;
wire n_524;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_751;
wire n_449;
wire n_749;
wire n_1208;
wire n_798;
wire n_1164;
wire n_509;
wire n_1209;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_1151;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_1100;
wire n_1214;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_1128;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_1204;
wire n_1160;
wire n_883;
wire n_823;
wire n_557;
wire n_1132;
wire n_643;
wire n_898;
wire n_617;
wire n_698;
wire n_1074;
wire n_1032;
wire n_845;
wire n_807;
wire n_1036;
wire n_739;
wire n_400;
wire n_955;
wire n_865;
wire n_1138;
wire n_893;
wire n_925;
wire n_485;
wire n_1099;
wire n_1026;
wire n_443;
wire n_1101;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_935;
wire n_1192;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_1130;
wire n_1127;
wire n_1095;
wire n_573;
wire n_769;
wire n_639;
wire n_676;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_1120;
wire n_685;
wire n_597;
wire n_832;
wire n_1187;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_605;
wire n_461;
wire n_873;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_1139;
wire n_718;
wire n_517;
wire n_1018;
wire n_1172;
wire n_747;
wire n_852;
wire n_667;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_1206;
wire n_621;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_691;
wire n_535;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_1140;
wire n_413;
wire n_1196;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_601;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1057;
wire n_1147;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_1143;
wire n_536;
wire n_895;
wire n_1126;
wire n_866;
wire n_622;
wire n_710;
wire n_1108;
wire n_387;
wire n_1182;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_1119;
wire n_761;
wire n_428;
wire n_581;
wire n_785;
wire n_746;
wire n_1205;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_720;
wire n_758;
wire n_516;
wire n_842;
wire n_525;
wire n_1163;
wire n_1173;
wire n_1180;
wire n_1116;
wire n_611;
wire n_943;
wire n_1168;
wire n_491;
wire n_843;
wire n_656;
wire n_772;
wire n_989;
wire n_1174;
wire n_797;
wire n_666;
wire n_1016;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_1035;
wire n_838;
wire n_499;
wire n_705;
wire n_647;
wire n_844;
wire n_448;
wire n_886;
wire n_1017;
wire n_1004;
wire n_953;
wire n_1094;
wire n_1176;
wire n_1190;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_1112;
wire n_454;
wire n_1213;
wire n_638;
wire n_1181;
wire n_910;
wire n_1211;
wire n_486;
wire n_911;
wire n_947;
wire n_653;
wire n_887;
wire n_1117;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_809;
wire n_1043;
wire n_1011;
wire n_926;
wire n_927;
wire n_1215;
wire n_986;
wire n_839;
wire n_734;
wire n_1088;
wire n_708;
wire n_919;
wire n_1081;
wire n_402;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_800;
wire n_779;
wire n_574;
wire n_929;
wire n_460;
wire n_1084;
wire n_1171;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_1122;
wire n_870;
wire n_659;
wire n_709;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_526;
wire n_1109;
wire n_921;
wire n_712;
wire n_1183;
wire n_711;
wire n_579;
wire n_937;
wire n_390;
wire n_473;
wire n_1193;
wire n_1148;
wire n_1054;
wire n_559;
wire n_1161;
wire n_458;
wire n_1070;
wire n_1085;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_1145;
wire n_771;
wire n_1121;
wire n_1152;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_492;
wire n_972;
wire n_699;
wire n_551;
wire n_456;
wire n_1149;
wire n_564;
wire n_1178;
wire n_624;
wire n_451;
wire n_1184;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_686;
wire n_796;
wire n_1041;
wire n_757;
wire n_594;
wire n_719;
wire n_565;
wire n_1195;
wire n_577;
wire n_936;
wire n_552;
wire n_1186;
wire n_1062;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_829;
wire n_1156;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_1142;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_1123;
wire n_884;
wire n_1201;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_645;
wire n_916;
wire n_1078;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_934;
wire n_482;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_608;
wire n_683;
wire n_527;
wire n_620;
wire n_420;
wire n_630;
wire n_394;
wire n_878;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_469;
wire n_1137;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_543;
wire n_1144;
wire n_889;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_1162;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_600;
wire n_464;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_1198;
wire n_584;
wire n_1110;
wire n_399;
wire n_979;
wire n_548;
wire n_905;
wire n_436;
wire n_833;
wire n_523;
wire n_707;
wire n_993;
wire n_689;
wire n_409;
wire n_799;
wire n_505;
wire n_1155;
wire n_756;
wire n_547;
wire n_537;
wire n_558;
wire n_810;
wire n_1133;
wire n_635;
wire n_787;
wire n_1194;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_1141;
wire n_1146;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_1158;
wire n_754;
wire n_1136;
wire n_941;
wire n_975;
wire n_1031;
wire n_550;
wire n_487;
wire n_1125;
wire n_652;
wire n_849;
wire n_553;
wire n_970;
wire n_1107;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_1159;
wire n_569;
wire n_1092;
wire n_441;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_1207;
wire n_1111;
wire n_511;
wire n_715;
wire n_467;
wire n_973;
wire n_416;
wire n_1053;
wire n_530;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_1106;
wire n_582;
wire n_1167;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_651;
wire n_404;
wire n_439;
wire n_1153;
wire n_518;
wire n_1210;
wire n_679;
wire n_1069;
wire n_1185;
wire n_612;
wire n_453;
wire n_633;
wire n_1170;
wire n_665;
wire n_902;
wire n_588;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_1165;
wire n_426;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_1166;
wire n_431;
wire n_812;
wire n_459;
wire n_1131;
wire n_502;
wire n_1175;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_1012;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_834;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1089;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_766;
wire n_743;
wire n_816;
wire n_1157;
wire n_430;
wire n_1002;
wire n_463;
wire n_1188;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_1019;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_438;
wire n_1124;
wire n_784;
wire n_515;
wire n_434;
wire n_983;
wire n_427;
wire n_1200;
wire n_1059;
wire n_1197;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_869;
wire n_1154;
wire n_437;
wire n_1082;
wire n_1113;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_1098;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_960;
wire n_956;
wire n_827;
wire n_531;
wire n_1001;
wire n_663;
wire n_508;
wire n_856;
wire n_1050;
wire n_778;
wire n_1025;
wire n_1134;
wire n_1177;
wire n_891;
wire n_1150;
wire n_398;
wire n_410;
wire n_1129;
wire n_1191;
wire n_566;
wire n_554;
wire n_602;
wire n_1023;
wire n_1013;
wire n_1076;
wire n_1118;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;

INVx1_ASAP7_75t_L g387 ( 
.A(n_111),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g388 ( 
.A(n_373),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_11),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_91),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_280),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_315),
.Y(n_392)
);

CKINVDCx14_ASAP7_75t_R g393 ( 
.A(n_367),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_335),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_381),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_249),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_259),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_192),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_245),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_326),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_329),
.Y(n_401)
);

BUFx2_ASAP7_75t_SL g402 ( 
.A(n_141),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_99),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_352),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_289),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_274),
.Y(n_406)
);

BUFx10_ASAP7_75t_L g407 ( 
.A(n_59),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_152),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_65),
.Y(n_409)
);

INVx1_ASAP7_75t_SL g410 ( 
.A(n_231),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_382),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_212),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_328),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_286),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_324),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_133),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_268),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_140),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_278),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_333),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_386),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_331),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_308),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_380),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_309),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_338),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_139),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_68),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_385),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_287),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_251),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_258),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_83),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_208),
.Y(n_434)
);

BUFx5_ASAP7_75t_L g435 ( 
.A(n_64),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_108),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_240),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_168),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_137),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_237),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_242),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_158),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_248),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_250),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_119),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_125),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_246),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_307),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_127),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_216),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_155),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_55),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_58),
.Y(n_453)
);

BUFx5_ASAP7_75t_L g454 ( 
.A(n_304),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_285),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_342),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_383),
.Y(n_457)
);

BUFx10_ASAP7_75t_L g458 ( 
.A(n_164),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_273),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_37),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_277),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_67),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_205),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_379),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_2),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_359),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_265),
.Y(n_467)
);

BUFx6f_ASAP7_75t_L g468 ( 
.A(n_196),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_305),
.Y(n_469)
);

INVx2_ASAP7_75t_SL g470 ( 
.A(n_377),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_43),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_330),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_244),
.Y(n_473)
);

CKINVDCx16_ASAP7_75t_R g474 ( 
.A(n_106),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_130),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_371),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_225),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_115),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_255),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_108),
.Y(n_480)
);

INVx1_ASAP7_75t_SL g481 ( 
.A(n_166),
.Y(n_481)
);

BUFx2_ASAP7_75t_L g482 ( 
.A(n_83),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_51),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_332),
.Y(n_484)
);

INVx2_ASAP7_75t_SL g485 ( 
.A(n_368),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_220),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_219),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_150),
.Y(n_488)
);

BUFx5_ASAP7_75t_L g489 ( 
.A(n_197),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_306),
.Y(n_490)
);

CKINVDCx16_ASAP7_75t_R g491 ( 
.A(n_365),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_366),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_213),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_238),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_316),
.Y(n_495)
);

BUFx10_ASAP7_75t_L g496 ( 
.A(n_131),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_122),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_294),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_378),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_295),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_193),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_296),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_61),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_90),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_87),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_63),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_33),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_370),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_88),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_228),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_247),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_170),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_136),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_110),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_301),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_214),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_72),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_18),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_375),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_120),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_269),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_354),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_256),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_356),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_185),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_310),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_116),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_303),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_257),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_369),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_243),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_293),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_227),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_267),
.Y(n_534)
);

BUFx2_ASAP7_75t_SL g535 ( 
.A(n_337),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_291),
.Y(n_536)
);

BUFx2_ASAP7_75t_L g537 ( 
.A(n_345),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_229),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_148),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_26),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_71),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_126),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_142),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_173),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_25),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_226),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_167),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_343),
.Y(n_548)
);

CKINVDCx16_ASAP7_75t_R g549 ( 
.A(n_46),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_112),
.Y(n_550)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_239),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_384),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_172),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_361),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_106),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_151),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_49),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_28),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_372),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g560 ( 
.A(n_241),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_145),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_36),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_374),
.Y(n_563)
);

INVxp67_ASAP7_75t_L g564 ( 
.A(n_147),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_49),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_92),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_175),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_138),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_190),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_376),
.Y(n_570)
);

BUFx5_ASAP7_75t_L g571 ( 
.A(n_191),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_143),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_38),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_255),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_178),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_109),
.Y(n_576)
);

BUFx5_ASAP7_75t_L g577 ( 
.A(n_320),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_327),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_254),
.Y(n_579)
);

CKINVDCx20_ASAP7_75t_R g580 ( 
.A(n_314),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_206),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_166),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_73),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_14),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_253),
.Y(n_585)
);

BUFx2_ASAP7_75t_L g586 ( 
.A(n_17),
.Y(n_586)
);

BUFx10_ASAP7_75t_L g587 ( 
.A(n_252),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_132),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_134),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_2),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_172),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_79),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_74),
.Y(n_593)
);

BUFx2_ASAP7_75t_L g594 ( 
.A(n_358),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_288),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_189),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_321),
.Y(n_597)
);

CKINVDCx20_ASAP7_75t_R g598 ( 
.A(n_102),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_216),
.Y(n_599)
);

INVxp67_ASAP7_75t_L g600 ( 
.A(n_482),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_537),
.B(n_1),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_422),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_391),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_392),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_394),
.Y(n_605)
);

INVxp67_ASAP7_75t_SL g606 ( 
.A(n_424),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_395),
.Y(n_607)
);

CKINVDCx20_ASAP7_75t_R g608 ( 
.A(n_426),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_435),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_405),
.Y(n_610)
);

CKINVDCx20_ASAP7_75t_R g611 ( 
.A(n_429),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_406),
.Y(n_612)
);

HB1xp67_ASAP7_75t_L g613 ( 
.A(n_474),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_435),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g615 ( 
.A(n_495),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_489),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_489),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_489),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_571),
.Y(n_619)
);

INVxp67_ASAP7_75t_SL g620 ( 
.A(n_528),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_411),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_571),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_571),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_413),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_414),
.Y(n_625)
);

NAND2xp33_ASAP7_75t_R g626 ( 
.A(n_594),
.B(n_0),
.Y(n_626)
);

INVxp33_ASAP7_75t_L g627 ( 
.A(n_586),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_444),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_415),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_417),
.Y(n_630)
);

CKINVDCx16_ASAP7_75t_R g631 ( 
.A(n_549),
.Y(n_631)
);

HB1xp67_ASAP7_75t_L g632 ( 
.A(n_387),
.Y(n_632)
);

INVxp67_ASAP7_75t_L g633 ( 
.A(n_407),
.Y(n_633)
);

INVxp67_ASAP7_75t_SL g634 ( 
.A(n_388),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_420),
.Y(n_635)
);

INVxp67_ASAP7_75t_L g636 ( 
.A(n_407),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_423),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_468),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_638),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_628),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_634),
.B(n_393),
.Y(n_641)
);

BUFx2_ASAP7_75t_L g642 ( 
.A(n_613),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_606),
.B(n_408),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_622),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_620),
.B(n_469),
.Y(n_645)
);

INVxp67_ASAP7_75t_L g646 ( 
.A(n_632),
.Y(n_646)
);

NAND2xp33_ASAP7_75t_SL g647 ( 
.A(n_626),
.B(n_497),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_609),
.Y(n_648)
);

INVx3_ASAP7_75t_L g649 ( 
.A(n_614),
.Y(n_649)
);

BUFx8_ASAP7_75t_L g650 ( 
.A(n_616),
.Y(n_650)
);

INVxp67_ASAP7_75t_L g651 ( 
.A(n_632),
.Y(n_651)
);

BUFx6f_ASAP7_75t_L g652 ( 
.A(n_617),
.Y(n_652)
);

INVx4_ASAP7_75t_L g653 ( 
.A(n_603),
.Y(n_653)
);

INVx3_ASAP7_75t_L g654 ( 
.A(n_618),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_619),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_623),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_600),
.B(n_428),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_604),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_605),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_607),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_601),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_610),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_612),
.Y(n_663)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_621),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_624),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_625),
.B(n_491),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_629),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_630),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_635),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_637),
.B(n_450),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_633),
.Y(n_671)
);

INVxp67_ASAP7_75t_L g672 ( 
.A(n_636),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_627),
.Y(n_673)
);

AND2x6_ASAP7_75t_L g674 ( 
.A(n_663),
.B(n_400),
.Y(n_674)
);

BUFx3_ASAP7_75t_L g675 ( 
.A(n_664),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_652),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_661),
.B(n_631),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_639),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_644),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_641),
.B(n_470),
.Y(n_680)
);

BUFx3_ASAP7_75t_L g681 ( 
.A(n_664),
.Y(n_681)
);

INVx5_ASAP7_75t_L g682 ( 
.A(n_658),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_673),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_641),
.B(n_485),
.Y(n_684)
);

NAND2xp33_ASAP7_75t_SL g685 ( 
.A(n_661),
.B(n_398),
.Y(n_685)
);

INVx4_ASAP7_75t_L g686 ( 
.A(n_665),
.Y(n_686)
);

INVx4_ASAP7_75t_L g687 ( 
.A(n_652),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_666),
.B(n_659),
.Y(n_688)
);

OR2x6_ASAP7_75t_L g689 ( 
.A(n_642),
.B(n_402),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_640),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_655),
.Y(n_691)
);

BUFx3_ASAP7_75t_L g692 ( 
.A(n_649),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_656),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_660),
.B(n_602),
.Y(n_694)
);

AND2x4_ASAP7_75t_L g695 ( 
.A(n_670),
.B(n_580),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_653),
.Y(n_696)
);

OR2x2_ASAP7_75t_L g697 ( 
.A(n_646),
.B(n_410),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_662),
.B(n_608),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g699 ( 
.A(n_648),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_654),
.Y(n_700)
);

AND2x4_ASAP7_75t_L g701 ( 
.A(n_645),
.B(n_437),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_671),
.B(n_430),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_643),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_657),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_667),
.B(n_611),
.Y(n_705)
);

BUFx3_ASAP7_75t_L g706 ( 
.A(n_650),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_657),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_669),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_668),
.Y(n_709)
);

OR2x2_ASAP7_75t_L g710 ( 
.A(n_651),
.B(n_647),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_672),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_665),
.Y(n_712)
);

OR2x2_ASAP7_75t_L g713 ( 
.A(n_673),
.B(n_481),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_678),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_688),
.B(n_691),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_693),
.B(n_401),
.Y(n_716)
);

A2O1A1Ixp33_ASAP7_75t_L g717 ( 
.A1(n_703),
.A2(n_419),
.B(n_421),
.C(n_404),
.Y(n_717)
);

OR2x6_ASAP7_75t_L g718 ( 
.A(n_675),
.B(n_535),
.Y(n_718)
);

NAND2x1p5_ASAP7_75t_L g719 ( 
.A(n_681),
.B(n_425),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_682),
.B(n_615),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_680),
.B(n_459),
.Y(n_721)
);

OAI221xp5_ASAP7_75t_L g722 ( 
.A1(n_707),
.A2(n_564),
.B1(n_475),
.B2(n_399),
.C(n_403),
.Y(n_722)
);

NAND2x1p5_ASAP7_75t_L g723 ( 
.A(n_682),
.B(n_464),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_704),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_683),
.Y(n_725)
);

INVxp67_ASAP7_75t_L g726 ( 
.A(n_713),
.Y(n_726)
);

AO22x2_ASAP7_75t_L g727 ( 
.A1(n_710),
.A2(n_440),
.B1(n_483),
.B2(n_431),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_684),
.B(n_466),
.Y(n_728)
);

BUFx3_ASAP7_75t_L g729 ( 
.A(n_692),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_712),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_699),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_708),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_700),
.Y(n_733)
);

NAND2x1p5_ASAP7_75t_L g734 ( 
.A(n_686),
.B(n_476),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_699),
.Y(n_735)
);

BUFx8_ASAP7_75t_L g736 ( 
.A(n_711),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_676),
.Y(n_737)
);

AO22x2_ASAP7_75t_L g738 ( 
.A1(n_695),
.A2(n_473),
.B1(n_503),
.B2(n_451),
.Y(n_738)
);

INVx4_ASAP7_75t_L g739 ( 
.A(n_690),
.Y(n_739)
);

AO22x2_ASAP7_75t_L g740 ( 
.A1(n_677),
.A2(n_477),
.B1(n_517),
.B2(n_438),
.Y(n_740)
);

AND2x4_ASAP7_75t_L g741 ( 
.A(n_701),
.B(n_709),
.Y(n_741)
);

AND2x4_ASAP7_75t_L g742 ( 
.A(n_689),
.B(n_501),
.Y(n_742)
);

NAND2x1p5_ASAP7_75t_L g743 ( 
.A(n_687),
.B(n_498),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_689),
.B(n_458),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_694),
.B(n_698),
.Y(n_745)
);

AO22x2_ASAP7_75t_L g746 ( 
.A1(n_685),
.A2(n_436),
.B1(n_465),
.B2(n_418),
.Y(n_746)
);

NAND2x1p5_ASAP7_75t_L g747 ( 
.A(n_702),
.B(n_502),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_674),
.Y(n_748)
);

AO22x2_ASAP7_75t_L g749 ( 
.A1(n_705),
.A2(n_523),
.B1(n_541),
.B2(n_513),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_674),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_674),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_696),
.B(n_389),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_679),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_678),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_679),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_678),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_688),
.B(n_519),
.Y(n_757)
);

AND2x4_ASAP7_75t_L g758 ( 
.A(n_675),
.B(n_520),
.Y(n_758)
);

NAND2x1p5_ASAP7_75t_L g759 ( 
.A(n_675),
.B(n_521),
.Y(n_759)
);

HB1xp67_ASAP7_75t_L g760 ( 
.A(n_695),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_688),
.A2(n_455),
.B1(n_457),
.B2(n_456),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_678),
.Y(n_762)
);

AND2x6_ASAP7_75t_L g763 ( 
.A(n_708),
.B(n_524),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_682),
.B(n_467),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_678),
.Y(n_765)
);

INVxp67_ASAP7_75t_L g766 ( 
.A(n_697),
.Y(n_766)
);

OAI221xp5_ASAP7_75t_L g767 ( 
.A1(n_703),
.A2(n_486),
.B1(n_518),
.B2(n_510),
.C(n_505),
.Y(n_767)
);

NAND2xp33_ASAP7_75t_L g768 ( 
.A(n_708),
.B(n_472),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_688),
.B(n_526),
.Y(n_769)
);

BUFx6f_ASAP7_75t_SL g770 ( 
.A(n_706),
.Y(n_770)
);

NAND2x1p5_ASAP7_75t_L g771 ( 
.A(n_675),
.B(n_530),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_688),
.B(n_390),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_675),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_679),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_678),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_678),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_745),
.B(n_496),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_772),
.B(n_532),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_766),
.B(n_725),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_757),
.B(n_534),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_769),
.B(n_490),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_724),
.B(n_492),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_752),
.B(n_499),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_773),
.B(n_500),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_741),
.B(n_508),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_721),
.B(n_552),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_728),
.B(n_554),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_732),
.B(n_515),
.Y(n_788)
);

NAND2xp33_ASAP7_75t_SL g789 ( 
.A(n_760),
.B(n_445),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_761),
.B(n_522),
.Y(n_790)
);

NAND2xp33_ASAP7_75t_SL g791 ( 
.A(n_739),
.B(n_478),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_734),
.B(n_536),
.Y(n_792)
);

NAND2xp33_ASAP7_75t_SL g793 ( 
.A(n_748),
.B(n_488),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_753),
.B(n_559),
.Y(n_794)
);

NAND2xp33_ASAP7_75t_SL g795 ( 
.A(n_750),
.B(n_507),
.Y(n_795)
);

NAND2xp33_ASAP7_75t_SL g796 ( 
.A(n_751),
.B(n_525),
.Y(n_796)
);

NAND2xp33_ASAP7_75t_SL g797 ( 
.A(n_744),
.B(n_527),
.Y(n_797)
);

NAND2xp33_ASAP7_75t_SL g798 ( 
.A(n_720),
.B(n_544),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_755),
.B(n_774),
.Y(n_799)
);

NAND2xp33_ASAP7_75t_SL g800 ( 
.A(n_733),
.B(n_764),
.Y(n_800)
);

AND2x4_ASAP7_75t_L g801 ( 
.A(n_735),
.B(n_540),
.Y(n_801)
);

NAND2xp33_ASAP7_75t_SL g802 ( 
.A(n_770),
.B(n_551),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_714),
.B(n_563),
.Y(n_803)
);

NAND2xp33_ASAP7_75t_SL g804 ( 
.A(n_737),
.B(n_582),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_754),
.B(n_776),
.Y(n_805)
);

NAND2xp33_ASAP7_75t_SL g806 ( 
.A(n_716),
.B(n_742),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_756),
.B(n_570),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_762),
.B(n_578),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_765),
.B(n_775),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_747),
.B(n_758),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_729),
.B(n_448),
.Y(n_811)
);

NOR2x1_ASAP7_75t_L g812 ( 
.A(n_718),
.B(n_768),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_740),
.B(n_746),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_736),
.B(n_461),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_743),
.B(n_461),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_727),
.B(n_763),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_SL g817 ( 
.A(n_719),
.B(n_461),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_771),
.B(n_484),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_759),
.B(n_484),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_723),
.B(n_484),
.Y(n_820)
);

NAND2xp33_ASAP7_75t_SL g821 ( 
.A(n_738),
.B(n_598),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_717),
.B(n_548),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_749),
.B(n_595),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_722),
.B(n_597),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_767),
.B(n_454),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_715),
.B(n_454),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_726),
.B(n_587),
.Y(n_827)
);

NAND2xp33_ASAP7_75t_SL g828 ( 
.A(n_730),
.B(n_396),
.Y(n_828)
);

NAND2xp33_ASAP7_75t_SL g829 ( 
.A(n_730),
.B(n_397),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_772),
.B(n_577),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_715),
.B(n_512),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_715),
.B(n_550),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_772),
.B(n_550),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_715),
.B(n_560),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_715),
.B(n_560),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_715),
.B(n_560),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_715),
.B(n_409),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_772),
.B(n_412),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_715),
.B(n_416),
.Y(n_839)
);

NAND2xp33_ASAP7_75t_SL g840 ( 
.A(n_730),
.B(n_427),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_715),
.B(n_432),
.Y(n_841)
);

NAND2xp33_ASAP7_75t_SL g842 ( 
.A(n_730),
.B(n_433),
.Y(n_842)
);

NAND2xp33_ASAP7_75t_SL g843 ( 
.A(n_730),
.B(n_434),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_715),
.B(n_439),
.Y(n_844)
);

NAND2xp33_ASAP7_75t_SL g845 ( 
.A(n_730),
.B(n_441),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_715),
.B(n_442),
.Y(n_846)
);

NAND2xp33_ASAP7_75t_SL g847 ( 
.A(n_730),
.B(n_443),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_715),
.B(n_446),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_772),
.B(n_447),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_715),
.B(n_449),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_715),
.B(n_452),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_715),
.B(n_453),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_715),
.B(n_460),
.Y(n_853)
);

AND2x4_ASAP7_75t_L g854 ( 
.A(n_731),
.B(n_546),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_715),
.B(n_462),
.Y(n_855)
);

A2O1A1Ixp33_ASAP7_75t_L g856 ( 
.A1(n_778),
.A2(n_561),
.B(n_565),
.C(n_558),
.Y(n_856)
);

A2O1A1Ixp33_ASAP7_75t_L g857 ( 
.A1(n_838),
.A2(n_579),
.B(n_581),
.C(n_576),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_854),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_849),
.B(n_471),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_801),
.Y(n_860)
);

AO31x2_ASAP7_75t_L g861 ( 
.A1(n_830),
.A2(n_591),
.A3(n_592),
.B(n_583),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_801),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_799),
.Y(n_863)
);

OAI21xp33_ASAP7_75t_L g864 ( 
.A1(n_777),
.A2(n_480),
.B(n_479),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_826),
.A2(n_593),
.B(n_463),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_780),
.B(n_833),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_805),
.Y(n_867)
);

A2O1A1Ixp33_ASAP7_75t_L g868 ( 
.A1(n_813),
.A2(n_806),
.B(n_800),
.C(n_795),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_837),
.B(n_487),
.Y(n_869)
);

AOI221xp5_ASAP7_75t_L g870 ( 
.A1(n_821),
.A2(n_798),
.B1(n_797),
.B2(n_804),
.C(n_789),
.Y(n_870)
);

O2A1O1Ixp5_ASAP7_75t_SL g871 ( 
.A1(n_823),
.A2(n_831),
.B(n_834),
.C(n_832),
.Y(n_871)
);

BUFx10_ASAP7_75t_L g872 ( 
.A(n_828),
.Y(n_872)
);

AND3x4_ASAP7_75t_L g873 ( 
.A(n_812),
.B(n_567),
.C(n_562),
.Y(n_873)
);

A2O1A1Ixp33_ASAP7_75t_L g874 ( 
.A1(n_793),
.A2(n_572),
.B(n_589),
.C(n_568),
.Y(n_874)
);

OAI21x1_ASAP7_75t_L g875 ( 
.A1(n_809),
.A2(n_261),
.B(n_260),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_825),
.Y(n_876)
);

NAND3x1_ASAP7_75t_L g877 ( 
.A(n_816),
.B(n_494),
.C(n_493),
.Y(n_877)
);

OAI22xp5_ASAP7_75t_L g878 ( 
.A1(n_839),
.A2(n_506),
.B1(n_509),
.B2(n_504),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_810),
.A2(n_263),
.B(n_262),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_796),
.B(n_511),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_782),
.A2(n_266),
.B(n_264),
.Y(n_881)
);

NAND3xp33_ASAP7_75t_L g882 ( 
.A(n_829),
.B(n_516),
.C(n_514),
.Y(n_882)
);

INVx8_ASAP7_75t_L g883 ( 
.A(n_827),
.Y(n_883)
);

AO31x2_ASAP7_75t_L g884 ( 
.A1(n_786),
.A2(n_271),
.A3(n_272),
.B(n_270),
.Y(n_884)
);

OAI22xp5_ASAP7_75t_L g885 ( 
.A1(n_841),
.A2(n_531),
.B1(n_533),
.B2(n_529),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_787),
.Y(n_886)
);

HB1xp67_ASAP7_75t_L g887 ( 
.A(n_779),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_844),
.B(n_538),
.Y(n_888)
);

OR2x2_ASAP7_75t_L g889 ( 
.A(n_846),
.B(n_539),
.Y(n_889)
);

A2O1A1Ixp33_ASAP7_75t_L g890 ( 
.A1(n_848),
.A2(n_543),
.B(n_545),
.C(n_542),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_850),
.B(n_547),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_794),
.A2(n_276),
.B(n_275),
.Y(n_892)
);

INVx4_ASAP7_75t_L g893 ( 
.A(n_791),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_851),
.B(n_553),
.Y(n_894)
);

OAI22xp5_ASAP7_75t_L g895 ( 
.A1(n_852),
.A2(n_556),
.B1(n_557),
.B2(n_555),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_814),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_853),
.B(n_566),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_855),
.B(n_569),
.Y(n_898)
);

OAI21x1_ASAP7_75t_L g899 ( 
.A1(n_788),
.A2(n_281),
.B(n_279),
.Y(n_899)
);

O2A1O1Ixp5_ASAP7_75t_SL g900 ( 
.A1(n_835),
.A2(n_599),
.B(n_596),
.C(n_574),
.Y(n_900)
);

AND3x4_ASAP7_75t_L g901 ( 
.A(n_802),
.B(n_575),
.C(n_573),
.Y(n_901)
);

OAI21x1_ASAP7_75t_L g902 ( 
.A1(n_803),
.A2(n_283),
.B(n_282),
.Y(n_902)
);

AND2x4_ASAP7_75t_L g903 ( 
.A(n_785),
.B(n_284),
.Y(n_903)
);

OAI22xp5_ASAP7_75t_L g904 ( 
.A1(n_781),
.A2(n_585),
.B1(n_588),
.B2(n_584),
.Y(n_904)
);

AOI21x1_ASAP7_75t_L g905 ( 
.A1(n_807),
.A2(n_292),
.B(n_290),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_783),
.B(n_590),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_836),
.Y(n_907)
);

AO31x2_ASAP7_75t_L g908 ( 
.A1(n_822),
.A2(n_298),
.A3(n_299),
.B(n_297),
.Y(n_908)
);

OAI21x1_ASAP7_75t_L g909 ( 
.A1(n_808),
.A2(n_302),
.B(n_300),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_824),
.Y(n_910)
);

INVx1_ASAP7_75t_SL g911 ( 
.A(n_840),
.Y(n_911)
);

AOI21xp33_ASAP7_75t_L g912 ( 
.A1(n_790),
.A2(n_3),
.B(n_4),
.Y(n_912)
);

OAI21x1_ASAP7_75t_L g913 ( 
.A1(n_784),
.A2(n_312),
.B(n_311),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_866),
.A2(n_792),
.B(n_815),
.Y(n_914)
);

O2A1O1Ixp33_ASAP7_75t_SL g915 ( 
.A1(n_868),
.A2(n_811),
.B(n_820),
.C(n_818),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_867),
.Y(n_916)
);

OAI21x1_ASAP7_75t_L g917 ( 
.A1(n_875),
.A2(n_819),
.B(n_817),
.Y(n_917)
);

INVx3_ASAP7_75t_L g918 ( 
.A(n_883),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_859),
.B(n_842),
.Y(n_919)
);

AO22x1_ASAP7_75t_L g920 ( 
.A1(n_873),
.A2(n_845),
.B1(n_847),
.B2(n_843),
.Y(n_920)
);

INVxp67_ASAP7_75t_L g921 ( 
.A(n_887),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_886),
.Y(n_922)
);

AND2x6_ASAP7_75t_L g923 ( 
.A(n_903),
.B(n_313),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_872),
.Y(n_924)
);

OAI221xp5_ASAP7_75t_L g925 ( 
.A1(n_870),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.C(n_8),
.Y(n_925)
);

OAI21xp5_ASAP7_75t_L g926 ( 
.A1(n_871),
.A2(n_876),
.B(n_900),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_860),
.B(n_317),
.Y(n_927)
);

NOR3xp33_ASAP7_75t_L g928 ( 
.A(n_893),
.B(n_9),
.C(n_10),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_858),
.Y(n_929)
);

OAI21x1_ASAP7_75t_L g930 ( 
.A1(n_899),
.A2(n_319),
.B(n_318),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_862),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_910),
.Y(n_932)
);

OAI21x1_ASAP7_75t_L g933 ( 
.A1(n_902),
.A2(n_323),
.B(n_322),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_896),
.Y(n_934)
);

OR2x6_ASAP7_75t_L g935 ( 
.A(n_879),
.B(n_325),
.Y(n_935)
);

BUFx2_ASAP7_75t_SL g936 ( 
.A(n_911),
.Y(n_936)
);

HB1xp67_ASAP7_75t_L g937 ( 
.A(n_907),
.Y(n_937)
);

INVx3_ASAP7_75t_L g938 ( 
.A(n_877),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_861),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_856),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_864),
.B(n_12),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_865),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_905),
.Y(n_943)
);

BUFx12f_ASAP7_75t_L g944 ( 
.A(n_889),
.Y(n_944)
);

OA21x2_ASAP7_75t_L g945 ( 
.A1(n_909),
.A2(n_336),
.B(n_334),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_857),
.Y(n_946)
);

OR2x2_ASAP7_75t_L g947 ( 
.A(n_869),
.B(n_13),
.Y(n_947)
);

CKINVDCx16_ASAP7_75t_R g948 ( 
.A(n_891),
.Y(n_948)
);

AO32x2_ASAP7_75t_L g949 ( 
.A1(n_878),
.A2(n_895),
.A3(n_885),
.B1(n_904),
.B2(n_912),
.Y(n_949)
);

BUFx6f_ASAP7_75t_L g950 ( 
.A(n_913),
.Y(n_950)
);

CKINVDCx8_ASAP7_75t_R g951 ( 
.A(n_901),
.Y(n_951)
);

AND2x4_ASAP7_75t_L g952 ( 
.A(n_880),
.B(n_339),
.Y(n_952)
);

OAI21x1_ASAP7_75t_L g953 ( 
.A1(n_892),
.A2(n_341),
.B(n_340),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_906),
.B(n_15),
.Y(n_954)
);

BUFx6f_ASAP7_75t_SL g955 ( 
.A(n_874),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_882),
.B(n_344),
.Y(n_956)
);

OA21x2_ASAP7_75t_L g957 ( 
.A1(n_881),
.A2(n_347),
.B(n_346),
.Y(n_957)
);

AOI21x1_ASAP7_75t_L g958 ( 
.A1(n_888),
.A2(n_349),
.B(n_348),
.Y(n_958)
);

OAI21x1_ASAP7_75t_L g959 ( 
.A1(n_894),
.A2(n_351),
.B(n_350),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_897),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_898),
.B(n_16),
.Y(n_961)
);

BUFx4f_ASAP7_75t_SL g962 ( 
.A(n_884),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_908),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_890),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_863),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_922),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_916),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_965),
.Y(n_968)
);

OA21x2_ASAP7_75t_L g969 ( 
.A1(n_926),
.A2(n_355),
.B(n_353),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_924),
.Y(n_970)
);

INVx4_ASAP7_75t_L g971 ( 
.A(n_934),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_934),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_929),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_932),
.Y(n_974)
);

BUFx3_ASAP7_75t_L g975 ( 
.A(n_918),
.Y(n_975)
);

OR2x6_ASAP7_75t_L g976 ( 
.A(n_936),
.B(n_357),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_931),
.Y(n_977)
);

HB1xp67_ASAP7_75t_L g978 ( 
.A(n_921),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_937),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_939),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_940),
.Y(n_981)
);

INVx3_ASAP7_75t_L g982 ( 
.A(n_944),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_942),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_961),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_954),
.Y(n_985)
);

A2O1A1Ixp33_ASAP7_75t_L g986 ( 
.A1(n_919),
.A2(n_21),
.B(n_19),
.C(n_20),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_927),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_946),
.Y(n_988)
);

BUFx4f_ASAP7_75t_L g989 ( 
.A(n_923),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_949),
.B(n_360),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_960),
.B(n_21),
.Y(n_991)
);

AOI22xp33_ASAP7_75t_L g992 ( 
.A1(n_941),
.A2(n_24),
.B1(n_22),
.B2(n_23),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_947),
.Y(n_993)
);

INVx6_ASAP7_75t_L g994 ( 
.A(n_948),
.Y(n_994)
);

INVx4_ASAP7_75t_L g995 ( 
.A(n_923),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_943),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_964),
.Y(n_997)
);

INVx3_ASAP7_75t_L g998 ( 
.A(n_951),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_958),
.Y(n_999)
);

BUFx2_ASAP7_75t_SL g1000 ( 
.A(n_955),
.Y(n_1000)
);

AO21x2_ASAP7_75t_L g1001 ( 
.A1(n_963),
.A2(n_363),
.B(n_362),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_R g1002 ( 
.A(n_970),
.B(n_998),
.Y(n_1002)
);

NAND2xp33_ASAP7_75t_R g1003 ( 
.A(n_982),
.B(n_956),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_984),
.B(n_985),
.Y(n_1004)
);

BUFx3_ASAP7_75t_L g1005 ( 
.A(n_972),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_980),
.Y(n_1006)
);

NAND2xp33_ASAP7_75t_R g1007 ( 
.A(n_976),
.B(n_938),
.Y(n_1007)
);

AND2x4_ASAP7_75t_L g1008 ( 
.A(n_995),
.B(n_952),
.Y(n_1008)
);

BUFx3_ASAP7_75t_L g1009 ( 
.A(n_972),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_R g1010 ( 
.A(n_989),
.B(n_962),
.Y(n_1010)
);

XNOR2xp5_ASAP7_75t_L g1011 ( 
.A(n_1000),
.B(n_920),
.Y(n_1011)
);

INVxp67_ASAP7_75t_L g1012 ( 
.A(n_978),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_979),
.B(n_959),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_993),
.B(n_928),
.Y(n_1014)
);

BUFx10_ASAP7_75t_L g1015 ( 
.A(n_994),
.Y(n_1015)
);

BUFx3_ASAP7_75t_L g1016 ( 
.A(n_975),
.Y(n_1016)
);

AND2x4_ASAP7_75t_L g1017 ( 
.A(n_987),
.B(n_935),
.Y(n_1017)
);

AND2x4_ASAP7_75t_L g1018 ( 
.A(n_973),
.B(n_935),
.Y(n_1018)
);

BUFx3_ASAP7_75t_L g1019 ( 
.A(n_971),
.Y(n_1019)
);

NAND2xp33_ASAP7_75t_R g1020 ( 
.A(n_990),
.B(n_945),
.Y(n_1020)
);

NAND2xp33_ASAP7_75t_R g1021 ( 
.A(n_990),
.B(n_957),
.Y(n_1021)
);

AND2x4_ASAP7_75t_L g1022 ( 
.A(n_977),
.B(n_950),
.Y(n_1022)
);

BUFx2_ASAP7_75t_L g1023 ( 
.A(n_997),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_1006),
.Y(n_1024)
);

OAI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_1011),
.A2(n_992),
.B1(n_925),
.B2(n_986),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_1022),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_1023),
.B(n_967),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_1012),
.B(n_974),
.Y(n_1028)
);

NAND2x1_ASAP7_75t_L g1029 ( 
.A(n_1013),
.B(n_983),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_1002),
.Y(n_1030)
);

AND2x4_ASAP7_75t_SL g1031 ( 
.A(n_1015),
.B(n_966),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_1004),
.B(n_968),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_1014),
.B(n_991),
.Y(n_1033)
);

AND2x4_ASAP7_75t_L g1034 ( 
.A(n_1018),
.B(n_996),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_1017),
.Y(n_1035)
);

INVx3_ASAP7_75t_L g1036 ( 
.A(n_1008),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_1005),
.Y(n_1037)
);

AND2x2_ASAP7_75t_L g1038 ( 
.A(n_1009),
.B(n_1016),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_1019),
.B(n_969),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_1010),
.B(n_999),
.Y(n_1040)
);

OAI211xp5_ASAP7_75t_L g1041 ( 
.A1(n_1003),
.A2(n_981),
.B(n_988),
.C(n_914),
.Y(n_1041)
);

AND2x4_ASAP7_75t_L g1042 ( 
.A(n_1007),
.B(n_1001),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1024),
.Y(n_1043)
);

HB1xp67_ASAP7_75t_L g1044 ( 
.A(n_1027),
.Y(n_1044)
);

BUFx3_ASAP7_75t_L g1045 ( 
.A(n_1038),
.Y(n_1045)
);

INVx4_ASAP7_75t_L g1046 ( 
.A(n_1030),
.Y(n_1046)
);

INVx4_ASAP7_75t_L g1047 ( 
.A(n_1031),
.Y(n_1047)
);

NAND3xp33_ASAP7_75t_L g1048 ( 
.A(n_1041),
.B(n_1020),
.C(n_1021),
.Y(n_1048)
);

INVx5_ASAP7_75t_L g1049 ( 
.A(n_1040),
.Y(n_1049)
);

BUFx3_ASAP7_75t_L g1050 ( 
.A(n_1037),
.Y(n_1050)
);

AOI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_1042),
.A2(n_915),
.B1(n_953),
.B2(n_917),
.Y(n_1051)
);

AOI222xp33_ASAP7_75t_L g1052 ( 
.A1(n_1028),
.A2(n_949),
.B1(n_34),
.B2(n_27),
.C1(n_39),
.C2(n_30),
.Y(n_1052)
);

AND2x4_ASAP7_75t_L g1053 ( 
.A(n_1026),
.B(n_930),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_1036),
.B(n_933),
.Y(n_1054)
);

AO21x2_ASAP7_75t_L g1055 ( 
.A1(n_1039),
.A2(n_1032),
.B(n_1034),
.Y(n_1055)
);

INVx5_ASAP7_75t_L g1056 ( 
.A(n_1034),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_1029),
.Y(n_1057)
);

INVx2_ASAP7_75t_L g1058 ( 
.A(n_1024),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_1033),
.B(n_29),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_1035),
.B(n_364),
.Y(n_1060)
);

OAI31xp33_ASAP7_75t_SL g1061 ( 
.A1(n_1025),
.A2(n_33),
.A3(n_31),
.B(n_32),
.Y(n_1061)
);

INVx3_ASAP7_75t_L g1062 ( 
.A(n_1047),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_1043),
.Y(n_1063)
);

INVxp33_ASAP7_75t_L g1064 ( 
.A(n_1046),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_1058),
.Y(n_1065)
);

AND2x2_ASAP7_75t_L g1066 ( 
.A(n_1045),
.B(n_35),
.Y(n_1066)
);

INVx3_ASAP7_75t_L g1067 ( 
.A(n_1050),
.Y(n_1067)
);

HB1xp67_ASAP7_75t_L g1068 ( 
.A(n_1057),
.Y(n_1068)
);

AND2x4_ASAP7_75t_L g1069 ( 
.A(n_1056),
.B(n_1054),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_1059),
.B(n_40),
.Y(n_1070)
);

OAI21xp33_ASAP7_75t_L g1071 ( 
.A1(n_1061),
.A2(n_41),
.B(n_42),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_1053),
.B(n_1051),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1052),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_1060),
.B(n_44),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1043),
.Y(n_1075)
);

AND2x4_ASAP7_75t_L g1076 ( 
.A(n_1049),
.B(n_45),
.Y(n_1076)
);

AND2x2_ASAP7_75t_L g1077 ( 
.A(n_1044),
.B(n_47),
.Y(n_1077)
);

NAND3xp33_ASAP7_75t_L g1078 ( 
.A(n_1048),
.B(n_48),
.C(n_50),
.Y(n_1078)
);

INVx1_ASAP7_75t_SL g1079 ( 
.A(n_1045),
.Y(n_1079)
);

BUFx2_ASAP7_75t_L g1080 ( 
.A(n_1055),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1063),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_1076),
.Y(n_1082)
);

NOR2x1_ASAP7_75t_L g1083 ( 
.A(n_1080),
.B(n_52),
.Y(n_1083)
);

NOR2xp33_ASAP7_75t_L g1084 ( 
.A(n_1070),
.B(n_53),
.Y(n_1084)
);

AO221x2_ASAP7_75t_L g1085 ( 
.A1(n_1078),
.A2(n_55),
.B1(n_57),
.B2(n_54),
.C(n_56),
.Y(n_1085)
);

BUFx3_ASAP7_75t_L g1086 ( 
.A(n_1067),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_1068),
.Y(n_1087)
);

AND2x4_ASAP7_75t_L g1088 ( 
.A(n_1075),
.B(n_60),
.Y(n_1088)
);

BUFx2_ASAP7_75t_L g1089 ( 
.A(n_1072),
.Y(n_1089)
);

OR2x2_ASAP7_75t_L g1090 ( 
.A(n_1065),
.B(n_62),
.Y(n_1090)
);

NAND2xp33_ASAP7_75t_R g1091 ( 
.A(n_1066),
.B(n_66),
.Y(n_1091)
);

AND2x2_ASAP7_75t_L g1092 ( 
.A(n_1069),
.B(n_69),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_1077),
.B(n_70),
.Y(n_1093)
);

BUFx6f_ASAP7_75t_L g1094 ( 
.A(n_1074),
.Y(n_1094)
);

AO221x2_ASAP7_75t_L g1095 ( 
.A1(n_1073),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.C(n_78),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_1064),
.B(n_77),
.Y(n_1096)
);

CKINVDCx20_ASAP7_75t_R g1097 ( 
.A(n_1079),
.Y(n_1097)
);

AOI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_1071),
.A2(n_82),
.B1(n_80),
.B2(n_81),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_1062),
.Y(n_1099)
);

BUFx2_ASAP7_75t_L g1100 ( 
.A(n_1097),
.Y(n_1100)
);

INVx3_ASAP7_75t_L g1101 ( 
.A(n_1086),
.Y(n_1101)
);

INVx3_ASAP7_75t_L g1102 ( 
.A(n_1094),
.Y(n_1102)
);

AOI22xp33_ASAP7_75t_L g1103 ( 
.A1(n_1095),
.A2(n_86),
.B1(n_84),
.B2(n_85),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_1092),
.B(n_86),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1090),
.Y(n_1105)
);

INVx1_ASAP7_75t_SL g1106 ( 
.A(n_1099),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_1088),
.Y(n_1107)
);

INVx4_ASAP7_75t_L g1108 ( 
.A(n_1082),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_1096),
.B(n_89),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_1084),
.B(n_91),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1093),
.Y(n_1111)
);

OAI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_1098),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.Y(n_1112)
);

AOI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_1085),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1081),
.Y(n_1114)
);

BUFx3_ASAP7_75t_L g1115 ( 
.A(n_1097),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_1089),
.B(n_100),
.Y(n_1116)
);

AND2x2_ASAP7_75t_L g1117 ( 
.A(n_1089),
.B(n_101),
.Y(n_1117)
);

OAI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_1083),
.A2(n_105),
.B1(n_103),
.B2(n_104),
.Y(n_1118)
);

CKINVDCx16_ASAP7_75t_R g1119 ( 
.A(n_1091),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1087),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1081),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_1119),
.B(n_107),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_1101),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_1102),
.Y(n_1124)
);

A2O1A1Ixp33_ASAP7_75t_SL g1125 ( 
.A1(n_1110),
.A2(n_115),
.B(n_113),
.C(n_114),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1114),
.Y(n_1126)
);

OAI21xp33_ASAP7_75t_L g1127 ( 
.A1(n_1103),
.A2(n_117),
.B(n_118),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1105),
.B(n_121),
.Y(n_1128)
);

INVx1_ASAP7_75t_SL g1129 ( 
.A(n_1100),
.Y(n_1129)
);

OAI321xp33_ASAP7_75t_L g1130 ( 
.A1(n_1112),
.A2(n_125),
.A3(n_127),
.B1(n_123),
.B2(n_124),
.C(n_126),
.Y(n_1130)
);

OAI21xp33_ASAP7_75t_L g1131 ( 
.A1(n_1113),
.A2(n_128),
.B(n_129),
.Y(n_1131)
);

NAND3xp33_ASAP7_75t_L g1132 ( 
.A(n_1118),
.B(n_128),
.C(n_130),
.Y(n_1132)
);

INVx2_ASAP7_75t_SL g1133 ( 
.A(n_1115),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1111),
.B(n_135),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_1107),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1120),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1121),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_1108),
.B(n_144),
.Y(n_1138)
);

HB1xp67_ASAP7_75t_L g1139 ( 
.A(n_1116),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1117),
.B(n_146),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_L g1141 ( 
.A(n_1129),
.B(n_1106),
.Y(n_1141)
);

HB1xp67_ASAP7_75t_L g1142 ( 
.A(n_1139),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1133),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1123),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1135),
.B(n_1109),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1126),
.Y(n_1146)
);

INVxp67_ASAP7_75t_L g1147 ( 
.A(n_1122),
.Y(n_1147)
);

AOI22xp33_ASAP7_75t_L g1148 ( 
.A1(n_1131),
.A2(n_1104),
.B1(n_151),
.B2(n_149),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1124),
.B(n_150),
.Y(n_1149)
);

AOI22xp33_ASAP7_75t_L g1150 ( 
.A1(n_1127),
.A2(n_155),
.B1(n_153),
.B2(n_154),
.Y(n_1150)
);

OR2x2_ASAP7_75t_L g1151 ( 
.A(n_1136),
.B(n_156),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_1128),
.B(n_157),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1151),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_1143),
.Y(n_1154)
);

INVxp67_ASAP7_75t_L g1155 ( 
.A(n_1141),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_1147),
.Y(n_1156)
);

INVx2_ASAP7_75t_SL g1157 ( 
.A(n_1149),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1146),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1144),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1145),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1152),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_1148),
.B(n_1138),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_1150),
.B(n_1134),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1142),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1142),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1156),
.B(n_1137),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1163),
.A2(n_1125),
.B(n_1132),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_SL g1168 ( 
.A(n_1155),
.B(n_1130),
.Y(n_1168)
);

NOR2x1_ASAP7_75t_L g1169 ( 
.A(n_1164),
.B(n_1140),
.Y(n_1169)
);

NAND4xp75_ASAP7_75t_L g1170 ( 
.A(n_1165),
.B(n_161),
.C(n_159),
.D(n_160),
.Y(n_1170)
);

NOR3x1_ASAP7_75t_L g1171 ( 
.A(n_1157),
.B(n_162),
.C(n_163),
.Y(n_1171)
);

NOR2x1_ASAP7_75t_L g1172 ( 
.A(n_1154),
.B(n_165),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1153),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1161),
.Y(n_1174)
);

AOI21x1_ASAP7_75t_L g1175 ( 
.A1(n_1162),
.A2(n_169),
.B(n_171),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_1159),
.B(n_174),
.Y(n_1176)
);

NAND3xp33_ASAP7_75t_SL g1177 ( 
.A(n_1160),
.B(n_176),
.C(n_177),
.Y(n_1177)
);

OAI322xp33_ASAP7_75t_L g1178 ( 
.A1(n_1158),
.A2(n_179),
.A3(n_180),
.B1(n_181),
.B2(n_182),
.C1(n_183),
.C2(n_184),
.Y(n_1178)
);

AOI211xp5_ASAP7_75t_L g1179 ( 
.A1(n_1167),
.A2(n_188),
.B(n_186),
.C(n_187),
.Y(n_1179)
);

INVx2_ASAP7_75t_SL g1180 ( 
.A(n_1172),
.Y(n_1180)
);

INVx1_ASAP7_75t_SL g1181 ( 
.A(n_1169),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1168),
.A2(n_194),
.B(n_195),
.Y(n_1182)
);

NOR2xp67_ASAP7_75t_SL g1183 ( 
.A(n_1170),
.B(n_195),
.Y(n_1183)
);

NAND4xp25_ASAP7_75t_L g1184 ( 
.A(n_1166),
.B(n_200),
.C(n_198),
.D(n_199),
.Y(n_1184)
);

NOR3xp33_ASAP7_75t_L g1185 ( 
.A(n_1173),
.B(n_201),
.C(n_202),
.Y(n_1185)
);

AOI321xp33_ASAP7_75t_L g1186 ( 
.A1(n_1174),
.A2(n_205),
.A3(n_207),
.B1(n_203),
.B2(n_204),
.C(n_206),
.Y(n_1186)
);

NOR2x1_ASAP7_75t_L g1187 ( 
.A(n_1177),
.B(n_204),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_1175),
.Y(n_1188)
);

AOI221xp5_ASAP7_75t_L g1189 ( 
.A1(n_1178),
.A2(n_211),
.B1(n_209),
.B2(n_210),
.C(n_212),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1171),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1176),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1180),
.Y(n_1192)
);

NAND4xp75_ASAP7_75t_L g1193 ( 
.A(n_1187),
.B(n_218),
.C(n_215),
.D(n_217),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1190),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1188),
.Y(n_1195)
);

AND2x4_ASAP7_75t_L g1196 ( 
.A(n_1181),
.B(n_217),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1188),
.Y(n_1197)
);

INVxp67_ASAP7_75t_L g1198 ( 
.A(n_1183),
.Y(n_1198)
);

AND2x4_ASAP7_75t_L g1199 ( 
.A(n_1191),
.B(n_221),
.Y(n_1199)
);

NAND4xp75_ASAP7_75t_L g1200 ( 
.A(n_1182),
.B(n_224),
.C(n_222),
.D(n_223),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_R g1201 ( 
.A(n_1192),
.B(n_1186),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_R g1202 ( 
.A(n_1194),
.B(n_1179),
.Y(n_1202)
);

NOR2xp33_ASAP7_75t_R g1203 ( 
.A(n_1198),
.B(n_1195),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_R g1204 ( 
.A(n_1197),
.B(n_1184),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_1196),
.B(n_1189),
.Y(n_1205)
);

INVx4_ASAP7_75t_L g1206 ( 
.A(n_1203),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1205),
.B(n_1199),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1206),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1207),
.Y(n_1209)
);

AND2x4_ASAP7_75t_SL g1210 ( 
.A(n_1208),
.B(n_1209),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1210),
.A2(n_1201),
.B1(n_1202),
.B2(n_1204),
.Y(n_1211)
);

OAI22xp5_ASAP7_75t_SL g1212 ( 
.A1(n_1211),
.A2(n_1193),
.B1(n_1200),
.B2(n_1185),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1212),
.A2(n_231),
.B1(n_229),
.B2(n_230),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1213),
.Y(n_1214)
);

OAI221xp5_ASAP7_75t_R g1215 ( 
.A1(n_1214),
.A2(n_234),
.B1(n_232),
.B2(n_233),
.C(n_235),
.Y(n_1215)
);

AOI211xp5_ASAP7_75t_L g1216 ( 
.A1(n_1215),
.A2(n_236),
.B(n_234),
.C(n_235),
.Y(n_1216)
);


endmodule