module fake_aes_1737_n_40 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_40);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_40;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_30;
wire n_13;
wire n_26;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
wire n_39;
INVx1_ASAP7_75t_L g11 ( .A(n_0), .Y(n_11) );
BUFx8_ASAP7_75t_L g12 ( .A(n_7), .Y(n_12) );
NOR2xp33_ASAP7_75t_L g13 ( .A(n_9), .B(n_8), .Y(n_13) );
NOR2xp33_ASAP7_75t_R g14 ( .A(n_9), .B(n_1), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_7), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_10), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_1), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_15), .B(n_8), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_17), .Y(n_19) );
INVx2_ASAP7_75t_SL g20 ( .A(n_17), .Y(n_20) );
HB1xp67_ASAP7_75t_L g21 ( .A(n_12), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_17), .Y(n_22) );
OAI22xp33_ASAP7_75t_L g23 ( .A1(n_21), .A2(n_11), .B1(n_13), .B2(n_12), .Y(n_23) );
NAND2xp33_ASAP7_75t_SL g24 ( .A(n_18), .B(n_14), .Y(n_24) );
INVx2_ASAP7_75t_L g25 ( .A(n_22), .Y(n_25) );
OAI22xp33_ASAP7_75t_L g26 ( .A1(n_20), .A2(n_11), .B1(n_12), .B2(n_16), .Y(n_26) );
AND2x2_ASAP7_75t_L g27 ( .A(n_25), .B(n_20), .Y(n_27) );
NAND4xp25_ASAP7_75t_L g28 ( .A(n_24), .B(n_19), .C(n_22), .D(n_12), .Y(n_28) );
AOI221xp5_ASAP7_75t_L g29 ( .A1(n_23), .A2(n_19), .B1(n_22), .B2(n_3), .C(n_4), .Y(n_29) );
AND2x2_ASAP7_75t_L g30 ( .A(n_27), .B(n_25), .Y(n_30) );
INVx2_ASAP7_75t_L g31 ( .A(n_28), .Y(n_31) );
INVx2_ASAP7_75t_L g32 ( .A(n_30), .Y(n_32) );
NAND2xp5_ASAP7_75t_SL g33 ( .A(n_31), .B(n_26), .Y(n_33) );
OAI221xp5_ASAP7_75t_L g34 ( .A1(n_33), .A2(n_29), .B1(n_31), .B2(n_3), .C(n_4), .Y(n_34) );
NAND2xp5_ASAP7_75t_L g35 ( .A(n_32), .B(n_0), .Y(n_35) );
INVxp67_ASAP7_75t_L g36 ( .A(n_32), .Y(n_36) );
AND2x4_ASAP7_75t_L g37 ( .A(n_36), .B(n_6), .Y(n_37) );
INVx1_ASAP7_75t_SL g38 ( .A(n_35), .Y(n_38) );
NOR3xp33_ASAP7_75t_SL g39 ( .A(n_38), .B(n_34), .C(n_5), .Y(n_39) );
AOI322xp5_ASAP7_75t_L g40 ( .A1(n_39), .A2(n_2), .A3(n_5), .B1(n_37), .B2(n_13), .C1(n_23), .C2(n_38), .Y(n_40) );
endmodule