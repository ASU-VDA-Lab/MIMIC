module real_jpeg_23687_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_37;
wire n_21;
wire n_35;
wire n_38;
wire n_33;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_23;
wire n_11;
wire n_14;
wire n_25;
wire n_7;
wire n_22;
wire n_18;
wire n_36;
wire n_39;
wire n_40;
wire n_41;
wire n_27;
wire n_26;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_0),
.B(n_4),
.Y(n_36)
);

HAxp5_ASAP7_75t_SL g40 ( 
.A(n_0),
.B(n_27),
.CON(n_40),
.SN(n_40)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g9 ( 
.A(n_2),
.B(n_4),
.Y(n_9)
);

AOI22xp5_ASAP7_75t_SL g12 ( 
.A1(n_2),
.A2(n_13),
.B1(n_14),
.B2(n_19),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_3),
.B(n_22),
.Y(n_31)
);

OR2x2_ASAP7_75t_SL g37 ( 
.A(n_3),
.B(n_22),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_4),
.B(n_12),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_4),
.B(n_19),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_4),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_4),
.B(n_5),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_5),
.B(n_16),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_5),
.B(n_16),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

AOI221xp5_ASAP7_75t_L g6 ( 
.A1(n_7),
.A2(n_20),
.B1(n_24),
.B2(n_28),
.C(n_29),
.Y(n_6)
);

NAND2xp5_ASAP7_75t_L g7 ( 
.A(n_8),
.B(n_10),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_9),
.Y(n_8)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_11),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_12),
.B(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g13 ( 
.A(n_14),
.Y(n_13)
);

OR2x2_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_17),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_23),
.Y(n_21)
);

AND2x2_ASAP7_75t_SL g28 ( 
.A(n_22),
.B(n_23),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_32),
.B1(n_37),
.B2(n_38),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_41),
.Y(n_39)
);

BUFx24_ASAP7_75t_SL g42 ( 
.A(n_40),
.Y(n_42)
);


endmodule