module fake_jpeg_30974_n_263 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_263);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_263;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_33;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_118;
wire n_155;
wire n_82;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx6_ASAP7_75t_SL g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_17),
.B(n_6),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_38),
.B(n_40),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_41),
.Y(n_61)
);

HAxp5_ASAP7_75t_SL g40 ( 
.A(n_18),
.B(n_0),
.CON(n_40),
.SN(n_40)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_18),
.B(n_6),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_42),
.Y(n_100)
);

BUFx12_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_50),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_44),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx8_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_17),
.A2(n_14),
.B1(n_5),
.B2(n_7),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_54),
.A2(n_27),
.B1(n_35),
.B2(n_24),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_34),
.Y(n_56)
);

NAND2xp33_ASAP7_75t_SL g89 ( 
.A(n_56),
.B(n_57),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx16f_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_40),
.A2(n_22),
.B1(n_29),
.B2(n_21),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_60),
.A2(n_91),
.B1(n_93),
.B2(n_25),
.Y(n_114)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_65),
.B(n_69),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_71),
.B(n_72),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_38),
.B(n_30),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_41),
.B(n_27),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_74),
.B(n_88),
.Y(n_112)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_75),
.B(n_78),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_76),
.A2(n_24),
.B1(n_23),
.B2(n_19),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_43),
.B(n_30),
.Y(n_78)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_53),
.A2(n_22),
.B1(n_29),
.B2(n_32),
.Y(n_79)
);

OA22x2_ASAP7_75t_L g110 ( 
.A1(n_79),
.A2(n_90),
.B1(n_91),
.B2(n_93),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_83),
.Y(n_117)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_51),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_86),
.B(n_87),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_43),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_45),
.B(n_19),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_45),
.A2(n_22),
.B1(n_29),
.B2(n_21),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_50),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_103),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_48),
.A2(n_21),
.B1(n_26),
.B2(n_16),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_50),
.A2(n_36),
.B(n_15),
.C(n_32),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_95),
.A2(n_97),
.B(n_25),
.C(n_15),
.Y(n_108)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_40),
.A2(n_36),
.B(n_15),
.C(n_32),
.Y(n_97)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_38),
.B(n_35),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_105),
.Y(n_121)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_51),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_47),
.Y(n_104)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_104),
.Y(n_107)
);

INVx6_ASAP7_75t_SL g105 ( 
.A(n_58),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_108),
.B(n_62),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_61),
.A2(n_25),
.B1(n_33),
.B2(n_31),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_109),
.A2(n_114),
.B1(n_63),
.B2(n_94),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_122),
.B1(n_90),
.B2(n_85),
.Y(n_135)
);

AND2x2_ASAP7_75t_SL g115 ( 
.A(n_68),
.B(n_0),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_115),
.B(n_134),
.C(n_63),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_99),
.B(n_33),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_120),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_31),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_77),
.B(n_23),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_129),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_79),
.A2(n_76),
.B1(n_84),
.B2(n_70),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_124),
.A2(n_125),
.B1(n_67),
.B2(n_80),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_79),
.A2(n_84),
.B1(n_70),
.B2(n_73),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_97),
.B(n_0),
.Y(n_129)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

NAND2x1_ASAP7_75t_SL g131 ( 
.A(n_95),
.B(n_1),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_131),
.A2(n_1),
.B(n_2),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_89),
.B(n_1),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_135),
.A2(n_140),
.B1(n_110),
.B2(n_115),
.Y(n_169)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_133),
.Y(n_136)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_138),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_127),
.B(n_66),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_147),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_110),
.A2(n_60),
.B1(n_73),
.B2(n_94),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_141),
.A2(n_143),
.B1(n_158),
.B2(n_160),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_108),
.A2(n_100),
.B1(n_80),
.B2(n_96),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_120),
.B(n_14),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_144),
.B(n_157),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_100),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_149),
.Y(n_175)
);

OAI21xp33_ASAP7_75t_L g181 ( 
.A1(n_146),
.A2(n_148),
.B(n_118),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_112),
.B(n_64),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_107),
.Y(n_150)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_150),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_129),
.B(n_3),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_151),
.B(n_152),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_64),
.Y(n_152)
);

MAJx2_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_64),
.C(n_62),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_118),
.C(n_121),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_67),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_154),
.B(n_156),
.Y(n_186)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_155),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_109),
.B(n_62),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_119),
.B(n_13),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_110),
.A2(n_123),
.B1(n_122),
.B2(n_117),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_161),
.B(n_162),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_128),
.B(n_8),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_111),
.B(n_116),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_163),
.B(n_164),
.Y(n_176)
);

NOR3xp33_ASAP7_75t_L g164 ( 
.A(n_116),
.B(n_82),
.C(n_81),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_142),
.B(n_115),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_168),
.B(n_188),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_169),
.A2(n_173),
.B1(n_184),
.B2(n_141),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_159),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_171),
.B(n_179),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_140),
.A2(n_134),
.B1(n_117),
.B2(n_107),
.Y(n_173)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_136),
.Y(n_178)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_178),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_159),
.Y(n_179)
);

AND2x6_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_121),
.Y(n_180)
);

AOI221xp5_ASAP7_75t_L g207 ( 
.A1(n_180),
.A2(n_162),
.B1(n_150),
.B2(n_4),
.C(n_7),
.Y(n_207)
);

HAxp5_ASAP7_75t_SL g202 ( 
.A(n_181),
.B(n_146),
.CON(n_202),
.SN(n_202)
);

INVx13_ASAP7_75t_L g182 ( 
.A(n_155),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_182),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_135),
.A2(n_121),
.B1(n_113),
.B2(n_106),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_138),
.Y(n_185)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_185),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_187),
.B(n_161),
.C(n_153),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_142),
.B(n_126),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_190),
.B(n_187),
.C(n_166),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_193),
.B(n_195),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_184),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_174),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_177),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_169),
.A2(n_173),
.B1(n_160),
.B2(n_183),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_197),
.A2(n_167),
.B1(n_132),
.B2(n_182),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_186),
.A2(n_183),
.B(n_175),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_198),
.A2(n_199),
.B(n_200),
.Y(n_210)
);

A2O1A1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_186),
.A2(n_145),
.B(n_154),
.C(n_156),
.Y(n_199)
);

AOI32xp33_ASAP7_75t_L g200 ( 
.A1(n_180),
.A2(n_163),
.A3(n_152),
.B1(n_149),
.B2(n_153),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_202),
.A2(n_207),
.B(n_189),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_188),
.A2(n_158),
.B1(n_151),
.B2(n_157),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_203),
.A2(n_189),
.B1(n_172),
.B2(n_167),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_175),
.A2(n_137),
.B(n_144),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_204),
.B(n_172),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_176),
.B(n_137),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_205),
.B(n_177),
.Y(n_211)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_165),
.Y(n_206)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_206),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_209),
.B(n_211),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_218),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_192),
.A2(n_165),
.B1(n_185),
.B2(n_178),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_213),
.A2(n_217),
.B1(n_220),
.B2(n_224),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_214),
.B(n_219),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_193),
.A2(n_179),
.B1(n_171),
.B2(n_170),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_190),
.B(n_166),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_168),
.C(n_170),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_222),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_126),
.C(n_106),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_198),
.B(n_197),
.C(n_200),
.Y(n_223)
);

MAJx2_ASAP7_75t_L g232 ( 
.A(n_223),
.B(n_199),
.C(n_204),
.Y(n_232)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_215),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_227),
.Y(n_237)
);

BUFx12_ASAP7_75t_L g227 ( 
.A(n_217),
.Y(n_227)
);

NAND2xp33_ASAP7_75t_SL g230 ( 
.A(n_216),
.B(n_199),
.Y(n_230)
);

NOR3xp33_ASAP7_75t_L g235 ( 
.A(n_230),
.B(n_229),
.C(n_223),
.Y(n_235)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_222),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_231),
.B(n_228),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_232),
.B(n_221),
.Y(n_239)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_235),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_226),
.B(n_205),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_238),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_228),
.B(n_218),
.C(n_212),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_239),
.B(n_242),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_233),
.A2(n_225),
.B1(n_231),
.B2(n_234),
.Y(n_240)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_240),
.Y(n_248)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_241),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_210),
.C(n_219),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_237),
.A2(n_207),
.B(n_208),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_245),
.A2(n_247),
.B(n_203),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_239),
.A2(n_227),
.B1(n_230),
.B2(n_242),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_253),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_249),
.B(n_208),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_251),
.B(n_252),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_194),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_246),
.B(n_238),
.C(n_227),
.Y(n_253)
);

AOI21x1_ASAP7_75t_L g254 ( 
.A1(n_247),
.A2(n_227),
.B(n_206),
.Y(n_254)
);

AO21x2_ASAP7_75t_L g257 ( 
.A1(n_254),
.A2(n_248),
.B(n_191),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_253),
.B(n_246),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_256),
.A2(n_257),
.B1(n_244),
.B2(n_194),
.Y(n_259)
);

AOI322xp5_ASAP7_75t_L g261 ( 
.A1(n_259),
.A2(n_260),
.A3(n_257),
.B1(n_258),
.B2(n_182),
.C1(n_167),
.C2(n_8),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_255),
.B(n_192),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_261),
.B(n_132),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_262),
.B(n_132),
.Y(n_263)
);


endmodule