module fake_netlist_5_1512_n_1351 (n_137, n_294, n_318, n_82, n_194, n_316, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_127, n_75, n_235, n_226, n_74, n_57, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_17, n_254, n_33, n_23, n_302, n_265, n_293, n_244, n_47, n_173, n_198, n_247, n_314, n_8, n_292, n_100, n_212, n_119, n_275, n_252, n_26, n_295, n_133, n_2, n_6, n_39, n_147, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_204, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_10, n_24, n_132, n_90, n_101, n_281, n_240, n_189, n_220, n_291, n_231, n_257, n_31, n_13, n_152, n_317, n_9, n_195, n_42, n_227, n_45, n_271, n_94, n_123, n_167, n_234, n_308, n_267, n_297, n_156, n_5, n_225, n_219, n_157, n_131, n_192, n_223, n_158, n_138, n_264, n_109, n_163, n_276, n_95, n_183, n_185, n_243, n_169, n_59, n_255, n_215, n_196, n_211, n_218, n_181, n_3, n_290, n_221, n_178, n_287, n_72, n_104, n_41, n_56, n_141, n_15, n_145, n_48, n_50, n_313, n_88, n_216, n_168, n_164, n_311, n_208, n_142, n_214, n_140, n_299, n_303, n_296, n_241, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_98, n_197, n_107, n_69, n_236, n_1, n_249, n_304, n_203, n_274, n_80, n_35, n_73, n_277, n_92, n_19, n_149, n_309, n_30, n_14, n_84, n_130, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_170, n_27, n_77, n_102, n_161, n_273, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_210, n_91, n_176, n_182, n_143, n_83, n_237, n_180, n_207, n_37, n_229, n_108, n_66, n_177, n_60, n_16, n_0, n_58, n_18, n_117, n_233, n_205, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_175, n_262, n_238, n_99, n_319, n_20, n_121, n_242, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_199, n_187, n_32, n_103, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_1351);

input n_137;
input n_294;
input n_318;
input n_82;
input n_194;
input n_316;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_17;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_8;
input n_292;
input n_100;
input n_212;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_2;
input n_6;
input n_39;
input n_147;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_204;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_10;
input n_24;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_31;
input n_13;
input n_152;
input n_317;
input n_9;
input n_195;
input n_42;
input n_227;
input n_45;
input n_271;
input n_94;
input n_123;
input n_167;
input n_234;
input n_308;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_158;
input n_138;
input n_264;
input n_109;
input n_163;
input n_276;
input n_95;
input n_183;
input n_185;
input n_243;
input n_169;
input n_59;
input n_255;
input n_215;
input n_196;
input n_211;
input n_218;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_287;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_15;
input n_145;
input n_48;
input n_50;
input n_313;
input n_88;
input n_216;
input n_168;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_140;
input n_299;
input n_303;
input n_296;
input n_241;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_98;
input n_197;
input n_107;
input n_69;
input n_236;
input n_1;
input n_249;
input n_304;
input n_203;
input n_274;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_149;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_170;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_210;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_237;
input n_180;
input n_207;
input n_37;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_16;
input n_0;
input n_58;
input n_18;
input n_117;
input n_233;
input n_205;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_175;
input n_262;
input n_238;
input n_99;
input n_319;
input n_20;
input n_121;
input n_242;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_199;
input n_187;
input n_32;
input n_103;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1351;

wire n_924;
wire n_1263;
wire n_977;
wire n_611;
wire n_1126;
wire n_1166;
wire n_469;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_667;
wire n_790;
wire n_1055;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1292;
wire n_1198;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_688;
wire n_800;
wire n_1347;
wire n_671;
wire n_819;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_625;
wire n_854;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_929;
wire n_1124;
wire n_902;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_731;
wire n_371;
wire n_1314;
wire n_709;
wire n_1236;
wire n_569;
wire n_920;
wire n_1289;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_1078;
wire n_775;
wire n_600;
wire n_1328;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_350;
wire n_798;
wire n_646;
wire n_436;
wire n_1216;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1284;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1069;
wire n_1075;
wire n_1322;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_907;
wire n_989;
wire n_1039;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_647;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_561;
wire n_1319;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_596;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_728;
wire n_1162;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_409;
wire n_887;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_759;
wire n_806;
wire n_324;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_649;
wire n_547;
wire n_1191;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1233;
wire n_526;
wire n_372;
wire n_677;
wire n_1333;
wire n_1121;
wire n_368;
wire n_604;
wire n_433;
wire n_949;
wire n_1008;
wire n_946;
wire n_1001;
wire n_498;
wire n_689;
wire n_738;
wire n_640;
wire n_624;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1054;
wire n_1269;
wire n_1095;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_374;
wire n_396;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_1336;
wire n_473;
wire n_1309;
wire n_1043;
wire n_355;
wire n_486;
wire n_614;
wire n_337;
wire n_1286;
wire n_1177;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1132;
wire n_388;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1006;
wire n_329;
wire n_1270;
wire n_582;
wire n_1332;
wire n_512;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1304;
wire n_1324;
wire n_987;
wire n_767;
wire n_993;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_513;
wire n_1094;
wire n_560;
wire n_340;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_960;
wire n_1290;
wire n_1123;
wire n_1047;
wire n_634;
wire n_1252;
wire n_348;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_950;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_389;
wire n_418;
wire n_912;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_376;
wire n_967;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_1343;
wire n_1203;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_507;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1329;
wire n_1312;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_943;
wire n_341;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1214;
wire n_1342;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1077;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1350;
wire n_1096;
wire n_833;
wire n_1307;
wire n_988;
wire n_814;
wire n_1201;
wire n_1114;
wire n_655;
wire n_669;
wire n_472;
wire n_1176;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_830;
wire n_1296;
wire n_801;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1019;
wire n_1105;
wire n_1338;
wire n_577;
wire n_338;
wire n_693;
wire n_836;
wire n_990;
wire n_975;
wire n_1256;
wire n_567;
wire n_778;
wire n_1122;
wire n_770;
wire n_458;
wire n_1102;
wire n_711;
wire n_1187;
wire n_1164;
wire n_489;
wire n_1174;
wire n_617;
wire n_1303;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_1116;
wire n_1212;
wire n_726;
wire n_982;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_774;
wire n_1335;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_557;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_393;
wire n_487;
wire n_665;
wire n_421;
wire n_910;
wire n_768;
wire n_1302;
wire n_1136;
wire n_1313;
wire n_754;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_1310;
wire n_427;
wire n_791;
wire n_732;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_676;
wire n_653;
wire n_642;
wire n_855;
wire n_1178;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_467;
wire n_1227;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_725;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_714;
wire n_909;
wire n_997;
wire n_932;
wire n_612;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_733;
wire n_941;
wire n_981;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_752;
wire n_905;
wire n_1108;
wire n_782;
wire n_1100;
wire n_862;
wire n_760;
wire n_381;
wire n_390;
wire n_1330;
wire n_481;
wire n_769;
wire n_1046;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_1225;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1344;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_432;
wire n_839;
wire n_1210;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_772;
wire n_499;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1012;
wire n_1348;
wire n_903;
wire n_740;
wire n_384;
wire n_1315;
wire n_1061;
wire n_333;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_632;
wire n_699;
wire n_979;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_1321;
wire n_585;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1076;
wire n_1091;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1220;
wire n_437;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_1042;
wire n_412;
wire n_657;
wire n_644;
wire n_1160;
wire n_491;
wire n_1258;
wire n_1074;
wire n_566;
wire n_565;
wire n_597;
wire n_1181;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1251;

INVx1_ASAP7_75t_L g321 ( 
.A(n_159),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_247),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_3),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_129),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_220),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_83),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_264),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_149),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_198),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_76),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_66),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_36),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_200),
.Y(n_333)
);

BUFx2_ASAP7_75t_L g334 ( 
.A(n_167),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_294),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_4),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_302),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_187),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_212),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_319),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_106),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_228),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_183),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_22),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_5),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_191),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_23),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_77),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_69),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_282),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_39),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_56),
.Y(n_352)
);

INVx1_ASAP7_75t_SL g353 ( 
.A(n_300),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_46),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_280),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_172),
.Y(n_356)
);

BUFx2_ASAP7_75t_L g357 ( 
.A(n_75),
.Y(n_357)
);

BUFx10_ASAP7_75t_L g358 ( 
.A(n_153),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_139),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_25),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_131),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_90),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_165),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_166),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_119),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_41),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_174),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_6),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_45),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_259),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_52),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_312),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_0),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_291),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_313),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_46),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_168),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_289),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_225),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_147),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_78),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_251),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_47),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_134),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_130),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_11),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_161),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_67),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_265),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_162),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_72),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_235),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_310),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_4),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_315),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_246),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_231),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_184),
.Y(n_398)
);

BUFx10_ASAP7_75t_L g399 ( 
.A(n_68),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_260),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_63),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_99),
.Y(n_402)
);

BUFx8_ASAP7_75t_SL g403 ( 
.A(n_136),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_62),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_226),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_135),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_39),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_124),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_317),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_108),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_70),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g412 ( 
.A(n_237),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_164),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_305),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_80),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_208),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_113),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_105),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_45),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_272),
.Y(n_420)
);

BUFx10_ASAP7_75t_L g421 ( 
.A(n_102),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_141),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_8),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_273),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_155),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_290),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_71),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_182),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_104),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_23),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_33),
.Y(n_431)
);

BUFx3_ASAP7_75t_L g432 ( 
.A(n_6),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_292),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_221),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_179),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_277),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_47),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_297),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_263),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_91),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_301),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_85),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_36),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_34),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_25),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_158),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_117),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_271),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_148),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_137),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_318),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g452 ( 
.A(n_107),
.Y(n_452)
);

BUFx10_ASAP7_75t_L g453 ( 
.A(n_173),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_24),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_311),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_216),
.Y(n_456)
);

INVx2_ASAP7_75t_SL g457 ( 
.A(n_195),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_215),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_30),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_110),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_248),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_94),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_283),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_253),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_230),
.Y(n_465)
);

CKINVDCx14_ASAP7_75t_R g466 ( 
.A(n_43),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_190),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_125),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_285),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_128),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_59),
.Y(n_471)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_258),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_10),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_304),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_95),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_43),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_177),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_87),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_81),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_140),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_232),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_204),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_199),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_194),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_22),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_14),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_73),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_267),
.Y(n_488)
);

BUFx8_ASAP7_75t_SL g489 ( 
.A(n_245),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_261),
.Y(n_490)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_252),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_266),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_288),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_154),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_206),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_144),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_202),
.Y(n_497)
);

INVxp33_ASAP7_75t_SL g498 ( 
.A(n_332),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_368),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_432),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_432),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_369),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_340),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_386),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_322),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_394),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_324),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_407),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_325),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_R g510 ( 
.A(n_466),
.B(n_60),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_437),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_329),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_335),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_338),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_372),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_445),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_486),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_340),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_497),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_339),
.Y(n_520)
);

INVxp33_ASAP7_75t_L g521 ( 
.A(n_491),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_372),
.Y(n_522)
);

INVxp67_ASAP7_75t_SL g523 ( 
.A(n_334),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_343),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_497),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_321),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_327),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_358),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_326),
.Y(n_529)
);

CKINVDCx16_ASAP7_75t_R g530 ( 
.A(n_380),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_346),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_328),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_349),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_332),
.Y(n_534)
);

INVxp67_ASAP7_75t_L g535 ( 
.A(n_376),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_350),
.Y(n_536)
);

INVxp33_ASAP7_75t_L g537 ( 
.A(n_403),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_357),
.B(n_0),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_356),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_430),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_330),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_359),
.Y(n_542)
);

CKINVDCx16_ASAP7_75t_R g543 ( 
.A(n_380),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_452),
.B(n_1),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_430),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_418),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_331),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_418),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_333),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_337),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_326),
.Y(n_551)
);

INVxp33_ASAP7_75t_L g552 ( 
.A(n_403),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_367),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_361),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_376),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_363),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_428),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_342),
.Y(n_558)
);

NOR2xp67_ASAP7_75t_L g559 ( 
.A(n_457),
.B(n_1),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_428),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_364),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_429),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_348),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_355),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_429),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_362),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_365),
.Y(n_567)
);

INVxp67_ASAP7_75t_SL g568 ( 
.A(n_341),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_381),
.Y(n_569)
);

INVxp67_ASAP7_75t_SL g570 ( 
.A(n_472),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_370),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_367),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_382),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_448),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_358),
.B(n_2),
.Y(n_575)
);

CKINVDCx16_ASAP7_75t_R g576 ( 
.A(n_448),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_375),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_390),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_377),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_378),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_385),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_387),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_391),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g584 ( 
.A(n_323),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_455),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_455),
.Y(n_586)
);

HB1xp67_ASAP7_75t_L g587 ( 
.A(n_336),
.Y(n_587)
);

CKINVDCx20_ASAP7_75t_R g588 ( 
.A(n_489),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_392),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_393),
.Y(n_590)
);

INVxp67_ASAP7_75t_SL g591 ( 
.A(n_395),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_401),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_402),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_396),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_489),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_405),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_397),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_413),
.Y(n_598)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_344),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_529),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_529),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_551),
.Y(n_602)
);

OA21x2_ASAP7_75t_L g603 ( 
.A1(n_551),
.A2(n_379),
.B(n_374),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_499),
.Y(n_604)
);

HB1xp67_ASAP7_75t_L g605 ( 
.A(n_584),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_572),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_499),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_572),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_553),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_553),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_526),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_553),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_516),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_527),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_516),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_532),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_521),
.B(n_457),
.Y(n_617)
);

OAI21x1_ASAP7_75t_L g618 ( 
.A1(n_541),
.A2(n_379),
.B(n_374),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_505),
.Y(n_619)
);

NAND2xp33_ASAP7_75t_R g620 ( 
.A(n_498),
.B(n_490),
.Y(n_620)
);

XNOR2xp5_ASAP7_75t_L g621 ( 
.A(n_546),
.B(n_345),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_547),
.Y(n_622)
);

BUFx2_ASAP7_75t_L g623 ( 
.A(n_588),
.Y(n_623)
);

INVxp67_ASAP7_75t_L g624 ( 
.A(n_587),
.Y(n_624)
);

BUFx2_ASAP7_75t_L g625 ( 
.A(n_588),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_507),
.B(n_384),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_549),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_502),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_550),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_558),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_563),
.Y(n_631)
);

AND2x4_ASAP7_75t_L g632 ( 
.A(n_591),
.B(n_384),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_535),
.B(n_358),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_509),
.B(n_388),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_534),
.Y(n_635)
);

INVx4_ASAP7_75t_L g636 ( 
.A(n_512),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_564),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_513),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_566),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_514),
.B(n_388),
.Y(n_640)
);

AND2x4_ASAP7_75t_L g641 ( 
.A(n_559),
.B(n_389),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_520),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_567),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_524),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_531),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_546),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_571),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_533),
.Y(n_648)
);

BUFx2_ASAP7_75t_L g649 ( 
.A(n_599),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_536),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_577),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_521),
.B(n_353),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_579),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_539),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_580),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_581),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_542),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_582),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_583),
.Y(n_659)
);

CKINVDCx20_ASAP7_75t_R g660 ( 
.A(n_548),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_554),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_589),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_590),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_592),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_593),
.Y(n_665)
);

CKINVDCx20_ASAP7_75t_R g666 ( 
.A(n_548),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_556),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_596),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_561),
.B(n_412),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_598),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_504),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_506),
.Y(n_672)
);

CKINVDCx16_ASAP7_75t_R g673 ( 
.A(n_530),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_569),
.B(n_490),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_573),
.Y(n_675)
);

CKINVDCx20_ASAP7_75t_R g676 ( 
.A(n_560),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_508),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_511),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_517),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_500),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_578),
.B(n_389),
.Y(n_681)
);

OAI21x1_ASAP7_75t_L g682 ( 
.A1(n_575),
.A2(n_414),
.B(n_400),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_501),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_518),
.Y(n_684)
);

OR2x6_ASAP7_75t_L g685 ( 
.A(n_649),
.B(n_555),
.Y(n_685)
);

OR2x2_ASAP7_75t_L g686 ( 
.A(n_635),
.B(n_543),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_608),
.B(n_568),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_608),
.B(n_570),
.Y(n_688)
);

BUFx3_ASAP7_75t_L g689 ( 
.A(n_684),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_603),
.B(n_519),
.Y(n_690)
);

BUFx3_ASAP7_75t_L g691 ( 
.A(n_680),
.Y(n_691)
);

AND2x6_ASAP7_75t_L g692 ( 
.A(n_632),
.B(n_400),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_L g693 ( 
.A1(n_632),
.A2(n_544),
.B1(n_538),
.B2(n_414),
.Y(n_693)
);

OR2x2_ASAP7_75t_L g694 ( 
.A(n_626),
.B(n_576),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_652),
.B(n_427),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_683),
.B(n_503),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_632),
.B(n_427),
.Y(n_697)
);

INVx3_ASAP7_75t_L g698 ( 
.A(n_604),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_671),
.Y(n_699)
);

AND2x4_ASAP7_75t_L g700 ( 
.A(n_672),
.B(n_503),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_604),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_619),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_603),
.B(n_525),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_604),
.Y(n_704)
);

INVx5_ASAP7_75t_L g705 ( 
.A(n_604),
.Y(n_705)
);

INVx4_ASAP7_75t_L g706 ( 
.A(n_628),
.Y(n_706)
);

NOR2x1p5_ASAP7_75t_L g707 ( 
.A(n_636),
.B(n_528),
.Y(n_707)
);

INVx4_ASAP7_75t_SL g708 ( 
.A(n_641),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_617),
.B(n_523),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_607),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_607),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_607),
.Y(n_712)
);

INVx3_ASAP7_75t_L g713 ( 
.A(n_607),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_624),
.B(n_594),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_628),
.Y(n_715)
);

INVx3_ASAP7_75t_L g716 ( 
.A(n_628),
.Y(n_716)
);

OAI22xp33_ASAP7_75t_L g717 ( 
.A1(n_620),
.A2(n_351),
.B1(n_352),
.B2(n_347),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_603),
.B(n_434),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_641),
.B(n_434),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_600),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_677),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_641),
.B(n_612),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_669),
.B(n_597),
.Y(n_723)
);

INVx6_ASAP7_75t_L g724 ( 
.A(n_628),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_634),
.B(n_475),
.Y(n_725)
);

INVx3_ASAP7_75t_L g726 ( 
.A(n_612),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_600),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_618),
.Y(n_728)
);

BUFx2_ASAP7_75t_L g729 ( 
.A(n_621),
.Y(n_729)
);

BUFx6f_ASAP7_75t_L g730 ( 
.A(n_618),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_678),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_633),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_640),
.B(n_475),
.Y(n_733)
);

AND2x6_ASAP7_75t_L g734 ( 
.A(n_681),
.B(n_435),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_611),
.Y(n_735)
);

BUFx6f_ASAP7_75t_L g736 ( 
.A(n_682),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_636),
.B(n_510),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_614),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_674),
.B(n_528),
.Y(n_739)
);

OR2x2_ASAP7_75t_L g740 ( 
.A(n_605),
.B(n_537),
.Y(n_740)
);

BUFx10_ASAP7_75t_L g741 ( 
.A(n_638),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_682),
.A2(n_447),
.B1(n_451),
.B2(n_436),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_638),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_600),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_612),
.Y(n_745)
);

CKINVDCx16_ASAP7_75t_R g746 ( 
.A(n_673),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_644),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_602),
.Y(n_748)
);

INVx4_ASAP7_75t_L g749 ( 
.A(n_639),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_622),
.Y(n_750)
);

NAND2x1p5_ASAP7_75t_L g751 ( 
.A(n_636),
.B(n_460),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_645),
.B(n_537),
.Y(n_752)
);

NAND2xp33_ASAP7_75t_L g753 ( 
.A(n_642),
.B(n_398),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_629),
.Y(n_754)
);

AND2x6_ASAP7_75t_L g755 ( 
.A(n_630),
.B(n_470),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_648),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_654),
.B(n_552),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_616),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_602),
.B(n_601),
.Y(n_759)
);

INVxp67_ASAP7_75t_L g760 ( 
.A(n_637),
.Y(n_760)
);

NAND2x1p5_ASAP7_75t_L g761 ( 
.A(n_639),
.B(n_482),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_643),
.Y(n_762)
);

AO22x2_ASAP7_75t_L g763 ( 
.A1(n_647),
.A2(n_487),
.B1(n_5),
.B2(n_2),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_642),
.B(n_552),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_602),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_615),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_653),
.Y(n_767)
);

INVx4_ASAP7_75t_L g768 ( 
.A(n_639),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_650),
.B(n_599),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_616),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_615),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_655),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_606),
.B(n_404),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_650),
.B(n_406),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_699),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_732),
.B(n_657),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_720),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_SL g778 ( 
.A(n_702),
.B(n_657),
.Y(n_778)
);

INVx3_ASAP7_75t_L g779 ( 
.A(n_726),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_721),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_718),
.B(n_656),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_758),
.Y(n_782)
);

BUFx8_ASAP7_75t_L g783 ( 
.A(n_743),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_727),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_718),
.B(n_658),
.Y(n_785)
);

NAND2x1p5_ASAP7_75t_L g786 ( 
.A(n_749),
.B(n_659),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_731),
.Y(n_787)
);

OR2x6_ASAP7_75t_SL g788 ( 
.A(n_747),
.B(n_661),
.Y(n_788)
);

AOI22xp5_ASAP7_75t_L g789 ( 
.A1(n_709),
.A2(n_667),
.B1(n_675),
.B2(n_661),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_722),
.B(n_667),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_744),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_722),
.B(n_675),
.Y(n_792)
);

NAND2xp33_ASAP7_75t_L g793 ( 
.A(n_692),
.B(n_408),
.Y(n_793)
);

O2A1O1Ixp33_ASAP7_75t_L g794 ( 
.A1(n_695),
.A2(n_664),
.B(n_665),
.C(n_663),
.Y(n_794)
);

NOR3xp33_ASAP7_75t_L g795 ( 
.A(n_769),
.B(n_625),
.C(n_623),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_739),
.B(n_409),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_735),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_714),
.B(n_515),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_738),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_739),
.B(n_410),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_749),
.B(n_768),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_748),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_768),
.B(n_668),
.Y(n_803)
);

INVx2_ASAP7_75t_SL g804 ( 
.A(n_696),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_708),
.B(n_411),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_750),
.Y(n_806)
);

AND2x4_ASAP7_75t_L g807 ( 
.A(n_700),
.B(n_670),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_754),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_690),
.B(n_627),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_690),
.B(n_627),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_703),
.B(n_631),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_726),
.B(n_631),
.Y(n_812)
);

NAND2x1_ASAP7_75t_L g813 ( 
.A(n_736),
.B(n_609),
.Y(n_813)
);

OAI22xp5_ASAP7_75t_L g814 ( 
.A1(n_693),
.A2(n_557),
.B1(n_522),
.B2(n_560),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_745),
.B(n_651),
.Y(n_815)
);

CKINVDCx20_ASAP7_75t_R g816 ( 
.A(n_746),
.Y(n_816)
);

OAI221xp5_ASAP7_75t_L g817 ( 
.A1(n_693),
.A2(n_662),
.B1(n_651),
.B2(n_679),
.C(n_354),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_723),
.B(n_562),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_745),
.B(n_662),
.Y(n_819)
);

AND2x6_ASAP7_75t_SL g820 ( 
.A(n_685),
.B(n_540),
.Y(n_820)
);

AND2x4_ASAP7_75t_L g821 ( 
.A(n_700),
.B(n_679),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_708),
.B(n_415),
.Y(n_822)
);

OAI22xp33_ASAP7_75t_L g823 ( 
.A1(n_694),
.A2(n_565),
.B1(n_574),
.B2(n_562),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_703),
.B(n_609),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_L g825 ( 
.A(n_737),
.B(n_565),
.Y(n_825)
);

NAND2xp33_ASAP7_75t_L g826 ( 
.A(n_692),
.B(n_416),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_765),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_736),
.B(n_742),
.Y(n_828)
);

AND2x4_ASAP7_75t_L g829 ( 
.A(n_689),
.B(n_613),
.Y(n_829)
);

INVxp67_ASAP7_75t_L g830 ( 
.A(n_686),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_736),
.B(n_610),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_696),
.B(n_574),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_708),
.B(n_417),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_742),
.B(n_610),
.Y(n_834)
);

AOI22xp5_ASAP7_75t_L g835 ( 
.A1(n_734),
.A2(n_420),
.B1(n_424),
.B2(n_422),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_762),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_695),
.A2(n_421),
.B1(n_453),
.B2(n_399),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_692),
.B(n_425),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_767),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_760),
.B(n_585),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_772),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_756),
.Y(n_842)
);

AOI22xp33_ASAP7_75t_L g843 ( 
.A1(n_692),
.A2(n_421),
.B1(n_453),
.B2(n_399),
.Y(n_843)
);

HB1xp67_ASAP7_75t_L g844 ( 
.A(n_685),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_691),
.Y(n_845)
);

INVx2_ASAP7_75t_SL g846 ( 
.A(n_740),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_766),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_759),
.Y(n_848)
);

INVx2_ASAP7_75t_SL g849 ( 
.A(n_687),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_719),
.B(n_613),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_719),
.B(n_613),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_725),
.B(n_426),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_771),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_759),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_L g855 ( 
.A1(n_725),
.A2(n_421),
.B1(n_453),
.B2(n_399),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_733),
.B(n_433),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_737),
.B(n_438),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_687),
.B(n_439),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_688),
.B(n_440),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_774),
.B(n_585),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_760),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_758),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_758),
.Y(n_863)
);

BUFx6f_ASAP7_75t_SL g864 ( 
.A(n_741),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_688),
.B(n_441),
.Y(n_865)
);

A2O1A1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_697),
.A2(n_446),
.B(n_449),
.C(n_442),
.Y(n_866)
);

BUFx2_ASAP7_75t_L g867 ( 
.A(n_832),
.Y(n_867)
);

INVx6_ASAP7_75t_L g868 ( 
.A(n_783),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_SL g869 ( 
.A1(n_860),
.A2(n_586),
.B1(n_545),
.B2(n_540),
.Y(n_869)
);

BUFx4f_ASAP7_75t_L g870 ( 
.A(n_846),
.Y(n_870)
);

BUFx2_ASAP7_75t_L g871 ( 
.A(n_840),
.Y(n_871)
);

BUFx6f_ASAP7_75t_L g872 ( 
.A(n_782),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_847),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_775),
.Y(n_874)
);

INVx2_ASAP7_75t_SL g875 ( 
.A(n_829),
.Y(n_875)
);

HB1xp67_ASAP7_75t_L g876 ( 
.A(n_830),
.Y(n_876)
);

NOR3xp33_ASAP7_75t_SL g877 ( 
.A(n_823),
.B(n_717),
.C(n_366),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_L g878 ( 
.A1(n_848),
.A2(n_854),
.B1(n_849),
.B2(n_785),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_858),
.B(n_859),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_782),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_790),
.B(n_741),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_858),
.B(n_733),
.Y(n_882)
);

INVx3_ASAP7_75t_L g883 ( 
.A(n_779),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_782),
.Y(n_884)
);

OR2x6_ASAP7_75t_L g885 ( 
.A(n_844),
.B(n_685),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_859),
.B(n_734),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_792),
.B(n_586),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_780),
.Y(n_888)
);

INVx2_ASAP7_75t_SL g889 ( 
.A(n_829),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_853),
.Y(n_890)
);

XOR2xp5_ASAP7_75t_L g891 ( 
.A(n_816),
.B(n_646),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_779),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_787),
.Y(n_893)
);

BUFx2_ASAP7_75t_L g894 ( 
.A(n_798),
.Y(n_894)
);

INVx1_ASAP7_75t_SL g895 ( 
.A(n_842),
.Y(n_895)
);

OAI22xp5_ASAP7_75t_L g896 ( 
.A1(n_828),
.A2(n_697),
.B1(n_763),
.B2(n_751),
.Y(n_896)
);

AOI211xp5_ASAP7_75t_L g897 ( 
.A1(n_825),
.A2(n_717),
.B(n_774),
.C(n_753),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_861),
.B(n_789),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_797),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_807),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_865),
.B(n_734),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_778),
.B(n_751),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_799),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_865),
.B(n_734),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_781),
.B(n_773),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_781),
.B(n_785),
.Y(n_906)
);

OR2x6_ASAP7_75t_L g907 ( 
.A(n_814),
.B(n_729),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_845),
.B(n_752),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_806),
.Y(n_909)
);

NOR2xp33_ASAP7_75t_L g910 ( 
.A(n_818),
.B(n_545),
.Y(n_910)
);

O2A1O1Ixp5_ASAP7_75t_L g911 ( 
.A1(n_796),
.A2(n_773),
.B(n_701),
.C(n_711),
.Y(n_911)
);

NOR3xp33_ASAP7_75t_SL g912 ( 
.A(n_776),
.B(n_371),
.C(n_360),
.Y(n_912)
);

AOI22xp5_ASAP7_75t_L g913 ( 
.A1(n_828),
.A2(n_755),
.B1(n_763),
.B2(n_770),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_809),
.B(n_770),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_809),
.A2(n_755),
.B1(n_763),
.B2(n_770),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_808),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_836),
.Y(n_917)
);

OR2x6_ASAP7_75t_L g918 ( 
.A(n_804),
.B(n_764),
.Y(n_918)
);

INVx5_ASAP7_75t_L g919 ( 
.A(n_807),
.Y(n_919)
);

INVx3_ASAP7_75t_L g920 ( 
.A(n_862),
.Y(n_920)
);

OR2x2_ASAP7_75t_L g921 ( 
.A(n_821),
.B(n_757),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_R g922 ( 
.A(n_864),
.B(n_646),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_839),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_810),
.B(n_755),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_821),
.B(n_715),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_810),
.B(n_755),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_811),
.B(n_716),
.Y(n_927)
);

INVx3_ASAP7_75t_L g928 ( 
.A(n_863),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_841),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_811),
.B(n_716),
.Y(n_930)
);

NAND2xp33_ASAP7_75t_SL g931 ( 
.A(n_864),
.B(n_707),
.Y(n_931)
);

BUFx2_ASAP7_75t_L g932 ( 
.A(n_783),
.Y(n_932)
);

OR2x2_ASAP7_75t_L g933 ( 
.A(n_800),
.B(n_660),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_R g934 ( 
.A(n_820),
.B(n_660),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_803),
.B(n_715),
.Y(n_935)
);

OAI21xp33_ASAP7_75t_SL g936 ( 
.A1(n_906),
.A2(n_834),
.B(n_824),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_879),
.B(n_878),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_914),
.A2(n_801),
.B(n_905),
.Y(n_938)
);

OAI21x1_ASAP7_75t_L g939 ( 
.A1(n_911),
.A2(n_831),
.B(n_813),
.Y(n_939)
);

OAI21x1_ASAP7_75t_L g940 ( 
.A1(n_927),
.A2(n_831),
.B(n_824),
.Y(n_940)
);

OAI22xp5_ASAP7_75t_L g941 ( 
.A1(n_897),
.A2(n_843),
.B1(n_834),
.B2(n_837),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_882),
.B(n_850),
.Y(n_942)
);

OAI21xp5_ASAP7_75t_L g943 ( 
.A1(n_924),
.A2(n_851),
.B(n_850),
.Y(n_943)
);

OAI21xp5_ASAP7_75t_L g944 ( 
.A1(n_924),
.A2(n_926),
.B(n_927),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_874),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_897),
.B(n_888),
.Y(n_946)
);

OAI21xp5_ASAP7_75t_L g947 ( 
.A1(n_926),
.A2(n_851),
.B(n_866),
.Y(n_947)
);

AO21x1_ASAP7_75t_L g948 ( 
.A1(n_886),
.A2(n_857),
.B(n_856),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_930),
.A2(n_786),
.B(n_793),
.Y(n_949)
);

OAI21x1_ASAP7_75t_SL g950 ( 
.A1(n_913),
.A2(n_794),
.B(n_812),
.Y(n_950)
);

OAI21x1_ASAP7_75t_L g951 ( 
.A1(n_920),
.A2(n_786),
.B(n_815),
.Y(n_951)
);

OAI21x1_ASAP7_75t_L g952 ( 
.A1(n_920),
.A2(n_819),
.B(n_784),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_883),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_893),
.B(n_852),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_899),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_871),
.B(n_795),
.Y(n_956)
);

OAI21x1_ASAP7_75t_L g957 ( 
.A1(n_928),
.A2(n_791),
.B(n_777),
.Y(n_957)
);

OAI22xp5_ASAP7_75t_L g958 ( 
.A1(n_915),
.A2(n_913),
.B1(n_896),
.B2(n_877),
.Y(n_958)
);

OAI21x1_ASAP7_75t_L g959 ( 
.A1(n_928),
.A2(n_827),
.B(n_802),
.Y(n_959)
);

INVx3_ASAP7_75t_L g960 ( 
.A(n_883),
.Y(n_960)
);

O2A1O1Ixp5_ASAP7_75t_L g961 ( 
.A1(n_901),
.A2(n_838),
.B(n_822),
.C(n_833),
.Y(n_961)
);

NAND3xp33_ASAP7_75t_L g962 ( 
.A(n_910),
.B(n_855),
.C(n_595),
.Y(n_962)
);

OAI21xp5_ASAP7_75t_SL g963 ( 
.A1(n_869),
.A2(n_817),
.B(n_835),
.Y(n_963)
);

AOI21x1_ASAP7_75t_SL g964 ( 
.A1(n_904),
.A2(n_826),
.B(n_761),
.Y(n_964)
);

OAI21x1_ASAP7_75t_L g965 ( 
.A1(n_935),
.A2(n_712),
.B(n_710),
.Y(n_965)
);

OAI21x1_ASAP7_75t_L g966 ( 
.A1(n_892),
.A2(n_704),
.B(n_698),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_923),
.B(n_761),
.Y(n_967)
);

OAI21x1_ASAP7_75t_L g968 ( 
.A1(n_925),
.A2(n_704),
.B(n_698),
.Y(n_968)
);

OAI22x1_ASAP7_75t_L g969 ( 
.A1(n_887),
.A2(n_676),
.B1(n_666),
.B2(n_383),
.Y(n_969)
);

AOI21x1_ASAP7_75t_L g970 ( 
.A1(n_896),
.A2(n_805),
.B(n_730),
.Y(n_970)
);

CKINVDCx20_ASAP7_75t_R g971 ( 
.A(n_922),
.Y(n_971)
);

OAI21xp33_ASAP7_75t_L g972 ( 
.A1(n_898),
.A2(n_676),
.B(n_666),
.Y(n_972)
);

OAI21xp5_ASAP7_75t_L g973 ( 
.A1(n_915),
.A2(n_713),
.B(n_706),
.Y(n_973)
);

INVx4_ASAP7_75t_L g974 ( 
.A(n_872),
.Y(n_974)
);

OR2x2_ASAP7_75t_L g975 ( 
.A(n_894),
.B(n_933),
.Y(n_975)
);

O2A1O1Ixp5_ASAP7_75t_L g976 ( 
.A1(n_902),
.A2(n_713),
.B(n_706),
.C(n_728),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_919),
.B(n_715),
.Y(n_977)
);

OAI21x1_ASAP7_75t_L g978 ( 
.A1(n_873),
.A2(n_730),
.B(n_728),
.Y(n_978)
);

AO31x2_ASAP7_75t_L g979 ( 
.A1(n_903),
.A2(n_728),
.A3(n_730),
.B(n_724),
.Y(n_979)
);

OAI22x1_ASAP7_75t_L g980 ( 
.A1(n_891),
.A2(n_419),
.B1(n_423),
.B2(n_373),
.Y(n_980)
);

OAI22xp5_ASAP7_75t_L g981 ( 
.A1(n_929),
.A2(n_788),
.B1(n_443),
.B2(n_444),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_909),
.B(n_724),
.Y(n_982)
);

OAI21x1_ASAP7_75t_L g983 ( 
.A1(n_890),
.A2(n_917),
.B(n_916),
.Y(n_983)
);

AND2x2_ASAP7_75t_L g984 ( 
.A(n_908),
.B(n_431),
.Y(n_984)
);

OAI21x1_ASAP7_75t_SL g985 ( 
.A1(n_875),
.A2(n_64),
.B(n_61),
.Y(n_985)
);

OAI21xp5_ASAP7_75t_L g986 ( 
.A1(n_921),
.A2(n_456),
.B(n_450),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_867),
.B(n_454),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_907),
.A2(n_459),
.B1(n_473),
.B2(n_471),
.Y(n_988)
);

OAI21xp5_ASAP7_75t_L g989 ( 
.A1(n_912),
.A2(n_461),
.B(n_458),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_872),
.Y(n_990)
);

AND2x2_ASAP7_75t_L g991 ( 
.A(n_895),
.B(n_476),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_889),
.B(n_724),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_872),
.Y(n_993)
);

BUFx8_ASAP7_75t_L g994 ( 
.A(n_975),
.Y(n_994)
);

OAI21x1_ASAP7_75t_L g995 ( 
.A1(n_978),
.A2(n_881),
.B(n_880),
.Y(n_995)
);

AND2x4_ASAP7_75t_L g996 ( 
.A(n_945),
.B(n_919),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_955),
.Y(n_997)
);

OAI21xp33_ASAP7_75t_SL g998 ( 
.A1(n_946),
.A2(n_918),
.B(n_907),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_937),
.B(n_895),
.Y(n_999)
);

AOI22xp33_ASAP7_75t_L g1000 ( 
.A1(n_941),
.A2(n_907),
.B1(n_900),
.B2(n_918),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_983),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_954),
.Y(n_1002)
);

OAI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_936),
.A2(n_870),
.B(n_918),
.Y(n_1003)
);

OAI21x1_ASAP7_75t_L g1004 ( 
.A1(n_939),
.A2(n_884),
.B(n_880),
.Y(n_1004)
);

OAI21x1_ASAP7_75t_SL g1005 ( 
.A1(n_950),
.A2(n_931),
.B(n_884),
.Y(n_1005)
);

BUFx3_ASAP7_75t_L g1006 ( 
.A(n_971),
.Y(n_1006)
);

O2A1O1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_963),
.A2(n_876),
.B(n_885),
.C(n_932),
.Y(n_1007)
);

OAI21x1_ASAP7_75t_L g1008 ( 
.A1(n_964),
.A2(n_884),
.B(n_880),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_942),
.B(n_900),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_972),
.B(n_900),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_942),
.B(n_919),
.Y(n_1011)
);

OAI21x1_ASAP7_75t_L g1012 ( 
.A1(n_951),
.A2(n_705),
.B(n_870),
.Y(n_1012)
);

OAI21x1_ASAP7_75t_SL g1013 ( 
.A1(n_985),
.A2(n_74),
.B(n_65),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_982),
.Y(n_1014)
);

OAI21x1_ASAP7_75t_L g1015 ( 
.A1(n_952),
.A2(n_705),
.B(n_82),
.Y(n_1015)
);

INVx3_ASAP7_75t_L g1016 ( 
.A(n_979),
.Y(n_1016)
);

INVx1_ASAP7_75t_SL g1017 ( 
.A(n_991),
.Y(n_1017)
);

OAI21x1_ASAP7_75t_L g1018 ( 
.A1(n_966),
.A2(n_705),
.B(n_84),
.Y(n_1018)
);

OAI21x1_ASAP7_75t_L g1019 ( 
.A1(n_957),
.A2(n_705),
.B(n_86),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_977),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_959),
.Y(n_1021)
);

OAI21x1_ASAP7_75t_SL g1022 ( 
.A1(n_970),
.A2(n_885),
.B(n_88),
.Y(n_1022)
);

CKINVDCx8_ASAP7_75t_R g1023 ( 
.A(n_977),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_979),
.Y(n_1024)
);

OAI21x1_ASAP7_75t_L g1025 ( 
.A1(n_940),
.A2(n_89),
.B(n_79),
.Y(n_1025)
);

OAI21x1_ASAP7_75t_L g1026 ( 
.A1(n_965),
.A2(n_93),
.B(n_92),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_979),
.Y(n_1027)
);

OAI21x1_ASAP7_75t_L g1028 ( 
.A1(n_968),
.A2(n_97),
.B(n_96),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_953),
.Y(n_1029)
);

AOI221xp5_ASAP7_75t_L g1030 ( 
.A1(n_988),
.A2(n_934),
.B1(n_485),
.B2(n_481),
.C(n_496),
.Y(n_1030)
);

OAI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_938),
.A2(n_885),
.B(n_463),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_958),
.B(n_462),
.Y(n_1032)
);

NOR2xp67_ASAP7_75t_L g1033 ( 
.A(n_962),
.B(n_98),
.Y(n_1033)
);

BUFx3_ASAP7_75t_L g1034 ( 
.A(n_990),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_953),
.Y(n_1035)
);

OA21x2_ASAP7_75t_L g1036 ( 
.A1(n_944),
.A2(n_465),
.B(n_464),
.Y(n_1036)
);

OAI21x1_ASAP7_75t_L g1037 ( 
.A1(n_949),
.A2(n_101),
.B(n_100),
.Y(n_1037)
);

OAI21x1_ASAP7_75t_L g1038 ( 
.A1(n_944),
.A2(n_109),
.B(n_103),
.Y(n_1038)
);

AND2x4_ASAP7_75t_L g1039 ( 
.A(n_960),
.B(n_993),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_960),
.Y(n_1040)
);

AOI22xp33_ASAP7_75t_L g1041 ( 
.A1(n_941),
.A2(n_480),
.B1(n_495),
.B2(n_494),
.Y(n_1041)
);

OAI21x1_ASAP7_75t_L g1042 ( 
.A1(n_961),
.A2(n_112),
.B(n_111),
.Y(n_1042)
);

AO31x2_ASAP7_75t_L g1043 ( 
.A1(n_948),
.A2(n_3),
.A3(n_7),
.B(n_8),
.Y(n_1043)
);

OAI21x1_ASAP7_75t_L g1044 ( 
.A1(n_943),
.A2(n_115),
.B(n_114),
.Y(n_1044)
);

AOI22xp33_ASAP7_75t_L g1045 ( 
.A1(n_958),
.A2(n_479),
.B1(n_493),
.B2(n_492),
.Y(n_1045)
);

OAI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_963),
.A2(n_868),
.B1(n_488),
.B2(n_484),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_L g1047 ( 
.A1(n_943),
.A2(n_118),
.B(n_116),
.Y(n_1047)
);

HB1xp67_ASAP7_75t_L g1048 ( 
.A(n_1017),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_1009),
.B(n_984),
.Y(n_1049)
);

AOI22xp33_ASAP7_75t_SL g1050 ( 
.A1(n_1032),
.A2(n_988),
.B1(n_986),
.B2(n_1046),
.Y(n_1050)
);

AOI22xp33_ASAP7_75t_L g1051 ( 
.A1(n_1032),
.A2(n_969),
.B1(n_986),
.B2(n_956),
.Y(n_1051)
);

INVx4_ASAP7_75t_L g1052 ( 
.A(n_1020),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_997),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1009),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_999),
.A2(n_967),
.B1(n_987),
.B2(n_973),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_1002),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_1006),
.Y(n_1057)
);

OAI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_1023),
.A2(n_973),
.B1(n_981),
.B2(n_989),
.Y(n_1058)
);

AOI22xp33_ASAP7_75t_L g1059 ( 
.A1(n_1030),
.A2(n_980),
.B1(n_989),
.B2(n_981),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_1006),
.Y(n_1060)
);

BUFx10_ASAP7_75t_L g1061 ( 
.A(n_996),
.Y(n_1061)
);

AOI22xp33_ASAP7_75t_L g1062 ( 
.A1(n_1045),
.A2(n_947),
.B1(n_992),
.B2(n_868),
.Y(n_1062)
);

AOI221xp5_ASAP7_75t_L g1063 ( 
.A1(n_1007),
.A2(n_947),
.B1(n_467),
.B2(n_477),
.C(n_483),
.Y(n_1063)
);

OAI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_1000),
.A2(n_974),
.B1(n_478),
.B2(n_474),
.Y(n_1064)
);

AND2x4_ASAP7_75t_L g1065 ( 
.A(n_996),
.B(n_974),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_1020),
.Y(n_1066)
);

OAI22xp33_ASAP7_75t_L g1067 ( 
.A1(n_1011),
.A2(n_469),
.B1(n_468),
.B2(n_976),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1040),
.Y(n_1068)
);

OAI221xp5_ASAP7_75t_L g1069 ( 
.A1(n_998),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.C(n_11),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_1010),
.B(n_9),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_994),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_1031),
.A2(n_320),
.B(n_121),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1029),
.Y(n_1073)
);

OAI22xp5_ASAP7_75t_L g1074 ( 
.A1(n_1023),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_1074)
);

INVxp67_ASAP7_75t_L g1075 ( 
.A(n_994),
.Y(n_1075)
);

AOI22xp33_ASAP7_75t_SL g1076 ( 
.A1(n_994),
.A2(n_1003),
.B1(n_1005),
.B2(n_996),
.Y(n_1076)
);

INVxp67_ASAP7_75t_L g1077 ( 
.A(n_1034),
.Y(n_1077)
);

AOI22xp33_ASAP7_75t_L g1078 ( 
.A1(n_1041),
.A2(n_12),
.B1(n_13),
.B2(n_15),
.Y(n_1078)
);

AOI22xp33_ASAP7_75t_L g1079 ( 
.A1(n_1033),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_1036),
.A2(n_316),
.B(n_122),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_1014),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_1081)
);

AOI21xp33_ASAP7_75t_L g1082 ( 
.A1(n_1036),
.A2(n_18),
.B(n_19),
.Y(n_1082)
);

OAI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_1034),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_1029),
.Y(n_1084)
);

HB1xp67_ASAP7_75t_L g1085 ( 
.A(n_1039),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_1039),
.B(n_20),
.Y(n_1086)
);

AOI22xp33_ASAP7_75t_SL g1087 ( 
.A1(n_1005),
.A2(n_21),
.B1(n_24),
.B2(n_26),
.Y(n_1087)
);

CKINVDCx6p67_ASAP7_75t_R g1088 ( 
.A(n_1020),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_1039),
.B(n_26),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1020),
.B(n_27),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_1035),
.Y(n_1091)
);

AND2x4_ASAP7_75t_L g1092 ( 
.A(n_1035),
.B(n_120),
.Y(n_1092)
);

AOI221x1_ASAP7_75t_L g1093 ( 
.A1(n_1022),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.C(n_30),
.Y(n_1093)
);

OAI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_1036),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_1094)
);

BUFx6f_ASAP7_75t_L g1095 ( 
.A(n_995),
.Y(n_1095)
);

AOI22xp33_ASAP7_75t_L g1096 ( 
.A1(n_1013),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_1096)
);

INVx1_ASAP7_75t_SL g1097 ( 
.A(n_1024),
.Y(n_1097)
);

AOI22xp33_ASAP7_75t_L g1098 ( 
.A1(n_1022),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_1043),
.B(n_35),
.Y(n_1099)
);

INVxp67_ASAP7_75t_SL g1100 ( 
.A(n_995),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1043),
.Y(n_1101)
);

AOI22xp33_ASAP7_75t_L g1102 ( 
.A1(n_1044),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_1001),
.B(n_37),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1043),
.Y(n_1104)
);

INVx6_ASAP7_75t_L g1105 ( 
.A(n_1008),
.Y(n_1105)
);

OR2x6_ASAP7_75t_L g1106 ( 
.A(n_1038),
.B(n_123),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_1044),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_1107)
);

CKINVDCx6p67_ASAP7_75t_R g1108 ( 
.A(n_1043),
.Y(n_1108)
);

BUFx3_ASAP7_75t_L g1109 ( 
.A(n_1057),
.Y(n_1109)
);

AOI22xp33_ASAP7_75t_SL g1110 ( 
.A1(n_1058),
.A2(n_1038),
.B1(n_1047),
.B2(n_1037),
.Y(n_1110)
);

AOI22xp33_ASAP7_75t_L g1111 ( 
.A1(n_1050),
.A2(n_1047),
.B1(n_1037),
.B2(n_1001),
.Y(n_1111)
);

OAI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_1059),
.A2(n_1024),
.B1(n_1027),
.B2(n_1016),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1072),
.A2(n_1042),
.B(n_1019),
.Y(n_1113)
);

AOI22xp33_ASAP7_75t_L g1114 ( 
.A1(n_1058),
.A2(n_1021),
.B1(n_1025),
.B2(n_1042),
.Y(n_1114)
);

INVx2_ASAP7_75t_SL g1115 ( 
.A(n_1060),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1053),
.Y(n_1116)
);

OAI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_1051),
.A2(n_1027),
.B1(n_1016),
.B2(n_1021),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_1080),
.A2(n_1015),
.B(n_1012),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_1049),
.B(n_1043),
.Y(n_1119)
);

INVx4_ASAP7_75t_L g1120 ( 
.A(n_1066),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1056),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1068),
.Y(n_1122)
);

OAI221xp5_ASAP7_75t_L g1123 ( 
.A1(n_1063),
.A2(n_1016),
.B1(n_44),
.B2(n_48),
.C(n_49),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_1071),
.Y(n_1124)
);

OR2x2_ASAP7_75t_L g1125 ( 
.A(n_1054),
.B(n_1008),
.Y(n_1125)
);

AOI22xp33_ASAP7_75t_SL g1126 ( 
.A1(n_1069),
.A2(n_1025),
.B1(n_1026),
.B2(n_1028),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_1062),
.A2(n_1028),
.B1(n_1026),
.B2(n_1019),
.Y(n_1127)
);

AOI22xp33_ASAP7_75t_SL g1128 ( 
.A1(n_1074),
.A2(n_1070),
.B1(n_1094),
.B2(n_1083),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_1086),
.B(n_1004),
.Y(n_1129)
);

AOI22xp33_ASAP7_75t_L g1130 ( 
.A1(n_1078),
.A2(n_1004),
.B1(n_1015),
.B2(n_1018),
.Y(n_1130)
);

INVx4_ASAP7_75t_L g1131 ( 
.A(n_1066),
.Y(n_1131)
);

AOI22xp33_ASAP7_75t_SL g1132 ( 
.A1(n_1074),
.A2(n_1018),
.B1(n_1012),
.B2(n_48),
.Y(n_1132)
);

AND2x4_ASAP7_75t_L g1133 ( 
.A(n_1085),
.B(n_126),
.Y(n_1133)
);

OAI22xp33_ASAP7_75t_L g1134 ( 
.A1(n_1093),
.A2(n_42),
.B1(n_44),
.B2(n_49),
.Y(n_1134)
);

AOI22xp33_ASAP7_75t_L g1135 ( 
.A1(n_1079),
.A2(n_42),
.B1(n_50),
.B2(n_51),
.Y(n_1135)
);

OR2x2_ASAP7_75t_L g1136 ( 
.A(n_1048),
.B(n_50),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1073),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1055),
.A2(n_219),
.B(n_314),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1084),
.Y(n_1139)
);

BUFx4f_ASAP7_75t_SL g1140 ( 
.A(n_1088),
.Y(n_1140)
);

AOI22xp33_ASAP7_75t_SL g1141 ( 
.A1(n_1083),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_1141)
);

AOI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_1087),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_1142)
);

NAND3xp33_ASAP7_75t_L g1143 ( 
.A(n_1098),
.B(n_54),
.C(n_55),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1091),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_1066),
.Y(n_1145)
);

AOI22xp33_ASAP7_75t_L g1146 ( 
.A1(n_1096),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1097),
.Y(n_1147)
);

OR2x2_ASAP7_75t_L g1148 ( 
.A(n_1090),
.B(n_57),
.Y(n_1148)
);

AOI22xp33_ASAP7_75t_L g1149 ( 
.A1(n_1102),
.A2(n_58),
.B1(n_59),
.B2(n_127),
.Y(n_1149)
);

OAI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_1077),
.A2(n_132),
.B1(n_133),
.B2(n_138),
.Y(n_1150)
);

AOI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_1075),
.A2(n_142),
.B1(n_143),
.B2(n_145),
.Y(n_1151)
);

AOI22xp33_ASAP7_75t_L g1152 ( 
.A1(n_1107),
.A2(n_1081),
.B1(n_1099),
.B2(n_1103),
.Y(n_1152)
);

OAI322xp33_ASAP7_75t_L g1153 ( 
.A1(n_1081),
.A2(n_146),
.A3(n_150),
.B1(n_151),
.B2(n_152),
.C1(n_156),
.C2(n_157),
.Y(n_1153)
);

AOI221x1_ASAP7_75t_SL g1154 ( 
.A1(n_1082),
.A2(n_160),
.B1(n_163),
.B2(n_169),
.C(n_170),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_L g1155 ( 
.A(n_1089),
.B(n_171),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1092),
.B(n_175),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_1076),
.A2(n_176),
.B1(n_178),
.B2(n_180),
.Y(n_1157)
);

NAND3xp33_ASAP7_75t_L g1158 ( 
.A(n_1106),
.B(n_181),
.C(n_185),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1065),
.B(n_1092),
.Y(n_1159)
);

OAI21xp5_ASAP7_75t_SL g1160 ( 
.A1(n_1064),
.A2(n_1067),
.B(n_1065),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1052),
.Y(n_1161)
);

AOI21xp33_ASAP7_75t_L g1162 ( 
.A1(n_1106),
.A2(n_186),
.B(n_188),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1106),
.A2(n_189),
.B1(n_192),
.B2(n_193),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_1061),
.Y(n_1164)
);

OAI211xp5_ASAP7_75t_SL g1165 ( 
.A1(n_1101),
.A2(n_196),
.B(n_197),
.C(n_201),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1097),
.Y(n_1166)
);

AOI22xp33_ASAP7_75t_L g1167 ( 
.A1(n_1108),
.A2(n_203),
.B1(n_205),
.B2(n_207),
.Y(n_1167)
);

AOI22xp33_ASAP7_75t_SL g1168 ( 
.A1(n_1061),
.A2(n_209),
.B1(n_210),
.B2(n_211),
.Y(n_1168)
);

OAI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1052),
.A2(n_213),
.B1(n_214),
.B2(n_217),
.Y(n_1169)
);

AND2x4_ASAP7_75t_L g1170 ( 
.A(n_1095),
.B(n_218),
.Y(n_1170)
);

OA21x2_ASAP7_75t_L g1171 ( 
.A1(n_1104),
.A2(n_222),
.B(n_223),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1116),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1122),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1121),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1137),
.Y(n_1175)
);

INVxp67_ASAP7_75t_SL g1176 ( 
.A(n_1147),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1125),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1119),
.B(n_1129),
.Y(n_1178)
);

AOI22xp33_ASAP7_75t_L g1179 ( 
.A1(n_1143),
.A2(n_1095),
.B1(n_1105),
.B2(n_1100),
.Y(n_1179)
);

AO21x1_ASAP7_75t_L g1180 ( 
.A1(n_1134),
.A2(n_1105),
.B(n_1095),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1166),
.Y(n_1181)
);

BUFx2_ASAP7_75t_L g1182 ( 
.A(n_1118),
.Y(n_1182)
);

AND2x2_ASAP7_75t_L g1183 ( 
.A(n_1139),
.B(n_224),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1144),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1171),
.Y(n_1185)
);

OR2x2_ASAP7_75t_L g1186 ( 
.A(n_1117),
.B(n_227),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1148),
.B(n_229),
.Y(n_1187)
);

HB1xp67_ASAP7_75t_L g1188 ( 
.A(n_1112),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1171),
.Y(n_1189)
);

AND2x2_ASAP7_75t_L g1190 ( 
.A(n_1110),
.B(n_1111),
.Y(n_1190)
);

OR2x2_ASAP7_75t_L g1191 ( 
.A(n_1136),
.B(n_233),
.Y(n_1191)
);

HB1xp67_ASAP7_75t_L g1192 ( 
.A(n_1145),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1127),
.Y(n_1193)
);

BUFx3_ASAP7_75t_L g1194 ( 
.A(n_1164),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1158),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1152),
.B(n_234),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1128),
.B(n_236),
.Y(n_1197)
);

OR2x2_ASAP7_75t_L g1198 ( 
.A(n_1114),
.B(n_1159),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1161),
.Y(n_1199)
);

AND2x4_ASAP7_75t_L g1200 ( 
.A(n_1170),
.B(n_238),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1154),
.B(n_239),
.Y(n_1201)
);

OR2x2_ASAP7_75t_L g1202 ( 
.A(n_1130),
.B(n_1158),
.Y(n_1202)
);

OAI211xp5_ASAP7_75t_SL g1203 ( 
.A1(n_1141),
.A2(n_240),
.B(n_241),
.C(n_242),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1170),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1132),
.B(n_243),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1126),
.B(n_244),
.Y(n_1206)
);

INVxp67_ASAP7_75t_L g1207 ( 
.A(n_1115),
.Y(n_1207)
);

AND2x2_ASAP7_75t_L g1208 ( 
.A(n_1156),
.B(n_249),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_1154),
.B(n_250),
.Y(n_1209)
);

OR2x2_ASAP7_75t_L g1210 ( 
.A(n_1113),
.B(n_254),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1165),
.Y(n_1211)
);

AND2x2_ASAP7_75t_L g1212 ( 
.A(n_1120),
.B(n_1131),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1164),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1178),
.B(n_1120),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1180),
.A2(n_1143),
.B1(n_1123),
.B2(n_1142),
.Y(n_1215)
);

OAI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1197),
.A2(n_1146),
.B1(n_1135),
.B2(n_1149),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1172),
.Y(n_1217)
);

AOI22xp5_ASAP7_75t_SL g1218 ( 
.A1(n_1195),
.A2(n_1124),
.B1(n_1109),
.B2(n_1138),
.Y(n_1218)
);

OAI211xp5_ASAP7_75t_L g1219 ( 
.A1(n_1195),
.A2(n_1163),
.B(n_1151),
.C(n_1162),
.Y(n_1219)
);

AOI211xp5_ASAP7_75t_L g1220 ( 
.A1(n_1180),
.A2(n_1153),
.B(n_1157),
.C(n_1150),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1178),
.B(n_1131),
.Y(n_1221)
);

AOI33xp33_ASAP7_75t_L g1222 ( 
.A1(n_1193),
.A2(n_1168),
.A3(n_1167),
.B1(n_1133),
.B2(n_1153),
.B3(n_1160),
.Y(n_1222)
);

BUFx2_ASAP7_75t_L g1223 ( 
.A(n_1177),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1172),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1176),
.B(n_1160),
.Y(n_1225)
);

OAI221xp5_ASAP7_75t_L g1226 ( 
.A1(n_1202),
.A2(n_1155),
.B1(n_1169),
.B2(n_1164),
.C(n_1140),
.Y(n_1226)
);

INVx3_ASAP7_75t_L g1227 ( 
.A(n_1172),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1174),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1174),
.Y(n_1229)
);

INVxp67_ASAP7_75t_L g1230 ( 
.A(n_1192),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1174),
.Y(n_1231)
);

AOI211xp5_ASAP7_75t_L g1232 ( 
.A1(n_1202),
.A2(n_1133),
.B(n_256),
.C(n_257),
.Y(n_1232)
);

OAI211xp5_ASAP7_75t_L g1233 ( 
.A1(n_1201),
.A2(n_255),
.B(n_262),
.C(n_268),
.Y(n_1233)
);

AOI22xp5_ASAP7_75t_L g1234 ( 
.A1(n_1211),
.A2(n_269),
.B1(n_270),
.B2(n_274),
.Y(n_1234)
);

OAI221xp5_ASAP7_75t_L g1235 ( 
.A1(n_1187),
.A2(n_275),
.B1(n_276),
.B2(n_278),
.C(n_279),
.Y(n_1235)
);

INVx1_ASAP7_75t_SL g1236 ( 
.A(n_1212),
.Y(n_1236)
);

INVx3_ASAP7_75t_L g1237 ( 
.A(n_1199),
.Y(n_1237)
);

OR2x2_ASAP7_75t_L g1238 ( 
.A(n_1223),
.B(n_1193),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1236),
.B(n_1190),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1223),
.B(n_1214),
.Y(n_1240)
);

BUFx2_ASAP7_75t_L g1241 ( 
.A(n_1227),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_1237),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1228),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1214),
.B(n_1190),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1227),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1221),
.B(n_1177),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1228),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_1221),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1230),
.B(n_1181),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1231),
.Y(n_1250)
);

AND2x4_ASAP7_75t_L g1251 ( 
.A(n_1227),
.B(n_1177),
.Y(n_1251)
);

INVx3_ASAP7_75t_R g1252 ( 
.A(n_1232),
.Y(n_1252)
);

NOR2xp67_ASAP7_75t_L g1253 ( 
.A(n_1237),
.B(n_1231),
.Y(n_1253)
);

NAND2x1_ASAP7_75t_L g1254 ( 
.A(n_1253),
.B(n_1241),
.Y(n_1254)
);

INVx1_ASAP7_75t_SL g1255 ( 
.A(n_1238),
.Y(n_1255)
);

AND2x4_ASAP7_75t_L g1256 ( 
.A(n_1248),
.B(n_1213),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1243),
.Y(n_1257)
);

NAND2x1p5_ASAP7_75t_L g1258 ( 
.A(n_1248),
.B(n_1194),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1243),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1247),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1247),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1250),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1250),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1244),
.B(n_1239),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1238),
.B(n_1239),
.Y(n_1265)
);

AND2x2_ASAP7_75t_SL g1266 ( 
.A(n_1252),
.B(n_1225),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1266),
.A2(n_1218),
.B(n_1252),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1264),
.B(n_1244),
.Y(n_1268)
);

INVx1_ASAP7_75t_SL g1269 ( 
.A(n_1256),
.Y(n_1269)
);

HB1xp67_ASAP7_75t_L g1270 ( 
.A(n_1255),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1257),
.Y(n_1271)
);

AOI221xp5_ASAP7_75t_L g1272 ( 
.A1(n_1255),
.A2(n_1215),
.B1(n_1216),
.B2(n_1249),
.C(n_1220),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1259),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1260),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1265),
.B(n_1246),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_SL g1276 ( 
.A(n_1258),
.B(n_1222),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1265),
.B(n_1246),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1256),
.B(n_1240),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1261),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1262),
.B(n_1240),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1270),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1278),
.B(n_1263),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_SL g1283 ( 
.A1(n_1267),
.A2(n_1196),
.B1(n_1219),
.B2(n_1205),
.Y(n_1283)
);

A2O1A1Ixp33_ASAP7_75t_L g1284 ( 
.A1(n_1272),
.A2(n_1222),
.B(n_1254),
.C(n_1205),
.Y(n_1284)
);

NAND4xp25_ASAP7_75t_L g1285 ( 
.A(n_1276),
.B(n_1196),
.C(n_1179),
.D(n_1209),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1270),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1271),
.Y(n_1287)
);

AND2x2_ASAP7_75t_L g1288 ( 
.A(n_1268),
.B(n_1242),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1269),
.B(n_1251),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1274),
.Y(n_1290)
);

AOI222xp33_ASAP7_75t_L g1291 ( 
.A1(n_1284),
.A2(n_1276),
.B1(n_1206),
.B2(n_1273),
.C1(n_1279),
.C2(n_1235),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1283),
.B(n_1280),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_SL g1293 ( 
.A1(n_1281),
.A2(n_1226),
.B1(n_1206),
.B2(n_1233),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1282),
.B(n_1289),
.Y(n_1294)
);

OAI21xp33_ASAP7_75t_L g1295 ( 
.A1(n_1283),
.A2(n_1277),
.B(n_1275),
.Y(n_1295)
);

AOI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1285),
.A2(n_1286),
.B1(n_1287),
.B2(n_1290),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1294),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1296),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1292),
.B(n_1274),
.Y(n_1299)
);

XOR2x2_ASAP7_75t_L g1300 ( 
.A(n_1291),
.B(n_1285),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1295),
.B(n_1288),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1293),
.B(n_1207),
.Y(n_1302)
);

INVx1_ASAP7_75t_SL g1303 ( 
.A(n_1297),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1299),
.Y(n_1304)
);

NAND3xp33_ASAP7_75t_SL g1305 ( 
.A(n_1298),
.B(n_1234),
.C(n_1191),
.Y(n_1305)
);

INVxp67_ASAP7_75t_SL g1306 ( 
.A(n_1299),
.Y(n_1306)
);

NOR3xp33_ASAP7_75t_L g1307 ( 
.A(n_1301),
.B(n_1302),
.C(n_1300),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1297),
.Y(n_1308)
);

NAND3xp33_ASAP7_75t_L g1309 ( 
.A(n_1298),
.B(n_1210),
.C(n_1191),
.Y(n_1309)
);

AOI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1307),
.A2(n_1213),
.B1(n_1211),
.B2(n_1200),
.Y(n_1310)
);

OAI21xp33_ASAP7_75t_L g1311 ( 
.A1(n_1303),
.A2(n_1198),
.B(n_1208),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1308),
.B(n_1245),
.Y(n_1312)
);

OAI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1305),
.A2(n_1210),
.B1(n_1188),
.B2(n_1186),
.Y(n_1313)
);

NOR3xp33_ASAP7_75t_L g1314 ( 
.A(n_1306),
.B(n_1203),
.C(n_1208),
.Y(n_1314)
);

AOI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1309),
.A2(n_1200),
.B1(n_1212),
.B2(n_1194),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1310),
.A2(n_1304),
.B1(n_1200),
.B2(n_1198),
.Y(n_1316)
);

AOI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1311),
.A2(n_1200),
.B1(n_1194),
.B2(n_1199),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_1315),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1312),
.B(n_1241),
.Y(n_1319)
);

A2O1A1Ixp33_ASAP7_75t_L g1320 ( 
.A1(n_1314),
.A2(n_1313),
.B(n_1186),
.C(n_1185),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_1318),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1316),
.B(n_1245),
.Y(n_1322)
);

INVxp33_ASAP7_75t_L g1323 ( 
.A(n_1319),
.Y(n_1323)
);

HB1xp67_ASAP7_75t_L g1324 ( 
.A(n_1320),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1317),
.B(n_1251),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1323),
.A2(n_1183),
.B(n_1182),
.Y(n_1326)
);

AO22x2_ASAP7_75t_L g1327 ( 
.A1(n_1321),
.A2(n_1183),
.B1(n_1181),
.B2(n_1251),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1324),
.B(n_1237),
.Y(n_1328)
);

NAND3xp33_ASAP7_75t_L g1329 ( 
.A(n_1322),
.B(n_1173),
.C(n_1182),
.Y(n_1329)
);

AOI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1325),
.A2(n_1204),
.B1(n_1173),
.B2(n_1175),
.Y(n_1330)
);

NOR3xp33_ASAP7_75t_L g1331 ( 
.A(n_1328),
.B(n_1204),
.C(n_1184),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1327),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1329),
.Y(n_1333)
);

HB1xp67_ASAP7_75t_L g1334 ( 
.A(n_1326),
.Y(n_1334)
);

OR2x6_ASAP7_75t_L g1335 ( 
.A(n_1330),
.B(n_1184),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_1328),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1328),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1336),
.B(n_1175),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1337),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_SL g1340 ( 
.A(n_1339),
.B(n_1332),
.Y(n_1340)
);

AOI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1338),
.A2(n_1333),
.B1(n_1334),
.B2(n_1331),
.Y(n_1341)
);

CKINVDCx20_ASAP7_75t_R g1342 ( 
.A(n_1340),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1341),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1342),
.B(n_1335),
.Y(n_1344)
);

AOI21xp33_ASAP7_75t_L g1345 ( 
.A1(n_1343),
.A2(n_281),
.B(n_284),
.Y(n_1345)
);

AOI222xp33_ASAP7_75t_L g1346 ( 
.A1(n_1344),
.A2(n_1345),
.B1(n_1185),
.B2(n_1189),
.C1(n_1217),
.C2(n_1224),
.Y(n_1346)
);

AOI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1344),
.A2(n_1189),
.B(n_1185),
.Y(n_1347)
);

AOI22xp5_ASAP7_75t_SL g1348 ( 
.A1(n_1347),
.A2(n_286),
.B1(n_287),
.B2(n_293),
.Y(n_1348)
);

AOI322xp5_ASAP7_75t_L g1349 ( 
.A1(n_1346),
.A2(n_1229),
.A3(n_1184),
.B1(n_296),
.B2(n_298),
.C1(n_299),
.C2(n_303),
.Y(n_1349)
);

AOI221xp5_ASAP7_75t_L g1350 ( 
.A1(n_1348),
.A2(n_1229),
.B1(n_295),
.B2(n_306),
.C(n_307),
.Y(n_1350)
);

AOI211xp5_ASAP7_75t_L g1351 ( 
.A1(n_1350),
.A2(n_1349),
.B(n_308),
.C(n_309),
.Y(n_1351)
);


endmodule