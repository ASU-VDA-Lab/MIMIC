module fake_netlist_1_12401_n_29 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_29);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_29;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
INVx1_ASAP7_75t_L g12 ( .A(n_1), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_2), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_0), .Y(n_14) );
NAND2xp5_ASAP7_75t_SL g15 ( .A(n_1), .B(n_4), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_10), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_9), .Y(n_17) );
NOR2xp33_ASAP7_75t_L g18 ( .A(n_16), .B(n_0), .Y(n_18) );
OAI22xp5_ASAP7_75t_SL g19 ( .A1(n_12), .A2(n_13), .B1(n_14), .B2(n_17), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_18), .Y(n_20) );
OAI221xp5_ASAP7_75t_L g21 ( .A1(n_20), .A2(n_19), .B1(n_15), .B2(n_4), .C(n_3), .Y(n_21) );
OR2x2_ASAP7_75t_L g22 ( .A(n_21), .B(n_15), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
INVx2_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
NOR2xp33_ASAP7_75t_R g25 ( .A(n_23), .B(n_2), .Y(n_25) );
HB1xp67_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
XNOR2xp5_ASAP7_75t_L g27 ( .A(n_24), .B(n_3), .Y(n_27) );
HB1xp67_ASAP7_75t_L g28 ( .A(n_26), .Y(n_28) );
AOI322xp5_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_27), .A3(n_5), .B1(n_6), .B2(n_7), .C1(n_8), .C2(n_11), .Y(n_29) );
endmodule