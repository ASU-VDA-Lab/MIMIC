module fake_jpeg_26535_n_323 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_323);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_323;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx8_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_7),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_38),
.Y(n_58)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_33),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx4f_ASAP7_75t_SL g57 ( 
.A(n_37),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_27),
.B(n_7),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_8),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_43),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx5_ASAP7_75t_SL g56 ( 
.A(n_44),
.Y(n_56)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_45),
.B(n_50),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_31),
.C(n_29),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_37),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_16),
.B1(n_31),
.B2(n_29),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_48),
.A2(n_61),
.B1(n_30),
.B2(n_28),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_21),
.Y(n_73)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_18),
.B1(n_32),
.B2(n_22),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_55),
.A2(n_59),
.B1(n_28),
.B2(n_24),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_39),
.A2(n_33),
.B1(n_31),
.B2(n_29),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_36),
.A2(n_17),
.B1(n_23),
.B2(n_27),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_17),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_62),
.B(n_63),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_41),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_42),
.A2(n_16),
.B1(n_31),
.B2(n_29),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_64),
.A2(n_40),
.B1(n_28),
.B2(n_24),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_58),
.B(n_23),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_66),
.B(n_71),
.Y(n_126)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_68),
.A2(n_94),
.B1(n_98),
.B2(n_99),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_70),
.A2(n_96),
.B1(n_56),
.B2(n_53),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_61),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_57),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_72),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_74),
.B(n_82),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_57),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_76),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_59),
.A2(n_26),
.B1(n_18),
.B2(n_22),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_78),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_60),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_21),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_63),
.A2(n_26),
.B(n_18),
.C(n_32),
.Y(n_81)
);

AO21x1_ASAP7_75t_L g114 ( 
.A1(n_81),
.A2(n_85),
.B(n_86),
.Y(n_114)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_44),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_57),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_87),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_42),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_93),
.C(n_44),
.Y(n_112)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_90),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_54),
.Y(n_115)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_46),
.B(n_42),
.Y(n_93)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_L g107 ( 
.A1(n_95),
.A2(n_93),
.B1(n_83),
.B2(n_88),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_58),
.A2(n_26),
.B(n_32),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_97),
.A2(n_22),
.B(n_24),
.Y(n_110)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_47),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_54),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_104),
.B(n_124),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_74),
.A2(n_53),
.B1(n_40),
.B2(n_56),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_105),
.A2(n_107),
.B1(n_115),
.B2(n_117),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_108),
.A2(n_110),
.B(n_122),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_112),
.A2(n_67),
.B(n_86),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_113),
.A2(n_112),
.B1(n_124),
.B2(n_111),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_82),
.A2(n_53),
.B1(n_56),
.B2(n_50),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_91),
.A2(n_45),
.B1(n_44),
.B2(n_37),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_120),
.A2(n_99),
.B1(n_89),
.B2(n_98),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_37),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_83),
.B(n_37),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_106),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_129),
.B(n_134),
.Y(n_170)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_131),
.B(n_132),
.Y(n_164)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_77),
.Y(n_133)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_114),
.B(n_88),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_135),
.B(n_139),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_67),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_143),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_122),
.Y(n_160)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_108),
.A2(n_76),
.B(n_97),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_140),
.Y(n_185)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_141),
.B(n_142),
.Y(n_189)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_120),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_119),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_127),
.A2(n_96),
.B1(n_81),
.B2(n_78),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_144),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_123),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_145),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_114),
.B(n_25),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_146),
.B(n_149),
.Y(n_173)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_147),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_148),
.A2(n_156),
.B1(n_157),
.B2(n_116),
.Y(n_183)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_115),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_115),
.B(n_85),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_152),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_110),
.B(n_65),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_103),
.Y(n_153)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_153),
.Y(n_163)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_113),
.Y(n_154)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_154),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_126),
.B(n_127),
.Y(n_155)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_155),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_128),
.A2(n_68),
.B1(n_94),
.B2(n_65),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_126),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_158),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_122),
.B(n_90),
.Y(n_159)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_159),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_160),
.B(n_178),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_108),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g210 ( 
.A1(n_166),
.A2(n_176),
.B(n_183),
.Y(n_210)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_129),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_175),
.B(n_181),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_134),
.B(n_108),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_138),
.B(n_122),
.C(n_118),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_177),
.B(n_159),
.C(n_136),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_150),
.B(n_156),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_140),
.B(n_100),
.Y(n_179)
);

FAx1_ASAP7_75t_SL g205 ( 
.A(n_179),
.B(n_177),
.CI(n_186),
.CON(n_205),
.SN(n_205)
);

AND2x6_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_11),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_182),
.Y(n_194)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_145),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_148),
.Y(n_182)
);

AOI21x1_ASAP7_75t_L g184 ( 
.A1(n_151),
.A2(n_43),
.B(n_69),
.Y(n_184)
);

OAI21xp33_ASAP7_75t_L g217 ( 
.A1(n_184),
.A2(n_186),
.B(n_170),
.Y(n_217)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_143),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_187),
.B(n_190),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_154),
.A2(n_128),
.B1(n_125),
.B2(n_109),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_188),
.A2(n_142),
.B1(n_132),
.B2(n_141),
.Y(n_195)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_147),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_153),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_191),
.Y(n_197)
);

AND2x6_ASAP7_75t_L g193 ( 
.A(n_155),
.B(n_137),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_193),
.B(n_12),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_195),
.A2(n_215),
.B1(n_183),
.B2(n_166),
.Y(n_226)
);

OAI32xp33_ASAP7_75t_L g198 ( 
.A1(n_170),
.A2(n_149),
.A3(n_135),
.B1(n_139),
.B2(n_131),
.Y(n_198)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_198),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_212),
.C(n_179),
.Y(n_222)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_189),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_202),
.Y(n_238)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_164),
.Y(n_202)
);

XNOR2x1_ASAP7_75t_L g203 ( 
.A(n_178),
.B(n_136),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_203),
.A2(n_205),
.B(n_209),
.Y(n_235)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_165),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_207),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_162),
.B(n_146),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_172),
.B(n_144),
.Y(n_208)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_208),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_161),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_185),
.A2(n_130),
.B(n_121),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_211),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_160),
.B(n_130),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_188),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_213),
.B(n_214),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_167),
.A2(n_109),
.B1(n_103),
.B2(n_125),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_172),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_218),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_184),
.Y(n_233)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_174),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_169),
.B(n_101),
.Y(n_219)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_219),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_163),
.Y(n_220)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_220),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_173),
.B(n_101),
.Y(n_221)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_221),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_222),
.B(n_238),
.C(n_230),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_176),
.C(n_166),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_236),
.C(n_243),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_201),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_225),
.B(n_9),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_226),
.A2(n_228),
.B1(n_231),
.B2(n_244),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_211),
.A2(n_192),
.B1(n_185),
.B2(n_193),
.Y(n_227)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_227),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_213),
.A2(n_192),
.B1(n_176),
.B2(n_168),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_218),
.A2(n_173),
.B1(n_180),
.B2(n_171),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_233),
.A2(n_210),
.B(n_221),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_208),
.A2(n_171),
.B1(n_92),
.B2(n_84),
.Y(n_234)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_234),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_75),
.C(n_37),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_199),
.B(n_37),
.C(n_43),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_195),
.A2(n_216),
.B1(n_200),
.B2(n_194),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_229),
.B(n_196),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_246),
.Y(n_276)
);

XNOR2x1_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_203),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_247),
.A2(n_233),
.B1(n_223),
.B2(n_234),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_249),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_222),
.B(n_212),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_210),
.C(n_202),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_253),
.C(n_258),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_198),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_255),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_219),
.C(n_209),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_235),
.B(n_205),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_227),
.B(n_205),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_262),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_239),
.A2(n_197),
.B1(n_204),
.B2(n_215),
.Y(n_257)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_257),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_25),
.C(n_43),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_30),
.C(n_20),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_263),
.Y(n_266)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_260),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_228),
.B(n_21),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_238),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_20),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_254),
.A2(n_223),
.B1(n_230),
.B2(n_237),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_268),
.A2(n_269),
.B1(n_278),
.B2(n_19),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_245),
.A2(n_241),
.B(n_233),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_270),
.A2(n_263),
.B(n_256),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_261),
.A2(n_226),
.B(n_242),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_271),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_253),
.A2(n_240),
.B(n_225),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_273),
.Y(n_290)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_277),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_247),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_258),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_280),
.B(n_8),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_281),
.A2(n_288),
.B(n_10),
.Y(n_297)
);

AO22x1_ASAP7_75t_L g282 ( 
.A1(n_271),
.A2(n_251),
.B1(n_250),
.B2(n_249),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_289),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_250),
.C(n_259),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_287),
.C(n_291),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_276),
.A2(n_267),
.B1(n_279),
.B2(n_268),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_284),
.A2(n_293),
.B1(n_14),
.B2(n_13),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_269),
.A2(n_20),
.B1(n_19),
.B2(n_9),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_14),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_265),
.B(n_19),
.C(n_8),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_266),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_273),
.B(n_19),
.C(n_6),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_290),
.B(n_272),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_296),
.Y(n_306)
);

NAND3xp33_ASAP7_75t_L g296 ( 
.A(n_289),
.B(n_278),
.C(n_272),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_299),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_283),
.B(n_275),
.C(n_274),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_285),
.B(n_274),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_300),
.B(n_304),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_275),
.C(n_10),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_301),
.B(n_302),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_303),
.B(n_291),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_13),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_308),
.B(n_309),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_298),
.A2(n_290),
.B(n_286),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_296),
.A2(n_282),
.B1(n_1),
.B2(n_2),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_311),
.Y(n_314)
);

AOI322xp5_ASAP7_75t_L g312 ( 
.A1(n_295),
.A2(n_12),
.A3(n_11),
.B1(n_10),
.B2(n_4),
.C1(n_0),
.C2(n_3),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_312),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_299),
.C(n_295),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_313),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_316),
.A2(n_317),
.B(n_310),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_5),
.C(n_3),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_318),
.B(n_308),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_320),
.A2(n_315),
.B(n_319),
.Y(n_321)
);

AOI321xp33_ASAP7_75t_L g322 ( 
.A1(n_321),
.A2(n_311),
.A3(n_314),
.B1(n_307),
.B2(n_4),
.C(n_5),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_4),
.Y(n_323)
);


endmodule