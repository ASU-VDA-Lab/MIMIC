module real_jpeg_30321_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_578;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_605;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_611;
wire n_393;
wire n_489;
wire n_221;
wire n_104;
wire n_153;
wire n_599;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_325;
wire n_594;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_586;
wire n_572;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_613;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_608;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_597;
wire n_42;
wire n_268;
wire n_313;
wire n_609;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_568;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g163 ( 
.A(n_0),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_0),
.Y(n_267)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_0),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_1),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_2),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_2),
.B(n_154),
.Y(n_254)
);

NAND2x1_ASAP7_75t_L g273 ( 
.A(n_2),
.B(n_274),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_2),
.B(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_2),
.B(n_354),
.Y(n_353)
);

NAND3xp33_ASAP7_75t_L g459 ( 
.A(n_2),
.B(n_162),
.C(n_460),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_2),
.B(n_465),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_2),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_2),
.B(n_460),
.Y(n_480)
);

NAND3xp33_ASAP7_75t_SL g543 ( 
.A(n_2),
.B(n_162),
.C(n_460),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_3),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_4),
.Y(n_75)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_4),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_5),
.A2(n_19),
.B(n_20),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_6),
.Y(n_128)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_6),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g462 ( 
.A(n_6),
.Y(n_462)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_6),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_7),
.B(n_213),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_7),
.B(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_7),
.B(n_311),
.Y(n_310)
);

AND2x2_ASAP7_75t_SL g332 ( 
.A(n_7),
.B(n_333),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_7),
.B(n_422),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g450 ( 
.A(n_7),
.B(n_216),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_7),
.B(n_478),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_7),
.B(n_518),
.Y(n_517)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_8),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_8),
.B(n_356),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_8),
.B(n_427),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_8),
.B(n_448),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_8),
.B(n_494),
.Y(n_493)
);

BUFx2_ASAP7_75t_R g33 ( 
.A(n_9),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_9),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_9),
.B(n_78),
.Y(n_77)
);

AND2x2_ASAP7_75t_SL g101 ( 
.A(n_9),
.B(n_102),
.Y(n_101)
);

AND2x4_ASAP7_75t_L g140 ( 
.A(n_9),
.B(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_9),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_9),
.B(n_228),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_9),
.B(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_10),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_10),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_10),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_11),
.Y(n_337)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_12),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_13),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_13),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_13),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_14),
.B(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

BUFx24_ASAP7_75t_L g96 ( 
.A(n_14),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_14),
.B(n_216),
.Y(n_215)
);

AOI22x1_ASAP7_75t_L g338 ( 
.A1(n_14),
.A2(n_15),
.B1(n_339),
.B2(n_342),
.Y(n_338)
);

NAND2x1_ASAP7_75t_L g263 ( 
.A(n_15),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_15),
.B(n_387),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_15),
.B(n_396),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_15),
.B(n_419),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_15),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_15),
.B(n_489),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_15),
.B(n_521),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g29 ( 
.A(n_16),
.B(n_30),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_16),
.B(n_41),
.Y(n_40)
);

AND2x2_ASAP7_75t_SL g72 ( 
.A(n_16),
.B(n_73),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_16),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_16),
.B(n_121),
.Y(n_120)
);

AND2x2_ASAP7_75t_SL g125 ( 
.A(n_16),
.B(n_126),
.Y(n_125)
);

AND2x4_ASAP7_75t_L g152 ( 
.A(n_16),
.B(n_109),
.Y(n_152)
);

AND2x2_ASAP7_75t_SL g162 ( 
.A(n_16),
.B(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_17),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_17),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_17),
.B(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_17),
.B(n_317),
.Y(n_316)
);

AND2x2_ASAP7_75t_SL g327 ( 
.A(n_17),
.B(n_328),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_17),
.B(n_380),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_614),
.Y(n_20)
);

A2O1A1O1Ixp25_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_129),
.B(n_286),
.C(n_594),
.D(n_613),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_181),
.Y(n_22)
);

OAI211xp5_ASAP7_75t_L g594 ( 
.A1(n_23),
.A2(n_595),
.B(n_598),
.C(n_600),
.Y(n_594)
);

NOR2xp67_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_113),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_88),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g599 ( 
.A(n_25),
.B(n_88),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_54),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g612 ( 
.A(n_26),
.B(n_54),
.C(n_88),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_44),
.C(n_49),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_27),
.B(n_91),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_32),
.C(n_40),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_28),
.A2(n_29),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_28),
.A2(n_29),
.B1(n_32),
.B2(n_176),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_28),
.B(n_125),
.C(n_129),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_28),
.A2(n_29),
.B1(n_301),
.B2(n_414),
.Y(n_413)
);

CKINVDCx11_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_29),
.B(n_301),
.C(n_304),
.Y(n_300)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_31),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_31),
.Y(n_515)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_32),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g606 ( 
.A1(n_32),
.A2(n_176),
.B1(n_607),
.B2(n_608),
.Y(n_606)
);

NAND2x1_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_34),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_38),
.Y(n_165)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_38),
.Y(n_356)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_39),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_40),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_40),
.A2(n_61),
.B1(n_70),
.B2(n_71),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_40),
.A2(n_61),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_40),
.A2(n_61),
.B1(n_310),
.B2(n_315),
.Y(n_309)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_44),
.B(n_49),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_46),
.Y(n_44)
);

NOR2x1_ASAP7_75t_R g105 ( 
.A(n_45),
.B(n_106),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g223 ( 
.A(n_45),
.B(n_224),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_45),
.B(n_224),
.Y(n_232)
);

INVx4_ASAP7_75t_SL g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_52),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_53),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_53),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_76),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_60),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_56),
.B(n_76),
.C(n_611),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_58),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

HB1xp67_ASAP7_75t_L g611 ( 
.A(n_60),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.C(n_70),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_61),
.B(n_310),
.C(n_316),
.Y(n_357)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_63),
.B(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_64),
.B(n_125),
.C(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_65),
.B(n_133),
.Y(n_204)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_69),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_69),
.Y(n_429)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_70),
.A2(n_71),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_70),
.A2(n_71),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_71),
.B(n_82),
.C(n_86),
.Y(n_605)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_72),
.Y(n_71)
);

MAJx2_ASAP7_75t_L g262 ( 
.A(n_72),
.B(n_263),
.C(n_265),
.Y(n_262)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_73),
.Y(n_449)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx4_ASAP7_75t_L g354 ( 
.A(n_74),
.Y(n_354)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_75),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_75),
.Y(n_420)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_80),
.B1(n_86),
.B2(n_87),
.Y(n_76)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_77),
.Y(n_86)
);

XOR2x2_ASAP7_75t_L g138 ( 
.A(n_77),
.B(n_139),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_77),
.B(n_144),
.C(n_146),
.Y(n_177)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

MAJx2_ASAP7_75t_L g209 ( 
.A(n_81),
.B(n_210),
.C(n_214),
.Y(n_209)
);

OAI22xp33_ASAP7_75t_SL g608 ( 
.A1(n_81),
.A2(n_82),
.B1(n_151),
.B2(n_152),
.Y(n_608)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_82),
.B(n_258),
.Y(n_257)
);

NOR3xp33_ASAP7_75t_SL g613 ( 
.A(n_82),
.B(n_152),
.C(n_176),
.Y(n_613)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_85),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_92),
.C(n_110),
.Y(n_88)
);

INVxp33_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XOR2x1_ASAP7_75t_L g179 ( 
.A(n_90),
.B(n_180),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_93),
.B(n_111),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_101),
.C(n_105),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_94),
.A2(n_95),
.B1(n_101),
.B2(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

AND2x4_ASAP7_75t_L g133 ( 
.A(n_96),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_96),
.B(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_96),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_96),
.B(n_393),
.Y(n_392)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_101),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_101),
.B(n_162),
.C(n_227),
.Y(n_226)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_102),
.Y(n_303)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_103),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

XOR2x1_ASAP7_75t_L g168 ( 
.A(n_105),
.B(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_113),
.B(n_599),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_171),
.C(n_179),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_114),
.B(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI21xp33_ASAP7_75t_L g187 ( 
.A1(n_115),
.A2(n_172),
.B(n_179),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_148),
.C(n_167),
.Y(n_115)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_116),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_131),
.C(n_138),
.Y(n_116)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_117),
.Y(n_283)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_125),
.B1(n_129),
.B2(n_130),
.Y(n_119)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_120),
.Y(n_129)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_122),
.Y(n_264)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_125),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_125),
.B(n_265),
.Y(n_377)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_130),
.B(n_204),
.Y(n_203)
);

XOR2x2_ASAP7_75t_L g456 ( 
.A(n_130),
.B(n_265),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_131),
.A2(n_132),
.B1(n_138),
.B2(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_136),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g282 ( 
.A(n_138),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_144),
.B1(n_146),
.B2(n_147),
.Y(n_139)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_140),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_140),
.A2(n_146),
.B1(n_253),
.B2(n_254),
.Y(n_350)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_142),
.Y(n_424)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_143),
.Y(n_307)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_144),
.Y(n_147)
);

NOR3xp33_ASAP7_75t_L g247 ( 
.A(n_146),
.B(n_248),
.C(n_252),
.Y(n_247)
);

OAI21xp33_ASAP7_75t_L g255 ( 
.A1(n_146),
.A2(n_248),
.B(n_252),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_148),
.A2(n_149),
.B1(n_168),
.B2(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

OA21x2_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_157),
.B(n_166),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_153),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_153),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_151),
.A2(n_152),
.B1(n_153),
.B2(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_151),
.B(n_232),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_151),
.A2(n_152),
.B1(n_223),
.B2(n_232),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

A2O1A1Ixp33_ASAP7_75t_SL g222 ( 
.A1(n_152),
.A2(n_223),
.B(n_226),
.C(n_231),
.Y(n_222)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_153),
.Y(n_221)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_157),
.B(n_220),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_162),
.C(n_164),
.Y(n_157)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_158),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g402 ( 
.A1(n_158),
.A2(n_206),
.B1(n_352),
.B2(n_353),
.Y(n_402)
);

OR2x2_ASAP7_75t_SL g158 ( 
.A(n_159),
.B(n_161),
.Y(n_158)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_159),
.Y(n_466)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx4_ASAP7_75t_L g492 ( 
.A(n_160),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_162),
.B(n_164),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_162),
.A2(n_227),
.B1(n_242),
.B2(n_243),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_162),
.Y(n_243)
);

XNOR2x2_ASAP7_75t_L g479 ( 
.A(n_162),
.B(n_480),
.Y(n_479)
);

INVx8_ASAP7_75t_L g394 ( 
.A(n_163),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_168),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_170),
.A2(n_241),
.B(n_244),
.Y(n_240)
);

OAI211xp5_ASAP7_75t_L g244 ( 
.A1(n_170),
.A2(n_227),
.B(n_243),
.C(n_245),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_172),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_172),
.A2(n_179),
.B1(n_185),
.B2(n_186),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_177),
.C(n_178),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_178),
.Y(n_198)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_179),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_233),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g595 ( 
.A1(n_182),
.A2(n_596),
.B(n_597),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_190),
.Y(n_182)
);

NOR2xp67_ASAP7_75t_L g597 ( 
.A(n_183),
.B(n_190),
.Y(n_597)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_187),
.B(n_188),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_196),
.C(n_199),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_192),
.B(n_197),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_195),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVxp67_ASAP7_75t_SL g199 ( 
.A(n_200),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_200),
.B(n_235),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_219),
.C(n_222),
.Y(n_200)
);

XOR2x1_ASAP7_75t_SL g284 ( 
.A(n_201),
.B(n_285),
.Y(n_284)
);

MAJx2_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_205),
.C(n_208),
.Y(n_201)
);

INVxp33_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g568 ( 
.A(n_203),
.B(n_209),
.Y(n_568)
);

XOR2xp5_ASAP7_75t_L g567 ( 
.A(n_205),
.B(n_568),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

MAJx2_ASAP7_75t_L g351 ( 
.A(n_206),
.B(n_352),
.C(n_355),
.Y(n_351)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_211),
.A2(n_212),
.B1(n_214),
.B2(n_215),
.Y(n_258)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g331 ( 
.A(n_218),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_219),
.B(n_222),
.Y(n_285)
);

INVx5_ASAP7_75t_SL g224 ( 
.A(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_226),
.B(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_227),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_227),
.B(n_243),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_227),
.B(n_296),
.Y(n_295)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_230),
.Y(n_251)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_230),
.Y(n_318)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_230),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

NOR2xp67_ASAP7_75t_L g596 ( 
.A(n_234),
.B(n_236),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_279),
.C(n_284),
.Y(n_236)
);

INVxp33_ASAP7_75t_SL g237 ( 
.A(n_238),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g576 ( 
.A(n_238),
.B(n_280),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_259),
.C(n_276),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g564 ( 
.A(n_239),
.B(n_565),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_246),
.C(n_256),
.Y(n_239)
);

INVxp67_ASAP7_75t_SL g366 ( 
.A(n_240),
.Y(n_366)
);

XNOR2x1_ASAP7_75t_L g415 ( 
.A(n_242),
.B(n_296),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_246),
.B(n_257),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_253),
.B(n_255),
.Y(n_246)
);

NOR2xp67_ASAP7_75t_L g349 ( 
.A(n_248),
.B(n_252),
.Y(n_349)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_249),
.Y(n_248)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g565 ( 
.A(n_260),
.B(n_277),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_268),
.C(n_273),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XNOR2x1_ASAP7_75t_L g362 ( 
.A(n_262),
.B(n_363),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_263),
.B(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_265),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_266),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g341 ( 
.A(n_267),
.Y(n_341)
);

INVxp67_ASAP7_75t_SL g268 ( 
.A(n_269),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_269),
.A2(n_270),
.B1(n_273),
.B2(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g364 ( 
.A(n_273),
.Y(n_364)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_275),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_283),
.Y(n_280)
);

XNOR2x1_ASAP7_75t_L g575 ( 
.A(n_284),
.B(n_576),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_585),
.Y(n_286)
);

NAND3xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_435),
.C(n_560),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_407),
.Y(n_288)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_289),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_369),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g589 ( 
.A(n_290),
.B(n_369),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_345),
.B2(n_368),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_291),
.B(n_579),
.C(n_580),
.Y(n_578)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_292),
.Y(n_291)
);

MAJx2_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_320),
.C(n_324),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_293),
.B(n_371),
.Y(n_370)
);

AO21x1_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_308),
.B(n_319),
.Y(n_293)
);

NAND2xp33_ASAP7_75t_SL g294 ( 
.A(n_295),
.B(n_300),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_295),
.B(n_300),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_295),
.B(n_300),
.Y(n_432)
);

NOR2x1_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_297),
.B(n_505),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_297),
.B(n_512),
.Y(n_511)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_301),
.Y(n_414)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

XNOR2x1_ASAP7_75t_SL g412 ( 
.A(n_304),
.B(n_413),
.Y(n_412)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_SL g306 ( 
.A(n_307),
.Y(n_306)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_307),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_308),
.B(n_432),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_309),
.B(n_316),
.Y(n_308)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_310),
.Y(n_315)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

BUFx4f_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_320),
.B(n_324),
.Y(n_371)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_326),
.B1(n_338),
.B2(n_344),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_332),
.Y(n_326)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_327),
.Y(n_360)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx6_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_332),
.Y(n_361)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx5_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_338),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_338),
.B(n_360),
.C(n_361),
.Y(n_359)
);

INVx3_ASAP7_75t_SL g339 ( 
.A(n_340),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_340),
.B(n_475),
.Y(n_474)
);

INVx8_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

BUFx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_344),
.A2(n_392),
.B(n_395),
.Y(n_391)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_345),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_365),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_346),
.Y(n_580)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_358),
.Y(n_346)
);

INVxp33_ASAP7_75t_SL g570 ( 
.A(n_347),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_351),
.C(n_357),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_348),
.B(n_351),
.Y(n_406)
);

XNOR2x1_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_355),
.Y(n_401)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_357),
.Y(n_405)
);

XNOR2x1_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_362),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_359),
.Y(n_571)
);

INVxp33_ASAP7_75t_L g572 ( 
.A(n_362),
.Y(n_572)
);

HB1xp67_ASAP7_75t_L g579 ( 
.A(n_365),
.Y(n_579)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_367),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_372),
.C(n_403),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_370),
.B(n_434),
.Y(n_433)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_373),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_373),
.B(n_404),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_391),
.C(n_399),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_375),
.B(n_410),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_376),
.B(n_378),
.C(n_384),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g544 ( 
.A1(n_376),
.A2(n_377),
.B1(n_545),
.B2(n_546),
.Y(n_544)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_378),
.A2(n_379),
.B1(n_385),
.B2(n_386),
.Y(n_546)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_383),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_SL g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx2_ASAP7_75t_SL g389 ( 
.A(n_390),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_391),
.B(n_400),
.Y(n_410)
);

INVx5_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_402),
.Y(n_400)
);

INVxp33_ASAP7_75t_SL g403 ( 
.A(n_404),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_406),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_433),
.Y(n_407)
);

OR2x2_ASAP7_75t_L g588 ( 
.A(n_408),
.B(n_433),
.Y(n_588)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_411),
.C(n_430),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_409),
.B(n_553),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_L g553 ( 
.A1(n_411),
.A2(n_431),
.B1(n_554),
.B2(n_555),
.Y(n_553)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_411),
.Y(n_555)
);

MAJx2_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_415),
.C(n_416),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_412),
.B(n_537),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_L g537 ( 
.A1(n_415),
.A2(n_416),
.B1(n_538),
.B2(n_539),
.Y(n_537)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_415),
.Y(n_539)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_416),
.Y(n_538)
);

MAJx2_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_421),
.C(n_425),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_417),
.A2(n_418),
.B1(n_425),
.B2(n_426),
.Y(n_444)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_421),
.B(n_444),
.Y(n_443)
);

INVx3_ASAP7_75t_SL g422 ( 
.A(n_423),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_431),
.Y(n_554)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_436),
.A2(n_550),
.B(n_559),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_438),
.A2(n_533),
.B(n_549),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_439),
.A2(n_481),
.B(n_532),
.Y(n_438)
);

NAND3xp33_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_467),
.C(n_468),
.Y(n_439)
);

AOI21xp33_ASAP7_75t_SL g532 ( 
.A1(n_440),
.A2(n_467),
.B(n_468),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_454),
.Y(n_440)
);

INVxp67_ASAP7_75t_SL g441 ( 
.A(n_442),
.Y(n_441)
);

NAND2xp33_ASAP7_75t_L g467 ( 
.A(n_442),
.B(n_455),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_445),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_443),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_445),
.B(n_454),
.C(n_548),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_450),
.C(n_451),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_446),
.A2(n_447),
.B1(n_450),
.B2(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

CKINVDCx16_ASAP7_75t_R g471 ( 
.A(n_450),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_451),
.B(n_470),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_453),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_452),
.B(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_457),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_456),
.B(n_463),
.C(n_543),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_R g558 ( 
.A(n_456),
.B(n_463),
.C(n_543),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_458),
.A2(n_459),
.B1(n_463),
.B2(n_464),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx4_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

BUFx2_ASAP7_75t_L g478 ( 
.A(n_462),
.Y(n_478)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_472),
.C(n_479),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_SL g495 ( 
.A(n_469),
.B(n_496),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_472),
.A2(n_473),
.B1(n_479),
.B2(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_476),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_474),
.A2(n_476),
.B1(n_477),
.B2(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_474),
.Y(n_486)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_479),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_L g481 ( 
.A1(n_482),
.A2(n_498),
.B(n_531),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_495),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_483),
.B(n_495),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_487),
.C(n_493),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_484),
.A2(n_485),
.B1(n_527),
.B2(n_528),
.Y(n_526)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_SL g527 ( 
.A(n_488),
.B(n_493),
.Y(n_527)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_499),
.A2(n_525),
.B(n_530),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_500),
.A2(n_510),
.B(n_524),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_504),
.Y(n_500)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_511),
.B(n_516),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_511),
.B(n_516),
.Y(n_524)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g516 ( 
.A1(n_517),
.A2(n_519),
.B1(n_520),
.B2(n_523),
.Y(n_516)
);

CKINVDCx14_ASAP7_75t_R g523 ( 
.A(n_517),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_519),
.B(n_523),
.Y(n_529)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_526),
.B(n_529),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_526),
.B(n_529),
.Y(n_530)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_527),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_534),
.B(n_547),
.Y(n_533)
);

NAND2xp33_ASAP7_75t_L g549 ( 
.A(n_534),
.B(n_547),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_535),
.A2(n_536),
.B1(n_540),
.B2(n_541),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_535),
.B(n_557),
.C(n_558),
.Y(n_556)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_542),
.B(n_544),
.Y(n_541)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_544),
.Y(n_557)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_552),
.B(n_556),
.Y(n_551)
);

OR2x2_ASAP7_75t_L g559 ( 
.A(n_552),
.B(n_556),
.Y(n_559)
);

AOI21xp5_ASAP7_75t_L g585 ( 
.A1(n_560),
.A2(n_586),
.B(n_590),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_561),
.A2(n_574),
.B1(n_577),
.B2(n_581),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_562),
.Y(n_561)
);

NOR2xp67_ASAP7_75t_L g591 ( 
.A(n_562),
.B(n_575),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_562),
.B(n_575),
.Y(n_593)
);

OAI22x1_ASAP7_75t_L g562 ( 
.A1(n_563),
.A2(n_566),
.B1(n_569),
.B2(n_573),
.Y(n_562)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_564),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g584 ( 
.A(n_564),
.B(n_567),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_567),
.B(n_569),
.Y(n_566)
);

HB1xp67_ASAP7_75t_L g573 ( 
.A(n_567),
.Y(n_573)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_569),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_570),
.B(n_571),
.C(n_572),
.Y(n_569)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_575),
.Y(n_574)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_578),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_578),
.B(n_582),
.Y(n_592)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_582),
.Y(n_581)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_583),
.B(n_584),
.Y(n_582)
);

OAI21x1_ASAP7_75t_L g586 ( 
.A1(n_587),
.A2(n_588),
.B(n_589),
.Y(n_586)
);

OAI21xp5_ASAP7_75t_L g590 ( 
.A1(n_591),
.A2(n_592),
.B(n_593),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_SL g600 ( 
.A(n_601),
.B(n_604),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_602),
.B(n_612),
.Y(n_601)
);

XOR2xp5_ASAP7_75t_L g602 ( 
.A(n_603),
.B(n_610),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_604),
.A2(n_605),
.B1(n_606),
.B2(n_609),
.Y(n_603)
);

CKINVDCx11_ASAP7_75t_R g604 ( 
.A(n_605),
.Y(n_604)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_606),
.Y(n_609)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_608),
.Y(n_607)
);

INVx5_ASAP7_75t_L g614 ( 
.A(n_615),
.Y(n_614)
);


endmodule