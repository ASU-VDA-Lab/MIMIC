module real_aes_15699_n_9 (n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_1, n_9);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_1;
output n_9;
wire n_17;
wire n_13;
wire n_12;
wire n_19;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_20;
wire n_18;
wire n_21;
wire n_10;
NOR3xp33_ASAP7_75t_SL g16 ( .A(n_0), .B(n_4), .C(n_17), .Y(n_16) );
NOR3xp33_ASAP7_75t_SL g10 ( .A(n_1), .B(n_6), .C(n_11), .Y(n_10) );
CKINVDCx5p33_ASAP7_75t_R g21 ( .A(n_2), .Y(n_21) );
CKINVDCx5p33_ASAP7_75t_R g18 ( .A(n_3), .Y(n_18) );
CKINVDCx5p33_ASAP7_75t_R g19 ( .A(n_5), .Y(n_19) );
CKINVDCx5p33_ASAP7_75t_R g20 ( .A(n_7), .Y(n_20) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_8), .Y(n_17) );
NAND2xp33_ASAP7_75t_R g9 ( .A(n_10), .B(n_21), .Y(n_9) );
NAND2xp33_ASAP7_75t_R g11 ( .A(n_12), .B(n_20), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_13), .Y(n_12) );
NAND2xp33_ASAP7_75t_R g13 ( .A(n_14), .B(n_19), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_15), .Y(n_14) );
NAND2xp33_ASAP7_75t_R g15 ( .A(n_16), .B(n_18), .Y(n_15) );
endmodule