module real_aes_7053_n_222 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_222);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_222;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_234;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_310;
wire n_725;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_236;
wire n_278;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_569;
wire n_303;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_498;
wire n_691;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_653;
wire n_290;
wire n_365;
wire n_637;
wire n_526;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_521;
wire n_418;
wire n_422;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_541;
wire n_224;
wire n_546;
wire n_639;
wire n_587;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g551 ( .A(n_0), .Y(n_551) );
AOI22xp5_ASAP7_75t_SL g579 ( .A1(n_1), .A2(n_187), .B1(n_542), .B2(n_580), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_2), .A2(n_35), .B1(n_296), .B2(n_335), .Y(n_722) );
AOI22xp33_ASAP7_75t_SL g600 ( .A1(n_3), .A2(n_11), .B1(n_504), .B2(n_519), .Y(n_600) );
AOI22xp5_ASAP7_75t_L g597 ( .A1(n_4), .A2(n_99), .B1(n_314), .B2(n_598), .Y(n_597) );
CKINVDCx20_ASAP7_75t_R g703 ( .A(n_5), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_6), .A2(n_12), .B1(n_455), .B2(n_488), .Y(n_487) );
AOI22xp33_ASAP7_75t_SL g721 ( .A1(n_7), .A2(n_214), .B1(n_390), .B2(n_575), .Y(n_721) );
INVx1_ASAP7_75t_L g538 ( .A(n_8), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g240 ( .A1(n_9), .A2(n_112), .B1(n_241), .B2(n_256), .Y(n_240) );
CKINVDCx20_ASAP7_75t_R g468 ( .A(n_10), .Y(n_468) );
CKINVDCx20_ASAP7_75t_R g705 ( .A(n_13), .Y(n_705) );
AOI221xp5_ASAP7_75t_L g454 ( .A1(n_14), .A2(n_95), .B1(n_455), .B2(n_456), .C(n_458), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_15), .A2(n_61), .B1(n_376), .B2(n_378), .Y(n_375) );
CKINVDCx20_ASAP7_75t_R g584 ( .A(n_16), .Y(n_584) );
AOI22xp33_ASAP7_75t_SL g333 ( .A1(n_17), .A2(n_141), .B1(n_334), .B2(n_335), .Y(n_333) );
AOI222xp33_ASAP7_75t_L g503 ( .A1(n_18), .A2(n_71), .B1(n_120), .B2(n_406), .C1(n_504), .C2(n_505), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_19), .B(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g545 ( .A(n_20), .Y(n_545) );
CKINVDCx20_ASAP7_75t_R g619 ( .A(n_21), .Y(n_619) );
NAND2xp5_ASAP7_75t_SL g327 ( .A(n_22), .B(n_328), .Y(n_327) );
AO22x2_ASAP7_75t_L g253 ( .A1(n_23), .A2(n_76), .B1(n_245), .B2(n_250), .Y(n_253) );
INVx1_ASAP7_75t_L g665 ( .A(n_23), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_24), .A2(n_134), .B1(n_359), .B2(n_361), .Y(n_358) );
CKINVDCx20_ASAP7_75t_R g357 ( .A(n_25), .Y(n_357) );
AOI22xp33_ASAP7_75t_SL g588 ( .A1(n_26), .A2(n_169), .B1(n_308), .B2(n_519), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_27), .A2(n_221), .B1(n_293), .B2(n_338), .Y(n_526) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_28), .A2(n_139), .B1(n_340), .B2(n_457), .Y(n_683) );
INVx1_ASAP7_75t_L g544 ( .A(n_29), .Y(n_544) );
CKINVDCx20_ASAP7_75t_R g416 ( .A(n_30), .Y(n_416) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_31), .A2(n_614), .B1(n_645), .B2(n_646), .Y(n_613) );
INVx1_ASAP7_75t_L g645 ( .A(n_31), .Y(n_645) );
AOI22xp33_ASAP7_75t_SL g329 ( .A1(n_32), .A2(n_143), .B1(n_283), .B2(n_287), .Y(n_329) );
AO22x2_ASAP7_75t_L g255 ( .A1(n_33), .A2(n_80), .B1(n_245), .B2(n_246), .Y(n_255) );
INVx1_ASAP7_75t_L g666 ( .A(n_33), .Y(n_666) );
CKINVDCx20_ASAP7_75t_R g432 ( .A(n_34), .Y(n_432) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_36), .A2(n_135), .B1(n_423), .B2(n_542), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_37), .A2(n_208), .B1(n_279), .B2(n_466), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_38), .A2(n_138), .B1(n_296), .B2(n_457), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_39), .A2(n_72), .B1(n_496), .B2(n_497), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g323 ( .A(n_40), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_41), .A2(n_79), .B1(n_383), .B2(n_621), .Y(n_620) );
CKINVDCx20_ASAP7_75t_R g367 ( .A(n_42), .Y(n_367) );
AOI22xp5_ASAP7_75t_L g718 ( .A1(n_43), .A2(n_75), .B1(n_263), .B2(n_457), .Y(n_718) );
CKINVDCx20_ASAP7_75t_R g639 ( .A(n_44), .Y(n_639) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_45), .Y(n_708) );
AOI222xp33_ASAP7_75t_L g304 ( .A1(n_46), .A2(n_153), .B1(n_204), .B2(n_305), .C1(n_308), .C2(n_312), .Y(n_304) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_47), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g530 ( .A1(n_48), .A2(n_62), .B1(n_423), .B2(n_531), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g617 ( .A(n_49), .Y(n_617) );
AOI22xp5_ASAP7_75t_SL g576 ( .A1(n_50), .A2(n_137), .B1(n_340), .B2(n_577), .Y(n_576) );
CKINVDCx20_ASAP7_75t_R g428 ( .A(n_51), .Y(n_428) );
AOI22xp5_ASAP7_75t_L g444 ( .A1(n_52), .A2(n_445), .B1(n_446), .B2(n_481), .Y(n_444) );
INVx1_ASAP7_75t_L g481 ( .A(n_52), .Y(n_481) );
AOI221xp5_ASAP7_75t_L g464 ( .A1(n_53), .A2(n_87), .B1(n_279), .B2(n_465), .C(n_467), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g673 ( .A(n_54), .Y(n_673) );
CKINVDCx20_ASAP7_75t_R g680 ( .A(n_55), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_56), .A2(n_215), .B1(n_332), .B2(n_686), .Y(n_685) );
CKINVDCx20_ASAP7_75t_R g368 ( .A(n_57), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_58), .A2(n_157), .B1(n_334), .B2(n_426), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g292 ( .A1(n_59), .A2(n_149), .B1(n_293), .B2(n_296), .Y(n_292) );
AOI22xp33_ASAP7_75t_SL g331 ( .A1(n_60), .A2(n_161), .B1(n_293), .B2(n_332), .Y(n_331) );
AOI22xp5_ASAP7_75t_SL g574 ( .A1(n_63), .A2(n_121), .B1(n_261), .B2(n_575), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_64), .A2(n_177), .B1(n_280), .B2(n_466), .Y(n_589) );
CKINVDCx20_ASAP7_75t_R g676 ( .A(n_65), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_66), .A2(n_185), .B1(n_299), .B2(n_335), .Y(n_684) );
CKINVDCx20_ASAP7_75t_R g631 ( .A(n_67), .Y(n_631) );
CKINVDCx20_ASAP7_75t_R g408 ( .A(n_68), .Y(n_408) );
AOI211xp5_ASAP7_75t_L g405 ( .A1(n_69), .A2(n_406), .B(n_407), .C(n_412), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_70), .A2(n_179), .B1(n_465), .B2(n_501), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_73), .A2(n_125), .B1(n_241), .B2(n_338), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_74), .A2(n_163), .B1(n_424), .B2(n_686), .Y(n_719) );
AOI222xp33_ASAP7_75t_L g477 ( .A1(n_77), .A2(n_97), .B1(n_116), .B2(n_370), .C1(n_478), .C2(n_479), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g352 ( .A(n_78), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_81), .A2(n_166), .B1(n_297), .B2(n_302), .Y(n_610) );
CKINVDCx20_ASAP7_75t_R g317 ( .A(n_82), .Y(n_317) );
CKINVDCx20_ASAP7_75t_R g637 ( .A(n_83), .Y(n_637) );
INVx1_ASAP7_75t_L g230 ( .A(n_84), .Y(n_230) );
INVx1_ASAP7_75t_L g532 ( .A(n_85), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_86), .A2(n_119), .B1(n_421), .B2(n_424), .Y(n_498) );
AOI22xp5_ASAP7_75t_L g605 ( .A1(n_88), .A2(n_165), .B1(n_293), .B2(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_89), .B(n_561), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_90), .A2(n_114), .B1(n_456), .B2(n_609), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_91), .A2(n_167), .B1(n_421), .B2(n_424), .Y(n_420) );
INVx1_ASAP7_75t_L g228 ( .A(n_92), .Y(n_228) );
AOI22xp33_ASAP7_75t_SL g324 ( .A1(n_93), .A2(n_124), .B1(n_308), .B2(n_315), .Y(n_324) );
AOI22xp33_ASAP7_75t_SL g608 ( .A1(n_94), .A2(n_142), .B1(n_382), .B2(n_609), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g709 ( .A1(n_96), .A2(n_210), .B1(n_315), .B2(n_710), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g281 ( .A1(n_98), .A2(n_130), .B1(n_282), .B2(n_287), .Y(n_281) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_100), .A2(n_175), .B1(n_308), .B2(n_519), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g590 ( .A(n_101), .Y(n_590) );
CKINVDCx20_ASAP7_75t_R g644 ( .A(n_102), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_103), .B(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g553 ( .A(n_104), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_105), .A2(n_201), .B1(n_392), .B2(n_395), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_106), .A2(n_144), .B1(n_241), .B2(n_388), .Y(n_525) );
INVx1_ASAP7_75t_L g567 ( .A(n_107), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g534 ( .A1(n_108), .A2(n_535), .B1(n_568), .B2(n_569), .Y(n_534) );
CKINVDCx16_ASAP7_75t_R g568 ( .A(n_108), .Y(n_568) );
INVx1_ASAP7_75t_L g462 ( .A(n_109), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g633 ( .A(n_110), .Y(n_633) );
INVx1_ASAP7_75t_L g521 ( .A(n_111), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_113), .A2(n_192), .B1(n_386), .B2(n_390), .Y(n_385) );
AOI221xp5_ASAP7_75t_L g448 ( .A1(n_115), .A2(n_160), .B1(n_261), .B2(n_434), .C(n_449), .Y(n_448) );
AOI22xp5_ASAP7_75t_L g586 ( .A1(n_117), .A2(n_148), .B1(n_288), .B2(n_314), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g410 ( .A1(n_118), .A2(n_171), .B1(n_361), .B2(n_411), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_122), .B(n_275), .Y(n_409) );
INVx2_ASAP7_75t_L g231 ( .A(n_123), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_126), .A2(n_183), .B1(n_288), .B2(n_411), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g413 ( .A(n_127), .Y(n_413) );
CKINVDCx20_ASAP7_75t_R g624 ( .A(n_128), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_129), .A2(n_168), .B1(n_381), .B2(n_383), .Y(n_380) );
CKINVDCx16_ASAP7_75t_R g403 ( .A(n_131), .Y(n_403) );
AND2x6_ASAP7_75t_L g227 ( .A(n_132), .B(n_228), .Y(n_227) );
HB1xp67_ASAP7_75t_L g659 ( .A(n_132), .Y(n_659) );
AO22x2_ASAP7_75t_L g244 ( .A1(n_133), .A2(n_182), .B1(n_245), .B2(n_246), .Y(n_244) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_136), .A2(n_193), .B1(n_426), .B2(n_547), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g260 ( .A1(n_140), .A2(n_164), .B1(n_261), .B2(n_269), .Y(n_260) );
AOI22xp33_ASAP7_75t_SL g528 ( .A1(n_145), .A2(n_162), .B1(n_382), .B2(n_529), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g611 ( .A(n_146), .Y(n_611) );
AOI22xp5_ASAP7_75t_L g668 ( .A1(n_147), .A2(n_669), .B1(n_688), .B2(n_689), .Y(n_668) );
CKINVDCx20_ASAP7_75t_R g688 ( .A(n_147), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_150), .A2(n_205), .B1(n_256), .B2(n_388), .Y(n_687) );
AOI22xp33_ASAP7_75t_SL g337 ( .A1(n_151), .A2(n_197), .B1(n_241), .B2(n_338), .Y(n_337) );
AO22x1_ASAP7_75t_L g449 ( .A1(n_152), .A2(n_180), .B1(n_450), .B2(n_452), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g341 ( .A(n_154), .Y(n_341) );
AO22x2_ASAP7_75t_L g249 ( .A1(n_155), .A2(n_195), .B1(n_245), .B2(n_250), .Y(n_249) );
AOI22xp5_ASAP7_75t_L g522 ( .A1(n_156), .A2(n_209), .B1(n_287), .B2(n_314), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_158), .A2(n_199), .B1(n_312), .B2(n_558), .Y(n_678) );
INVx1_ASAP7_75t_L g435 ( .A(n_159), .Y(n_435) );
AOI22xp33_ASAP7_75t_SL g339 ( .A1(n_170), .A2(n_198), .B1(n_261), .B2(n_340), .Y(n_339) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_172), .A2(n_220), .B1(n_491), .B2(n_493), .Y(n_490) );
AOI22xp33_ASAP7_75t_L g298 ( .A1(n_173), .A2(n_196), .B1(n_299), .B2(n_302), .Y(n_298) );
INVx1_ASAP7_75t_L g559 ( .A(n_174), .Y(n_559) );
CKINVDCx20_ASAP7_75t_R g627 ( .A(n_176), .Y(n_627) );
CKINVDCx20_ASAP7_75t_R g681 ( .A(n_178), .Y(n_681) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_181), .Y(n_430) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_182), .B(n_664), .Y(n_663) );
NAND2xp5_ASAP7_75t_SL g326 ( .A(n_184), .B(n_279), .Y(n_326) );
AOI211xp5_ASAP7_75t_L g222 ( .A1(n_186), .A2(n_223), .B(n_232), .C(n_667), .Y(n_222) );
INVx1_ASAP7_75t_L g698 ( .A(n_188), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g274 ( .A1(n_189), .A2(n_202), .B1(n_275), .B2(n_279), .Y(n_274) );
CKINVDCx20_ASAP7_75t_R g674 ( .A(n_190), .Y(n_674) );
INVx1_ASAP7_75t_L g564 ( .A(n_191), .Y(n_564) );
INVx1_ASAP7_75t_L g459 ( .A(n_194), .Y(n_459) );
INVx1_ASAP7_75t_L g662 ( .A(n_195), .Y(n_662) );
CKINVDCx20_ASAP7_75t_R g372 ( .A(n_200), .Y(n_372) );
INVx1_ASAP7_75t_L g540 ( .A(n_203), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_206), .Y(n_471) );
INVx1_ASAP7_75t_L g245 ( .A(n_207), .Y(n_245) );
INVx1_ASAP7_75t_L g247 ( .A(n_207), .Y(n_247) );
CKINVDCx20_ASAP7_75t_R g642 ( .A(n_211), .Y(n_642) );
CKINVDCx20_ASAP7_75t_R g640 ( .A(n_212), .Y(n_640) );
INVx1_ASAP7_75t_L g556 ( .A(n_213), .Y(n_556) );
OA22x2_ASAP7_75t_L g483 ( .A1(n_216), .A2(n_484), .B1(n_485), .B2(n_506), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_216), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g596 ( .A(n_217), .Y(n_596) );
CKINVDCx20_ASAP7_75t_R g712 ( .A(n_218), .Y(n_712) );
AOI22xp5_ASAP7_75t_L g344 ( .A1(n_219), .A2(n_345), .B1(n_396), .B2(n_397), .Y(n_344) );
CKINVDCx20_ASAP7_75t_R g396 ( .A(n_219), .Y(n_396) );
CKINVDCx20_ASAP7_75t_R g223 ( .A(n_224), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_225), .Y(n_224) );
HB1xp67_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AND2x4_ASAP7_75t_L g226 ( .A(n_227), .B(n_229), .Y(n_226) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_228), .Y(n_658) );
OAI21xp5_ASAP7_75t_L g696 ( .A1(n_229), .A2(n_657), .B(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_231), .Y(n_229) );
AOI221xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_399), .B1(n_652), .B2(n_653), .C(n_654), .Y(n_232) );
INVx1_ASAP7_75t_L g653 ( .A(n_233), .Y(n_653) );
AOI22xp5_ASAP7_75t_SL g233 ( .A1(n_234), .A2(n_235), .B1(n_343), .B2(n_398), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AO22x2_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_237), .B1(n_318), .B2(n_342), .Y(n_235) );
INVx2_ASAP7_75t_SL g236 ( .A(n_237), .Y(n_236) );
XOR2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_317), .Y(n_237) );
NAND4xp75_ASAP7_75t_L g238 ( .A(n_239), .B(n_273), .C(n_291), .D(n_304), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_260), .Y(n_239) );
BUFx3_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
BUFx3_ASAP7_75t_L g394 ( .A(n_242), .Y(n_394) );
BUFx3_ASAP7_75t_L g457 ( .A(n_242), .Y(n_457) );
AND2x2_ASAP7_75t_L g242 ( .A(n_243), .B(n_251), .Y(n_242) );
AND2x2_ASAP7_75t_L g301 ( .A(n_243), .B(n_272), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_243), .B(n_251), .Y(n_438) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_243), .B(n_272), .Y(n_461) );
AND2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_248), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_244), .B(n_249), .Y(n_259) );
INVx2_ASAP7_75t_L g267 ( .A(n_244), .Y(n_267) );
AND2x2_ASAP7_75t_L g286 ( .A(n_244), .B(n_253), .Y(n_286) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx1_ASAP7_75t_L g250 ( .A(n_247), .Y(n_250) );
INVx1_ASAP7_75t_L g289 ( .A(n_248), .Y(n_289) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g268 ( .A(n_249), .Y(n_268) );
AND2x2_ASAP7_75t_L g278 ( .A(n_249), .B(n_267), .Y(n_278) );
INVx1_ASAP7_75t_L g311 ( .A(n_249), .Y(n_311) );
AND2x4_ASAP7_75t_L g257 ( .A(n_251), .B(n_258), .Y(n_257) );
AND2x2_ASAP7_75t_L g295 ( .A(n_251), .B(n_266), .Y(n_295) );
AND2x4_ASAP7_75t_L g297 ( .A(n_251), .B(n_278), .Y(n_297) );
AND2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_254), .Y(n_251) );
OR2x2_ASAP7_75t_L g265 ( .A(n_252), .B(n_255), .Y(n_265) );
AND2x2_ASAP7_75t_L g272 ( .A(n_252), .B(n_255), .Y(n_272) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g290 ( .A(n_253), .B(n_255), .Y(n_290) );
AND2x2_ASAP7_75t_L g310 ( .A(n_254), .B(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g470 ( .A(n_254), .Y(n_470) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g285 ( .A(n_255), .Y(n_285) );
BUFx3_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
BUFx3_ASAP7_75t_L g338 ( .A(n_257), .Y(n_338) );
BUFx2_ASAP7_75t_L g424 ( .A(n_257), .Y(n_424) );
BUFx3_ASAP7_75t_L g453 ( .A(n_257), .Y(n_453) );
BUFx3_ASAP7_75t_L g542 ( .A(n_257), .Y(n_542) );
AND2x2_ASAP7_75t_L g580 ( .A(n_258), .B(n_470), .Y(n_580) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
OR2x6_ASAP7_75t_L g303 ( .A(n_259), .B(n_285), .Y(n_303) );
INVx1_ASAP7_75t_L g429 ( .A(n_261), .Y(n_429) );
INVx3_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
INVx2_ASAP7_75t_SL g497 ( .A(n_262), .Y(n_497) );
OAI221xp5_ASAP7_75t_SL g616 ( .A1(n_262), .A2(n_617), .B1(n_618), .B2(n_619), .C(n_620), .Y(n_616) );
INVx11_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx11_ASAP7_75t_L g389 ( .A(n_263), .Y(n_389) );
AND2x6_ASAP7_75t_L g263 ( .A(n_264), .B(n_266), .Y(n_263) );
AND2x4_ASAP7_75t_L g277 ( .A(n_264), .B(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g350 ( .A(n_265), .B(n_351), .Y(n_350) );
AND2x4_ASAP7_75t_L g271 ( .A(n_266), .B(n_272), .Y(n_271) );
AND2x6_ASAP7_75t_L g307 ( .A(n_266), .B(n_290), .Y(n_307) );
AND2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g390 ( .A(n_270), .Y(n_390) );
OAI22xp5_ASAP7_75t_L g427 ( .A1(n_270), .A2(n_428), .B1(n_429), .B2(n_430), .Y(n_427) );
INVx2_ASAP7_75t_L g455 ( .A(n_270), .Y(n_455) );
OAI221xp5_ASAP7_75t_SL g543 ( .A1(n_270), .A2(n_436), .B1(n_544), .B2(n_545), .C(n_546), .Y(n_543) );
INVx3_ASAP7_75t_L g609 ( .A(n_270), .Y(n_609) );
INVx6_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
BUFx3_ASAP7_75t_L g340 ( .A(n_271), .Y(n_340) );
BUFx3_ASAP7_75t_L g529 ( .A(n_271), .Y(n_529) );
AND2x6_ASAP7_75t_L g280 ( .A(n_272), .B(n_278), .Y(n_280) );
NAND2x1p5_ASAP7_75t_L g356 ( .A(n_272), .B(n_278), .Y(n_356) );
AND2x2_ASAP7_75t_SL g273 ( .A(n_274), .B(n_281), .Y(n_273) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g328 ( .A(n_276), .Y(n_328) );
INVx5_ASAP7_75t_L g466 ( .A(n_276), .Y(n_466) );
INVx2_ASAP7_75t_L g517 ( .A(n_276), .Y(n_517) );
INVx4_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g351 ( .A(n_278), .Y(n_351) );
BUFx4f_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
BUFx2_ASAP7_75t_L g501 ( .A(n_280), .Y(n_501) );
BUFx2_ASAP7_75t_L g515 ( .A(n_280), .Y(n_515) );
BUFx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx1_ASAP7_75t_L g360 ( .A(n_283), .Y(n_360) );
BUFx2_ASAP7_75t_L g411 ( .A(n_283), .Y(n_411) );
BUFx3_ASAP7_75t_L g519 ( .A(n_283), .Y(n_519) );
AND2x4_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x4_ASAP7_75t_L g309 ( .A(n_286), .B(n_310), .Y(n_309) );
AND2x4_ASAP7_75t_L g315 ( .A(n_286), .B(n_316), .Y(n_315) );
NAND2x1p5_ASAP7_75t_L g469 ( .A(n_286), .B(n_470), .Y(n_469) );
BUFx3_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
BUFx6f_ASAP7_75t_L g363 ( .A(n_288), .Y(n_363) );
BUFx2_ASAP7_75t_SL g598 ( .A(n_288), .Y(n_598) );
BUFx2_ASAP7_75t_SL g710 ( .A(n_288), .Y(n_710) );
AND2x4_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
INVx1_ASAP7_75t_L g476 ( .A(n_289), .Y(n_476) );
INVx1_ASAP7_75t_L g475 ( .A(n_290), .Y(n_475) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_298), .Y(n_291) );
INVx3_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx3_ASAP7_75t_L g686 ( .A(n_294), .Y(n_686) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
BUFx6f_ASAP7_75t_L g377 ( .A(n_295), .Y(n_377) );
BUFx2_ASAP7_75t_SL g577 ( .A(n_295), .Y(n_577) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_296), .Y(n_626) );
BUFx3_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
BUFx3_ASAP7_75t_L g332 ( .A(n_297), .Y(n_332) );
INVx2_ASAP7_75t_L g379 ( .A(n_297), .Y(n_379) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_297), .Y(n_423) );
BUFx3_ASAP7_75t_L g451 ( .A(n_297), .Y(n_451) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_299), .Y(n_621) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx1_ASAP7_75t_L g334 ( .A(n_300), .Y(n_334) );
INVx5_ASAP7_75t_L g382 ( .A(n_300), .Y(n_382) );
INVx4_ASAP7_75t_L g492 ( .A(n_300), .Y(n_492) );
BUFx3_ASAP7_75t_L g548 ( .A(n_300), .Y(n_548) );
INVx3_ASAP7_75t_L g575 ( .A(n_300), .Y(n_575) );
INVx8_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
BUFx2_ASAP7_75t_L g335 ( .A(n_302), .Y(n_335) );
BUFx4f_ASAP7_75t_SL g383 ( .A(n_302), .Y(n_383) );
BUFx2_ASAP7_75t_L g493 ( .A(n_302), .Y(n_493) );
INVx6_ASAP7_75t_SL g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_SL g426 ( .A(n_303), .Y(n_426) );
INVx1_ASAP7_75t_SL g531 ( .A(n_303), .Y(n_531) );
INVx4_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OAI21xp5_ASAP7_75t_SL g707 ( .A1(n_306), .A2(n_708), .B(n_709), .Y(n_707) );
INVx4_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g322 ( .A(n_307), .Y(n_322) );
BUFx3_ASAP7_75t_L g406 ( .A(n_307), .Y(n_406) );
BUFx6f_ASAP7_75t_L g478 ( .A(n_307), .Y(n_478) );
INVx2_ASAP7_75t_L g585 ( .A(n_307), .Y(n_585) );
INVx4_ASAP7_75t_L g480 ( .A(n_308), .Y(n_480) );
BUFx6f_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_309), .Y(n_366) );
BUFx6f_ASAP7_75t_L g415 ( .A(n_309), .Y(n_415) );
BUFx4f_ASAP7_75t_SL g504 ( .A(n_309), .Y(n_504) );
BUFx2_ASAP7_75t_L g558 ( .A(n_309), .Y(n_558) );
INVx1_ASAP7_75t_L g316 ( .A(n_311), .Y(n_316) );
INVx1_ASAP7_75t_L g417 ( .A(n_312), .Y(n_417) );
INVx3_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
BUFx4f_ASAP7_75t_SL g505 ( .A(n_314), .Y(n_505) );
BUFx12f_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
BUFx6f_ASAP7_75t_L g371 ( .A(n_315), .Y(n_371) );
BUFx6f_ASAP7_75t_L g562 ( .A(n_315), .Y(n_562) );
INVx4_ASAP7_75t_SL g342 ( .A(n_318), .Y(n_342) );
XOR2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_341), .Y(n_318) );
NAND3x1_ASAP7_75t_L g319 ( .A(n_320), .B(n_330), .C(n_336), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g320 ( .A(n_321), .B(n_325), .Y(n_320) );
OAI21xp5_ASAP7_75t_SL g321 ( .A1(n_322), .A2(n_323), .B(n_324), .Y(n_321) );
OAI222xp33_ASAP7_75t_L g364 ( .A1(n_322), .A2(n_365), .B1(n_367), .B2(n_368), .C1(n_369), .C2(n_372), .Y(n_364) );
OAI21xp5_ASAP7_75t_SL g520 ( .A1(n_322), .A2(n_521), .B(n_522), .Y(n_520) );
OAI21xp5_ASAP7_75t_L g595 ( .A1(n_322), .A2(n_596), .B(n_597), .Y(n_595) );
NAND3xp33_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .C(n_329), .Y(n_325) );
AND2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_333), .Y(n_330) );
AND2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_339), .Y(n_336) );
BUFx2_ASAP7_75t_L g395 ( .A(n_338), .Y(n_395) );
INVx1_ASAP7_75t_L g398 ( .A(n_343), .Y(n_398) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_SL g397 ( .A(n_345), .Y(n_397) );
AND2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_373), .Y(n_345) );
NOR2xp33_ASAP7_75t_SL g346 ( .A(n_347), .B(n_364), .Y(n_346) );
OAI221xp5_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_352), .B1(n_353), .B2(n_357), .C(n_358), .Y(n_347) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_348), .A2(n_634), .B1(n_673), .B2(n_674), .Y(n_672) );
INVx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_SL g552 ( .A(n_349), .Y(n_552) );
INVx2_ASAP7_75t_L g632 ( .A(n_349), .Y(n_632) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
BUFx3_ASAP7_75t_L g704 ( .A(n_350), .Y(n_704) );
OAI211xp5_ASAP7_75t_L g407 ( .A1(n_353), .A2(n_408), .B(n_409), .C(n_410), .Y(n_407) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_355), .A2(n_551), .B1(n_552), .B2(n_553), .Y(n_550) );
BUFx3_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g635 ( .A(n_356), .Y(n_635) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
OAI222xp33_ASAP7_75t_L g636 ( .A1(n_365), .A2(n_369), .B1(n_637), .B2(n_638), .C1(n_639), .C2(n_640), .Y(n_636) );
CKINVDCx20_ASAP7_75t_R g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx3_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g373 ( .A(n_374), .B(n_384), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_375), .B(n_380), .Y(n_374) );
BUFx3_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_377), .Y(n_434) );
BUFx3_ASAP7_75t_L g496 ( .A(n_377), .Y(n_496) );
INVx3_ASAP7_75t_L g623 ( .A(n_377), .Y(n_623) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
BUFx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
CKINVDCx20_ASAP7_75t_R g463 ( .A(n_383), .Y(n_463) );
NAND2xp5_ASAP7_75t_SL g384 ( .A(n_385), .B(n_391), .Y(n_384) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx2_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
INVx5_ASAP7_75t_SL g606 ( .A(n_389), .Y(n_606) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g652 ( .A(n_399), .Y(n_652) );
AOI22xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_439), .B1(n_650), .B2(n_651), .Y(n_399) );
INVx1_ASAP7_75t_SL g650 ( .A(n_400), .Y(n_650) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
XNOR2xp5_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
AND2x2_ASAP7_75t_L g404 ( .A(n_405), .B(n_418), .Y(n_404) );
INVx3_ASAP7_75t_L g677 ( .A(n_406), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_414), .B1(n_416), .B2(n_417), .Y(n_412) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
BUFx6f_ASAP7_75t_L g714 ( .A(n_415), .Y(n_714) );
NOR3xp33_ASAP7_75t_L g418 ( .A(n_419), .B(n_427), .C(n_431), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_420), .B(n_425), .Y(n_419) );
INVx3_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx4_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_433), .B1(n_435), .B2(n_436), .Y(n_431) );
OAI221xp5_ASAP7_75t_SL g537 ( .A1(n_433), .A2(n_538), .B1(n_539), .B2(n_540), .C(n_541), .Y(n_537) );
INVx1_ASAP7_75t_SL g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g651 ( .A(n_439), .Y(n_651) );
XOR2xp5_ASAP7_75t_L g439 ( .A(n_440), .B(n_570), .Y(n_439) );
OAI22xp5_ASAP7_75t_SL g440 ( .A1(n_441), .A2(n_442), .B1(n_507), .B2(n_508), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
OAI22xp5_ASAP7_75t_SL g442 ( .A1(n_443), .A2(n_444), .B1(n_482), .B2(n_483), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
AND4x1_ASAP7_75t_L g447 ( .A(n_448), .B(n_454), .C(n_464), .D(n_477), .Y(n_447) );
BUFx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g618 ( .A(n_453), .Y(n_618) );
BUFx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g489 ( .A(n_457), .Y(n_489) );
OAI22xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_460), .B1(n_462), .B2(n_463), .Y(n_458) );
BUFx2_ASAP7_75t_R g460 ( .A(n_461), .Y(n_460) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OAI22xp5_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_469), .B1(n_471), .B2(n_472), .Y(n_467) );
INVx4_ASAP7_75t_L g566 ( .A(n_469), .Y(n_566) );
BUFx3_ASAP7_75t_L g643 ( .A(n_469), .Y(n_643) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_469), .A2(n_712), .B1(n_713), .B2(n_715), .Y(n_711) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_472), .A2(n_564), .B1(n_565), .B2(n_567), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g641 ( .A1(n_472), .A2(n_642), .B1(n_643), .B2(n_644), .Y(n_641) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
CKINVDCx16_ASAP7_75t_R g473 ( .A(n_474), .Y(n_473) );
OAI22xp5_ASAP7_75t_L g679 ( .A1(n_474), .A2(n_565), .B1(n_680), .B2(n_681), .Y(n_679) );
OR2x6_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
INVx2_ASAP7_75t_SL g555 ( .A(n_478), .Y(n_555) );
INVx2_ASAP7_75t_L g638 ( .A(n_478), .Y(n_638) );
INVx3_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_SL g506 ( .A(n_485), .Y(n_506) );
NAND4xp75_ASAP7_75t_L g485 ( .A(n_486), .B(n_494), .C(n_499), .D(n_503), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_490), .Y(n_486) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
BUFx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_498), .Y(n_494) );
INVx1_ASAP7_75t_L g539 ( .A(n_497), .Y(n_539) );
AND2x2_ASAP7_75t_SL g499 ( .A(n_500), .B(n_502), .Y(n_499) );
INVx1_ASAP7_75t_SL g507 ( .A(n_508), .Y(n_507) );
XOR2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_533), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
XOR2x2_ASAP7_75t_SL g510 ( .A(n_511), .B(n_532), .Y(n_510) );
NAND2x1p5_ASAP7_75t_L g511 ( .A(n_512), .B(n_523), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_513), .B(n_520), .Y(n_512) );
NAND3xp33_ASAP7_75t_L g513 ( .A(n_514), .B(n_516), .C(n_518), .Y(n_513) );
NOR2x1_ASAP7_75t_L g523 ( .A(n_524), .B(n_527), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_525), .B(n_526), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_528), .B(n_530), .Y(n_527) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g569 ( .A(n_535), .Y(n_569) );
AND2x2_ASAP7_75t_SL g535 ( .A(n_536), .B(n_549), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_537), .B(n_543), .Y(n_536) );
INVx3_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
NOR3xp33_ASAP7_75t_L g549 ( .A(n_550), .B(n_554), .C(n_563), .Y(n_549) );
OAI221xp5_ASAP7_75t_SL g554 ( .A1(n_555), .A2(n_556), .B1(n_557), .B2(n_559), .C(n_560), .Y(n_554) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
BUFx4f_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AOI22xp5_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_572), .B1(n_591), .B2(n_649), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
XOR2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_590), .Y(n_572) );
NAND4xp75_ASAP7_75t_SL g573 ( .A(n_574), .B(n_576), .C(n_578), .D(n_582), .Y(n_573) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g582 ( .A(n_583), .B(n_587), .Y(n_582) );
OAI21xp5_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_585), .B(n_586), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
INVx1_ASAP7_75t_L g649 ( .A(n_591), .Y(n_649) );
AOI22xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_612), .B1(n_647), .B2(n_648), .Y(n_591) );
INVx3_ASAP7_75t_SL g647 ( .A(n_592), .Y(n_647) );
XOR2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_611), .Y(n_592) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_594), .B(n_602), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_595), .B(n_599), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_600), .B(n_601), .Y(n_599) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_603), .B(n_607), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_610), .Y(n_607) );
INVx3_ASAP7_75t_L g648 ( .A(n_612), .Y(n_648) );
BUFx3_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g646 ( .A(n_614), .Y(n_646) );
AND2x2_ASAP7_75t_SL g614 ( .A(n_615), .B(n_629), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g615 ( .A(n_616), .B(n_622), .Y(n_615) );
OAI221xp5_ASAP7_75t_SL g622 ( .A1(n_623), .A2(n_624), .B1(n_625), .B2(n_627), .C(n_628), .Y(n_622) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
NOR3xp33_ASAP7_75t_L g629 ( .A(n_630), .B(n_636), .C(n_641), .Y(n_629) );
OAI22xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_632), .B1(n_633), .B2(n_634), .Y(n_630) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g706 ( .A(n_635), .Y(n_706) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NOR2x1_ASAP7_75t_L g655 ( .A(n_656), .B(n_660), .Y(n_655) );
OR2x2_ASAP7_75t_SL g725 ( .A(n_656), .B(n_661), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_657), .B(n_659), .Y(n_656) );
CKINVDCx20_ASAP7_75t_R g691 ( .A(n_657), .Y(n_691) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_658), .B(n_694), .Y(n_697) );
CKINVDCx16_ASAP7_75t_R g694 ( .A(n_659), .Y(n_694) );
CKINVDCx20_ASAP7_75t_R g660 ( .A(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
OAI322xp33_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_690), .A3(n_692), .B1(n_695), .B2(n_698), .C1(n_699), .C2(n_723), .Y(n_667) );
CKINVDCx20_ASAP7_75t_R g689 ( .A(n_669), .Y(n_689) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_SL g670 ( .A(n_671), .B(n_682), .Y(n_670) );
NOR3xp33_ASAP7_75t_L g671 ( .A(n_672), .B(n_675), .C(n_679), .Y(n_671) );
OAI21xp33_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_677), .B(n_678), .Y(n_675) );
AND4x1_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .C(n_685), .D(n_687), .Y(n_682) );
HB1xp67_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
HB1xp67_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
CKINVDCx20_ASAP7_75t_R g695 ( .A(n_696), .Y(n_695) );
XOR2x2_ASAP7_75t_L g699 ( .A(n_698), .B(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_701), .B(n_716), .Y(n_700) );
NOR3xp33_ASAP7_75t_L g701 ( .A(n_702), .B(n_707), .C(n_711), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g702 ( .A1(n_703), .A2(n_704), .B1(n_705), .B2(n_706), .Y(n_702) );
INVx2_ASAP7_75t_SL g713 ( .A(n_714), .Y(n_713) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_717), .B(n_720), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_718), .B(n_719), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_721), .B(n_722), .Y(n_720) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_724), .Y(n_723) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_725), .Y(n_724) );
endmodule