module fake_netlist_6_2063_n_1766 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1766);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1766;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1627;
wire n_1295;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g165 ( 
.A(n_160),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_27),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_48),
.Y(n_167)
);

INVxp67_ASAP7_75t_SL g168 ( 
.A(n_110),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_143),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_122),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_108),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_40),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_1),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_61),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_159),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_26),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_58),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_89),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_68),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_93),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_115),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_11),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_76),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_114),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_66),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_141),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_163),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_42),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_153),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_82),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_131),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_41),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_3),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_100),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_21),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_49),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_57),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_137),
.Y(n_199)
);

BUFx10_ASAP7_75t_L g200 ( 
.A(n_132),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_28),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_162),
.Y(n_202)
);

BUFx10_ASAP7_75t_L g203 ( 
.A(n_18),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_16),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_154),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_83),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_164),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_2),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_147),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_142),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_49),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_148),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_134),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_69),
.Y(n_214)
);

BUFx8_ASAP7_75t_SL g215 ( 
.A(n_5),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_38),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_71),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_118),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_50),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_4),
.Y(n_220)
);

BUFx10_ASAP7_75t_L g221 ( 
.A(n_25),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_1),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_59),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_102),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_12),
.Y(n_225)
);

INVx2_ASAP7_75t_SL g226 ( 
.A(n_111),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_125),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_70),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_38),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_67),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_62),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_50),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_126),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_138),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_80),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_107),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_81),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_17),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_53),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_5),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_84),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_22),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_29),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_44),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_116),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_21),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_105),
.Y(n_247)
);

BUFx2_ASAP7_75t_SL g248 ( 
.A(n_39),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_22),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_74),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_146),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_106),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_29),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_3),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_44),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_129),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_43),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_99),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_25),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_9),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_34),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_109),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_11),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_72),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_36),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_4),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_53),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_48),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_63),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_119),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_161),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_117),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_158),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_91),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_52),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_34),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_27),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_37),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_156),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_140),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_133),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_130),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_14),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_52),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_78),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_37),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_0),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_92),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_88),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_75),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_0),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_55),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_101),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_8),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_46),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_150),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_56),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_19),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_23),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_103),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_120),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_124),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_6),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_86),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g305 ( 
.A(n_35),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_149),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_35),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_46),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_155),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_55),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_64),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_112),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_13),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_12),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_56),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_65),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_36),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_95),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_157),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_51),
.Y(n_320)
);

BUFx8_ASAP7_75t_SL g321 ( 
.A(n_15),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_18),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_14),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_127),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_45),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_145),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_123),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_175),
.B(n_2),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_215),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_321),
.Y(n_330)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_169),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_174),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_202),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_196),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_209),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_206),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_310),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_207),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_210),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_212),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_224),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_213),
.Y(n_342)
);

INVxp33_ASAP7_75t_L g343 ( 
.A(n_314),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_205),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_217),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_218),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_223),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_228),
.Y(n_348)
);

INVxp33_ASAP7_75t_SL g349 ( 
.A(n_166),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_196),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_230),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_231),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_216),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_233),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_196),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_196),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_196),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_203),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_203),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_241),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_169),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_245),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_226),
.B(n_6),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_325),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_283),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_242),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_247),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g368 ( 
.A(n_305),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_250),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_205),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_251),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_203),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_242),
.B(n_7),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_172),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_252),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_256),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_169),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_242),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_226),
.B(n_7),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_242),
.Y(n_380)
);

INVxp67_ASAP7_75t_SL g381 ( 
.A(n_170),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_181),
.B(n_8),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_242),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_254),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_254),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_258),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_200),
.Y(n_387)
);

NOR2xp67_ASAP7_75t_L g388 ( 
.A(n_181),
.B(n_9),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_262),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_272),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_273),
.Y(n_391)
);

NOR2xp67_ASAP7_75t_L g392 ( 
.A(n_167),
.B(n_10),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_254),
.Y(n_393)
);

NOR2xp67_ASAP7_75t_L g394 ( 
.A(n_193),
.B(n_10),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_274),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_254),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_221),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_279),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_254),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_190),
.B(n_13),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_303),
.Y(n_401)
);

INVxp67_ASAP7_75t_SL g402 ( 
.A(n_303),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_303),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_280),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_235),
.B(n_15),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_333),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_332),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_336),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_402),
.B(n_303),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_338),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_373),
.B(n_303),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_339),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_361),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_334),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_340),
.B(n_177),
.Y(n_415)
);

AND2x4_ASAP7_75t_L g416 ( 
.A(n_373),
.B(n_165),
.Y(n_416)
);

HB1xp67_ASAP7_75t_L g417 ( 
.A(n_365),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_335),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_334),
.Y(n_419)
);

OAI21x1_ASAP7_75t_L g420 ( 
.A1(n_331),
.A2(n_180),
.B(n_171),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_341),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_350),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_361),
.Y(n_423)
);

AND2x6_ASAP7_75t_L g424 ( 
.A(n_331),
.B(n_169),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_350),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_355),
.Y(n_426)
);

NOR2x1_ASAP7_75t_L g427 ( 
.A(n_331),
.B(n_388),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_361),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_355),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_344),
.B(n_370),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_365),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_363),
.B(n_177),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_342),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_377),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_347),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_356),
.B(n_184),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_356),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_377),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_387),
.B(n_200),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_357),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_345),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_377),
.Y(n_442)
);

CKINVDCx16_ASAP7_75t_R g443 ( 
.A(n_364),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_357),
.B(n_186),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_354),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_366),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_331),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_366),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_367),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_R g450 ( 
.A(n_346),
.B(n_281),
.Y(n_450)
);

OA21x2_ASAP7_75t_L g451 ( 
.A1(n_378),
.A2(n_219),
.B(n_204),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_378),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_380),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_368),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_368),
.A2(n_286),
.B1(n_225),
.B2(n_183),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_380),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_383),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_383),
.Y(n_458)
);

INVx3_ASAP7_75t_L g459 ( 
.A(n_384),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_384),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_387),
.B(n_200),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_369),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_337),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_385),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_385),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_393),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_376),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_386),
.B(n_178),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_390),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_391),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_393),
.Y(n_471)
);

NAND3xp33_ASAP7_75t_L g472 ( 
.A(n_382),
.B(n_211),
.C(n_208),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_379),
.B(n_178),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_396),
.B(n_179),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_396),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_399),
.B(n_179),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_404),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_399),
.Y(n_478)
);

OR2x6_ASAP7_75t_L g479 ( 
.A(n_392),
.B(n_248),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_432),
.B(n_381),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_415),
.B(n_349),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_431),
.B(n_364),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_432),
.B(n_401),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_448),
.Y(n_484)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_417),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_419),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_430),
.B(n_401),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_452),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_452),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_419),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_411),
.Y(n_491)
);

INVx4_ASAP7_75t_L g492 ( 
.A(n_452),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_431),
.B(n_403),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_419),
.Y(n_494)
);

BUFx4f_ASAP7_75t_L g495 ( 
.A(n_451),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_468),
.B(n_430),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_448),
.Y(n_497)
);

INVx8_ASAP7_75t_L g498 ( 
.A(n_416),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_417),
.B(n_403),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_448),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_411),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_454),
.B(n_343),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_411),
.B(n_288),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_454),
.B(n_353),
.Y(n_504)
);

AND2x2_ASAP7_75t_SL g505 ( 
.A(n_473),
.B(n_328),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_452),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_439),
.A2(n_352),
.B1(n_371),
.B2(n_398),
.Y(n_507)
);

NOR2x1p5_ASAP7_75t_L g508 ( 
.A(n_406),
.B(n_329),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_452),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_414),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_452),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_414),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_422),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_416),
.B(n_168),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_473),
.B(n_348),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_453),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_408),
.B(n_351),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_422),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_410),
.B(n_360),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_409),
.Y(n_520)
);

BUFx4f_ASAP7_75t_L g521 ( 
.A(n_451),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_409),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_425),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_458),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_458),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_453),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_412),
.B(n_362),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_425),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_426),
.Y(n_529)
);

INVx5_ASAP7_75t_L g530 ( 
.A(n_424),
.Y(n_530)
);

NAND2xp33_ASAP7_75t_L g531 ( 
.A(n_472),
.B(n_169),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_453),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_463),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_433),
.B(n_375),
.Y(n_534)
);

BUFx10_ASAP7_75t_L g535 ( 
.A(n_435),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_416),
.B(n_474),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_436),
.B(n_353),
.Y(n_537)
);

INVx4_ASAP7_75t_L g538 ( 
.A(n_453),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_426),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_436),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_416),
.B(n_188),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_458),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_445),
.B(n_389),
.Y(n_543)
);

INVx4_ASAP7_75t_L g544 ( 
.A(n_453),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_429),
.Y(n_545)
);

NAND3xp33_ASAP7_75t_L g546 ( 
.A(n_472),
.B(n_405),
.C(n_400),
.Y(n_546)
);

INVx4_ASAP7_75t_L g547 ( 
.A(n_453),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_474),
.B(n_199),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_460),
.Y(n_549)
);

BUFx10_ASAP7_75t_L g550 ( 
.A(n_449),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_462),
.B(n_395),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_436),
.B(n_392),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_476),
.B(n_214),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_467),
.B(n_330),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_460),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_456),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_469),
.B(n_374),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_429),
.Y(n_558)
);

BUFx2_ASAP7_75t_L g559 ( 
.A(n_463),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_437),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_470),
.B(n_397),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_437),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_440),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_476),
.B(n_227),
.Y(n_564)
);

AND2x4_ASAP7_75t_L g565 ( 
.A(n_479),
.B(n_444),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_477),
.B(n_358),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_444),
.B(n_427),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_461),
.B(n_359),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_450),
.B(n_443),
.Y(n_569)
);

BUFx4_ASAP7_75t_L g570 ( 
.A(n_443),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_456),
.Y(n_571)
);

NAND2xp33_ASAP7_75t_L g572 ( 
.A(n_424),
.B(n_444),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_479),
.B(n_372),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_456),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_456),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_427),
.B(n_234),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_479),
.A2(n_388),
.B1(n_394),
.B2(n_222),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_L g578 ( 
.A1(n_479),
.A2(n_394),
.B1(n_232),
.B2(n_322),
.Y(n_578)
);

BUFx4f_ASAP7_75t_L g579 ( 
.A(n_451),
.Y(n_579)
);

BUFx4f_ASAP7_75t_L g580 ( 
.A(n_451),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_440),
.B(n_236),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_460),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_446),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_466),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_479),
.B(n_182),
.Y(n_585)
);

INVx4_ASAP7_75t_L g586 ( 
.A(n_456),
.Y(n_586)
);

INVx4_ASAP7_75t_L g587 ( 
.A(n_456),
.Y(n_587)
);

INVx2_ASAP7_75t_SL g588 ( 
.A(n_479),
.Y(n_588)
);

OR2x2_ASAP7_75t_L g589 ( 
.A(n_455),
.B(n_240),
.Y(n_589)
);

BUFx10_ASAP7_75t_L g590 ( 
.A(n_424),
.Y(n_590)
);

OAI22xp33_ASAP7_75t_L g591 ( 
.A1(n_455),
.A2(n_239),
.B1(n_244),
.B2(n_243),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_466),
.Y(n_592)
);

AND2x6_ASAP7_75t_L g593 ( 
.A(n_446),
.B(n_237),
.Y(n_593)
);

OAI22xp33_ASAP7_75t_SL g594 ( 
.A1(n_464),
.A2(n_315),
.B1(n_295),
.B2(n_287),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_466),
.Y(n_595)
);

INVxp67_ASAP7_75t_SL g596 ( 
.A(n_457),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_464),
.B(n_264),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_465),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_451),
.B(n_249),
.Y(n_599)
);

INVx4_ASAP7_75t_L g600 ( 
.A(n_457),
.Y(n_600)
);

AND2x6_ASAP7_75t_L g601 ( 
.A(n_465),
.B(n_269),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_475),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_475),
.B(n_182),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_441),
.B(n_185),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_459),
.Y(n_605)
);

NAND2xp33_ASAP7_75t_SL g606 ( 
.A(n_459),
.B(n_323),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_478),
.Y(n_607)
);

OA22x2_ASAP7_75t_L g608 ( 
.A1(n_420),
.A2(n_266),
.B1(n_320),
.B2(n_253),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_457),
.Y(n_609)
);

AND2x4_ASAP7_75t_L g610 ( 
.A(n_420),
.B(n_270),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_407),
.Y(n_611)
);

BUFx8_ASAP7_75t_SL g612 ( 
.A(n_418),
.Y(n_612)
);

OAI22xp5_ASAP7_75t_L g613 ( 
.A1(n_459),
.A2(n_275),
.B1(n_220),
.B2(n_229),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_478),
.B(n_255),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_457),
.B(n_185),
.Y(n_615)
);

NAND3xp33_ASAP7_75t_L g616 ( 
.A(n_459),
.B(n_278),
.C(n_268),
.Y(n_616)
);

AND3x2_ASAP7_75t_L g617 ( 
.A(n_478),
.B(n_327),
.C(n_311),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_471),
.Y(n_618)
);

AND3x1_ASAP7_75t_L g619 ( 
.A(n_471),
.B(n_263),
.C(n_257),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g620 ( 
.A(n_420),
.B(n_271),
.Y(n_620)
);

AND2x4_ASAP7_75t_L g621 ( 
.A(n_447),
.B(n_282),
.Y(n_621)
);

INVx1_ASAP7_75t_SL g622 ( 
.A(n_421),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_471),
.B(n_285),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_471),
.B(n_187),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_424),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_447),
.B(n_291),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_413),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_457),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_447),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_413),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_502),
.B(n_221),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_496),
.B(n_187),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_491),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_480),
.B(n_191),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_498),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_520),
.B(n_457),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_522),
.B(n_293),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_627),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_491),
.Y(n_639)
);

BUFx3_ASAP7_75t_L g640 ( 
.A(n_612),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_501),
.B(n_296),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_481),
.B(n_191),
.Y(n_642)
);

INVx2_ASAP7_75t_SL g643 ( 
.A(n_502),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_L g644 ( 
.A1(n_599),
.A2(n_308),
.B1(n_302),
.B2(n_306),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_515),
.B(n_565),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_L g646 ( 
.A(n_568),
.B(n_192),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_501),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_565),
.B(n_192),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_505),
.B(n_195),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_552),
.B(n_301),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_486),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_552),
.B(n_423),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_490),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_494),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_536),
.B(n_423),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_505),
.B(n_195),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_493),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_565),
.B(n_198),
.Y(n_658)
);

AOI22xp5_ASAP7_75t_L g659 ( 
.A1(n_546),
.A2(n_290),
.B1(n_304),
.B2(n_326),
.Y(n_659)
);

OAI22xp5_ASAP7_75t_L g660 ( 
.A1(n_588),
.A2(n_198),
.B1(n_290),
.B2(n_289),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_573),
.B(n_289),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_540),
.B(n_423),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_599),
.A2(n_166),
.B1(n_173),
.B2(n_176),
.Y(n_663)
);

AOI22xp5_ASAP7_75t_L g664 ( 
.A1(n_585),
.A2(n_312),
.B1(n_309),
.B2(n_326),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_493),
.B(n_300),
.Y(n_665)
);

AOI22xp33_ASAP7_75t_L g666 ( 
.A1(n_608),
.A2(n_297),
.B1(n_176),
.B2(n_189),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_499),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_588),
.A2(n_318),
.B1(n_304),
.B2(n_309),
.Y(n_668)
);

NAND3xp33_ASAP7_75t_L g669 ( 
.A(n_606),
.B(n_238),
.C(n_259),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_537),
.B(n_300),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_626),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_485),
.B(n_221),
.Y(n_672)
);

INVx8_ASAP7_75t_L g673 ( 
.A(n_498),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_627),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_540),
.B(n_423),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_483),
.B(n_442),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_630),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_608),
.A2(n_297),
.B1(n_189),
.B2(n_194),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_630),
.Y(n_679)
);

AND2x6_ASAP7_75t_SL g680 ( 
.A(n_557),
.B(n_173),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_567),
.B(n_442),
.Y(n_681)
);

AOI22xp33_ASAP7_75t_L g682 ( 
.A1(n_608),
.A2(n_299),
.B1(n_197),
.B2(n_201),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_484),
.Y(n_683)
);

NAND3xp33_ASAP7_75t_L g684 ( 
.A(n_606),
.B(n_260),
.C(n_261),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_487),
.B(n_442),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_484),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_537),
.B(n_312),
.Y(n_687)
);

A2O1A1Ixp33_ASAP7_75t_L g688 ( 
.A1(n_495),
.A2(n_324),
.B(n_316),
.C(n_318),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_531),
.A2(n_299),
.B1(n_197),
.B2(n_201),
.Y(n_689)
);

AOI22xp33_ASAP7_75t_L g690 ( 
.A1(n_531),
.A2(n_307),
.B1(n_246),
.B2(n_292),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_497),
.Y(n_691)
);

INVxp67_ASAP7_75t_L g692 ( 
.A(n_504),
.Y(n_692)
);

OR2x2_ASAP7_75t_L g693 ( 
.A(n_504),
.B(n_194),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_495),
.A2(n_580),
.B1(n_521),
.B2(n_579),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_503),
.B(n_324),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_499),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_577),
.B(n_578),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_624),
.B(n_442),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_612),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_497),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_548),
.B(n_553),
.Y(n_701)
);

OAI22xp5_ASAP7_75t_L g702 ( 
.A1(n_514),
.A2(n_319),
.B1(n_316),
.B2(n_276),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_564),
.B(n_319),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_528),
.B(n_438),
.Y(n_704)
);

NAND3xp33_ASAP7_75t_SL g705 ( 
.A(n_507),
.B(n_246),
.C(n_317),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_589),
.B(n_265),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_529),
.B(n_438),
.Y(n_707)
);

OR2x2_ASAP7_75t_L g708 ( 
.A(n_559),
.B(n_482),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_561),
.B(n_267),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_558),
.B(n_438),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_626),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_560),
.B(n_434),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_510),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_495),
.A2(n_521),
.B1(n_579),
.B2(n_580),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_510),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_512),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_583),
.B(n_434),
.Y(n_717)
);

INVxp67_ASAP7_75t_L g718 ( 
.A(n_559),
.Y(n_718)
);

OR2x2_ASAP7_75t_L g719 ( 
.A(n_533),
.B(n_298),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_512),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_598),
.B(n_602),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_498),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_L g723 ( 
.A1(n_521),
.A2(n_307),
.B1(n_292),
.B2(n_294),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_513),
.Y(n_724)
);

NAND3xp33_ASAP7_75t_L g725 ( 
.A(n_616),
.B(n_277),
.C(n_284),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_513),
.B(n_434),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_518),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_518),
.B(n_428),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_500),
.Y(n_729)
);

INVx4_ASAP7_75t_L g730 ( 
.A(n_498),
.Y(n_730)
);

NAND3xp33_ASAP7_75t_L g731 ( 
.A(n_589),
.B(n_317),
.C(n_313),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_523),
.B(n_428),
.Y(n_732)
);

O2A1O1Ixp5_ASAP7_75t_L g733 ( 
.A1(n_579),
.A2(n_428),
.B(n_413),
.C(n_424),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_523),
.B(n_424),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_591),
.B(n_535),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_541),
.B(n_603),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_539),
.B(n_424),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_539),
.B(n_294),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_535),
.B(n_313),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_545),
.B(n_298),
.Y(n_740)
);

AOI22xp5_ASAP7_75t_L g741 ( 
.A1(n_615),
.A2(n_424),
.B1(n_60),
.B2(n_73),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_545),
.Y(n_742)
);

HB1xp67_ASAP7_75t_L g743 ( 
.A(n_619),
.Y(n_743)
);

BUFx5_ASAP7_75t_L g744 ( 
.A(n_590),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_562),
.B(n_152),
.Y(n_745)
);

OAI22xp5_ASAP7_75t_L g746 ( 
.A1(n_580),
.A2(n_151),
.B1(n_139),
.B2(n_136),
.Y(n_746)
);

OR2x6_ASAP7_75t_L g747 ( 
.A(n_569),
.B(n_16),
.Y(n_747)
);

INVx2_ASAP7_75t_SL g748 ( 
.A(n_570),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_535),
.B(n_17),
.Y(n_749)
);

INVx2_ASAP7_75t_SL g750 ( 
.A(n_570),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_562),
.Y(n_751)
);

AOI21x1_ASAP7_75t_L g752 ( 
.A1(n_623),
.A2(n_135),
.B(n_128),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_550),
.B(n_594),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_563),
.B(n_19),
.Y(n_754)
);

NOR2xp67_ASAP7_75t_L g755 ( 
.A(n_519),
.B(n_121),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_550),
.B(n_20),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_550),
.B(n_20),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_566),
.B(n_23),
.Y(n_758)
);

AOI22xp33_ASAP7_75t_L g759 ( 
.A1(n_610),
.A2(n_24),
.B1(n_26),
.B2(n_28),
.Y(n_759)
);

A2O1A1Ixp33_ASAP7_75t_L g760 ( 
.A1(n_563),
.A2(n_24),
.B(n_30),
.C(n_31),
.Y(n_760)
);

AND2x6_ASAP7_75t_SL g761 ( 
.A(n_527),
.B(n_30),
.Y(n_761)
);

AOI21xp5_ASAP7_75t_L g762 ( 
.A1(n_596),
.A2(n_113),
.B(n_104),
.Y(n_762)
);

INVx1_ASAP7_75t_SL g763 ( 
.A(n_611),
.Y(n_763)
);

OAI22xp5_ASAP7_75t_L g764 ( 
.A1(n_576),
.A2(n_98),
.B1(n_97),
.B2(n_96),
.Y(n_764)
);

INVxp67_ASAP7_75t_L g765 ( 
.A(n_534),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_618),
.B(n_94),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_614),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_614),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_500),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_625),
.B(n_31),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_625),
.B(n_32),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_618),
.B(n_605),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_524),
.Y(n_773)
);

AOI22xp33_ASAP7_75t_L g774 ( 
.A1(n_610),
.A2(n_32),
.B1(n_33),
.B2(n_39),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_613),
.B(n_33),
.Y(n_775)
);

OR2x2_ASAP7_75t_L g776 ( 
.A(n_622),
.B(n_40),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_488),
.B(n_556),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_604),
.B(n_41),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_590),
.B(n_530),
.Y(n_779)
);

OAI22xp33_ASAP7_75t_L g780 ( 
.A1(n_581),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_488),
.B(n_79),
.Y(n_781)
);

INVx2_ASAP7_75t_SL g782 ( 
.A(n_611),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_524),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_488),
.B(n_77),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_554),
.B(n_597),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_572),
.A2(n_85),
.B1(n_87),
.B2(n_90),
.Y(n_786)
);

NOR3xp33_ASAP7_75t_L g787 ( 
.A(n_517),
.B(n_47),
.C(n_51),
.Y(n_787)
);

AOI22xp5_ASAP7_75t_L g788 ( 
.A1(n_572),
.A2(n_47),
.B1(n_54),
.B2(n_593),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_621),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_590),
.B(n_54),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_489),
.B(n_571),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_489),
.B(n_571),
.Y(n_792)
);

AO22x1_ASAP7_75t_L g793 ( 
.A1(n_610),
.A2(n_620),
.B1(n_593),
.B2(n_601),
.Y(n_793)
);

NOR2xp67_ASAP7_75t_L g794 ( 
.A(n_543),
.B(n_551),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_489),
.B(n_574),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_530),
.B(n_621),
.Y(n_796)
);

BUFx6f_ASAP7_75t_L g797 ( 
.A(n_506),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_511),
.B(n_574),
.Y(n_798)
);

OAI22xp33_ASAP7_75t_L g799 ( 
.A1(n_629),
.A2(n_595),
.B1(n_542),
.B2(n_592),
.Y(n_799)
);

INVx5_ASAP7_75t_L g800 ( 
.A(n_593),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_617),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_511),
.B(n_571),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_631),
.B(n_508),
.Y(n_803)
);

OAI21xp5_ASAP7_75t_L g804 ( 
.A1(n_733),
.A2(n_620),
.B(n_549),
.Y(n_804)
);

AOI21x1_ASAP7_75t_L g805 ( 
.A1(n_796),
.A2(n_629),
.B(n_620),
.Y(n_805)
);

A2O1A1Ixp33_ASAP7_75t_L g806 ( 
.A1(n_632),
.A2(n_556),
.B(n_609),
.C(n_574),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_701),
.B(n_516),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_701),
.B(n_516),
.Y(n_808)
);

INVx3_ASAP7_75t_L g809 ( 
.A(n_797),
.Y(n_809)
);

OAI21xp5_ASAP7_75t_L g810 ( 
.A1(n_694),
.A2(n_555),
.B(n_549),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_789),
.Y(n_811)
);

INVx3_ASAP7_75t_SL g812 ( 
.A(n_699),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_655),
.A2(n_492),
.B(n_600),
.Y(n_813)
);

A2O1A1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_632),
.A2(n_556),
.B(n_609),
.C(n_575),
.Y(n_814)
);

BUFx12f_ASAP7_75t_L g815 ( 
.A(n_748),
.Y(n_815)
);

OAI21xp5_ASAP7_75t_L g816 ( 
.A1(n_694),
.A2(n_555),
.B(n_582),
.Y(n_816)
);

OR2x2_ASAP7_75t_L g817 ( 
.A(n_692),
.B(n_525),
.Y(n_817)
);

OAI21xp5_ASAP7_75t_L g818 ( 
.A1(n_714),
.A2(n_652),
.B(n_697),
.Y(n_818)
);

OR2x6_ASAP7_75t_SL g819 ( 
.A(n_708),
.B(n_669),
.Y(n_819)
);

INVx4_ASAP7_75t_L g820 ( 
.A(n_635),
.Y(n_820)
);

OAI21xp5_ASAP7_75t_L g821 ( 
.A1(n_714),
.A2(n_582),
.B(n_584),
.Y(n_821)
);

AO32x1_ASAP7_75t_L g822 ( 
.A1(n_746),
.A2(n_607),
.A3(n_595),
.B1(n_592),
.B2(n_584),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_634),
.B(n_609),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_681),
.A2(n_492),
.B(n_600),
.Y(n_824)
);

AOI22xp5_ASAP7_75t_L g825 ( 
.A1(n_645),
.A2(n_601),
.B1(n_593),
.B2(n_628),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_633),
.Y(n_826)
);

A2O1A1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_646),
.A2(n_575),
.B(n_511),
.C(n_516),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_718),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_639),
.Y(n_829)
);

BUFx4f_ASAP7_75t_L g830 ( 
.A(n_750),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_634),
.B(n_642),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_785),
.B(n_530),
.Y(n_832)
);

NOR2xp67_ASAP7_75t_L g833 ( 
.A(n_765),
.B(n_525),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_642),
.B(n_628),
.Y(n_834)
);

AND2x4_ASAP7_75t_L g835 ( 
.A(n_647),
.B(n_492),
.Y(n_835)
);

AND2x2_ASAP7_75t_SL g836 ( 
.A(n_759),
.B(n_544),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_703),
.B(n_601),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_793),
.A2(n_544),
.B(n_600),
.Y(n_838)
);

INVxp67_ASAP7_75t_L g839 ( 
.A(n_672),
.Y(n_839)
);

A2O1A1Ixp33_ASAP7_75t_L g840 ( 
.A1(n_736),
.A2(n_703),
.B(n_656),
.C(n_649),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_636),
.A2(n_544),
.B(n_587),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_683),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_695),
.B(n_601),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_736),
.A2(n_601),
.B1(n_593),
.B2(n_538),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_695),
.B(n_657),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_686),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_640),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_671),
.B(n_601),
.Y(n_848)
);

AND2x4_ASAP7_75t_L g849 ( 
.A(n_667),
.B(n_696),
.Y(n_849)
);

A2O1A1Ixp33_ASAP7_75t_L g850 ( 
.A1(n_706),
.A2(n_709),
.B(n_785),
.C(n_778),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_L g851 ( 
.A1(n_644),
.A2(n_593),
.B1(n_509),
.B2(n_526),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_662),
.A2(n_587),
.B(n_586),
.Y(n_852)
);

O2A1O1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_775),
.A2(n_530),
.B(n_509),
.C(n_526),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_711),
.B(n_586),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_643),
.B(n_587),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_675),
.A2(n_586),
.B(n_547),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_698),
.A2(n_547),
.B(n_538),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_767),
.B(n_538),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_691),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_768),
.B(n_547),
.Y(n_860)
);

AOI22xp5_ASAP7_75t_L g861 ( 
.A1(n_735),
.A2(n_650),
.B1(n_794),
.B2(n_706),
.Y(n_861)
);

A2O1A1Ixp33_ASAP7_75t_L g862 ( 
.A1(n_738),
.A2(n_740),
.B(n_754),
.C(n_644),
.Y(n_862)
);

AOI21xp5_ASAP7_75t_L g863 ( 
.A1(n_777),
.A2(n_530),
.B(n_509),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_791),
.A2(n_506),
.B(n_509),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_713),
.Y(n_865)
);

INVx4_ASAP7_75t_L g866 ( 
.A(n_635),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_705),
.B(n_506),
.Y(n_867)
);

AO22x1_ASAP7_75t_L g868 ( 
.A1(n_787),
.A2(n_506),
.B1(n_509),
.B2(n_526),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_792),
.A2(n_506),
.B(n_526),
.Y(n_869)
);

BUFx2_ASAP7_75t_L g870 ( 
.A(n_747),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_693),
.B(n_670),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_743),
.B(n_526),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_797),
.Y(n_873)
);

OAI22xp5_ASAP7_75t_L g874 ( 
.A1(n_759),
.A2(n_532),
.B1(n_774),
.B2(n_663),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_776),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_795),
.A2(n_532),
.B(n_802),
.Y(n_876)
);

OAI22xp5_ASAP7_75t_L g877 ( 
.A1(n_774),
.A2(n_532),
.B1(n_663),
.B2(n_682),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_685),
.A2(n_532),
.B(n_676),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_715),
.B(n_532),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_779),
.A2(n_800),
.B(n_798),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_800),
.A2(n_798),
.B(n_772),
.Y(n_881)
);

AND2x2_ASAP7_75t_SL g882 ( 
.A(n_723),
.B(n_666),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_716),
.B(n_720),
.Y(n_883)
);

NOR2xp67_ASAP7_75t_L g884 ( 
.A(n_782),
.B(n_725),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_724),
.B(n_727),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_687),
.B(n_738),
.Y(n_886)
);

OAI22xp5_ASAP7_75t_L g887 ( 
.A1(n_666),
.A2(n_682),
.B1(n_678),
.B2(n_723),
.Y(n_887)
);

INVx5_ASAP7_75t_L g888 ( 
.A(n_635),
.Y(n_888)
);

A2O1A1Ixp33_ASAP7_75t_L g889 ( 
.A1(n_740),
.A2(n_754),
.B(n_742),
.C(n_751),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_R g890 ( 
.A(n_763),
.B(n_719),
.Y(n_890)
);

AO32x2_ASAP7_75t_L g891 ( 
.A1(n_660),
.A2(n_764),
.A3(n_702),
.B1(n_678),
.B2(n_801),
.Y(n_891)
);

NAND2x1_ASAP7_75t_L g892 ( 
.A(n_730),
.B(n_635),
.Y(n_892)
);

AOI21xp33_ASAP7_75t_L g893 ( 
.A1(n_661),
.A2(n_664),
.B(n_684),
.Y(n_893)
);

OAI21xp5_ASAP7_75t_L g894 ( 
.A1(n_688),
.A2(n_799),
.B(n_637),
.Y(n_894)
);

O2A1O1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_770),
.A2(n_771),
.B(n_790),
.C(n_760),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_651),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_800),
.A2(n_721),
.B(n_797),
.Y(n_897)
);

INVx1_ASAP7_75t_SL g898 ( 
.A(n_743),
.Y(n_898)
);

NAND2xp33_ASAP7_75t_L g899 ( 
.A(n_722),
.B(n_744),
.Y(n_899)
);

O2A1O1Ixp33_ASAP7_75t_L g900 ( 
.A1(n_641),
.A2(n_758),
.B(n_665),
.C(n_780),
.Y(n_900)
);

O2A1O1Ixp5_ASAP7_75t_L g901 ( 
.A1(n_799),
.A2(n_745),
.B(n_653),
.C(n_654),
.Y(n_901)
);

OAI21x1_ASAP7_75t_L g902 ( 
.A1(n_781),
.A2(n_784),
.B(n_734),
.Y(n_902)
);

O2A1O1Ixp33_ASAP7_75t_SL g903 ( 
.A1(n_766),
.A2(n_737),
.B(n_788),
.C(n_658),
.Y(n_903)
);

AOI22xp5_ASAP7_75t_L g904 ( 
.A1(n_755),
.A2(n_648),
.B1(n_753),
.B2(n_731),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_700),
.B(n_773),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_797),
.Y(n_906)
);

OAI22xp5_ASAP7_75t_L g907 ( 
.A1(n_689),
.A2(n_690),
.B1(n_747),
.B2(n_659),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_729),
.B(n_783),
.Y(n_908)
);

INVx3_ASAP7_75t_L g909 ( 
.A(n_769),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_800),
.A2(n_730),
.B(n_673),
.Y(n_910)
);

OR2x2_ASAP7_75t_L g911 ( 
.A(n_739),
.B(n_668),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_673),
.A2(n_722),
.B(n_732),
.Y(n_912)
);

INVx1_ASAP7_75t_SL g913 ( 
.A(n_747),
.Y(n_913)
);

AOI22xp33_ASAP7_75t_L g914 ( 
.A1(n_689),
.A2(n_690),
.B1(n_638),
.B2(n_674),
.Y(n_914)
);

OAI21xp5_ASAP7_75t_L g915 ( 
.A1(n_726),
.A2(n_728),
.B(n_704),
.Y(n_915)
);

BUFx2_ASAP7_75t_L g916 ( 
.A(n_680),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_677),
.B(n_679),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_707),
.Y(n_918)
);

AO22x1_ASAP7_75t_L g919 ( 
.A1(n_780),
.A2(n_761),
.B1(n_756),
.B2(n_749),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_710),
.B(n_712),
.Y(n_920)
);

OAI21xp5_ASAP7_75t_L g921 ( 
.A1(n_717),
.A2(n_786),
.B(n_741),
.Y(n_921)
);

OAI22xp5_ASAP7_75t_L g922 ( 
.A1(n_722),
.A2(n_673),
.B1(n_757),
.B2(n_762),
.Y(n_922)
);

OAI22xp5_ASAP7_75t_L g923 ( 
.A1(n_722),
.A2(n_774),
.B1(n_759),
.B2(n_644),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_744),
.B(n_752),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_744),
.A2(n_498),
.B(n_655),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_744),
.A2(n_498),
.B(n_655),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_744),
.B(n_701),
.Y(n_927)
);

NOR2xp33_ASAP7_75t_L g928 ( 
.A(n_744),
.B(n_642),
.Y(n_928)
);

O2A1O1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_632),
.A2(n_531),
.B(n_697),
.C(n_775),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_655),
.A2(n_498),
.B(n_652),
.Y(n_930)
);

INVx3_ASAP7_75t_L g931 ( 
.A(n_797),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_797),
.Y(n_932)
);

HB1xp67_ASAP7_75t_L g933 ( 
.A(n_718),
.Y(n_933)
);

BUFx3_ASAP7_75t_L g934 ( 
.A(n_640),
.Y(n_934)
);

CKINVDCx10_ASAP7_75t_R g935 ( 
.A(n_699),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_701),
.B(n_632),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_633),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_655),
.A2(n_498),
.B(n_652),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_789),
.Y(n_939)
);

OR2x2_ASAP7_75t_L g940 ( 
.A(n_692),
.B(n_431),
.Y(n_940)
);

O2A1O1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_632),
.A2(n_531),
.B(n_697),
.C(n_775),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_631),
.B(n_431),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_655),
.A2(n_498),
.B(n_652),
.Y(n_943)
);

NAND2x1p5_ASAP7_75t_L g944 ( 
.A(n_635),
.B(n_722),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_655),
.A2(n_498),
.B(n_652),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_642),
.B(n_765),
.Y(n_946)
);

AO21x2_ASAP7_75t_L g947 ( 
.A1(n_799),
.A2(n_645),
.B(n_688),
.Y(n_947)
);

O2A1O1Ixp33_ASAP7_75t_SL g948 ( 
.A1(n_688),
.A2(n_745),
.B(n_775),
.C(n_766),
.Y(n_948)
);

OAI21xp5_ASAP7_75t_L g949 ( 
.A1(n_733),
.A2(n_521),
.B(n_495),
.Y(n_949)
);

OAI21xp33_ASAP7_75t_L g950 ( 
.A1(n_646),
.A2(n_632),
.B(n_642),
.Y(n_950)
);

NOR2x1_ASAP7_75t_L g951 ( 
.A(n_755),
.B(n_508),
.Y(n_951)
);

OAI22xp5_ASAP7_75t_L g952 ( 
.A1(n_759),
.A2(n_774),
.B1(n_644),
.B2(n_632),
.Y(n_952)
);

A2O1A1Ixp33_ASAP7_75t_L g953 ( 
.A1(n_632),
.A2(n_701),
.B(n_646),
.C(n_496),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_701),
.B(n_632),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_655),
.A2(n_498),
.B(n_652),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_701),
.B(n_632),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_642),
.B(n_765),
.Y(n_957)
);

NAND3xp33_ASAP7_75t_L g958 ( 
.A(n_632),
.B(n_646),
.C(n_642),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_701),
.B(n_632),
.Y(n_959)
);

INVx3_ASAP7_75t_L g960 ( 
.A(n_797),
.Y(n_960)
);

AOI22xp33_ASAP7_75t_L g961 ( 
.A1(n_632),
.A2(n_505),
.B1(n_701),
.B2(n_697),
.Y(n_961)
);

INVx3_ASAP7_75t_L g962 ( 
.A(n_797),
.Y(n_962)
);

A2O1A1Ixp33_ASAP7_75t_L g963 ( 
.A1(n_632),
.A2(n_701),
.B(n_646),
.C(n_496),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_789),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_655),
.A2(n_498),
.B(n_652),
.Y(n_965)
);

NOR3xp33_ASAP7_75t_L g966 ( 
.A(n_646),
.B(n_642),
.C(n_443),
.Y(n_966)
);

A2O1A1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_632),
.A2(n_701),
.B(n_646),
.C(n_496),
.Y(n_967)
);

BUFx3_ASAP7_75t_L g968 ( 
.A(n_640),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_655),
.A2(n_498),
.B(n_652),
.Y(n_969)
);

OAI21xp33_ASAP7_75t_L g970 ( 
.A1(n_646),
.A2(n_632),
.B(n_642),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_655),
.A2(n_498),
.B(n_652),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_655),
.A2(n_498),
.B(n_652),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_633),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_701),
.B(n_632),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_631),
.B(n_431),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_655),
.A2(n_498),
.B(n_652),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_701),
.B(n_632),
.Y(n_977)
);

INVx3_ASAP7_75t_L g978 ( 
.A(n_797),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_701),
.B(n_632),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_797),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_789),
.Y(n_981)
);

AOI22xp5_ASAP7_75t_L g982 ( 
.A1(n_632),
.A2(n_701),
.B1(n_645),
.B2(n_642),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_633),
.B(n_639),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_642),
.B(n_765),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_701),
.B(n_632),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_655),
.A2(n_498),
.B(n_652),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_SL g987 ( 
.A(n_701),
.B(n_632),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_797),
.Y(n_988)
);

BUFx2_ASAP7_75t_L g989 ( 
.A(n_890),
.Y(n_989)
);

INVx2_ASAP7_75t_SL g990 ( 
.A(n_828),
.Y(n_990)
);

OAI21x1_ASAP7_75t_L g991 ( 
.A1(n_876),
.A2(n_804),
.B(n_864),
.Y(n_991)
);

BUFx8_ASAP7_75t_L g992 ( 
.A(n_815),
.Y(n_992)
);

AOI21x1_ASAP7_75t_L g993 ( 
.A1(n_924),
.A2(n_832),
.B(n_823),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_936),
.B(n_954),
.Y(n_994)
);

NAND2xp33_ASAP7_75t_L g995 ( 
.A(n_952),
.B(n_923),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_956),
.B(n_959),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_950),
.B(n_970),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_974),
.A2(n_979),
.B1(n_985),
.B2(n_963),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_952),
.A2(n_967),
.B(n_953),
.C(n_850),
.Y(n_999)
);

A2O1A1Ixp33_ASAP7_75t_L g1000 ( 
.A1(n_923),
.A2(n_840),
.B(n_862),
.C(n_958),
.Y(n_1000)
);

OAI21x1_ASAP7_75t_L g1001 ( 
.A1(n_804),
.A2(n_869),
.B(n_816),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_831),
.B(n_946),
.Y(n_1002)
);

OAI21x1_ASAP7_75t_L g1003 ( 
.A1(n_810),
.A2(n_821),
.B(n_816),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_957),
.B(n_984),
.Y(n_1004)
);

A2O1A1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_874),
.A2(n_982),
.B(n_887),
.C(n_977),
.Y(n_1005)
);

OAI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_987),
.A2(n_941),
.B(n_929),
.Y(n_1006)
);

BUFx8_ASAP7_75t_L g1007 ( 
.A(n_870),
.Y(n_1007)
);

OR2x2_ASAP7_75t_L g1008 ( 
.A(n_940),
.B(n_942),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_899),
.A2(n_927),
.B(n_928),
.Y(n_1009)
);

AOI21x1_ASAP7_75t_L g1010 ( 
.A1(n_930),
.A2(n_943),
.B(n_938),
.Y(n_1010)
);

OAI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_961),
.A2(n_836),
.B1(n_861),
.B2(n_882),
.Y(n_1011)
);

OAI21x1_ASAP7_75t_L g1012 ( 
.A1(n_810),
.A2(n_821),
.B(n_852),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_983),
.B(n_811),
.Y(n_1013)
);

AOI21x1_ASAP7_75t_L g1014 ( 
.A1(n_945),
.A2(n_965),
.B(n_955),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_845),
.B(n_975),
.Y(n_1015)
);

OAI21x1_ASAP7_75t_L g1016 ( 
.A1(n_856),
.A2(n_926),
.B(n_925),
.Y(n_1016)
);

OAI21x1_ASAP7_75t_L g1017 ( 
.A1(n_838),
.A2(n_805),
.B(n_841),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_969),
.A2(n_972),
.B(n_971),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_976),
.A2(n_986),
.B(n_843),
.Y(n_1019)
);

OAI21x1_ASAP7_75t_L g1020 ( 
.A1(n_912),
.A2(n_878),
.B(n_824),
.Y(n_1020)
);

OAI21xp33_ASAP7_75t_L g1021 ( 
.A1(n_886),
.A2(n_907),
.B(n_887),
.Y(n_1021)
);

OAI21x1_ASAP7_75t_L g1022 ( 
.A1(n_813),
.A2(n_857),
.B(n_902),
.Y(n_1022)
);

A2O1A1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_874),
.A2(n_877),
.B(n_907),
.C(n_900),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_920),
.A2(n_837),
.B(n_949),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_949),
.A2(n_807),
.B(n_808),
.Y(n_1025)
);

OR2x2_ASAP7_75t_L g1026 ( 
.A(n_898),
.B(n_933),
.Y(n_1026)
);

OAI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_818),
.A2(n_894),
.B(n_901),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_881),
.A2(n_888),
.B(n_834),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_888),
.A2(n_903),
.B(n_915),
.Y(n_1029)
);

OAI21x1_ASAP7_75t_L g1030 ( 
.A1(n_880),
.A2(n_863),
.B(n_897),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_820),
.Y(n_1031)
);

AOI221xp5_ASAP7_75t_SL g1032 ( 
.A1(n_877),
.A2(n_889),
.B1(n_839),
.B2(n_865),
.C(n_883),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_817),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_871),
.B(n_898),
.Y(n_1034)
);

BUFx4f_ASAP7_75t_L g1035 ( 
.A(n_812),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_888),
.A2(n_915),
.B(n_851),
.Y(n_1036)
);

OAI21x1_ASAP7_75t_L g1037 ( 
.A1(n_910),
.A2(n_879),
.B(n_944),
.Y(n_1037)
);

INVx4_ASAP7_75t_L g1038 ( 
.A(n_888),
.Y(n_1038)
);

AOI21xp33_ASAP7_75t_L g1039 ( 
.A1(n_911),
.A2(n_895),
.B(n_893),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_939),
.Y(n_1040)
);

AND3x4_ASAP7_75t_L g1041 ( 
.A(n_966),
.B(n_849),
.C(n_884),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_921),
.A2(n_948),
.B(n_848),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_918),
.B(n_833),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_885),
.B(n_872),
.Y(n_1044)
);

CKINVDCx20_ASAP7_75t_R g1045 ( 
.A(n_847),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_875),
.B(n_913),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_854),
.A2(n_858),
.B(n_860),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_964),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_906),
.Y(n_1049)
);

NAND3xp33_ASAP7_75t_SL g1050 ( 
.A(n_904),
.B(n_803),
.C(n_913),
.Y(n_1050)
);

AO31x2_ASAP7_75t_L g1051 ( 
.A1(n_806),
.A2(n_814),
.A3(n_827),
.B(n_867),
.Y(n_1051)
);

OAI21x1_ASAP7_75t_L g1052 ( 
.A1(n_944),
.A2(n_892),
.B(n_908),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_844),
.A2(n_914),
.B1(n_825),
.B2(n_896),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_981),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_849),
.B(n_937),
.Y(n_1055)
);

CKINVDCx20_ASAP7_75t_R g1056 ( 
.A(n_934),
.Y(n_1056)
);

OAI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_905),
.A2(n_917),
.B(n_853),
.Y(n_1057)
);

INVx3_ASAP7_75t_L g1058 ( 
.A(n_820),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_855),
.A2(n_922),
.B(n_835),
.Y(n_1059)
);

CKINVDCx20_ASAP7_75t_R g1060 ( 
.A(n_968),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_973),
.B(n_829),
.Y(n_1061)
);

OAI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_842),
.A2(n_859),
.B(n_846),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_835),
.A2(n_947),
.B(n_866),
.Y(n_1063)
);

AO21x1_ASAP7_75t_L g1064 ( 
.A1(n_826),
.A2(n_983),
.B(n_866),
.Y(n_1064)
);

AOI21xp33_ASAP7_75t_L g1065 ( 
.A1(n_951),
.A2(n_947),
.B(n_909),
.Y(n_1065)
);

NAND2x1p5_ASAP7_75t_L g1066 ( 
.A(n_906),
.B(n_988),
.Y(n_1066)
);

OAI21x1_ASAP7_75t_L g1067 ( 
.A1(n_809),
.A2(n_960),
.B(n_931),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_906),
.A2(n_988),
.B(n_980),
.Y(n_1068)
);

OAI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_909),
.A2(n_809),
.B(n_962),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_932),
.A2(n_980),
.B(n_988),
.Y(n_1070)
);

AOI21x1_ASAP7_75t_L g1071 ( 
.A1(n_868),
.A2(n_919),
.B(n_822),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_932),
.A2(n_980),
.B(n_931),
.Y(n_1072)
);

OAI21x1_ASAP7_75t_L g1073 ( 
.A1(n_978),
.A2(n_962),
.B(n_960),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_932),
.B(n_978),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_873),
.A2(n_822),
.B(n_891),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_819),
.B(n_873),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_822),
.A2(n_830),
.B(n_891),
.Y(n_1077)
);

A2O1A1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_830),
.A2(n_891),
.B(n_916),
.C(n_935),
.Y(n_1078)
);

OAI21x1_ASAP7_75t_L g1079 ( 
.A1(n_876),
.A2(n_804),
.B(n_864),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_L g1080 ( 
.A(n_936),
.B(n_954),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_SL g1081 ( 
.A1(n_923),
.A2(n_952),
.B(n_730),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_982),
.B(n_950),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_936),
.B(n_954),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_865),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_899),
.A2(n_714),
.B(n_694),
.Y(n_1085)
);

AND2x2_ASAP7_75t_L g1086 ( 
.A(n_942),
.B(n_975),
.Y(n_1086)
);

AOI21x1_ASAP7_75t_L g1087 ( 
.A1(n_924),
.A2(n_832),
.B(n_823),
.Y(n_1087)
);

HB1xp67_ASAP7_75t_L g1088 ( 
.A(n_828),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_L g1089 ( 
.A1(n_876),
.A2(n_804),
.B(n_864),
.Y(n_1089)
);

OAI21x1_ASAP7_75t_L g1090 ( 
.A1(n_876),
.A2(n_804),
.B(n_864),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_936),
.B(n_954),
.Y(n_1091)
);

NAND2x1p5_ASAP7_75t_L g1092 ( 
.A(n_888),
.B(n_820),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_936),
.B(n_954),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_876),
.A2(n_804),
.B(n_864),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_942),
.B(n_975),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_899),
.A2(n_714),
.B(n_694),
.Y(n_1096)
);

BUFx2_ASAP7_75t_SL g1097 ( 
.A(n_934),
.Y(n_1097)
);

AND2x4_ASAP7_75t_L g1098 ( 
.A(n_983),
.B(n_939),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_935),
.Y(n_1099)
);

OAI21xp5_ASAP7_75t_SL g1100 ( 
.A1(n_946),
.A2(n_568),
.B(n_515),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_906),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_942),
.B(n_975),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_899),
.A2(n_714),
.B(n_694),
.Y(n_1103)
);

BUFx2_ASAP7_75t_L g1104 ( 
.A(n_890),
.Y(n_1104)
);

A2O1A1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_952),
.A2(n_963),
.B(n_967),
.C(n_953),
.Y(n_1105)
);

OAI21x1_ASAP7_75t_L g1106 ( 
.A1(n_876),
.A2(n_804),
.B(n_864),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_936),
.B(n_954),
.Y(n_1107)
);

OAI21x1_ASAP7_75t_L g1108 ( 
.A1(n_876),
.A2(n_804),
.B(n_864),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_936),
.B(n_954),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_899),
.A2(n_714),
.B(n_694),
.Y(n_1110)
);

AOI21xp33_ASAP7_75t_L g1111 ( 
.A1(n_950),
.A2(n_970),
.B(n_831),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_SL g1112 ( 
.A1(n_895),
.A2(n_952),
.B(n_923),
.Y(n_1112)
);

AOI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_882),
.A2(n_952),
.B1(n_887),
.B2(n_950),
.Y(n_1113)
);

AOI21xp5_ASAP7_75t_L g1114 ( 
.A1(n_899),
.A2(n_714),
.B(n_694),
.Y(n_1114)
);

AO21x1_ASAP7_75t_L g1115 ( 
.A1(n_952),
.A2(n_954),
.B(n_936),
.Y(n_1115)
);

BUFx2_ASAP7_75t_L g1116 ( 
.A(n_890),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_935),
.Y(n_1117)
);

OAI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_953),
.A2(n_967),
.B(n_963),
.Y(n_1118)
);

O2A1O1Ixp33_ASAP7_75t_SL g1119 ( 
.A1(n_953),
.A2(n_963),
.B(n_967),
.C(n_952),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_876),
.A2(n_804),
.B(n_864),
.Y(n_1120)
);

AOI221xp5_ASAP7_75t_L g1121 ( 
.A1(n_887),
.A2(n_907),
.B1(n_952),
.B2(n_591),
.C(n_706),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_876),
.A2(n_804),
.B(n_864),
.Y(n_1122)
);

OAI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_953),
.A2(n_967),
.B(n_963),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_876),
.A2(n_804),
.B(n_864),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_936),
.B(n_954),
.Y(n_1125)
);

NAND2x1p5_ASAP7_75t_L g1126 ( 
.A(n_888),
.B(n_820),
.Y(n_1126)
);

INVx2_ASAP7_75t_SL g1127 ( 
.A(n_828),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_899),
.A2(n_714),
.B(n_694),
.Y(n_1128)
);

INVxp67_ASAP7_75t_L g1129 ( 
.A(n_942),
.Y(n_1129)
);

OAI22xp5_ASAP7_75t_L g1130 ( 
.A1(n_936),
.A2(n_956),
.B1(n_959),
.B2(n_954),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_865),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_SL g1132 ( 
.A1(n_923),
.A2(n_952),
.B(n_730),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_876),
.A2(n_804),
.B(n_864),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_950),
.B(n_970),
.Y(n_1134)
);

OAI22xp5_ASAP7_75t_L g1135 ( 
.A1(n_936),
.A2(n_956),
.B1(n_959),
.B2(n_954),
.Y(n_1135)
);

INVx3_ASAP7_75t_L g1136 ( 
.A(n_820),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1130),
.B(n_1135),
.Y(n_1137)
);

OR2x6_ASAP7_75t_L g1138 ( 
.A(n_1097),
.B(n_1081),
.Y(n_1138)
);

INVxp67_ASAP7_75t_L g1139 ( 
.A(n_1088),
.Y(n_1139)
);

BUFx10_ASAP7_75t_L g1140 ( 
.A(n_1099),
.Y(n_1140)
);

HB1xp67_ASAP7_75t_L g1141 ( 
.A(n_1088),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_1017),
.A2(n_1022),
.B(n_1030),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1009),
.A2(n_1024),
.B(n_1029),
.Y(n_1143)
);

BUFx2_ASAP7_75t_SL g1144 ( 
.A(n_1056),
.Y(n_1144)
);

CKINVDCx20_ASAP7_75t_R g1145 ( 
.A(n_1045),
.Y(n_1145)
);

BUFx6f_ASAP7_75t_L g1146 ( 
.A(n_1049),
.Y(n_1146)
);

CKINVDCx20_ASAP7_75t_R g1147 ( 
.A(n_1045),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_1086),
.B(n_1095),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_994),
.B(n_996),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_1099),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1080),
.B(n_1083),
.Y(n_1151)
);

AO21x2_ASAP7_75t_L g1152 ( 
.A1(n_1027),
.A2(n_1123),
.B(n_1118),
.Y(n_1152)
);

INVx3_ASAP7_75t_L g1153 ( 
.A(n_1038),
.Y(n_1153)
);

AND2x4_ASAP7_75t_L g1154 ( 
.A(n_1013),
.B(n_1098),
.Y(n_1154)
);

O2A1O1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_1100),
.A2(n_1002),
.B(n_1004),
.C(n_1039),
.Y(n_1155)
);

BUFx3_ASAP7_75t_L g1156 ( 
.A(n_1056),
.Y(n_1156)
);

A2O1A1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_1121),
.A2(n_1134),
.B(n_997),
.C(n_1021),
.Y(n_1157)
);

BUFx6f_ASAP7_75t_L g1158 ( 
.A(n_1049),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1091),
.B(n_1093),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_1102),
.B(n_1008),
.Y(n_1160)
);

BUFx6f_ASAP7_75t_L g1161 ( 
.A(n_1049),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1107),
.B(n_1109),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1042),
.A2(n_1019),
.B(n_1059),
.Y(n_1163)
);

BUFx10_ASAP7_75t_L g1164 ( 
.A(n_1117),
.Y(n_1164)
);

AND2x4_ASAP7_75t_L g1165 ( 
.A(n_1013),
.B(n_1098),
.Y(n_1165)
);

AND2x2_ASAP7_75t_SL g1166 ( 
.A(n_995),
.B(n_1113),
.Y(n_1166)
);

INVx2_ASAP7_75t_SL g1167 ( 
.A(n_990),
.Y(n_1167)
);

AND2x2_ASAP7_75t_L g1168 ( 
.A(n_1034),
.B(n_1004),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1125),
.B(n_1002),
.Y(n_1169)
);

BUFx3_ASAP7_75t_L g1170 ( 
.A(n_1060),
.Y(n_1170)
);

INVxp67_ASAP7_75t_L g1171 ( 
.A(n_1026),
.Y(n_1171)
);

BUFx2_ASAP7_75t_SL g1172 ( 
.A(n_1060),
.Y(n_1172)
);

INVx3_ASAP7_75t_L g1173 ( 
.A(n_1038),
.Y(n_1173)
);

A2O1A1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_997),
.A2(n_1134),
.B(n_1111),
.C(n_1023),
.Y(n_1174)
);

OR2x6_ASAP7_75t_L g1175 ( 
.A(n_1132),
.B(n_1092),
.Y(n_1175)
);

AND2x4_ASAP7_75t_L g1176 ( 
.A(n_1013),
.B(n_1098),
.Y(n_1176)
);

A2O1A1Ixp33_ASAP7_75t_SL g1177 ( 
.A1(n_1006),
.A2(n_1076),
.B(n_1113),
.C(n_1018),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_1049),
.Y(n_1178)
);

INVx3_ASAP7_75t_SL g1179 ( 
.A(n_1117),
.Y(n_1179)
);

BUFx4f_ASAP7_75t_L g1180 ( 
.A(n_1041),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1131),
.Y(n_1181)
);

INVx3_ASAP7_75t_SL g1182 ( 
.A(n_1127),
.Y(n_1182)
);

AND2x2_ASAP7_75t_SL g1183 ( 
.A(n_995),
.B(n_1035),
.Y(n_1183)
);

AOI221x1_ASAP7_75t_L g1184 ( 
.A1(n_1105),
.A2(n_999),
.B1(n_1011),
.B2(n_1023),
.C(n_1000),
.Y(n_1184)
);

OA21x2_ASAP7_75t_L g1185 ( 
.A1(n_1012),
.A2(n_1025),
.B(n_1001),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1105),
.A2(n_999),
.B1(n_1005),
.B2(n_998),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1040),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1085),
.A2(n_1114),
.B(n_1096),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1129),
.B(n_1015),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_1129),
.B(n_1055),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1115),
.B(n_1082),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1033),
.B(n_1046),
.Y(n_1192)
);

HB1xp67_ASAP7_75t_L g1193 ( 
.A(n_1046),
.Y(n_1193)
);

NAND3xp33_ASAP7_75t_L g1194 ( 
.A(n_1000),
.B(n_1005),
.C(n_1082),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1044),
.B(n_1119),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1119),
.B(n_1112),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_SL g1197 ( 
.A1(n_1053),
.A2(n_1110),
.B(n_1128),
.Y(n_1197)
);

NOR2xp67_ASAP7_75t_SL g1198 ( 
.A(n_989),
.B(n_1104),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1048),
.Y(n_1199)
);

BUFx4f_ASAP7_75t_SL g1200 ( 
.A(n_992),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1043),
.B(n_1032),
.Y(n_1201)
);

CKINVDCx11_ASAP7_75t_R g1202 ( 
.A(n_1116),
.Y(n_1202)
);

INVx4_ASAP7_75t_L g1203 ( 
.A(n_1101),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1050),
.A2(n_1041),
.B1(n_1076),
.B2(n_1054),
.Y(n_1204)
);

AOI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1050),
.A2(n_1078),
.B1(n_1064),
.B2(n_1061),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1078),
.B(n_1036),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1035),
.B(n_1062),
.Y(n_1207)
);

O2A1O1Ixp5_ASAP7_75t_SL g1208 ( 
.A1(n_1065),
.A2(n_1074),
.B(n_1057),
.C(n_1069),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_1007),
.A2(n_1103),
.B1(n_1074),
.B2(n_1077),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1101),
.B(n_1066),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1101),
.B(n_1066),
.Y(n_1211)
);

INVx5_ASAP7_75t_L g1212 ( 
.A(n_1101),
.Y(n_1212)
);

OR2x6_ASAP7_75t_L g1213 ( 
.A(n_1092),
.B(n_1126),
.Y(n_1213)
);

INVx2_ASAP7_75t_SL g1214 ( 
.A(n_1007),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_992),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1047),
.B(n_1003),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1136),
.B(n_1031),
.Y(n_1217)
);

BUFx6f_ASAP7_75t_L g1218 ( 
.A(n_1126),
.Y(n_1218)
);

AND2x4_ASAP7_75t_L g1219 ( 
.A(n_1031),
.B(n_1058),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1028),
.A2(n_1063),
.B(n_1133),
.Y(n_1220)
);

BUFx2_ASAP7_75t_L g1221 ( 
.A(n_1007),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1072),
.B(n_1136),
.Y(n_1222)
);

AOI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1058),
.A2(n_1052),
.B1(n_1068),
.B2(n_1070),
.Y(n_1223)
);

AND2x4_ASAP7_75t_L g1224 ( 
.A(n_1037),
.B(n_1073),
.Y(n_1224)
);

OR2x2_ASAP7_75t_L g1225 ( 
.A(n_1051),
.B(n_1075),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_991),
.A2(n_1124),
.B(n_1106),
.Y(n_1226)
);

AOI221xp5_ASAP7_75t_L g1227 ( 
.A1(n_1071),
.A2(n_1051),
.B1(n_1087),
.B2(n_993),
.C(n_1122),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1051),
.B(n_1089),
.Y(n_1228)
);

OR2x6_ASAP7_75t_L g1229 ( 
.A(n_1067),
.B(n_1079),
.Y(n_1229)
);

BUFx2_ASAP7_75t_L g1230 ( 
.A(n_1051),
.Y(n_1230)
);

A2O1A1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1090),
.A2(n_1120),
.B(n_1094),
.C(n_1108),
.Y(n_1231)
);

A2O1A1Ixp33_ASAP7_75t_SL g1232 ( 
.A1(n_1010),
.A2(n_1014),
.B(n_1016),
.C(n_1020),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1130),
.B(n_936),
.Y(n_1233)
);

NAND3xp33_ASAP7_75t_L g1234 ( 
.A(n_1100),
.B(n_963),
.C(n_953),
.Y(n_1234)
);

NOR4xp25_ASAP7_75t_L g1235 ( 
.A(n_1121),
.B(n_953),
.C(n_967),
.D(n_963),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1130),
.B(n_936),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_1099),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1086),
.B(n_942),
.Y(n_1238)
);

INVx3_ASAP7_75t_L g1239 ( 
.A(n_1038),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1130),
.B(n_936),
.Y(n_1240)
);

AND2x4_ASAP7_75t_L g1241 ( 
.A(n_1013),
.B(n_1098),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1121),
.A2(n_950),
.B1(n_970),
.B2(n_958),
.Y(n_1242)
);

HB1xp67_ASAP7_75t_L g1243 ( 
.A(n_1088),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1084),
.Y(n_1244)
);

AND2x4_ASAP7_75t_L g1245 ( 
.A(n_1013),
.B(n_1098),
.Y(n_1245)
);

AOI221xp5_ASAP7_75t_L g1246 ( 
.A1(n_1100),
.A2(n_1121),
.B1(n_1004),
.B2(n_1002),
.C(n_706),
.Y(n_1246)
);

CKINVDCx6p67_ASAP7_75t_R g1247 ( 
.A(n_1045),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1084),
.Y(n_1248)
);

INVx3_ASAP7_75t_L g1249 ( 
.A(n_1038),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_994),
.A2(n_952),
.B1(n_954),
.B2(n_936),
.Y(n_1250)
);

AND2x2_ASAP7_75t_L g1251 ( 
.A(n_1086),
.B(n_942),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1130),
.B(n_936),
.Y(n_1252)
);

AND2x4_ASAP7_75t_L g1253 ( 
.A(n_1013),
.B(n_1098),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1121),
.A2(n_950),
.B1(n_970),
.B2(n_958),
.Y(n_1254)
);

OR2x2_ASAP7_75t_L g1255 ( 
.A(n_1008),
.B(n_1015),
.Y(n_1255)
);

BUFx6f_ASAP7_75t_SL g1256 ( 
.A(n_990),
.Y(n_1256)
);

INVx3_ASAP7_75t_SL g1257 ( 
.A(n_1099),
.Y(n_1257)
);

NAND2x1p5_ASAP7_75t_L g1258 ( 
.A(n_1038),
.B(n_888),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1084),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1009),
.A2(n_928),
.B(n_927),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1009),
.A2(n_928),
.B(n_927),
.Y(n_1261)
);

OAI21xp33_ASAP7_75t_L g1262 ( 
.A1(n_1100),
.A2(n_431),
.B(n_417),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_SL g1263 ( 
.A(n_1086),
.B(n_850),
.Y(n_1263)
);

NAND3xp33_ASAP7_75t_L g1264 ( 
.A(n_1100),
.B(n_963),
.C(n_953),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_SL g1265 ( 
.A1(n_1112),
.A2(n_1064),
.B(n_1036),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_L g1266 ( 
.A(n_1100),
.B(n_946),
.Y(n_1266)
);

AND2x4_ASAP7_75t_L g1267 ( 
.A(n_1013),
.B(n_1098),
.Y(n_1267)
);

AND2x4_ASAP7_75t_L g1268 ( 
.A(n_1013),
.B(n_1098),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1084),
.Y(n_1269)
);

BUFx4f_ASAP7_75t_L g1270 ( 
.A(n_1041),
.Y(n_1270)
);

HB1xp67_ASAP7_75t_L g1271 ( 
.A(n_1088),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_1099),
.Y(n_1272)
);

CKINVDCx8_ASAP7_75t_R g1273 ( 
.A(n_1097),
.Y(n_1273)
);

BUFx4_ASAP7_75t_SL g1274 ( 
.A(n_1056),
.Y(n_1274)
);

A2O1A1Ixp33_ASAP7_75t_SL g1275 ( 
.A1(n_1118),
.A2(n_632),
.B(n_642),
.C(n_481),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_L g1276 ( 
.A(n_1100),
.B(n_946),
.Y(n_1276)
);

AOI21xp33_ASAP7_75t_L g1277 ( 
.A1(n_1121),
.A2(n_970),
.B(n_950),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1009),
.A2(n_928),
.B(n_927),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1086),
.B(n_942),
.Y(n_1279)
);

OR2x2_ASAP7_75t_L g1280 ( 
.A(n_1152),
.B(n_1191),
.Y(n_1280)
);

OR2x2_ASAP7_75t_L g1281 ( 
.A(n_1152),
.B(n_1191),
.Y(n_1281)
);

BUFx10_ASAP7_75t_L g1282 ( 
.A(n_1256),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1166),
.B(n_1242),
.Y(n_1283)
);

CKINVDCx20_ASAP7_75t_R g1284 ( 
.A(n_1145),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1169),
.B(n_1149),
.Y(n_1285)
);

INVx8_ASAP7_75t_L g1286 ( 
.A(n_1212),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1181),
.Y(n_1287)
);

BUFx3_ASAP7_75t_L g1288 ( 
.A(n_1273),
.Y(n_1288)
);

INVx3_ASAP7_75t_L g1289 ( 
.A(n_1219),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1187),
.Y(n_1290)
);

AO21x1_ASAP7_75t_SL g1291 ( 
.A1(n_1206),
.A2(n_1137),
.B(n_1277),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1199),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1244),
.Y(n_1293)
);

AOI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1188),
.A2(n_1226),
.B(n_1260),
.Y(n_1294)
);

NOR2x1_ASAP7_75t_R g1295 ( 
.A(n_1150),
.B(n_1237),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1149),
.A2(n_1162),
.B1(n_1159),
.B2(n_1151),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1248),
.Y(n_1297)
);

BUFx2_ASAP7_75t_L g1298 ( 
.A(n_1141),
.Y(n_1298)
);

AOI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1246),
.A2(n_1277),
.B1(n_1254),
.B2(n_1276),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1259),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1269),
.Y(n_1301)
);

INVx3_ASAP7_75t_L g1302 ( 
.A(n_1219),
.Y(n_1302)
);

HB1xp67_ASAP7_75t_L g1303 ( 
.A(n_1243),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1189),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1190),
.Y(n_1305)
);

INVx3_ASAP7_75t_L g1306 ( 
.A(n_1175),
.Y(n_1306)
);

INVx1_ASAP7_75t_SL g1307 ( 
.A(n_1182),
.Y(n_1307)
);

AOI21x1_ASAP7_75t_L g1308 ( 
.A1(n_1261),
.A2(n_1278),
.B(n_1216),
.Y(n_1308)
);

BUFx10_ASAP7_75t_L g1309 ( 
.A(n_1256),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1271),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1255),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1142),
.A2(n_1220),
.B(n_1163),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1160),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1210),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1157),
.B(n_1174),
.Y(n_1315)
);

CKINVDCx11_ASAP7_75t_R g1316 ( 
.A(n_1179),
.Y(n_1316)
);

BUFx8_ASAP7_75t_L g1317 ( 
.A(n_1221),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1266),
.A2(n_1234),
.B1(n_1264),
.B2(n_1194),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1211),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1148),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1192),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1168),
.Y(n_1322)
);

OA21x2_ASAP7_75t_L g1323 ( 
.A1(n_1143),
.A2(n_1227),
.B(n_1231),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1196),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1228),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1196),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1201),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1201),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1265),
.Y(n_1329)
);

AOI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1183),
.A2(n_1262),
.B1(n_1204),
.B2(n_1251),
.Y(n_1330)
);

BUFx2_ASAP7_75t_L g1331 ( 
.A(n_1167),
.Y(n_1331)
);

OAI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1169),
.A2(n_1159),
.B1(n_1151),
.B2(n_1162),
.Y(n_1332)
);

AOI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1238),
.A2(n_1279),
.B1(n_1207),
.B2(n_1234),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1263),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1264),
.A2(n_1194),
.B1(n_1186),
.B2(n_1250),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1216),
.A2(n_1208),
.B(n_1223),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1222),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1155),
.B(n_1250),
.Y(n_1338)
);

INVx3_ASAP7_75t_L g1339 ( 
.A(n_1175),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1225),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1197),
.A2(n_1185),
.B(n_1186),
.Y(n_1341)
);

HB1xp67_ASAP7_75t_L g1342 ( 
.A(n_1171),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1230),
.Y(n_1343)
);

INVx11_ASAP7_75t_L g1344 ( 
.A(n_1274),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1217),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1235),
.B(n_1240),
.Y(n_1346)
);

CKINVDCx11_ASAP7_75t_R g1347 ( 
.A(n_1257),
.Y(n_1347)
);

HB1xp67_ASAP7_75t_L g1348 ( 
.A(n_1139),
.Y(n_1348)
);

BUFx2_ASAP7_75t_R g1349 ( 
.A(n_1272),
.Y(n_1349)
);

INVx1_ASAP7_75t_SL g1350 ( 
.A(n_1202),
.Y(n_1350)
);

INVx1_ASAP7_75t_SL g1351 ( 
.A(n_1144),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1235),
.B(n_1240),
.Y(n_1352)
);

BUFx2_ASAP7_75t_R g1353 ( 
.A(n_1215),
.Y(n_1353)
);

OAI22xp33_ASAP7_75t_SL g1354 ( 
.A1(n_1233),
.A2(n_1236),
.B1(n_1252),
.B2(n_1137),
.Y(n_1354)
);

BUFx3_ASAP7_75t_L g1355 ( 
.A(n_1154),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1233),
.A2(n_1206),
.B1(n_1270),
.B2(n_1180),
.Y(n_1356)
);

BUFx6f_ASAP7_75t_L g1357 ( 
.A(n_1146),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_1147),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1180),
.A2(n_1270),
.B1(n_1193),
.B2(n_1195),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1158),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1161),
.Y(n_1361)
);

AOI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1198),
.A2(n_1245),
.B1(n_1268),
.B2(n_1267),
.Y(n_1362)
);

OAI21x1_ASAP7_75t_L g1363 ( 
.A1(n_1185),
.A2(n_1195),
.B(n_1209),
.Y(n_1363)
);

OR2x6_ASAP7_75t_L g1364 ( 
.A(n_1138),
.B(n_1229),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1205),
.A2(n_1138),
.B1(n_1268),
.B2(n_1267),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1178),
.Y(n_1366)
);

CKINVDCx11_ASAP7_75t_R g1367 ( 
.A(n_1140),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_SL g1368 ( 
.A1(n_1203),
.A2(n_1214),
.B(n_1138),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1184),
.A2(n_1258),
.B(n_1232),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_1247),
.Y(n_1370)
);

OA21x2_ASAP7_75t_L g1371 ( 
.A1(n_1224),
.A2(n_1177),
.B(n_1275),
.Y(n_1371)
);

INVx2_ASAP7_75t_SL g1372 ( 
.A(n_1165),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1172),
.A2(n_1253),
.B1(n_1245),
.B2(n_1176),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1178),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1178),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1165),
.Y(n_1376)
);

HB1xp67_ASAP7_75t_L g1377 ( 
.A(n_1176),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1241),
.Y(n_1378)
);

CKINVDCx11_ASAP7_75t_R g1379 ( 
.A(n_1140),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1241),
.Y(n_1380)
);

BUFx4f_ASAP7_75t_SL g1381 ( 
.A(n_1156),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1229),
.Y(n_1382)
);

INVx4_ASAP7_75t_L g1383 ( 
.A(n_1213),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1253),
.Y(n_1384)
);

OAI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1229),
.A2(n_1224),
.B(n_1213),
.Y(n_1385)
);

BUFx6f_ASAP7_75t_L g1386 ( 
.A(n_1218),
.Y(n_1386)
);

AOI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1170),
.A2(n_1200),
.B1(n_1164),
.B2(n_1218),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_SL g1388 ( 
.A1(n_1153),
.A2(n_1173),
.B1(n_1239),
.B2(n_1249),
.Y(n_1388)
);

CKINVDCx11_ASAP7_75t_R g1389 ( 
.A(n_1164),
.Y(n_1389)
);

BUFx12f_ASAP7_75t_L g1390 ( 
.A(n_1215),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1169),
.B(n_1002),
.Y(n_1391)
);

OA21x2_ASAP7_75t_L g1392 ( 
.A1(n_1143),
.A2(n_1163),
.B(n_1188),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1296),
.B(n_1285),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1346),
.B(n_1352),
.Y(n_1394)
);

INVx3_ASAP7_75t_L g1395 ( 
.A(n_1364),
.Y(n_1395)
);

INVxp67_ASAP7_75t_SL g1396 ( 
.A(n_1303),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1325),
.Y(n_1397)
);

BUFx6f_ASAP7_75t_L g1398 ( 
.A(n_1364),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1346),
.B(n_1352),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1298),
.Y(n_1400)
);

NAND2x1p5_ASAP7_75t_L g1401 ( 
.A(n_1306),
.B(n_1339),
.Y(n_1401)
);

OAI21x1_ASAP7_75t_L g1402 ( 
.A1(n_1312),
.A2(n_1294),
.B(n_1308),
.Y(n_1402)
);

AND2x2_ASAP7_75t_L g1403 ( 
.A(n_1340),
.B(n_1283),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1280),
.B(n_1281),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1280),
.Y(n_1405)
);

BUFx3_ASAP7_75t_L g1406 ( 
.A(n_1368),
.Y(n_1406)
);

OR2x2_ASAP7_75t_L g1407 ( 
.A(n_1281),
.B(n_1343),
.Y(n_1407)
);

INVx3_ASAP7_75t_L g1408 ( 
.A(n_1364),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1382),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1382),
.Y(n_1410)
);

HB1xp67_ASAP7_75t_L g1411 ( 
.A(n_1298),
.Y(n_1411)
);

OAI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1336),
.A2(n_1341),
.B(n_1363),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1391),
.B(n_1332),
.Y(n_1413)
);

OR2x6_ASAP7_75t_L g1414 ( 
.A(n_1306),
.B(n_1339),
.Y(n_1414)
);

BUFx2_ASAP7_75t_L g1415 ( 
.A(n_1385),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1337),
.Y(n_1416)
);

OA21x2_ASAP7_75t_L g1417 ( 
.A1(n_1341),
.A2(n_1338),
.B(n_1369),
.Y(n_1417)
);

BUFx4f_ASAP7_75t_L g1418 ( 
.A(n_1286),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1324),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1392),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1326),
.Y(n_1421)
);

OAI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1392),
.A2(n_1323),
.B(n_1329),
.Y(n_1422)
);

AOI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1354),
.A2(n_1315),
.B(n_1335),
.Y(n_1423)
);

AO21x2_ASAP7_75t_L g1424 ( 
.A1(n_1327),
.A2(n_1328),
.B(n_1334),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_SL g1425 ( 
.A1(n_1318),
.A2(n_1383),
.B(n_1365),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1287),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1283),
.B(n_1318),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1371),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1311),
.B(n_1299),
.Y(n_1429)
);

AO21x2_ASAP7_75t_L g1430 ( 
.A1(n_1333),
.A2(n_1300),
.B(n_1297),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1290),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1299),
.B(n_1304),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1371),
.Y(n_1433)
);

AO21x2_ASAP7_75t_L g1434 ( 
.A1(n_1315),
.A2(n_1293),
.B(n_1292),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1301),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_1316),
.Y(n_1436)
);

OAI21xp5_ASAP7_75t_L g1437 ( 
.A1(n_1335),
.A2(n_1356),
.B(n_1330),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1322),
.B(n_1313),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1310),
.B(n_1320),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1291),
.B(n_1314),
.Y(n_1440)
);

OR2x2_ASAP7_75t_L g1441 ( 
.A(n_1356),
.B(n_1305),
.Y(n_1441)
);

BUFx3_ASAP7_75t_L g1442 ( 
.A(n_1286),
.Y(n_1442)
);

BUFx2_ASAP7_75t_L g1443 ( 
.A(n_1383),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1319),
.B(n_1345),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1321),
.B(n_1342),
.Y(n_1445)
);

CKINVDCx6p67_ASAP7_75t_R g1446 ( 
.A(n_1316),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1289),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1289),
.B(n_1302),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1289),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1302),
.Y(n_1450)
);

INVx1_ASAP7_75t_SL g1451 ( 
.A(n_1331),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1302),
.B(n_1359),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_L g1453 ( 
.A(n_1348),
.Y(n_1453)
);

OR2x2_ASAP7_75t_L g1454 ( 
.A(n_1359),
.B(n_1351),
.Y(n_1454)
);

INVxp67_ASAP7_75t_L g1455 ( 
.A(n_1307),
.Y(n_1455)
);

AND2x4_ASAP7_75t_L g1456 ( 
.A(n_1376),
.B(n_1378),
.Y(n_1456)
);

AO21x2_ASAP7_75t_L g1457 ( 
.A1(n_1360),
.A2(n_1366),
.B(n_1361),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1374),
.Y(n_1458)
);

OR2x2_ASAP7_75t_L g1459 ( 
.A(n_1404),
.B(n_1375),
.Y(n_1459)
);

AOI221xp5_ASAP7_75t_L g1460 ( 
.A1(n_1437),
.A2(n_1373),
.B1(n_1384),
.B2(n_1350),
.C(n_1288),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1404),
.B(n_1380),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1393),
.B(n_1388),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1394),
.B(n_1386),
.Y(n_1463)
);

INVx3_ASAP7_75t_L g1464 ( 
.A(n_1398),
.Y(n_1464)
);

AND2x2_ASAP7_75t_L g1465 ( 
.A(n_1394),
.B(n_1386),
.Y(n_1465)
);

OR2x2_ASAP7_75t_L g1466 ( 
.A(n_1434),
.B(n_1377),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1405),
.Y(n_1467)
);

INVx3_ASAP7_75t_L g1468 ( 
.A(n_1398),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1399),
.B(n_1372),
.Y(n_1469)
);

HB1xp67_ASAP7_75t_L g1470 ( 
.A(n_1434),
.Y(n_1470)
);

AND2x4_ASAP7_75t_L g1471 ( 
.A(n_1395),
.B(n_1355),
.Y(n_1471)
);

INVx1_ASAP7_75t_SL g1472 ( 
.A(n_1400),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1417),
.B(n_1357),
.Y(n_1473)
);

BUFx2_ASAP7_75t_L g1474 ( 
.A(n_1414),
.Y(n_1474)
);

AND2x4_ASAP7_75t_L g1475 ( 
.A(n_1395),
.B(n_1355),
.Y(n_1475)
);

INVxp67_ASAP7_75t_L g1476 ( 
.A(n_1424),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1405),
.B(n_1357),
.Y(n_1477)
);

AOI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1423),
.A2(n_1420),
.B(n_1422),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1417),
.B(n_1362),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1397),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_L g1481 ( 
.A(n_1424),
.Y(n_1481)
);

NAND4xp25_ASAP7_75t_L g1482 ( 
.A(n_1413),
.B(n_1429),
.C(n_1432),
.D(n_1445),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1424),
.Y(n_1483)
);

OR2x2_ASAP7_75t_L g1484 ( 
.A(n_1407),
.B(n_1387),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1420),
.Y(n_1485)
);

BUFx2_ASAP7_75t_L g1486 ( 
.A(n_1414),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1428),
.B(n_1433),
.Y(n_1487)
);

BUFx3_ASAP7_75t_L g1488 ( 
.A(n_1398),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1407),
.Y(n_1489)
);

INVxp67_ASAP7_75t_L g1490 ( 
.A(n_1457),
.Y(n_1490)
);

OR2x2_ASAP7_75t_L g1491 ( 
.A(n_1430),
.B(n_1288),
.Y(n_1491)
);

NAND3xp33_ASAP7_75t_L g1492 ( 
.A(n_1482),
.B(n_1440),
.C(n_1454),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1472),
.B(n_1396),
.Y(n_1493)
);

HB1xp67_ASAP7_75t_L g1494 ( 
.A(n_1489),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1463),
.B(n_1415),
.Y(n_1495)
);

OAI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1482),
.A2(n_1454),
.B(n_1455),
.Y(n_1496)
);

OA21x2_ASAP7_75t_L g1497 ( 
.A1(n_1476),
.A2(n_1412),
.B(n_1402),
.Y(n_1497)
);

OAI21xp5_ASAP7_75t_SL g1498 ( 
.A1(n_1460),
.A2(n_1427),
.B(n_1452),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1463),
.B(n_1403),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1472),
.B(n_1411),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1465),
.B(n_1403),
.Y(n_1501)
);

OAI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1462),
.A2(n_1441),
.B1(n_1446),
.B2(n_1427),
.Y(n_1502)
);

NAND3xp33_ASAP7_75t_L g1503 ( 
.A(n_1491),
.B(n_1440),
.C(n_1441),
.Y(n_1503)
);

NAND3xp33_ASAP7_75t_L g1504 ( 
.A(n_1491),
.B(n_1452),
.C(n_1438),
.Y(n_1504)
);

NAND3xp33_ASAP7_75t_L g1505 ( 
.A(n_1491),
.B(n_1409),
.C(n_1410),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1480),
.Y(n_1506)
);

OAI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1462),
.A2(n_1460),
.B1(n_1484),
.B2(n_1446),
.Y(n_1507)
);

OAI21xp33_ASAP7_75t_L g1508 ( 
.A1(n_1484),
.A2(n_1453),
.B(n_1444),
.Y(n_1508)
);

NAND3xp33_ASAP7_75t_L g1509 ( 
.A(n_1478),
.B(n_1409),
.C(n_1410),
.Y(n_1509)
);

NAND3xp33_ASAP7_75t_L g1510 ( 
.A(n_1478),
.B(n_1416),
.C(n_1421),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1461),
.B(n_1416),
.Y(n_1511)
);

OAI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1484),
.A2(n_1451),
.B1(n_1418),
.B2(n_1370),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1461),
.B(n_1430),
.Y(n_1513)
);

OAI21xp33_ASAP7_75t_L g1514 ( 
.A1(n_1479),
.A2(n_1444),
.B(n_1439),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1471),
.A2(n_1425),
.B1(n_1398),
.B2(n_1408),
.Y(n_1515)
);

AOI21xp33_ASAP7_75t_L g1516 ( 
.A1(n_1466),
.A2(n_1430),
.B(n_1425),
.Y(n_1516)
);

NOR2xp33_ASAP7_75t_L g1517 ( 
.A(n_1461),
.B(n_1381),
.Y(n_1517)
);

NAND3xp33_ASAP7_75t_L g1518 ( 
.A(n_1490),
.B(n_1419),
.C(n_1421),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1469),
.B(n_1479),
.Y(n_1519)
);

NAND3xp33_ASAP7_75t_L g1520 ( 
.A(n_1490),
.B(n_1419),
.C(n_1447),
.Y(n_1520)
);

AOI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1469),
.A2(n_1456),
.B1(n_1398),
.B2(n_1448),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_L g1522 ( 
.A(n_1469),
.B(n_1436),
.Y(n_1522)
);

OAI21xp5_ASAP7_75t_SL g1523 ( 
.A1(n_1479),
.A2(n_1408),
.B(n_1474),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1474),
.B(n_1408),
.Y(n_1524)
);

OAI221xp5_ASAP7_75t_L g1525 ( 
.A1(n_1466),
.A2(n_1406),
.B1(n_1439),
.B2(n_1401),
.C(n_1358),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1459),
.B(n_1477),
.Y(n_1526)
);

OA211x2_ASAP7_75t_L g1527 ( 
.A1(n_1476),
.A2(n_1418),
.B(n_1442),
.C(n_1406),
.Y(n_1527)
);

NAND3xp33_ASAP7_75t_L g1528 ( 
.A(n_1481),
.B(n_1447),
.C(n_1449),
.Y(n_1528)
);

NAND3xp33_ASAP7_75t_L g1529 ( 
.A(n_1481),
.B(n_1449),
.C(n_1450),
.Y(n_1529)
);

NAND3xp33_ASAP7_75t_L g1530 ( 
.A(n_1483),
.B(n_1449),
.C(n_1450),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1519),
.B(n_1473),
.Y(n_1531)
);

NOR2xp33_ASAP7_75t_L g1532 ( 
.A(n_1492),
.B(n_1525),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1519),
.B(n_1473),
.Y(n_1533)
);

BUFx2_ASAP7_75t_L g1534 ( 
.A(n_1524),
.Y(n_1534)
);

AOI33xp33_ASAP7_75t_L g1535 ( 
.A1(n_1515),
.A2(n_1426),
.A3(n_1435),
.B1(n_1431),
.B2(n_1467),
.B3(n_1458),
.Y(n_1535)
);

OR2x2_ASAP7_75t_L g1536 ( 
.A(n_1513),
.B(n_1470),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1506),
.Y(n_1537)
);

AND2x4_ASAP7_75t_L g1538 ( 
.A(n_1506),
.B(n_1487),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1494),
.B(n_1526),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1497),
.Y(n_1540)
);

HB1xp67_ASAP7_75t_L g1541 ( 
.A(n_1505),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1497),
.Y(n_1542)
);

INVx2_ASAP7_75t_SL g1543 ( 
.A(n_1497),
.Y(n_1543)
);

INVx1_ASAP7_75t_SL g1544 ( 
.A(n_1493),
.Y(n_1544)
);

HB1xp67_ASAP7_75t_L g1545 ( 
.A(n_1520),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1504),
.B(n_1470),
.Y(n_1546)
);

BUFx3_ASAP7_75t_L g1547 ( 
.A(n_1509),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1514),
.B(n_1467),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1503),
.B(n_1483),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1511),
.Y(n_1550)
);

AOI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1498),
.A2(n_1456),
.B1(n_1475),
.B2(n_1471),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1518),
.Y(n_1552)
);

INVx3_ASAP7_75t_L g1553 ( 
.A(n_1499),
.Y(n_1553)
);

AND3x1_ASAP7_75t_L g1554 ( 
.A(n_1522),
.B(n_1468),
.C(n_1464),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1530),
.Y(n_1555)
);

AND2x4_ASAP7_75t_L g1556 ( 
.A(n_1521),
.B(n_1485),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1531),
.B(n_1499),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1540),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1531),
.B(n_1501),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1537),
.Y(n_1560)
);

INVx3_ASAP7_75t_L g1561 ( 
.A(n_1538),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1540),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1540),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1531),
.B(n_1501),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1533),
.B(n_1495),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1533),
.B(n_1495),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1537),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1533),
.B(n_1523),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1537),
.Y(n_1569)
);

AND2x4_ASAP7_75t_L g1570 ( 
.A(n_1556),
.B(n_1486),
.Y(n_1570)
);

INVx3_ASAP7_75t_R g1571 ( 
.A(n_1549),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1540),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1542),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1553),
.B(n_1514),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1542),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1552),
.B(n_1508),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1538),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1538),
.Y(n_1578)
);

HB1xp67_ASAP7_75t_L g1579 ( 
.A(n_1541),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1552),
.B(n_1508),
.Y(n_1580)
);

AOI21xp33_ASAP7_75t_L g1581 ( 
.A1(n_1532),
.A2(n_1507),
.B(n_1496),
.Y(n_1581)
);

INVxp67_ASAP7_75t_L g1582 ( 
.A(n_1545),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1546),
.B(n_1510),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1542),
.Y(n_1584)
);

NOR5xp2_ASAP7_75t_L g1585 ( 
.A(n_1545),
.B(n_1528),
.C(n_1529),
.D(n_1516),
.E(n_1527),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1552),
.B(n_1500),
.Y(n_1586)
);

INVxp67_ASAP7_75t_L g1587 ( 
.A(n_1541),
.Y(n_1587)
);

AND3x2_ASAP7_75t_L g1588 ( 
.A(n_1532),
.B(n_1517),
.C(n_1443),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1569),
.Y(n_1589)
);

NAND2x1_ASAP7_75t_L g1590 ( 
.A(n_1574),
.B(n_1534),
.Y(n_1590)
);

NOR2xp67_ASAP7_75t_L g1591 ( 
.A(n_1582),
.B(n_1553),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1583),
.B(n_1576),
.Y(n_1592)
);

INVx3_ASAP7_75t_L g1593 ( 
.A(n_1561),
.Y(n_1593)
);

OAI21xp33_ASAP7_75t_L g1594 ( 
.A1(n_1581),
.A2(n_1551),
.B(n_1547),
.Y(n_1594)
);

AND2x2_ASAP7_75t_SL g1595 ( 
.A(n_1585),
.B(n_1554),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1583),
.B(n_1555),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1569),
.Y(n_1597)
);

OAI322xp33_ASAP7_75t_L g1598 ( 
.A1(n_1582),
.A2(n_1546),
.A3(n_1549),
.B1(n_1555),
.B2(n_1536),
.C1(n_1548),
.C2(n_1544),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1586),
.B(n_1544),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1586),
.B(n_1547),
.Y(n_1600)
);

NAND2x1p5_ASAP7_75t_L g1601 ( 
.A(n_1583),
.B(n_1554),
.Y(n_1601)
);

AND2x4_ASAP7_75t_L g1602 ( 
.A(n_1568),
.B(n_1547),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1558),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1568),
.B(n_1534),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1560),
.Y(n_1605)
);

BUFx2_ASAP7_75t_L g1606 ( 
.A(n_1579),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1576),
.B(n_1539),
.Y(n_1607)
);

NOR2x1_ASAP7_75t_L g1608 ( 
.A(n_1580),
.B(n_1547),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1558),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1560),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1560),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1581),
.B(n_1550),
.Y(n_1612)
);

OAI21xp5_ASAP7_75t_L g1613 ( 
.A1(n_1587),
.A2(n_1555),
.B(n_1551),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1567),
.Y(n_1614)
);

NOR2x1p5_ASAP7_75t_SL g1615 ( 
.A(n_1558),
.B(n_1542),
.Y(n_1615)
);

AND2x4_ASAP7_75t_L g1616 ( 
.A(n_1568),
.B(n_1551),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1580),
.B(n_1550),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1558),
.Y(n_1618)
);

AND2x4_ASAP7_75t_L g1619 ( 
.A(n_1570),
.B(n_1556),
.Y(n_1619)
);

INVx2_ASAP7_75t_L g1620 ( 
.A(n_1562),
.Y(n_1620)
);

INVx1_ASAP7_75t_SL g1621 ( 
.A(n_1588),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1570),
.B(n_1556),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1579),
.B(n_1536),
.Y(n_1623)
);

NAND2x2_ASAP7_75t_L g1624 ( 
.A(n_1588),
.B(n_1488),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1587),
.B(n_1550),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1562),
.Y(n_1626)
);

BUFx2_ASAP7_75t_L g1627 ( 
.A(n_1565),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1567),
.Y(n_1628)
);

AND2x4_ASAP7_75t_L g1629 ( 
.A(n_1570),
.B(n_1556),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1567),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1557),
.B(n_1534),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1608),
.B(n_1557),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1604),
.B(n_1574),
.Y(n_1633)
);

NAND2x1p5_ASAP7_75t_L g1634 ( 
.A(n_1595),
.B(n_1585),
.Y(n_1634)
);

INVx1_ASAP7_75t_SL g1635 ( 
.A(n_1621),
.Y(n_1635)
);

INVxp67_ASAP7_75t_SL g1636 ( 
.A(n_1601),
.Y(n_1636)
);

NOR2x1_ASAP7_75t_L g1637 ( 
.A(n_1606),
.B(n_1284),
.Y(n_1637)
);

AOI22xp33_ASAP7_75t_L g1638 ( 
.A1(n_1594),
.A2(n_1502),
.B1(n_1570),
.B2(n_1512),
.Y(n_1638)
);

AOI22xp33_ASAP7_75t_L g1639 ( 
.A1(n_1595),
.A2(n_1570),
.B1(n_1574),
.B2(n_1475),
.Y(n_1639)
);

OR2x2_ASAP7_75t_L g1640 ( 
.A(n_1592),
.B(n_1596),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1605),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1612),
.B(n_1557),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1600),
.B(n_1592),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1610),
.Y(n_1644)
);

OR2x6_ASAP7_75t_L g1645 ( 
.A(n_1590),
.B(n_1286),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1602),
.B(n_1559),
.Y(n_1646)
);

INVxp67_ASAP7_75t_L g1647 ( 
.A(n_1602),
.Y(n_1647)
);

HB1xp67_ASAP7_75t_L g1648 ( 
.A(n_1604),
.Y(n_1648)
);

INVx1_ASAP7_75t_SL g1649 ( 
.A(n_1602),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1611),
.Y(n_1650)
);

AO21x2_ASAP7_75t_L g1651 ( 
.A1(n_1591),
.A2(n_1571),
.B(n_1563),
.Y(n_1651)
);

NAND2xp5_ASAP7_75t_L g1652 ( 
.A(n_1607),
.B(n_1559),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1616),
.B(n_1559),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1616),
.B(n_1564),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1627),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1596),
.B(n_1549),
.Y(n_1656)
);

INVxp67_ASAP7_75t_L g1657 ( 
.A(n_1625),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1614),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1628),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1616),
.B(n_1564),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1630),
.Y(n_1661)
);

OR2x6_ASAP7_75t_L g1662 ( 
.A(n_1613),
.B(n_1571),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1589),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1601),
.B(n_1564),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1623),
.B(n_1536),
.Y(n_1665)
);

AOI22xp33_ASAP7_75t_L g1666 ( 
.A1(n_1624),
.A2(n_1570),
.B1(n_1471),
.B2(n_1475),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1631),
.B(n_1565),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1635),
.B(n_1617),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1653),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1647),
.B(n_1599),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1653),
.Y(n_1671)
);

AOI21xp33_ASAP7_75t_SL g1672 ( 
.A1(n_1634),
.A2(n_1370),
.B(n_1358),
.Y(n_1672)
);

OAI22xp5_ASAP7_75t_L g1673 ( 
.A1(n_1634),
.A2(n_1662),
.B1(n_1637),
.B2(n_1638),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1649),
.B(n_1648),
.Y(n_1674)
);

OAI21xp5_ASAP7_75t_L g1675 ( 
.A1(n_1634),
.A2(n_1623),
.B(n_1571),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1657),
.B(n_1655),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1643),
.B(n_1347),
.Y(n_1677)
);

INVxp67_ASAP7_75t_L g1678 ( 
.A(n_1640),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1655),
.B(n_1631),
.Y(n_1679)
);

OAI21xp5_ASAP7_75t_L g1680 ( 
.A1(n_1662),
.A2(n_1546),
.B(n_1597),
.Y(n_1680)
);

OAI221xp5_ASAP7_75t_L g1681 ( 
.A1(n_1662),
.A2(n_1624),
.B1(n_1598),
.B2(n_1593),
.C(n_1561),
.Y(n_1681)
);

OAI32xp33_ASAP7_75t_L g1682 ( 
.A1(n_1632),
.A2(n_1593),
.A3(n_1561),
.B1(n_1577),
.B2(n_1578),
.Y(n_1682)
);

OAI21xp33_ASAP7_75t_L g1683 ( 
.A1(n_1662),
.A2(n_1615),
.B(n_1535),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1654),
.B(n_1660),
.Y(n_1684)
);

O2A1O1Ixp33_ASAP7_75t_SL g1685 ( 
.A1(n_1636),
.A2(n_1284),
.B(n_1593),
.C(n_1577),
.Y(n_1685)
);

OAI21xp33_ASAP7_75t_L g1686 ( 
.A1(n_1639),
.A2(n_1535),
.B(n_1619),
.Y(n_1686)
);

OR2x6_ASAP7_75t_L g1687 ( 
.A(n_1640),
.B(n_1390),
.Y(n_1687)
);

O2A1O1Ixp33_ASAP7_75t_L g1688 ( 
.A1(n_1651),
.A2(n_1543),
.B(n_1629),
.C(n_1619),
.Y(n_1688)
);

AOI221xp5_ASAP7_75t_L g1689 ( 
.A1(n_1646),
.A2(n_1629),
.B1(n_1622),
.B2(n_1619),
.C(n_1543),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1654),
.B(n_1565),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1641),
.Y(n_1691)
);

OAI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1664),
.A2(n_1629),
.B(n_1622),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1641),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1684),
.B(n_1660),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1678),
.B(n_1663),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1691),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1693),
.Y(n_1697)
);

OR2x2_ASAP7_75t_L g1698 ( 
.A(n_1674),
.B(n_1642),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1669),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1671),
.B(n_1633),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1673),
.B(n_1668),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1679),
.B(n_1652),
.Y(n_1702)
);

INVx2_ASAP7_75t_SL g1703 ( 
.A(n_1687),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1676),
.B(n_1633),
.Y(n_1704)
);

INVx2_ASAP7_75t_SL g1705 ( 
.A(n_1687),
.Y(n_1705)
);

AND2x4_ASAP7_75t_L g1706 ( 
.A(n_1687),
.B(n_1664),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1670),
.B(n_1677),
.Y(n_1707)
);

NOR2x1_ASAP7_75t_L g1708 ( 
.A(n_1675),
.B(n_1651),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1692),
.B(n_1667),
.Y(n_1709)
);

OR2x2_ASAP7_75t_L g1710 ( 
.A(n_1690),
.B(n_1667),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1692),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1686),
.B(n_1663),
.Y(n_1712)
);

OR2x2_ASAP7_75t_L g1713 ( 
.A(n_1675),
.B(n_1665),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1672),
.B(n_1644),
.Y(n_1714)
);

AOI21xp33_ASAP7_75t_L g1715 ( 
.A1(n_1708),
.A2(n_1713),
.B(n_1705),
.Y(n_1715)
);

AOI21xp5_ASAP7_75t_L g1716 ( 
.A1(n_1701),
.A2(n_1680),
.B(n_1683),
.Y(n_1716)
);

AOI211xp5_ASAP7_75t_L g1717 ( 
.A1(n_1712),
.A2(n_1681),
.B(n_1685),
.C(n_1688),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1699),
.Y(n_1718)
);

OAI22xp5_ASAP7_75t_L g1719 ( 
.A1(n_1712),
.A2(n_1666),
.B1(n_1645),
.B2(n_1689),
.Y(n_1719)
);

O2A1O1Ixp33_ASAP7_75t_L g1720 ( 
.A1(n_1714),
.A2(n_1651),
.B(n_1682),
.C(n_1656),
.Y(n_1720)
);

NOR3xp33_ASAP7_75t_SL g1721 ( 
.A(n_1707),
.B(n_1711),
.C(n_1714),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1700),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_SL g1723 ( 
.A(n_1706),
.B(n_1656),
.Y(n_1723)
);

AOI222xp33_ASAP7_75t_L g1724 ( 
.A1(n_1695),
.A2(n_1658),
.B1(n_1650),
.B2(n_1644),
.C1(n_1659),
.C2(n_1661),
.Y(n_1724)
);

AOI21xp5_ASAP7_75t_L g1725 ( 
.A1(n_1695),
.A2(n_1645),
.B(n_1650),
.Y(n_1725)
);

NOR3xp33_ASAP7_75t_L g1726 ( 
.A(n_1715),
.B(n_1703),
.C(n_1704),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1723),
.B(n_1706),
.Y(n_1727)
);

AOI211x1_ASAP7_75t_L g1728 ( 
.A1(n_1716),
.A2(n_1709),
.B(n_1694),
.C(n_1697),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1721),
.B(n_1698),
.Y(n_1729)
);

NOR2x1_ASAP7_75t_L g1730 ( 
.A(n_1718),
.B(n_1696),
.Y(n_1730)
);

NOR3x1_ASAP7_75t_L g1731 ( 
.A(n_1722),
.B(n_1702),
.C(n_1710),
.Y(n_1731)
);

NAND3xp33_ASAP7_75t_L g1732 ( 
.A(n_1720),
.B(n_1659),
.C(n_1658),
.Y(n_1732)
);

AOI22xp5_ASAP7_75t_L g1733 ( 
.A1(n_1717),
.A2(n_1645),
.B1(n_1661),
.B2(n_1622),
.Y(n_1733)
);

NOR2xp67_ASAP7_75t_L g1734 ( 
.A(n_1725),
.B(n_1390),
.Y(n_1734)
);

NAND4xp25_ASAP7_75t_L g1735 ( 
.A(n_1724),
.B(n_1665),
.C(n_1527),
.D(n_1620),
.Y(n_1735)
);

INVxp67_ASAP7_75t_L g1736 ( 
.A(n_1727),
.Y(n_1736)
);

NOR2x1_ASAP7_75t_L g1737 ( 
.A(n_1730),
.B(n_1719),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1728),
.B(n_1566),
.Y(n_1738)
);

NOR3xp33_ASAP7_75t_L g1739 ( 
.A(n_1726),
.B(n_1729),
.C(n_1734),
.Y(n_1739)
);

NAND4xp75_ASAP7_75t_L g1740 ( 
.A(n_1731),
.B(n_1347),
.C(n_1389),
.D(n_1379),
.Y(n_1740)
);

AOI22xp33_ASAP7_75t_SL g1741 ( 
.A1(n_1738),
.A2(n_1732),
.B1(n_1645),
.B2(n_1733),
.Y(n_1741)
);

AOI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1739),
.A2(n_1735),
.B1(n_1379),
.B2(n_1389),
.Y(n_1742)
);

INVx3_ASAP7_75t_L g1743 ( 
.A(n_1740),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1736),
.Y(n_1744)
);

INVxp67_ASAP7_75t_L g1745 ( 
.A(n_1737),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1736),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1744),
.Y(n_1747)
);

NOR4xp75_ASAP7_75t_L g1748 ( 
.A(n_1743),
.B(n_1367),
.C(n_1344),
.D(n_1353),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1746),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1745),
.Y(n_1750)
);

AOI211xp5_ASAP7_75t_L g1751 ( 
.A1(n_1742),
.A2(n_1295),
.B(n_1349),
.C(n_1367),
.Y(n_1751)
);

NOR3xp33_ASAP7_75t_L g1752 ( 
.A(n_1747),
.B(n_1741),
.C(n_1344),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1750),
.B(n_1561),
.Y(n_1753)
);

NAND5xp2_ASAP7_75t_L g1754 ( 
.A(n_1751),
.B(n_1317),
.C(n_1309),
.D(n_1282),
.E(n_1521),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1753),
.Y(n_1755)
);

NAND4xp25_ASAP7_75t_L g1756 ( 
.A(n_1755),
.B(n_1752),
.C(n_1749),
.D(n_1754),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1756),
.Y(n_1757)
);

AOI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1756),
.A2(n_1748),
.B1(n_1317),
.B2(n_1309),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1758),
.B(n_1282),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1757),
.Y(n_1760)
);

NAND3xp33_ASAP7_75t_L g1761 ( 
.A(n_1760),
.B(n_1317),
.C(n_1603),
.Y(n_1761)
);

AO221x2_ASAP7_75t_L g1762 ( 
.A1(n_1759),
.A2(n_1309),
.B1(n_1626),
.B2(n_1603),
.C(n_1620),
.Y(n_1762)
);

AOI221xp5_ASAP7_75t_L g1763 ( 
.A1(n_1761),
.A2(n_1626),
.B1(n_1618),
.B2(n_1609),
.C(n_1584),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1763),
.Y(n_1764)
);

OAI221xp5_ASAP7_75t_R g1765 ( 
.A1(n_1764),
.A2(n_1762),
.B1(n_1618),
.B2(n_1609),
.C(n_1572),
.Y(n_1765)
);

AOI211xp5_ASAP7_75t_L g1766 ( 
.A1(n_1765),
.A2(n_1573),
.B(n_1563),
.C(n_1575),
.Y(n_1766)
);


endmodule