module fake_ariane_1090_n_1876 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1876);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1876;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_899;
wire n_352;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_718;
wire n_329;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_101),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_104),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_113),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_52),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_156),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_109),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_46),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_36),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_106),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_179),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_89),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_75),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_91),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_126),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_74),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_33),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_30),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_64),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_11),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_8),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_170),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_163),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_151),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_6),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_61),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_161),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_142),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_39),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_178),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_45),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_27),
.Y(n_212)
);

BUFx10_ASAP7_75t_L g213 ( 
.A(n_48),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_6),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_77),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_57),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_132),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_150),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_177),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_24),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_2),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g222 ( 
.A(n_112),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_58),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_144),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_11),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_44),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_24),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_131),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_76),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_5),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_174),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_48),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_164),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_115),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_35),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_120),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_165),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_52),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_92),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_63),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_172),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_143),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_60),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_37),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_47),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_102),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_118),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_30),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_33),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_171),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_111),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_168),
.Y(n_252)
);

BUFx5_ASAP7_75t_L g253 ( 
.A(n_153),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_87),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_82),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_124),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_20),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_162),
.Y(n_258)
);

BUFx10_ASAP7_75t_L g259 ( 
.A(n_23),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_157),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_26),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_70),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_36),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_65),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_40),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_29),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_127),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_29),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_72),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_105),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_20),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_49),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_73),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_8),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_32),
.Y(n_275)
);

BUFx10_ASAP7_75t_L g276 ( 
.A(n_85),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_88),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_47),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_12),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_79),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_121),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_107),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_86),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_95),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_147),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_97),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_78),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_35),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g289 ( 
.A(n_49),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_119),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_56),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_44),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_176),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_166),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_128),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_17),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_66),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_54),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_149),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_158),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_122),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_4),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_154),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_58),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_3),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_167),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_46),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_145),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_38),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_67),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_125),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_19),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_25),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_51),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_61),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_18),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_96),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_2),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_116),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_155),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_173),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_117),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_37),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_110),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_57),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_169),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_175),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_51),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_108),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_93),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_100),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_99),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_21),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_80),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_17),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_41),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_41),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_69),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_4),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_98),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_50),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_25),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_60),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_56),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_34),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_3),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_53),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_53),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_45),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_1),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_1),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_137),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_103),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_39),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_10),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_28),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_9),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_59),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_42),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_134),
.Y(n_360)
);

INVxp67_ASAP7_75t_SL g361 ( 
.A(n_205),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_212),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_199),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_240),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_181),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_181),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_184),
.B(n_0),
.Y(n_367)
);

BUFx2_ASAP7_75t_L g368 ( 
.A(n_201),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_260),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_287),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_205),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_206),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_332),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_201),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_206),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_184),
.B(n_0),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_198),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_195),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_276),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_298),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_195),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_235),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_203),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_203),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_207),
.B(n_5),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_276),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_313),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_349),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_276),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_307),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_335),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_224),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_328),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_289),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_185),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_289),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_349),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_336),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_359),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_333),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_333),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_207),
.B(n_7),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_268),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_R g404 ( 
.A(n_182),
.B(n_130),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_256),
.B(n_7),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_209),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_209),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_211),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_211),
.Y(n_409)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_197),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_183),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_183),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_202),
.Y(n_413)
);

NOR2xp67_ASAP7_75t_L g414 ( 
.A(n_302),
.B(n_9),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_188),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_227),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_210),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_202),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_227),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_258),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_230),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_258),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_189),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_230),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_243),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_243),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_245),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_210),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_299),
.Y(n_429)
);

CKINVDCx16_ASAP7_75t_R g430 ( 
.A(n_213),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_299),
.Y(n_431)
);

CKINVDCx16_ASAP7_75t_R g432 ( 
.A(n_213),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_245),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_200),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_261),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_213),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_259),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_261),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_214),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_216),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_220),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_217),
.B(n_10),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_259),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_263),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_263),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_223),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_272),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_272),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_259),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_403),
.Y(n_450)
);

NAND2xp33_ASAP7_75t_L g451 ( 
.A(n_442),
.B(n_268),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_403),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_378),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_378),
.B(n_344),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_381),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_381),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_383),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_383),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_384),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_384),
.B(n_344),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_417),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_417),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_428),
.B(n_217),
.Y(n_463)
);

OR2x2_ASAP7_75t_L g464 ( 
.A(n_368),
.B(n_357),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_428),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_361),
.B(n_357),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_406),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_396),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_371),
.B(n_274),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_407),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_408),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_409),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_416),
.Y(n_473)
);

OR2x2_ASAP7_75t_L g474 ( 
.A(n_368),
.B(n_274),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_374),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_394),
.Y(n_476)
);

INVx3_ASAP7_75t_L g477 ( 
.A(n_419),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_421),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_424),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_425),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_426),
.B(n_268),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_427),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_433),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_372),
.B(n_291),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_392),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_375),
.B(n_291),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_435),
.Y(n_487)
);

AND2x4_ASAP7_75t_L g488 ( 
.A(n_444),
.B(n_268),
.Y(n_488)
);

AND2x4_ASAP7_75t_L g489 ( 
.A(n_445),
.B(n_268),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_447),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_448),
.Y(n_491)
);

INVx4_ASAP7_75t_L g492 ( 
.A(n_392),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_367),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_388),
.B(n_360),
.Y(n_494)
);

INVxp67_ASAP7_75t_L g495 ( 
.A(n_439),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_397),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_376),
.Y(n_497)
);

INVx4_ASAP7_75t_L g498 ( 
.A(n_379),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_385),
.Y(n_499)
);

INVx1_ASAP7_75t_SL g500 ( 
.A(n_411),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_405),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_402),
.B(n_218),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_438),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_412),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_401),
.B(n_305),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_414),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_404),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_413),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_379),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_386),
.B(n_218),
.Y(n_510)
);

AND2x4_ASAP7_75t_L g511 ( 
.A(n_400),
.B(n_305),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_410),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_410),
.B(n_309),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_386),
.B(n_360),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_389),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_418),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_389),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_420),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_395),
.Y(n_519)
);

OA21x2_ASAP7_75t_L g520 ( 
.A1(n_395),
.A2(n_237),
.B(n_234),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_370),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g522 ( 
.A(n_377),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_415),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_390),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_415),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_422),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_423),
.B(n_234),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_459),
.Y(n_528)
);

NAND2xp33_ASAP7_75t_R g529 ( 
.A(n_485),
.B(n_365),
.Y(n_529)
);

AND2x6_ASAP7_75t_L g530 ( 
.A(n_521),
.B(n_237),
.Y(n_530)
);

AND2x2_ASAP7_75t_SL g531 ( 
.A(n_520),
.B(n_228),
.Y(n_531)
);

AND2x4_ASAP7_75t_L g532 ( 
.A(n_503),
.B(n_429),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_459),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_459),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_459),
.Y(n_535)
);

INVx1_ASAP7_75t_SL g536 ( 
.A(n_500),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_459),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_501),
.B(n_365),
.Y(n_538)
);

NAND3xp33_ASAP7_75t_L g539 ( 
.A(n_507),
.B(n_434),
.C(n_423),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_498),
.B(n_366),
.Y(n_540)
);

BUFx4f_ASAP7_75t_L g541 ( 
.A(n_520),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_501),
.B(n_507),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_501),
.B(n_366),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_501),
.B(n_370),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_459),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_457),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_498),
.B(n_434),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_459),
.Y(n_548)
);

INVx5_ASAP7_75t_L g549 ( 
.A(n_459),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_498),
.B(n_440),
.Y(n_550)
);

INVxp67_ASAP7_75t_SL g551 ( 
.A(n_463),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_507),
.B(n_498),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_520),
.A2(n_431),
.B1(n_343),
.B2(n_341),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_459),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_498),
.B(n_440),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_522),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_459),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_461),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g559 ( 
.A1(n_493),
.A2(n_441),
.B1(n_446),
.B2(n_232),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_461),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_461),
.Y(n_561)
);

AND2x6_ASAP7_75t_L g562 ( 
.A(n_521),
.B(n_252),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_461),
.Y(n_563)
);

INVx5_ASAP7_75t_L g564 ( 
.A(n_461),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_461),
.Y(n_565)
);

AND3x1_ASAP7_75t_L g566 ( 
.A(n_519),
.B(n_315),
.C(n_309),
.Y(n_566)
);

INVx4_ASAP7_75t_L g567 ( 
.A(n_461),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_498),
.B(n_441),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_515),
.B(n_446),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_501),
.B(n_499),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_461),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_461),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_515),
.B(n_380),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_503),
.B(n_430),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_461),
.Y(n_575)
);

OR2x6_ASAP7_75t_L g576 ( 
.A(n_466),
.B(n_315),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_509),
.B(n_432),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_457),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_509),
.B(n_390),
.Y(n_579)
);

BUFx10_ASAP7_75t_L g580 ( 
.A(n_485),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_453),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_453),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_501),
.B(n_194),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_499),
.B(n_222),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_453),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_453),
.Y(n_586)
);

AOI22xp33_ASAP7_75t_L g587 ( 
.A1(n_520),
.A2(n_339),
.B1(n_316),
.B2(n_318),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_455),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_455),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_458),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_458),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_499),
.B(n_269),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_462),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_462),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_455),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_455),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_456),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_462),
.Y(n_598)
);

OAI22xp33_ASAP7_75t_L g599 ( 
.A1(n_514),
.A2(n_391),
.B1(n_221),
.B2(n_248),
.Y(n_599)
);

BUFx3_ASAP7_75t_L g600 ( 
.A(n_467),
.Y(n_600)
);

NAND2xp33_ASAP7_75t_L g601 ( 
.A(n_521),
.B(n_509),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_456),
.Y(n_602)
);

CKINVDCx6p67_ASAP7_75t_R g603 ( 
.A(n_504),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_456),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_499),
.B(n_311),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_456),
.Y(n_606)
);

INVx4_ASAP7_75t_L g607 ( 
.A(n_471),
.Y(n_607)
);

CKINVDCx20_ASAP7_75t_R g608 ( 
.A(n_522),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_465),
.Y(n_609)
);

NAND2xp33_ASAP7_75t_L g610 ( 
.A(n_521),
.B(n_253),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_465),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_515),
.B(n_391),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_503),
.B(n_316),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_465),
.Y(n_614)
);

AND2x6_ASAP7_75t_L g615 ( 
.A(n_521),
.B(n_252),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_465),
.Y(n_616)
);

INVx4_ASAP7_75t_L g617 ( 
.A(n_471),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_471),
.Y(n_618)
);

INVxp67_ASAP7_75t_SL g619 ( 
.A(n_463),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_493),
.B(n_267),
.Y(n_620)
);

INVxp67_ASAP7_75t_L g621 ( 
.A(n_475),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_517),
.B(n_362),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_517),
.B(n_436),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_L g624 ( 
.A1(n_493),
.A2(n_312),
.B1(n_226),
.B2(n_238),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_450),
.Y(n_625)
);

AND2x6_ASAP7_75t_L g626 ( 
.A(n_521),
.B(n_267),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_470),
.Y(n_627)
);

INVx5_ASAP7_75t_L g628 ( 
.A(n_470),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_471),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_450),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_471),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_471),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_477),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_470),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_477),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_450),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_470),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_452),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_452),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_452),
.Y(n_640)
);

AOI22xp33_ASAP7_75t_L g641 ( 
.A1(n_520),
.A2(n_354),
.B1(n_342),
.B2(n_341),
.Y(n_641)
);

OR2x6_ASAP7_75t_L g642 ( 
.A(n_466),
.B(n_318),
.Y(n_642)
);

INVxp67_ASAP7_75t_SL g643 ( 
.A(n_463),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_509),
.B(n_225),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_520),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_477),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_470),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_477),
.Y(n_648)
);

INVx1_ASAP7_75t_SL g649 ( 
.A(n_500),
.Y(n_649)
);

XNOR2x2_ASAP7_75t_R g650 ( 
.A(n_500),
.B(n_382),
.Y(n_650)
);

CKINVDCx6p67_ASAP7_75t_R g651 ( 
.A(n_504),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_520),
.A2(n_323),
.B1(n_342),
.B2(n_339),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_470),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_470),
.Y(n_654)
);

INVx2_ASAP7_75t_SL g655 ( 
.A(n_503),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_497),
.B(n_270),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_470),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_454),
.B(n_323),
.Y(n_658)
);

INVxp33_ASAP7_75t_L g659 ( 
.A(n_475),
.Y(n_659)
);

AND2x4_ASAP7_75t_L g660 ( 
.A(n_466),
.B(n_337),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_509),
.B(n_244),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_470),
.Y(n_662)
);

INVx2_ASAP7_75t_SL g663 ( 
.A(n_466),
.Y(n_663)
);

INVx6_ASAP7_75t_L g664 ( 
.A(n_470),
.Y(n_664)
);

BUFx3_ASAP7_75t_L g665 ( 
.A(n_467),
.Y(n_665)
);

INVx4_ASAP7_75t_L g666 ( 
.A(n_477),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_514),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_487),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_487),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_487),
.Y(n_670)
);

BUFx6f_ASAP7_75t_L g671 ( 
.A(n_487),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_517),
.B(n_519),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_514),
.Y(n_673)
);

INVx3_ASAP7_75t_L g674 ( 
.A(n_487),
.Y(n_674)
);

AO22x2_ASAP7_75t_L g675 ( 
.A1(n_511),
.A2(n_337),
.B1(n_343),
.B2(n_354),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_497),
.B(n_270),
.Y(n_676)
);

NAND2xp33_ASAP7_75t_L g677 ( 
.A(n_521),
.B(n_253),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_477),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_546),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_663),
.B(n_509),
.Y(n_680)
);

AOI22xp5_ASAP7_75t_L g681 ( 
.A1(n_667),
.A2(n_519),
.B1(n_525),
.B2(n_523),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_SL g682 ( 
.A(n_536),
.B(n_649),
.Y(n_682)
);

BUFx3_ASAP7_75t_L g683 ( 
.A(n_580),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_667),
.B(n_497),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_673),
.B(n_523),
.Y(n_685)
);

NAND3xp33_ASAP7_75t_L g686 ( 
.A(n_569),
.B(n_495),
.C(n_523),
.Y(n_686)
);

AND2x2_ASAP7_75t_SL g687 ( 
.A(n_531),
.B(n_502),
.Y(n_687)
);

INVxp67_ASAP7_75t_L g688 ( 
.A(n_574),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_673),
.B(n_525),
.Y(n_689)
);

BUFx8_ASAP7_75t_L g690 ( 
.A(n_574),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_542),
.B(n_525),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_546),
.Y(n_692)
);

AOI22xp5_ASAP7_75t_L g693 ( 
.A1(n_672),
.A2(n_521),
.B1(n_510),
.B2(n_502),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_529),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_551),
.B(n_510),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_619),
.B(n_527),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_556),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_643),
.B(n_527),
.Y(n_698)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_570),
.A2(n_451),
.B(n_478),
.Y(n_699)
);

O2A1O1Ixp5_ASAP7_75t_L g700 ( 
.A1(n_552),
.A2(n_492),
.B(n_478),
.C(n_483),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_532),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_538),
.B(n_521),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_532),
.B(n_476),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_590),
.Y(n_704)
);

OA22x2_ASAP7_75t_L g705 ( 
.A1(n_576),
.A2(n_511),
.B1(n_505),
.B2(n_512),
.Y(n_705)
);

AOI221xp5_ASAP7_75t_L g706 ( 
.A1(n_599),
.A2(n_511),
.B1(n_513),
.B2(n_512),
.C(n_476),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_532),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_590),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_543),
.B(n_521),
.Y(n_709)
);

INVx2_ASAP7_75t_SL g710 ( 
.A(n_580),
.Y(n_710)
);

BUFx6f_ASAP7_75t_L g711 ( 
.A(n_634),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_581),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_578),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_581),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_578),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_541),
.B(n_492),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_541),
.B(n_492),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_544),
.B(n_492),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_582),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_655),
.B(n_492),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_655),
.B(n_492),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_556),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_573),
.B(n_495),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_541),
.B(n_487),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_608),
.Y(n_725)
);

OAI22xp33_ASAP7_75t_L g726 ( 
.A1(n_576),
.A2(n_474),
.B1(n_464),
.B2(n_494),
.Y(n_726)
);

OAI22xp33_ASAP7_75t_L g727 ( 
.A1(n_576),
.A2(n_474),
.B1(n_464),
.B2(n_494),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_585),
.Y(n_728)
);

INVxp67_ASAP7_75t_L g729 ( 
.A(n_623),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_577),
.B(n_524),
.Y(n_730)
);

INVxp67_ASAP7_75t_L g731 ( 
.A(n_622),
.Y(n_731)
);

AOI22xp5_ASAP7_75t_L g732 ( 
.A1(n_675),
.A2(n_511),
.B1(n_506),
.B2(n_524),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_585),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_607),
.B(n_487),
.Y(n_734)
);

NAND2xp33_ASAP7_75t_L g735 ( 
.A(n_634),
.B(n_487),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_659),
.B(n_508),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_539),
.B(n_506),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_584),
.B(n_478),
.Y(n_738)
);

BUFx6f_ASAP7_75t_L g739 ( 
.A(n_634),
.Y(n_739)
);

BUFx3_ASAP7_75t_L g740 ( 
.A(n_580),
.Y(n_740)
);

OAI22xp5_ASAP7_75t_SL g741 ( 
.A1(n_608),
.A2(n_387),
.B1(n_399),
.B2(n_398),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_592),
.B(n_478),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_663),
.B(n_583),
.Y(n_743)
);

INVxp67_ASAP7_75t_L g744 ( 
.A(n_612),
.Y(n_744)
);

NAND3xp33_ASAP7_75t_L g745 ( 
.A(n_559),
.B(n_512),
.C(n_474),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_605),
.B(n_579),
.Y(n_746)
);

BUFx6f_ASAP7_75t_SL g747 ( 
.A(n_660),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_607),
.B(n_506),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_586),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_607),
.B(n_487),
.Y(n_750)
);

CKINVDCx20_ASAP7_75t_R g751 ( 
.A(n_603),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_617),
.B(n_511),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_555),
.B(n_478),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_568),
.B(n_511),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_621),
.B(n_511),
.Y(n_755)
);

OR2x6_ASAP7_75t_L g756 ( 
.A(n_576),
.B(n_504),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_586),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_617),
.B(n_505),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_617),
.B(n_666),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_588),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_588),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_591),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_L g763 ( 
.A(n_666),
.B(n_505),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_666),
.B(n_505),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_591),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_593),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_645),
.B(n_531),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_589),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_603),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_547),
.B(n_505),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_593),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_550),
.B(n_505),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_595),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_600),
.B(n_478),
.Y(n_774)
);

INVxp67_ASAP7_75t_L g775 ( 
.A(n_566),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_594),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_594),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_600),
.B(n_482),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_601),
.A2(n_677),
.B(n_610),
.Y(n_779)
);

OR2x2_ASAP7_75t_L g780 ( 
.A(n_642),
.B(n_468),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_540),
.B(n_505),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_642),
.B(n_482),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_595),
.Y(n_783)
);

INVx2_ASAP7_75t_SL g784 ( 
.A(n_613),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_651),
.B(n_508),
.Y(n_785)
);

OR2x6_ASAP7_75t_L g786 ( 
.A(n_642),
.B(n_504),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_665),
.B(n_482),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_665),
.B(n_482),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_645),
.B(n_487),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_598),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_613),
.B(n_482),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_642),
.B(n_644),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_675),
.A2(n_513),
.B1(n_490),
.B2(n_473),
.Y(n_793)
);

BUFx3_ASAP7_75t_L g794 ( 
.A(n_651),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_620),
.B(n_482),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_598),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_656),
.B(n_483),
.Y(n_797)
);

OAI22xp5_ASAP7_75t_SL g798 ( 
.A1(n_553),
.A2(n_393),
.B1(n_364),
.B2(n_369),
.Y(n_798)
);

BUFx6f_ASAP7_75t_SL g799 ( 
.A(n_660),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_660),
.B(n_483),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_676),
.B(n_483),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_618),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_661),
.B(n_483),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_L g804 ( 
.A1(n_675),
.A2(n_513),
.B1(n_490),
.B2(n_473),
.Y(n_804)
);

AOI22xp5_ASAP7_75t_L g805 ( 
.A1(n_675),
.A2(n_451),
.B1(n_479),
.B2(n_480),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_658),
.B(n_483),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_658),
.B(n_467),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_618),
.B(n_473),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_629),
.B(n_474),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_629),
.B(n_472),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_631),
.B(n_473),
.Y(n_811)
);

INVxp67_ASAP7_75t_L g812 ( 
.A(n_624),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_SL g813 ( 
.A(n_650),
.B(n_518),
.Y(n_813)
);

OR2x2_ASAP7_75t_L g814 ( 
.A(n_650),
.B(n_468),
.Y(n_814)
);

A2O1A1Ixp33_ASAP7_75t_L g815 ( 
.A1(n_631),
.A2(n_472),
.B(n_480),
.C(n_479),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_632),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_632),
.B(n_472),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_587),
.B(n_508),
.Y(n_818)
);

INVx3_ASAP7_75t_L g819 ( 
.A(n_596),
.Y(n_819)
);

OAI221xp5_ASAP7_75t_L g820 ( 
.A1(n_641),
.A2(n_479),
.B1(n_480),
.B2(n_491),
.C(n_464),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_633),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_596),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_633),
.B(n_491),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_635),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_635),
.B(n_646),
.Y(n_825)
);

INVx2_ASAP7_75t_SL g826 ( 
.A(n_625),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_646),
.B(n_648),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_648),
.B(n_491),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_678),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_678),
.B(n_490),
.Y(n_830)
);

OR2x6_ASAP7_75t_L g831 ( 
.A(n_597),
.B(n_518),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_652),
.B(n_454),
.Y(n_832)
);

INVx2_ASAP7_75t_SL g833 ( 
.A(n_625),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_634),
.B(n_513),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_597),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_602),
.B(n_454),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_602),
.B(n_454),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_609),
.B(n_614),
.Y(n_838)
);

INVx2_ASAP7_75t_SL g839 ( 
.A(n_630),
.Y(n_839)
);

INVx4_ASAP7_75t_L g840 ( 
.A(n_634),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_609),
.B(n_460),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_637),
.B(n_464),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_630),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_614),
.Y(n_844)
);

INVx3_ASAP7_75t_L g845 ( 
.A(n_840),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_819),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_744),
.B(n_508),
.Y(n_847)
);

BUFx2_ASAP7_75t_SL g848 ( 
.A(n_751),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_685),
.B(n_516),
.Y(n_849)
);

NAND3xp33_ASAP7_75t_L g850 ( 
.A(n_731),
.B(n_601),
.C(n_526),
.Y(n_850)
);

AOI21xp5_ASAP7_75t_L g851 ( 
.A1(n_759),
.A2(n_677),
.B(n_610),
.Y(n_851)
);

INVx2_ASAP7_75t_SL g852 ( 
.A(n_690),
.Y(n_852)
);

OAI22xp5_ASAP7_75t_L g853 ( 
.A1(n_687),
.A2(n_567),
.B1(n_606),
.B2(n_604),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_759),
.A2(n_557),
.B(n_533),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_703),
.B(n_518),
.Y(n_855)
);

NOR2xp67_ASAP7_75t_L g856 ( 
.A(n_694),
.B(n_516),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_712),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_685),
.B(n_516),
.Y(n_858)
);

A2O1A1Ixp33_ASAP7_75t_L g859 ( 
.A1(n_691),
.A2(n_606),
.B(n_611),
.C(n_604),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_789),
.A2(n_557),
.B(n_533),
.Y(n_860)
);

INVx3_ASAP7_75t_L g861 ( 
.A(n_840),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_729),
.B(n_518),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_714),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_687),
.B(n_637),
.Y(n_864)
);

AOI21xp5_ASAP7_75t_L g865 ( 
.A1(n_789),
.A2(n_560),
.B(n_558),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_753),
.A2(n_560),
.B(n_558),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_713),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_688),
.B(n_516),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_724),
.A2(n_563),
.B(n_561),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_696),
.B(n_526),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_724),
.A2(n_709),
.B(n_702),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_SL g872 ( 
.A1(n_767),
.A2(n_653),
.B(n_647),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_693),
.B(n_637),
.Y(n_873)
);

O2A1O1Ixp33_ASAP7_75t_L g874 ( 
.A1(n_754),
.A2(n_616),
.B(n_611),
.C(n_490),
.Y(n_874)
);

NAND3xp33_ASAP7_75t_L g875 ( 
.A(n_686),
.B(n_526),
.C(n_373),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_715),
.Y(n_876)
);

BUFx6f_ASAP7_75t_L g877 ( 
.A(n_711),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_698),
.B(n_526),
.Y(n_878)
);

HB1xp67_ASAP7_75t_L g879 ( 
.A(n_747),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_695),
.B(n_616),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_723),
.B(n_363),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_812),
.B(n_567),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_819),
.Y(n_883)
);

OAI22xp5_ASAP7_75t_L g884 ( 
.A1(n_752),
.A2(n_567),
.B1(n_534),
.B2(n_554),
.Y(n_884)
);

O2A1O1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_726),
.A2(n_494),
.B(n_563),
.C(n_565),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_719),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_702),
.A2(n_565),
.B(n_561),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_684),
.B(n_460),
.Y(n_888)
);

OAI21xp33_ASAP7_75t_L g889 ( 
.A1(n_691),
.A2(n_257),
.B(n_249),
.Y(n_889)
);

NAND3xp33_ASAP7_75t_SL g890 ( 
.A(n_706),
.B(n_443),
.C(n_437),
.Y(n_890)
);

A2O1A1Ixp33_ASAP7_75t_L g891 ( 
.A1(n_743),
.A2(n_460),
.B(n_638),
.C(n_636),
.Y(n_891)
);

BUFx3_ASAP7_75t_L g892 ( 
.A(n_794),
.Y(n_892)
);

AOI22xp5_ASAP7_75t_L g893 ( 
.A1(n_726),
.A2(n_562),
.B1(n_530),
.B2(n_626),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_681),
.B(n_637),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_689),
.B(n_627),
.Y(n_895)
);

INVx3_ASAP7_75t_L g896 ( 
.A(n_711),
.Y(n_896)
);

AOI21xp5_ASAP7_75t_L g897 ( 
.A1(n_709),
.A2(n_721),
.B(n_720),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_743),
.B(n_460),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_809),
.B(n_636),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_746),
.B(n_627),
.Y(n_900)
);

INVx1_ASAP7_75t_SL g901 ( 
.A(n_682),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_728),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_716),
.A2(n_535),
.B(n_528),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_716),
.A2(n_535),
.B(n_528),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_809),
.B(n_638),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_711),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_762),
.Y(n_907)
);

HB1xp67_ASAP7_75t_L g908 ( 
.A(n_747),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_717),
.A2(n_545),
.B(n_537),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_717),
.A2(n_545),
.B(n_537),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_765),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_734),
.A2(n_572),
.B(n_548),
.Y(n_912)
);

CKINVDCx12_ASAP7_75t_R g913 ( 
.A(n_741),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_734),
.A2(n_572),
.B(n_548),
.Y(n_914)
);

NOR2x1p5_ASAP7_75t_L g915 ( 
.A(n_683),
.B(n_469),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_766),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_746),
.A2(n_640),
.B(n_639),
.C(n_488),
.Y(n_917)
);

NOR2xp67_ASAP7_75t_L g918 ( 
.A(n_710),
.B(n_496),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_750),
.A2(n_825),
.B(n_742),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_784),
.B(n_639),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_843),
.B(n_640),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_733),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_750),
.A2(n_575),
.B(n_647),
.Y(n_923)
);

AOI33xp33_ASAP7_75t_L g924 ( 
.A1(n_727),
.A2(n_469),
.A3(n_484),
.B1(n_486),
.B2(n_489),
.B3(n_481),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_680),
.B(n_530),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_680),
.B(n_530),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_749),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_771),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_757),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_825),
.A2(n_575),
.B(n_653),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_752),
.B(n_530),
.Y(n_931)
);

NOR2xp67_ASAP7_75t_L g932 ( 
.A(n_769),
.B(n_496),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_738),
.A2(n_797),
.B(n_795),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_801),
.A2(n_657),
.B(n_654),
.Y(n_934)
);

OAI21xp5_ASAP7_75t_L g935 ( 
.A1(n_779),
.A2(n_657),
.B(n_654),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_748),
.B(n_530),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_748),
.B(n_530),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_727),
.B(n_530),
.Y(n_938)
);

OAI21xp5_ASAP7_75t_L g939 ( 
.A1(n_700),
.A2(n_670),
.B(n_669),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_776),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_818),
.B(n_562),
.Y(n_941)
);

AOI21x1_ASAP7_75t_L g942 ( 
.A1(n_808),
.A2(n_670),
.B(n_669),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_827),
.A2(n_554),
.B(n_534),
.Y(n_943)
);

OR2x6_ASAP7_75t_L g944 ( 
.A(n_756),
.B(n_496),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_730),
.B(n_627),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_737),
.B(n_562),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_838),
.A2(n_554),
.B(n_534),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_737),
.B(n_562),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_730),
.B(n_674),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_777),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_790),
.Y(n_951)
);

O2A1O1Ixp33_ASAP7_75t_L g952 ( 
.A1(n_755),
.A2(n_674),
.B(n_571),
.C(n_190),
.Y(n_952)
);

AOI22xp5_ASAP7_75t_L g953 ( 
.A1(n_792),
.A2(n_562),
.B1(n_615),
.B2(n_626),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_796),
.Y(n_954)
);

OAI21xp5_ASAP7_75t_L g955 ( 
.A1(n_699),
.A2(n_571),
.B(n_674),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_774),
.A2(n_571),
.B(n_637),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_807),
.B(n_782),
.Y(n_957)
);

OAI22xp5_ASAP7_75t_L g958 ( 
.A1(n_758),
.A2(n_664),
.B1(n_668),
.B2(n_671),
.Y(n_958)
);

OAI22xp5_ASAP7_75t_L g959 ( 
.A1(n_758),
.A2(n_664),
.B1(n_668),
.B2(n_671),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_778),
.A2(n_668),
.B(n_662),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_794),
.B(n_469),
.Y(n_961)
);

OR2x6_ASAP7_75t_L g962 ( 
.A(n_756),
.B(n_496),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_782),
.B(n_562),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_806),
.B(n_763),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_763),
.B(n_662),
.Y(n_965)
);

OR2x2_ASAP7_75t_L g966 ( 
.A(n_780),
.B(n_469),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_760),
.Y(n_967)
);

OAI21xp5_ASAP7_75t_L g968 ( 
.A1(n_764),
.A2(n_615),
.B(n_562),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_761),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_787),
.A2(n_668),
.B(n_662),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_788),
.A2(n_668),
.B(n_662),
.Y(n_971)
);

OAI321xp33_ASAP7_75t_L g972 ( 
.A1(n_732),
.A2(n_281),
.A3(n_334),
.B1(n_320),
.B2(n_273),
.C(n_293),
.Y(n_972)
);

INVx2_ASAP7_75t_L g973 ( 
.A(n_768),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_711),
.Y(n_974)
);

CKINVDCx10_ASAP7_75t_R g975 ( 
.A(n_799),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_764),
.B(n_615),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_802),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_793),
.B(n_615),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_793),
.B(n_615),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_816),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_718),
.A2(n_671),
.B(n_662),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_821),
.Y(n_982)
);

O2A1O1Ixp33_ASAP7_75t_L g983 ( 
.A1(n_842),
.A2(n_196),
.B(n_486),
.C(n_484),
.Y(n_983)
);

OAI21xp5_ASAP7_75t_L g984 ( 
.A1(n_808),
.A2(n_626),
.B(n_615),
.Y(n_984)
);

OAI21xp5_ASAP7_75t_L g985 ( 
.A1(n_811),
.A2(n_626),
.B(n_615),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_718),
.A2(n_671),
.B(n_564),
.Y(n_986)
);

HB1xp67_ASAP7_75t_L g987 ( 
.A(n_799),
.Y(n_987)
);

AND2x4_ASAP7_75t_L g988 ( 
.A(n_785),
.B(n_484),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_739),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_773),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_804),
.B(n_626),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_739),
.B(n_671),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_L g993 ( 
.A1(n_791),
.A2(n_664),
.B1(n_325),
.B2(n_351),
.Y(n_993)
);

INVx4_ASAP7_75t_L g994 ( 
.A(n_831),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_811),
.A2(n_564),
.B(n_549),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_830),
.A2(n_564),
.B(n_549),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_824),
.Y(n_997)
);

OAI21xp5_ASAP7_75t_L g998 ( 
.A1(n_830),
.A2(n_626),
.B(n_564),
.Y(n_998)
);

OAI22xp5_ASAP7_75t_L g999 ( 
.A1(n_679),
.A2(n_664),
.B1(n_356),
.B2(n_355),
.Y(n_999)
);

AOI21x1_ASAP7_75t_L g1000 ( 
.A1(n_810),
.A2(n_277),
.B(n_273),
.Y(n_1000)
);

OAI21xp33_ASAP7_75t_L g1001 ( 
.A1(n_770),
.A2(n_266),
.B(n_265),
.Y(n_1001)
);

OAI21xp33_ASAP7_75t_SL g1002 ( 
.A1(n_705),
.A2(n_486),
.B(n_484),
.Y(n_1002)
);

BUFx2_ASAP7_75t_L g1003 ( 
.A(n_697),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_817),
.A2(n_564),
.B(n_549),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_722),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_823),
.A2(n_549),
.B(n_628),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_828),
.A2(n_767),
.B(n_735),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_836),
.A2(n_549),
.B(n_628),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_804),
.B(n_701),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_837),
.A2(n_628),
.B(n_187),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_841),
.A2(n_628),
.B(n_191),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_783),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_707),
.B(n_626),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_829),
.A2(n_628),
.B(n_247),
.Y(n_1014)
);

OAI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_815),
.A2(n_486),
.B(n_489),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_803),
.A2(n_246),
.B(n_353),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_775),
.B(n_792),
.Y(n_1017)
);

AO21x1_ASAP7_75t_L g1018 ( 
.A1(n_803),
.A2(n_286),
.B(n_334),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_692),
.A2(n_296),
.B1(n_271),
.B2(n_275),
.Y(n_1019)
);

AOI22xp33_ASAP7_75t_L g1020 ( 
.A1(n_832),
.A2(n_489),
.B1(n_488),
.B2(n_481),
.Y(n_1020)
);

NOR3xp33_ASAP7_75t_L g1021 ( 
.A(n_745),
.B(n_304),
.C(n_288),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_844),
.A2(n_772),
.B(n_770),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_826),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_772),
.A2(n_290),
.B(n_215),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_833),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_822),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_800),
.B(n_481),
.Y(n_1027)
);

A2O1A1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_781),
.A2(n_489),
.B(n_488),
.C(n_481),
.Y(n_1028)
);

NAND2x1_ASAP7_75t_L g1029 ( 
.A(n_739),
.B(n_481),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_834),
.A2(n_208),
.B(n_204),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_839),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_690),
.B(n_449),
.Y(n_1032)
);

BUFx2_ASAP7_75t_L g1033 ( 
.A(n_1005),
.Y(n_1033)
);

CKINVDCx20_ASAP7_75t_R g1034 ( 
.A(n_913),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_867),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_876),
.Y(n_1036)
);

AND2x4_ASAP7_75t_L g1037 ( 
.A(n_892),
.B(n_756),
.Y(n_1037)
);

AND2x6_ASAP7_75t_L g1038 ( 
.A(n_877),
.B(n_805),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_957),
.B(n_708),
.Y(n_1039)
);

O2A1O1Ixp33_ASAP7_75t_SL g1040 ( 
.A1(n_964),
.A2(n_965),
.B(n_976),
.C(n_864),
.Y(n_1040)
);

OAI21xp33_ASAP7_75t_SL g1041 ( 
.A1(n_924),
.A2(n_705),
.B(n_781),
.Y(n_1041)
);

HB1xp67_ASAP7_75t_L g1042 ( 
.A(n_855),
.Y(n_1042)
);

AND2x4_ASAP7_75t_L g1043 ( 
.A(n_892),
.B(n_786),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_975),
.Y(n_1044)
);

OR2x6_ASAP7_75t_L g1045 ( 
.A(n_852),
.B(n_786),
.Y(n_1045)
);

O2A1O1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_1021),
.A2(n_683),
.B(n_740),
.C(n_704),
.Y(n_1046)
);

OA22x2_ASAP7_75t_L g1047 ( 
.A1(n_988),
.A2(n_798),
.B1(n_786),
.B2(n_725),
.Y(n_1047)
);

A2O1A1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_1022),
.A2(n_820),
.B(n_740),
.C(n_835),
.Y(n_1048)
);

O2A1O1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_1021),
.A2(n_814),
.B(n_831),
.C(n_736),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_862),
.B(n_813),
.Y(n_1050)
);

O2A1O1Ixp33_ASAP7_75t_L g1051 ( 
.A1(n_847),
.A2(n_831),
.B(n_320),
.C(n_284),
.Y(n_1051)
);

O2A1O1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_847),
.A2(n_338),
.B(n_293),
.C(n_286),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_877),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_857),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_1017),
.B(n_739),
.Y(n_1055)
);

BUFx3_ASAP7_75t_L g1056 ( 
.A(n_1003),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_898),
.B(n_481),
.Y(n_1057)
);

A2O1A1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_882),
.A2(n_338),
.B(n_277),
.C(n_281),
.Y(n_1058)
);

AOI22xp33_ASAP7_75t_L g1059 ( 
.A1(n_890),
.A2(n_488),
.B1(n_481),
.B2(n_489),
.Y(n_1059)
);

BUFx8_ASAP7_75t_L g1060 ( 
.A(n_961),
.Y(n_1060)
);

O2A1O1Ixp5_ASAP7_75t_L g1061 ( 
.A1(n_873),
.A2(n_489),
.B(n_488),
.C(n_284),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_1017),
.B(n_488),
.Y(n_1062)
);

BUFx2_ASAP7_75t_L g1063 ( 
.A(n_961),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_881),
.B(n_488),
.Y(n_1064)
);

O2A1O1Ixp33_ASAP7_75t_SL g1065 ( 
.A1(n_965),
.A2(n_864),
.B(n_931),
.C(n_891),
.Y(n_1065)
);

NOR3xp33_ASAP7_75t_SL g1066 ( 
.A(n_889),
.B(n_1019),
.C(n_279),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_881),
.B(n_966),
.Y(n_1067)
);

NOR2xp33_ASAP7_75t_L g1068 ( 
.A(n_988),
.B(n_278),
.Y(n_1068)
);

OAI22xp33_ASAP7_75t_L g1069 ( 
.A1(n_849),
.A2(n_346),
.B1(n_358),
.B2(n_350),
.Y(n_1069)
);

A2O1A1Ixp33_ASAP7_75t_L g1070 ( 
.A1(n_882),
.A2(n_949),
.B(n_945),
.C(n_900),
.Y(n_1070)
);

AOI22x1_ASAP7_75t_L g1071 ( 
.A1(n_933),
.A2(n_489),
.B1(n_348),
.B2(n_347),
.Y(n_1071)
);

BUFx4f_ASAP7_75t_L g1072 ( 
.A(n_944),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_897),
.A2(n_236),
.B(n_228),
.Y(n_1073)
);

INVx4_ASAP7_75t_L g1074 ( 
.A(n_994),
.Y(n_1074)
);

HB1xp67_ASAP7_75t_L g1075 ( 
.A(n_879),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_899),
.A2(n_345),
.B1(n_292),
.B2(n_314),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_877),
.Y(n_1077)
);

OR2x2_ASAP7_75t_L g1078 ( 
.A(n_868),
.B(n_236),
.Y(n_1078)
);

O2A1O1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_858),
.A2(n_12),
.B(n_13),
.C(n_14),
.Y(n_1079)
);

NOR2xp33_ASAP7_75t_L g1080 ( 
.A(n_875),
.B(n_186),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_857),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_877),
.Y(n_1082)
);

OAI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_871),
.A2(n_352),
.B(n_340),
.Y(n_1083)
);

AO21x1_ASAP7_75t_L g1084 ( 
.A1(n_946),
.A2(n_253),
.B(n_283),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_868),
.B(n_13),
.Y(n_1085)
);

NAND2x1p5_ASAP7_75t_L g1086 ( 
.A(n_994),
.B(n_283),
.Y(n_1086)
);

INVx4_ASAP7_75t_L g1087 ( 
.A(n_944),
.Y(n_1087)
);

NAND2x1p5_ASAP7_75t_L g1088 ( 
.A(n_845),
.B(n_283),
.Y(n_1088)
);

NAND2x1p5_ASAP7_75t_L g1089 ( 
.A(n_845),
.B(n_283),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_900),
.B(n_253),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_870),
.B(n_878),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_851),
.A2(n_981),
.B(n_986),
.Y(n_1092)
);

NAND3xp33_ASAP7_75t_SL g1093 ( 
.A(n_1001),
.B(n_331),
.C(n_330),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_1009),
.B(n_253),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_888),
.B(n_253),
.Y(n_1095)
);

BUFx3_ASAP7_75t_L g1096 ( 
.A(n_879),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_935),
.A2(n_942),
.B(n_904),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_921),
.B(n_1023),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_936),
.A2(n_937),
.B(n_854),
.Y(n_1099)
);

BUFx2_ASAP7_75t_SL g1100 ( 
.A(n_908),
.Y(n_1100)
);

HB1xp67_ASAP7_75t_L g1101 ( 
.A(n_908),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_945),
.B(n_192),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_905),
.B(n_253),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_924),
.B(n_949),
.Y(n_1104)
);

CKINVDCx20_ASAP7_75t_R g1105 ( 
.A(n_848),
.Y(n_1105)
);

AOI33xp33_ASAP7_75t_L g1106 ( 
.A1(n_907),
.A2(n_14),
.A3(n_15),
.B1(n_16),
.B2(n_18),
.B3(n_19),
.Y(n_1106)
);

OAI22xp5_ASAP7_75t_SL g1107 ( 
.A1(n_1032),
.A2(n_329),
.B1(n_327),
.B2(n_326),
.Y(n_1107)
);

OAI22x1_ASAP7_75t_L g1108 ( 
.A1(n_1032),
.A2(n_324),
.B1(n_322),
.B2(n_321),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_915),
.B(n_15),
.Y(n_1109)
);

HB1xp67_ASAP7_75t_L g1110 ( 
.A(n_987),
.Y(n_1110)
);

INVx1_ASAP7_75t_SL g1111 ( 
.A(n_901),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_911),
.B(n_253),
.Y(n_1112)
);

A2O1A1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_948),
.A2(n_319),
.B(n_317),
.C(n_310),
.Y(n_1113)
);

O2A1O1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_891),
.A2(n_16),
.B(n_21),
.C(n_22),
.Y(n_1114)
);

NOR2xp67_ASAP7_75t_L g1115 ( 
.A(n_987),
.B(n_193),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_916),
.Y(n_1116)
);

AND2x4_ASAP7_75t_L g1117 ( 
.A(n_944),
.B(n_22),
.Y(n_1117)
);

OR2x6_ASAP7_75t_L g1118 ( 
.A(n_962),
.B(n_283),
.Y(n_1118)
);

INVx3_ASAP7_75t_L g1119 ( 
.A(n_974),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_887),
.A2(n_308),
.B(n_306),
.Y(n_1120)
);

O2A1O1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_1002),
.A2(n_23),
.B(n_26),
.C(n_27),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_893),
.A2(n_938),
.B1(n_940),
.B2(n_954),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_974),
.Y(n_1123)
);

BUFx6f_ASAP7_75t_L g1124 ( 
.A(n_974),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_863),
.Y(n_1125)
);

BUFx2_ASAP7_75t_L g1126 ( 
.A(n_962),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_880),
.A2(n_303),
.B(n_301),
.Y(n_1127)
);

NAND3xp33_ASAP7_75t_L g1128 ( 
.A(n_850),
.B(n_300),
.C(n_297),
.Y(n_1128)
);

BUFx3_ASAP7_75t_L g1129 ( 
.A(n_962),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_873),
.A2(n_295),
.B(n_294),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_974),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_928),
.B(n_253),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_918),
.B(n_1025),
.Y(n_1133)
);

A2O1A1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_885),
.A2(n_285),
.B(n_282),
.C(n_280),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_950),
.B(n_28),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_1031),
.B(n_264),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_951),
.B(n_977),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_856),
.B(n_31),
.Y(n_1138)
);

AOI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_932),
.A2(n_262),
.B1(n_255),
.B2(n_254),
.Y(n_1139)
);

AOI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_963),
.A2(n_239),
.B1(n_250),
.B2(n_242),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_896),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_896),
.Y(n_1142)
);

INVx3_ASAP7_75t_L g1143 ( 
.A(n_861),
.Y(n_1143)
);

INVx3_ASAP7_75t_L g1144 ( 
.A(n_861),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_980),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_R g1146 ( 
.A(n_906),
.B(n_251),
.Y(n_1146)
);

HB1xp67_ASAP7_75t_L g1147 ( 
.A(n_982),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_997),
.B(n_241),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_SL g1149 ( 
.A(n_972),
.B(n_906),
.Y(n_1149)
);

O2A1O1Ixp33_ASAP7_75t_SL g1150 ( 
.A1(n_992),
.A2(n_31),
.B(n_32),
.C(n_34),
.Y(n_1150)
);

AOI21x1_ASAP7_75t_L g1151 ( 
.A1(n_1000),
.A2(n_233),
.B(n_231),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_989),
.Y(n_1152)
);

HB1xp67_ASAP7_75t_L g1153 ( 
.A(n_846),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_920),
.B(n_1020),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_886),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_989),
.B(n_229),
.Y(n_1156)
);

AND2x4_ASAP7_75t_L g1157 ( 
.A(n_1028),
.B(n_38),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_1029),
.Y(n_1158)
);

OAI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_859),
.A2(n_219),
.B(n_42),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1007),
.A2(n_114),
.B(n_160),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_1020),
.B(n_40),
.Y(n_1161)
);

NOR2xp33_ASAP7_75t_L g1162 ( 
.A(n_883),
.B(n_1027),
.Y(n_1162)
);

AOI221xp5_ASAP7_75t_L g1163 ( 
.A1(n_983),
.A2(n_43),
.B1(n_50),
.B2(n_54),
.C(n_55),
.Y(n_1163)
);

O2A1O1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_917),
.A2(n_43),
.B(n_55),
.C(n_59),
.Y(n_1164)
);

BUFx8_ASAP7_75t_L g1165 ( 
.A(n_902),
.Y(n_1165)
);

INVx4_ASAP7_75t_L g1166 ( 
.A(n_922),
.Y(n_1166)
);

INVx3_ASAP7_75t_L g1167 ( 
.A(n_967),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_958),
.A2(n_959),
.B(n_866),
.Y(n_1168)
);

OAI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_859),
.A2(n_917),
.B(n_919),
.Y(n_1169)
);

AND3x1_ASAP7_75t_SL g1170 ( 
.A(n_1030),
.B(n_180),
.C(n_68),
.Y(n_1170)
);

BUFx3_ASAP7_75t_L g1171 ( 
.A(n_927),
.Y(n_1171)
);

O2A1O1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_1028),
.A2(n_62),
.B(n_71),
.C(n_81),
.Y(n_1172)
);

BUFx2_ASAP7_75t_L g1173 ( 
.A(n_925),
.Y(n_1173)
);

AOI22xp33_ASAP7_75t_L g1174 ( 
.A1(n_929),
.A2(n_83),
.B1(n_84),
.B2(n_90),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_969),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_894),
.A2(n_94),
.B(n_123),
.C(n_129),
.Y(n_1176)
);

OAI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_968),
.A2(n_133),
.B1(n_135),
.B2(n_136),
.Y(n_1177)
);

BUFx2_ASAP7_75t_L g1178 ( 
.A(n_926),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_990),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_934),
.A2(n_138),
.B(n_139),
.Y(n_1180)
);

CKINVDCx11_ASAP7_75t_R g1181 ( 
.A(n_1012),
.Y(n_1181)
);

OAI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1015),
.A2(n_140),
.B1(n_141),
.B2(n_146),
.Y(n_1182)
);

OAI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_895),
.A2(n_148),
.B1(n_159),
.B2(n_953),
.Y(n_1183)
);

HB1xp67_ASAP7_75t_L g1184 ( 
.A(n_1026),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_973),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_1024),
.B(n_991),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_999),
.B(n_973),
.Y(n_1187)
);

AO31x2_ASAP7_75t_L g1188 ( 
.A1(n_1084),
.A2(n_1018),
.A3(n_853),
.B(n_1010),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_SL g1189 ( 
.A1(n_1159),
.A2(n_984),
.B(n_985),
.Y(n_1189)
);

AOI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_1067),
.A2(n_894),
.B1(n_978),
.B2(n_979),
.Y(n_1190)
);

AOI21xp33_ASAP7_75t_L g1191 ( 
.A1(n_1052),
.A2(n_952),
.B(n_941),
.Y(n_1191)
);

OAI22x1_ASAP7_75t_L g1192 ( 
.A1(n_1157),
.A2(n_992),
.B1(n_1013),
.B2(n_895),
.Y(n_1192)
);

O2A1O1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_1070),
.A2(n_993),
.B(n_1016),
.C(n_874),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1168),
.A2(n_970),
.B(n_971),
.Y(n_1194)
);

AO31x2_ASAP7_75t_L g1195 ( 
.A1(n_1122),
.A2(n_1011),
.A3(n_910),
.B(n_909),
.Y(n_1195)
);

INVx8_ASAP7_75t_L g1196 ( 
.A(n_1044),
.Y(n_1196)
);

AOI221x1_ASAP7_75t_L g1197 ( 
.A1(n_1182),
.A2(n_872),
.B1(n_903),
.B2(n_869),
.C(n_960),
.Y(n_1197)
);

OAI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1083),
.A2(n_1159),
.B(n_1055),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1063),
.B(n_884),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_1092),
.A2(n_955),
.B(n_947),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1097),
.A2(n_939),
.B(n_930),
.Y(n_1201)
);

INVx3_ASAP7_75t_L g1202 ( 
.A(n_1053),
.Y(n_1202)
);

O2A1O1Ixp5_ASAP7_75t_L g1203 ( 
.A1(n_1083),
.A2(n_998),
.B(n_1014),
.C(n_956),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1042),
.B(n_943),
.Y(n_1204)
);

NAND3xp33_ASAP7_75t_SL g1205 ( 
.A(n_1066),
.B(n_912),
.C(n_914),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1098),
.B(n_860),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1099),
.A2(n_923),
.B(n_865),
.Y(n_1207)
);

OAI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1048),
.A2(n_1008),
.B(n_1004),
.Y(n_1208)
);

OA21x2_ASAP7_75t_L g1209 ( 
.A1(n_1169),
.A2(n_1006),
.B(n_995),
.Y(n_1209)
);

AOI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1090),
.A2(n_996),
.B(n_1073),
.Y(n_1210)
);

NAND3xp33_ASAP7_75t_L g1211 ( 
.A(n_1163),
.B(n_1106),
.C(n_1114),
.Y(n_1211)
);

AOI221x1_ASAP7_75t_L g1212 ( 
.A1(n_1182),
.A2(n_1177),
.B1(n_1183),
.B2(n_1122),
.C(n_1157),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1169),
.A2(n_1040),
.B(n_1065),
.Y(n_1213)
);

OAI22x1_ASAP7_75t_L g1214 ( 
.A1(n_1117),
.A2(n_1050),
.B1(n_1161),
.B2(n_1043),
.Y(n_1214)
);

AOI22x1_ASAP7_75t_SL g1215 ( 
.A1(n_1034),
.A2(n_1105),
.B1(n_1142),
.B2(n_1152),
.Y(n_1215)
);

OAI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1058),
.A2(n_1076),
.B(n_1148),
.Y(n_1216)
);

NAND3xp33_ASAP7_75t_L g1217 ( 
.A(n_1164),
.B(n_1079),
.C(n_1076),
.Y(n_1217)
);

OAI22x1_ASAP7_75t_L g1218 ( 
.A1(n_1117),
.A2(n_1043),
.B1(n_1037),
.B2(n_1080),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1160),
.A2(n_1180),
.B(n_1094),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1094),
.A2(n_1186),
.B(n_1090),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1103),
.A2(n_1112),
.B(n_1132),
.Y(n_1221)
);

AO21x1_ASAP7_75t_L g1222 ( 
.A1(n_1177),
.A2(n_1183),
.B(n_1187),
.Y(n_1222)
);

AO32x2_ASAP7_75t_L g1223 ( 
.A1(n_1087),
.A2(n_1166),
.A3(n_1074),
.B1(n_1107),
.B2(n_1047),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1091),
.A2(n_1104),
.B(n_1085),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1081),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1185),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1103),
.A2(n_1132),
.B(n_1112),
.Y(n_1227)
);

OAI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1104),
.A2(n_1041),
.B(n_1061),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1088),
.A2(n_1089),
.B(n_1095),
.Y(n_1229)
);

NOR2xp67_ASAP7_75t_L g1230 ( 
.A(n_1147),
.B(n_1075),
.Y(n_1230)
);

OAI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1134),
.A2(n_1039),
.B(n_1113),
.Y(n_1231)
);

NOR2xp67_ASAP7_75t_L g1232 ( 
.A(n_1101),
.B(n_1110),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1039),
.A2(n_1102),
.B(n_1095),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1137),
.A2(n_1057),
.B(n_1172),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1088),
.A2(n_1089),
.B(n_1176),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1125),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1111),
.B(n_1137),
.Y(n_1237)
);

AND2x4_ASAP7_75t_L g1238 ( 
.A(n_1087),
.B(n_1037),
.Y(n_1238)
);

AO22x1_ASAP7_75t_L g1239 ( 
.A1(n_1165),
.A2(n_1060),
.B1(n_1109),
.B2(n_1068),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1057),
.A2(n_1046),
.B(n_1154),
.Y(n_1240)
);

A2O1A1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_1051),
.A2(n_1121),
.B(n_1049),
.C(n_1162),
.Y(n_1241)
);

O2A1O1Ixp33_ASAP7_75t_SL g1242 ( 
.A1(n_1135),
.A2(n_1156),
.B(n_1062),
.C(n_1136),
.Y(n_1242)
);

INVx4_ASAP7_75t_L g1243 ( 
.A(n_1056),
.Y(n_1243)
);

HB1xp67_ASAP7_75t_L g1244 ( 
.A(n_1153),
.Y(n_1244)
);

AO31x2_ASAP7_75t_L g1245 ( 
.A1(n_1166),
.A2(n_1155),
.A3(n_1175),
.B(n_1179),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1111),
.B(n_1064),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1128),
.A2(n_1149),
.B(n_1071),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1086),
.A2(n_1151),
.B(n_1119),
.Y(n_1248)
);

NOR2xp33_ASAP7_75t_L g1249 ( 
.A(n_1033),
.B(n_1096),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_L g1250 ( 
.A(n_1060),
.B(n_1181),
.Y(n_1250)
);

INVx5_ASAP7_75t_L g1251 ( 
.A(n_1118),
.Y(n_1251)
);

NAND2x1p5_ASAP7_75t_L g1252 ( 
.A(n_1072),
.B(n_1074),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1093),
.A2(n_1072),
.B(n_1078),
.Y(n_1253)
);

CKINVDCx6p67_ASAP7_75t_R g1254 ( 
.A(n_1100),
.Y(n_1254)
);

INVxp67_ASAP7_75t_SL g1255 ( 
.A(n_1167),
.Y(n_1255)
);

INVxp67_ASAP7_75t_L g1256 ( 
.A(n_1165),
.Y(n_1256)
);

INVx1_ASAP7_75t_SL g1257 ( 
.A(n_1146),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_1047),
.B(n_1045),
.Y(n_1258)
);

A2O1A1Ixp33_ASAP7_75t_L g1259 ( 
.A1(n_1135),
.A2(n_1138),
.B(n_1127),
.C(n_1059),
.Y(n_1259)
);

BUFx10_ASAP7_75t_L g1260 ( 
.A(n_1053),
.Y(n_1260)
);

INVx3_ASAP7_75t_L g1261 ( 
.A(n_1053),
.Y(n_1261)
);

INVxp67_ASAP7_75t_L g1262 ( 
.A(n_1184),
.Y(n_1262)
);

AO31x2_ASAP7_75t_L g1263 ( 
.A1(n_1035),
.A2(n_1036),
.A3(n_1145),
.B(n_1116),
.Y(n_1263)
);

AND2x6_ASAP7_75t_L g1264 ( 
.A(n_1129),
.B(n_1158),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_SL g1265 ( 
.A(n_1143),
.B(n_1144),
.Y(n_1265)
);

OAI21xp5_ASAP7_75t_SL g1266 ( 
.A1(n_1069),
.A2(n_1139),
.B(n_1140),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1143),
.A2(n_1144),
.B(n_1118),
.Y(n_1267)
);

AOI221xp5_ASAP7_75t_L g1268 ( 
.A1(n_1108),
.A2(n_1150),
.B1(n_1130),
.B2(n_1133),
.C(n_1120),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1171),
.Y(n_1269)
);

NOR2xp67_ASAP7_75t_L g1270 ( 
.A(n_1115),
.B(n_1131),
.Y(n_1270)
);

AO31x2_ASAP7_75t_L g1271 ( 
.A1(n_1173),
.A2(n_1178),
.A3(n_1126),
.B(n_1141),
.Y(n_1271)
);

AOI31xp67_ASAP7_75t_L g1272 ( 
.A1(n_1170),
.A2(n_1038),
.A3(n_1174),
.B(n_1077),
.Y(n_1272)
);

CKINVDCx8_ASAP7_75t_R g1273 ( 
.A(n_1045),
.Y(n_1273)
);

BUFx2_ASAP7_75t_L g1274 ( 
.A(n_1045),
.Y(n_1274)
);

AO21x1_ASAP7_75t_L g1275 ( 
.A1(n_1038),
.A2(n_1118),
.B(n_1082),
.Y(n_1275)
);

NOR2xp33_ASAP7_75t_L g1276 ( 
.A(n_1158),
.B(n_1077),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1077),
.A2(n_1082),
.B(n_1123),
.Y(n_1277)
);

AO31x2_ASAP7_75t_L g1278 ( 
.A1(n_1038),
.A2(n_1082),
.A3(n_1123),
.B(n_1124),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1123),
.A2(n_1131),
.B(n_1124),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1038),
.A2(n_1124),
.B(n_1131),
.Y(n_1280)
);

OA21x2_ASAP7_75t_L g1281 ( 
.A1(n_1097),
.A2(n_1092),
.B(n_1169),
.Y(n_1281)
);

INVxp67_ASAP7_75t_SL g1282 ( 
.A(n_1042),
.Y(n_1282)
);

CKINVDCx6p67_ASAP7_75t_R g1283 ( 
.A(n_1034),
.Y(n_1283)
);

OAI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1070),
.A2(n_744),
.B1(n_729),
.B2(n_731),
.Y(n_1284)
);

OAI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1070),
.A2(n_744),
.B1(n_729),
.B2(n_731),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1070),
.A2(n_601),
.B(n_1168),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1070),
.A2(n_601),
.B(n_1168),
.Y(n_1287)
);

AOI221xp5_ASAP7_75t_SL g1288 ( 
.A1(n_1163),
.A2(n_729),
.B1(n_731),
.B2(n_744),
.C(n_1076),
.Y(n_1288)
);

BUFx2_ASAP7_75t_SL g1289 ( 
.A(n_1105),
.Y(n_1289)
);

NOR2x1_ASAP7_75t_R g1290 ( 
.A(n_1044),
.B(n_697),
.Y(n_1290)
);

NAND3xp33_ASAP7_75t_L g1291 ( 
.A(n_1066),
.B(n_729),
.C(n_731),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1097),
.A2(n_1092),
.B(n_1099),
.Y(n_1292)
);

INVx5_ASAP7_75t_L g1293 ( 
.A(n_1118),
.Y(n_1293)
);

OAI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1070),
.A2(n_744),
.B(n_685),
.Y(n_1294)
);

A2O1A1Ixp33_ASAP7_75t_L g1295 ( 
.A1(n_1159),
.A2(n_731),
.B(n_729),
.C(n_744),
.Y(n_1295)
);

NOR3xp33_ASAP7_75t_L g1296 ( 
.A(n_1163),
.B(n_731),
.C(n_729),
.Y(n_1296)
);

NAND3xp33_ASAP7_75t_L g1297 ( 
.A(n_1066),
.B(n_729),
.C(n_731),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_SL g1298 ( 
.A(n_1055),
.B(n_957),
.Y(n_1298)
);

CKINVDCx20_ASAP7_75t_R g1299 ( 
.A(n_1044),
.Y(n_1299)
);

AOI221x1_ASAP7_75t_L g1300 ( 
.A1(n_1182),
.A2(n_1159),
.B1(n_1177),
.B2(n_1083),
.C(n_1183),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1070),
.A2(n_601),
.B(n_1168),
.Y(n_1301)
);

AOI22xp5_ASAP7_75t_L g1302 ( 
.A1(n_1067),
.A2(n_731),
.B1(n_729),
.B2(n_881),
.Y(n_1302)
);

AOI221xp5_ASAP7_75t_L g1303 ( 
.A1(n_1076),
.A2(n_731),
.B1(n_729),
.B2(n_623),
.C(n_599),
.Y(n_1303)
);

BUFx2_ASAP7_75t_L g1304 ( 
.A(n_1056),
.Y(n_1304)
);

OAI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1070),
.A2(n_744),
.B(n_685),
.Y(n_1305)
);

CKINVDCx11_ASAP7_75t_R g1306 ( 
.A(n_1105),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1067),
.B(n_731),
.Y(n_1307)
);

AO31x2_ASAP7_75t_L g1308 ( 
.A1(n_1084),
.A2(n_1018),
.A3(n_859),
.B(n_1122),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1185),
.Y(n_1309)
);

BUFx10_ASAP7_75t_L g1310 ( 
.A(n_1044),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1070),
.A2(n_601),
.B(n_1168),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1097),
.A2(n_1092),
.B(n_1099),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_L g1313 ( 
.A(n_1067),
.B(n_731),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1185),
.Y(n_1314)
);

CKINVDCx6p67_ASAP7_75t_R g1315 ( 
.A(n_1034),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1054),
.Y(n_1316)
);

INVxp67_ASAP7_75t_SL g1317 ( 
.A(n_1042),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1067),
.B(n_731),
.Y(n_1318)
);

INVx2_ASAP7_75t_SL g1319 ( 
.A(n_1165),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1070),
.A2(n_601),
.B(n_1168),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1185),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1147),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1067),
.B(n_731),
.Y(n_1323)
);

OAI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1070),
.A2(n_744),
.B(n_685),
.Y(n_1324)
);

OAI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1070),
.A2(n_744),
.B(n_685),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1147),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1067),
.B(n_731),
.Y(n_1327)
);

INVx1_ASAP7_75t_SL g1328 ( 
.A(n_1111),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1185),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1097),
.A2(n_1092),
.B(n_1099),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1097),
.A2(n_1092),
.B(n_1099),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_SL g1332 ( 
.A(n_1055),
.B(n_957),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1070),
.A2(n_601),
.B(n_1168),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1070),
.A2(n_601),
.B(n_1168),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1087),
.B(n_1037),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_SL g1336 ( 
.A1(n_1159),
.A2(n_1039),
.B(n_1046),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1070),
.A2(n_601),
.B(n_1168),
.Y(n_1337)
);

AOI221x1_ASAP7_75t_L g1338 ( 
.A1(n_1182),
.A2(n_1159),
.B1(n_1177),
.B2(n_1083),
.C(n_1183),
.Y(n_1338)
);

OR2x6_ASAP7_75t_L g1339 ( 
.A(n_1045),
.B(n_852),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1185),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1070),
.A2(n_601),
.B(n_1168),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1070),
.A2(n_601),
.B(n_1168),
.Y(n_1342)
);

AO31x2_ASAP7_75t_L g1343 ( 
.A1(n_1084),
.A2(n_1018),
.A3(n_859),
.B(n_1122),
.Y(n_1343)
);

INVxp67_ASAP7_75t_L g1344 ( 
.A(n_1075),
.Y(n_1344)
);

OR2x6_ASAP7_75t_L g1345 ( 
.A(n_1045),
.B(n_852),
.Y(n_1345)
);

A2O1A1Ixp33_ASAP7_75t_L g1346 ( 
.A1(n_1159),
.A2(n_731),
.B(n_729),
.C(n_744),
.Y(n_1346)
);

O2A1O1Ixp33_ASAP7_75t_SL g1347 ( 
.A1(n_1070),
.A2(n_957),
.B(n_964),
.C(n_1104),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_1044),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1097),
.A2(n_1092),
.B(n_1099),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1185),
.Y(n_1350)
);

CKINVDCx20_ASAP7_75t_R g1351 ( 
.A(n_1299),
.Y(n_1351)
);

CKINVDCx11_ASAP7_75t_R g1352 ( 
.A(n_1310),
.Y(n_1352)
);

NAND2xp5_ASAP7_75t_L g1353 ( 
.A(n_1237),
.B(n_1313),
.Y(n_1353)
);

INVx3_ASAP7_75t_L g1354 ( 
.A(n_1260),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1263),
.Y(n_1355)
);

OAI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1212),
.A2(n_1338),
.B1(n_1300),
.B2(n_1216),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1222),
.A2(n_1211),
.B1(n_1198),
.B2(n_1303),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1296),
.A2(n_1217),
.B1(n_1214),
.B2(n_1258),
.Y(n_1358)
);

INVx1_ASAP7_75t_SL g1359 ( 
.A(n_1257),
.Y(n_1359)
);

INVx4_ASAP7_75t_SL g1360 ( 
.A(n_1264),
.Y(n_1360)
);

BUFx10_ASAP7_75t_L g1361 ( 
.A(n_1348),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1224),
.A2(n_1218),
.B1(n_1269),
.B2(n_1297),
.Y(n_1362)
);

OAI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1295),
.A2(n_1346),
.B1(n_1302),
.B2(n_1266),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1284),
.A2(n_1285),
.B1(n_1294),
.B2(n_1325),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1307),
.B(n_1318),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1305),
.A2(n_1324),
.B1(n_1336),
.B2(n_1291),
.Y(n_1366)
);

AOI22xp5_ASAP7_75t_SL g1367 ( 
.A1(n_1239),
.A2(n_1250),
.B1(n_1256),
.B2(n_1319),
.Y(n_1367)
);

INVx8_ASAP7_75t_L g1368 ( 
.A(n_1264),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1231),
.A2(n_1189),
.B1(n_1327),
.B2(n_1323),
.Y(n_1369)
);

OAI22xp33_ASAP7_75t_L g1370 ( 
.A1(n_1190),
.A2(n_1251),
.B1(n_1293),
.B2(n_1282),
.Y(n_1370)
);

AND2x4_ASAP7_75t_L g1371 ( 
.A(n_1238),
.B(n_1335),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1236),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_SL g1373 ( 
.A1(n_1251),
.A2(n_1293),
.B1(n_1199),
.B2(n_1317),
.Y(n_1373)
);

BUFx2_ASAP7_75t_L g1374 ( 
.A(n_1243),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1322),
.A2(n_1326),
.B1(n_1298),
.B2(n_1332),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_1306),
.Y(n_1376)
);

INVx6_ASAP7_75t_L g1377 ( 
.A(n_1243),
.Y(n_1377)
);

HB1xp67_ASAP7_75t_L g1378 ( 
.A(n_1281),
.Y(n_1378)
);

CKINVDCx6p67_ASAP7_75t_R g1379 ( 
.A(n_1196),
.Y(n_1379)
);

BUFx2_ASAP7_75t_L g1380 ( 
.A(n_1339),
.Y(n_1380)
);

OAI22xp5_ASAP7_75t_L g1381 ( 
.A1(n_1241),
.A2(n_1259),
.B1(n_1344),
.B2(n_1228),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1275),
.A2(n_1225),
.B1(n_1316),
.B2(n_1253),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1226),
.A2(n_1350),
.B1(n_1329),
.B2(n_1321),
.Y(n_1383)
);

BUFx6f_ASAP7_75t_L g1384 ( 
.A(n_1264),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1309),
.A2(n_1350),
.B1(n_1340),
.B2(n_1329),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_1196),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_1283),
.Y(n_1387)
);

CKINVDCx11_ASAP7_75t_R g1388 ( 
.A(n_1310),
.Y(n_1388)
);

OAI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1251),
.A2(n_1293),
.B1(n_1246),
.B2(n_1206),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1314),
.Y(n_1390)
);

CKINVDCx16_ASAP7_75t_R g1391 ( 
.A(n_1215),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1244),
.B(n_1289),
.Y(n_1392)
);

BUFx12f_ASAP7_75t_L g1393 ( 
.A(n_1339),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1321),
.Y(n_1394)
);

BUFx10_ASAP7_75t_L g1395 ( 
.A(n_1249),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1340),
.A2(n_1328),
.B1(n_1264),
.B2(n_1274),
.Y(n_1396)
);

OAI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1213),
.A2(n_1345),
.B1(n_1230),
.B2(n_1240),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1245),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_SL g1399 ( 
.A1(n_1223),
.A2(n_1234),
.B1(n_1288),
.B2(n_1335),
.Y(n_1399)
);

BUFx6f_ASAP7_75t_L g1400 ( 
.A(n_1280),
.Y(n_1400)
);

OAI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1345),
.A2(n_1273),
.B1(n_1315),
.B2(n_1232),
.Y(n_1401)
);

CKINVDCx11_ASAP7_75t_R g1402 ( 
.A(n_1254),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1191),
.A2(n_1268),
.B1(n_1192),
.B2(n_1262),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1245),
.Y(n_1404)
);

BUFx2_ASAP7_75t_SL g1405 ( 
.A(n_1270),
.Y(n_1405)
);

CKINVDCx11_ASAP7_75t_R g1406 ( 
.A(n_1260),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1233),
.A2(n_1204),
.B1(n_1247),
.B2(n_1255),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1223),
.B(n_1252),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1286),
.A2(n_1334),
.B1(n_1342),
.B2(n_1287),
.Y(n_1409)
);

AOI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1242),
.A2(n_1276),
.B1(n_1265),
.B2(n_1267),
.Y(n_1410)
);

AOI22xp33_ASAP7_75t_SL g1411 ( 
.A1(n_1223),
.A2(n_1301),
.B1(n_1337),
.B2(n_1311),
.Y(n_1411)
);

CKINVDCx20_ASAP7_75t_R g1412 ( 
.A(n_1290),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1271),
.Y(n_1413)
);

BUFx10_ASAP7_75t_L g1414 ( 
.A(n_1202),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1261),
.B(n_1278),
.Y(n_1415)
);

BUFx12f_ASAP7_75t_L g1416 ( 
.A(n_1278),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1205),
.A2(n_1221),
.B1(n_1227),
.B2(n_1220),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1209),
.A2(n_1341),
.B1(n_1333),
.B2(n_1320),
.Y(n_1418)
);

BUFx12f_ASAP7_75t_L g1419 ( 
.A(n_1277),
.Y(n_1419)
);

INVx6_ASAP7_75t_L g1420 ( 
.A(n_1279),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1347),
.Y(n_1421)
);

NAND2x1p5_ASAP7_75t_L g1422 ( 
.A(n_1229),
.B(n_1235),
.Y(n_1422)
);

NAND2xp33_ASAP7_75t_SL g1423 ( 
.A(n_1208),
.B(n_1272),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1248),
.Y(n_1424)
);

INVx6_ASAP7_75t_L g1425 ( 
.A(n_1281),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_SL g1426 ( 
.A1(n_1209),
.A2(n_1219),
.B1(n_1308),
.B2(n_1343),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1207),
.A2(n_1200),
.B1(n_1194),
.B2(n_1201),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1308),
.A2(n_1343),
.B1(n_1193),
.B2(n_1349),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1343),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_SL g1430 ( 
.A1(n_1308),
.A2(n_1203),
.B1(n_1197),
.B2(n_1188),
.Y(n_1430)
);

AOI22xp33_ASAP7_75t_L g1431 ( 
.A1(n_1331),
.A2(n_1292),
.B1(n_1312),
.B2(n_1330),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_SL g1432 ( 
.A1(n_1188),
.A2(n_1047),
.B1(n_1216),
.B2(n_1157),
.Y(n_1432)
);

INVx1_ASAP7_75t_SL g1433 ( 
.A(n_1195),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1210),
.A2(n_1295),
.B1(n_1346),
.B2(n_1216),
.Y(n_1434)
);

AOI22xp5_ASAP7_75t_SL g1435 ( 
.A1(n_1195),
.A2(n_1047),
.B1(n_556),
.B2(n_608),
.Y(n_1435)
);

AOI22x1_ASAP7_75t_L g1436 ( 
.A1(n_1195),
.A2(n_1305),
.B1(n_1324),
.B2(n_1294),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_1348),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1313),
.B(n_1067),
.Y(n_1438)
);

BUFx12f_ASAP7_75t_L g1439 ( 
.A(n_1306),
.Y(n_1439)
);

OAI21xp5_ASAP7_75t_L g1440 ( 
.A1(n_1216),
.A2(n_744),
.B(n_729),
.Y(n_1440)
);

BUFx4f_ASAP7_75t_SL g1441 ( 
.A(n_1299),
.Y(n_1441)
);

INVx4_ASAP7_75t_L g1442 ( 
.A(n_1306),
.Y(n_1442)
);

CKINVDCx11_ASAP7_75t_R g1443 ( 
.A(n_1299),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1216),
.A2(n_1047),
.B1(n_890),
.B2(n_1222),
.Y(n_1444)
);

CKINVDCx16_ASAP7_75t_R g1445 ( 
.A(n_1299),
.Y(n_1445)
);

INVx6_ASAP7_75t_L g1446 ( 
.A(n_1243),
.Y(n_1446)
);

INVx5_ASAP7_75t_L g1447 ( 
.A(n_1264),
.Y(n_1447)
);

INVx4_ASAP7_75t_L g1448 ( 
.A(n_1306),
.Y(n_1448)
);

INVx1_ASAP7_75t_SL g1449 ( 
.A(n_1304),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1216),
.A2(n_1047),
.B1(n_890),
.B2(n_1222),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1237),
.B(n_1313),
.Y(n_1451)
);

NAND2x1p5_ASAP7_75t_L g1452 ( 
.A(n_1251),
.B(n_1293),
.Y(n_1452)
);

OAI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1212),
.A2(n_1338),
.B1(n_1300),
.B2(n_1216),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1216),
.A2(n_1047),
.B1(n_890),
.B2(n_1222),
.Y(n_1454)
);

CKINVDCx5p33_ASAP7_75t_R g1455 ( 
.A(n_1348),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1216),
.A2(n_1047),
.B1(n_890),
.B2(n_1222),
.Y(n_1456)
);

CKINVDCx11_ASAP7_75t_R g1457 ( 
.A(n_1299),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_SL g1458 ( 
.A1(n_1216),
.A2(n_1047),
.B1(n_1157),
.B2(n_364),
.Y(n_1458)
);

AOI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1303),
.A2(n_623),
.B1(n_731),
.B2(n_729),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1216),
.A2(n_1047),
.B1(n_890),
.B2(n_1222),
.Y(n_1460)
);

BUFx2_ASAP7_75t_SL g1461 ( 
.A(n_1299),
.Y(n_1461)
);

OAI21xp33_ASAP7_75t_L g1462 ( 
.A1(n_1303),
.A2(n_1216),
.B(n_1295),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1216),
.A2(n_798),
.B1(n_1047),
.B2(n_890),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1216),
.A2(n_798),
.B1(n_1047),
.B2(n_890),
.Y(n_1464)
);

OAI22xp5_ASAP7_75t_SL g1465 ( 
.A1(n_1291),
.A2(n_913),
.B1(n_731),
.B2(n_556),
.Y(n_1465)
);

HB1xp67_ASAP7_75t_L g1466 ( 
.A(n_1281),
.Y(n_1466)
);

INVx6_ASAP7_75t_L g1467 ( 
.A(n_1243),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1216),
.A2(n_1047),
.B1(n_890),
.B2(n_1222),
.Y(n_1468)
);

BUFx8_ASAP7_75t_SL g1469 ( 
.A(n_1299),
.Y(n_1469)
);

CKINVDCx9p33_ASAP7_75t_R g1470 ( 
.A(n_1215),
.Y(n_1470)
);

NAND2x1p5_ASAP7_75t_L g1471 ( 
.A(n_1251),
.B(n_1293),
.Y(n_1471)
);

BUFx6f_ASAP7_75t_L g1472 ( 
.A(n_1264),
.Y(n_1472)
);

INVx3_ASAP7_75t_L g1473 ( 
.A(n_1425),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1355),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1394),
.Y(n_1475)
);

AOI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1434),
.A2(n_1409),
.B(n_1378),
.Y(n_1476)
);

INVx3_ASAP7_75t_L g1477 ( 
.A(n_1425),
.Y(n_1477)
);

CKINVDCx20_ASAP7_75t_R g1478 ( 
.A(n_1469),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1390),
.B(n_1415),
.Y(n_1479)
);

OAI21x1_ASAP7_75t_L g1480 ( 
.A1(n_1427),
.A2(n_1431),
.B(n_1422),
.Y(n_1480)
);

INVx1_ASAP7_75t_SL g1481 ( 
.A(n_1359),
.Y(n_1481)
);

HB1xp67_ASAP7_75t_L g1482 ( 
.A(n_1381),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1378),
.B(n_1466),
.Y(n_1483)
);

BUFx6f_ASAP7_75t_L g1484 ( 
.A(n_1447),
.Y(n_1484)
);

AOI21x1_ASAP7_75t_L g1485 ( 
.A1(n_1466),
.A2(n_1363),
.B(n_1421),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1398),
.Y(n_1486)
);

INVx2_ASAP7_75t_SL g1487 ( 
.A(n_1377),
.Y(n_1487)
);

AND2x4_ASAP7_75t_L g1488 ( 
.A(n_1360),
.B(n_1447),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1426),
.B(n_1429),
.Y(n_1489)
);

AO21x2_ASAP7_75t_L g1490 ( 
.A1(n_1356),
.A2(n_1453),
.B(n_1404),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_1443),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1353),
.B(n_1451),
.Y(n_1492)
);

OR2x6_ASAP7_75t_L g1493 ( 
.A(n_1368),
.B(n_1384),
.Y(n_1493)
);

HB1xp67_ASAP7_75t_L g1494 ( 
.A(n_1449),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1372),
.Y(n_1495)
);

INVxp67_ASAP7_75t_L g1496 ( 
.A(n_1438),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1413),
.Y(n_1497)
);

OAI21x1_ASAP7_75t_L g1498 ( 
.A1(n_1431),
.A2(n_1422),
.B(n_1418),
.Y(n_1498)
);

OR2x6_ASAP7_75t_L g1499 ( 
.A(n_1368),
.B(n_1472),
.Y(n_1499)
);

INVx3_ASAP7_75t_L g1500 ( 
.A(n_1420),
.Y(n_1500)
);

INVx4_ASAP7_75t_L g1501 ( 
.A(n_1360),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1426),
.B(n_1428),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1375),
.Y(n_1503)
);

AOI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1462),
.A2(n_1458),
.B1(n_1454),
.B2(n_1468),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1383),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1365),
.B(n_1441),
.Y(n_1506)
);

INVx2_ASAP7_75t_SL g1507 ( 
.A(n_1377),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1385),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1428),
.B(n_1430),
.Y(n_1509)
);

BUFx2_ASAP7_75t_L g1510 ( 
.A(n_1424),
.Y(n_1510)
);

HB1xp67_ASAP7_75t_L g1511 ( 
.A(n_1375),
.Y(n_1511)
);

BUFx2_ASAP7_75t_L g1512 ( 
.A(n_1423),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1430),
.B(n_1432),
.Y(n_1513)
);

BUFx2_ASAP7_75t_L g1514 ( 
.A(n_1416),
.Y(n_1514)
);

OAI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1357),
.A2(n_1459),
.B1(n_1364),
.B2(n_1444),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1432),
.B(n_1369),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1369),
.B(n_1408),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1433),
.B(n_1411),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1411),
.B(n_1357),
.Y(n_1519)
);

OAI21x1_ASAP7_75t_L g1520 ( 
.A1(n_1417),
.A2(n_1436),
.B(n_1407),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1400),
.Y(n_1521)
);

INVx1_ASAP7_75t_SL g1522 ( 
.A(n_1395),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1392),
.B(n_1399),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1356),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1453),
.Y(n_1525)
);

AND2x2_ASAP7_75t_L g1526 ( 
.A(n_1399),
.B(n_1366),
.Y(n_1526)
);

AND2x4_ASAP7_75t_L g1527 ( 
.A(n_1360),
.B(n_1472),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1389),
.Y(n_1528)
);

HB1xp67_ASAP7_75t_L g1529 ( 
.A(n_1374),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1389),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1397),
.Y(n_1531)
);

AO21x2_ASAP7_75t_L g1532 ( 
.A1(n_1370),
.A2(n_1397),
.B(n_1410),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1458),
.A2(n_1463),
.B1(n_1464),
.B2(n_1460),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1366),
.B(n_1358),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1370),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1444),
.B(n_1450),
.Y(n_1536)
);

AO21x2_ASAP7_75t_L g1537 ( 
.A1(n_1440),
.A2(n_1401),
.B(n_1435),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1382),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1403),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1419),
.Y(n_1540)
);

BUFx2_ASAP7_75t_SL g1541 ( 
.A(n_1395),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1450),
.B(n_1468),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1454),
.B(n_1460),
.Y(n_1543)
);

OAI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1456),
.A2(n_1362),
.B1(n_1465),
.B2(n_1391),
.Y(n_1544)
);

OAI21x1_ASAP7_75t_L g1545 ( 
.A1(n_1452),
.A2(n_1471),
.B(n_1456),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1373),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1373),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1414),
.Y(n_1548)
);

OAI21x1_ASAP7_75t_L g1549 ( 
.A1(n_1452),
.A2(n_1396),
.B(n_1354),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1380),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1354),
.Y(n_1551)
);

OA21x2_ASAP7_75t_L g1552 ( 
.A1(n_1371),
.A2(n_1401),
.B(n_1387),
.Y(n_1552)
);

INVx2_ASAP7_75t_SL g1553 ( 
.A(n_1446),
.Y(n_1553)
);

INVx3_ASAP7_75t_L g1554 ( 
.A(n_1446),
.Y(n_1554)
);

AND2x4_ASAP7_75t_L g1555 ( 
.A(n_1479),
.B(n_1442),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1517),
.B(n_1367),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1524),
.B(n_1467),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_SL g1558 ( 
.A(n_1515),
.B(n_1393),
.Y(n_1558)
);

AO32x2_ASAP7_75t_L g1559 ( 
.A1(n_1544),
.A2(n_1448),
.A3(n_1442),
.B1(n_1470),
.B2(n_1467),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1524),
.B(n_1467),
.Y(n_1560)
);

OAI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1504),
.A2(n_1445),
.B1(n_1441),
.B2(n_1376),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1475),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1475),
.Y(n_1563)
);

OAI21xp5_ASAP7_75t_L g1564 ( 
.A1(n_1482),
.A2(n_1412),
.B(n_1351),
.Y(n_1564)
);

AND2x4_ASAP7_75t_L g1565 ( 
.A(n_1473),
.B(n_1386),
.Y(n_1565)
);

AND2x6_ASAP7_75t_L g1566 ( 
.A(n_1488),
.B(n_1470),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1496),
.B(n_1461),
.Y(n_1567)
);

AOI21xp5_ASAP7_75t_SL g1568 ( 
.A1(n_1552),
.A2(n_1455),
.B(n_1437),
.Y(n_1568)
);

INVx1_ASAP7_75t_SL g1569 ( 
.A(n_1541),
.Y(n_1569)
);

OAI211xp5_ASAP7_75t_L g1570 ( 
.A1(n_1504),
.A2(n_1519),
.B(n_1533),
.C(n_1526),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_SL g1571 ( 
.A(n_1519),
.B(n_1361),
.Y(n_1571)
);

A2O1A1Ixp33_ASAP7_75t_L g1572 ( 
.A1(n_1536),
.A2(n_1405),
.B(n_1402),
.C(n_1406),
.Y(n_1572)
);

OR2x6_ASAP7_75t_L g1573 ( 
.A(n_1488),
.B(n_1439),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1495),
.B(n_1379),
.Y(n_1574)
);

AND2x4_ASAP7_75t_L g1575 ( 
.A(n_1473),
.B(n_1352),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_1491),
.Y(n_1576)
);

NAND2x1_ASAP7_75t_L g1577 ( 
.A(n_1554),
.B(n_1388),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1523),
.B(n_1457),
.Y(n_1578)
);

A2O1A1Ixp33_ASAP7_75t_L g1579 ( 
.A1(n_1536),
.A2(n_1542),
.B(n_1516),
.C(n_1526),
.Y(n_1579)
);

OAI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1542),
.A2(n_1543),
.B1(n_1539),
.B2(n_1516),
.Y(n_1580)
);

AO32x2_ASAP7_75t_L g1581 ( 
.A1(n_1487),
.A2(n_1507),
.A3(n_1553),
.B1(n_1511),
.B2(n_1503),
.Y(n_1581)
);

NOR2xp33_ASAP7_75t_L g1582 ( 
.A(n_1534),
.B(n_1522),
.Y(n_1582)
);

OA21x2_ASAP7_75t_L g1583 ( 
.A1(n_1520),
.A2(n_1480),
.B(n_1498),
.Y(n_1583)
);

AOI21xp5_ASAP7_75t_SL g1584 ( 
.A1(n_1552),
.A2(n_1488),
.B(n_1532),
.Y(n_1584)
);

AO32x2_ASAP7_75t_L g1585 ( 
.A1(n_1487),
.A2(n_1553),
.A3(n_1507),
.B1(n_1490),
.B2(n_1501),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1529),
.B(n_1550),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1494),
.B(n_1506),
.Y(n_1587)
);

AOI21xp5_ASAP7_75t_L g1588 ( 
.A1(n_1532),
.A2(n_1531),
.B(n_1512),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1509),
.B(n_1502),
.Y(n_1589)
);

NOR2xp33_ASAP7_75t_L g1590 ( 
.A(n_1534),
.B(n_1541),
.Y(n_1590)
);

A2O1A1Ixp33_ASAP7_75t_L g1591 ( 
.A1(n_1513),
.A2(n_1539),
.B(n_1525),
.C(n_1518),
.Y(n_1591)
);

AO32x2_ASAP7_75t_L g1592 ( 
.A1(n_1490),
.A2(n_1501),
.A3(n_1525),
.B1(n_1513),
.B2(n_1483),
.Y(n_1592)
);

AO32x2_ASAP7_75t_L g1593 ( 
.A1(n_1490),
.A2(n_1501),
.A3(n_1483),
.B1(n_1489),
.B2(n_1505),
.Y(n_1593)
);

OA21x2_ASAP7_75t_L g1594 ( 
.A1(n_1476),
.A2(n_1530),
.B(n_1528),
.Y(n_1594)
);

NOR2xp33_ASAP7_75t_L g1595 ( 
.A(n_1485),
.B(n_1537),
.Y(n_1595)
);

BUFx12f_ASAP7_75t_L g1596 ( 
.A(n_1478),
.Y(n_1596)
);

AND2x4_ASAP7_75t_L g1597 ( 
.A(n_1473),
.B(n_1477),
.Y(n_1597)
);

OAI22xp5_ASAP7_75t_SL g1598 ( 
.A1(n_1552),
.A2(n_1540),
.B1(n_1492),
.B2(n_1481),
.Y(n_1598)
);

OAI21xp33_ASAP7_75t_L g1599 ( 
.A1(n_1485),
.A2(n_1476),
.B(n_1489),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1505),
.B(n_1508),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1497),
.Y(n_1601)
);

AND2x4_ASAP7_75t_L g1602 ( 
.A(n_1477),
.B(n_1514),
.Y(n_1602)
);

NOR2xp67_ASAP7_75t_SL g1603 ( 
.A(n_1484),
.B(n_1552),
.Y(n_1603)
);

HB1xp67_ASAP7_75t_L g1604 ( 
.A(n_1510),
.Y(n_1604)
);

OAI21x1_ASAP7_75t_L g1605 ( 
.A1(n_1545),
.A2(n_1549),
.B(n_1500),
.Y(n_1605)
);

O2A1O1Ixp33_ASAP7_75t_L g1606 ( 
.A1(n_1537),
.A2(n_1538),
.B(n_1528),
.C(n_1530),
.Y(n_1606)
);

A2O1A1Ixp33_ASAP7_75t_L g1607 ( 
.A1(n_1535),
.A2(n_1547),
.B(n_1546),
.C(n_1538),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1601),
.Y(n_1608)
);

INVx2_ASAP7_75t_L g1609 ( 
.A(n_1594),
.Y(n_1609)
);

HB1xp67_ASAP7_75t_L g1610 ( 
.A(n_1604),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1562),
.Y(n_1611)
);

INVxp67_ASAP7_75t_SL g1612 ( 
.A(n_1604),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1583),
.B(n_1521),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1588),
.B(n_1589),
.Y(n_1614)
);

BUFx2_ASAP7_75t_L g1615 ( 
.A(n_1585),
.Y(n_1615)
);

BUFx2_ASAP7_75t_L g1616 ( 
.A(n_1585),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1563),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_SL g1618 ( 
.A1(n_1570),
.A2(n_1537),
.B1(n_1546),
.B2(n_1547),
.Y(n_1618)
);

BUFx2_ASAP7_75t_L g1619 ( 
.A(n_1585),
.Y(n_1619)
);

AND2x4_ASAP7_75t_L g1620 ( 
.A(n_1597),
.B(n_1605),
.Y(n_1620)
);

INVxp67_ASAP7_75t_L g1621 ( 
.A(n_1590),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1586),
.B(n_1486),
.Y(n_1622)
);

AOI22xp33_ASAP7_75t_L g1623 ( 
.A1(n_1580),
.A2(n_1527),
.B1(n_1499),
.B2(n_1493),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1593),
.B(n_1592),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1592),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1592),
.Y(n_1626)
);

BUFx2_ASAP7_75t_L g1627 ( 
.A(n_1581),
.Y(n_1627)
);

BUFx2_ASAP7_75t_L g1628 ( 
.A(n_1581),
.Y(n_1628)
);

OAI22xp33_ASAP7_75t_L g1629 ( 
.A1(n_1558),
.A2(n_1561),
.B1(n_1580),
.B2(n_1582),
.Y(n_1629)
);

INVx1_ASAP7_75t_SL g1630 ( 
.A(n_1569),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1581),
.B(n_1474),
.Y(n_1631)
);

NAND3xp33_ASAP7_75t_L g1632 ( 
.A(n_1558),
.B(n_1551),
.C(n_1548),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1617),
.Y(n_1633)
);

INVx3_ASAP7_75t_L g1634 ( 
.A(n_1620),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1617),
.Y(n_1635)
);

BUFx2_ASAP7_75t_L g1636 ( 
.A(n_1610),
.Y(n_1636)
);

OAI31xp33_ASAP7_75t_L g1637 ( 
.A1(n_1629),
.A2(n_1570),
.A3(n_1579),
.B(n_1591),
.Y(n_1637)
);

BUFx3_ASAP7_75t_L g1638 ( 
.A(n_1630),
.Y(n_1638)
);

INVx5_ASAP7_75t_SL g1639 ( 
.A(n_1620),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1621),
.B(n_1555),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1608),
.Y(n_1641)
);

NAND3xp33_ASAP7_75t_L g1642 ( 
.A(n_1618),
.B(n_1561),
.C(n_1595),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1608),
.Y(n_1643)
);

A2O1A1Ixp33_ASAP7_75t_SL g1644 ( 
.A1(n_1612),
.A2(n_1548),
.B(n_1590),
.C(n_1564),
.Y(n_1644)
);

INVx3_ASAP7_75t_L g1645 ( 
.A(n_1620),
.Y(n_1645)
);

OAI33xp33_ASAP7_75t_L g1646 ( 
.A1(n_1629),
.A2(n_1606),
.A3(n_1598),
.B1(n_1599),
.B2(n_1560),
.B3(n_1557),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1608),
.Y(n_1647)
);

AOI33xp33_ASAP7_75t_L g1648 ( 
.A1(n_1624),
.A2(n_1578),
.A3(n_1587),
.B1(n_1569),
.B2(n_1606),
.B3(n_1556),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1621),
.B(n_1602),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1611),
.Y(n_1650)
);

OAI21xp33_ASAP7_75t_SL g1651 ( 
.A1(n_1624),
.A2(n_1568),
.B(n_1571),
.Y(n_1651)
);

INVx4_ASAP7_75t_L g1652 ( 
.A(n_1620),
.Y(n_1652)
);

AO22x1_ASAP7_75t_L g1653 ( 
.A1(n_1624),
.A2(n_1566),
.B1(n_1595),
.B2(n_1582),
.Y(n_1653)
);

NAND3xp33_ASAP7_75t_SL g1654 ( 
.A(n_1627),
.B(n_1564),
.C(n_1579),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1614),
.B(n_1557),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1611),
.Y(n_1656)
);

AND2x4_ASAP7_75t_L g1657 ( 
.A(n_1620),
.B(n_1573),
.Y(n_1657)
);

AO21x2_ASAP7_75t_L g1658 ( 
.A1(n_1609),
.A2(n_1591),
.B(n_1607),
.Y(n_1658)
);

AO21x2_ASAP7_75t_L g1659 ( 
.A1(n_1609),
.A2(n_1607),
.B(n_1560),
.Y(n_1659)
);

OAI31xp33_ASAP7_75t_L g1660 ( 
.A1(n_1627),
.A2(n_1572),
.A3(n_1559),
.B(n_1571),
.Y(n_1660)
);

OAI221xp5_ASAP7_75t_L g1661 ( 
.A1(n_1618),
.A2(n_1572),
.B1(n_1584),
.B2(n_1603),
.C(n_1574),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1614),
.B(n_1622),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1614),
.B(n_1600),
.Y(n_1663)
);

NAND4xp25_ASAP7_75t_L g1664 ( 
.A(n_1630),
.B(n_1567),
.C(n_1551),
.D(n_1565),
.Y(n_1664)
);

AND2x4_ASAP7_75t_L g1665 ( 
.A(n_1620),
.B(n_1573),
.Y(n_1665)
);

HB1xp67_ASAP7_75t_L g1666 ( 
.A(n_1610),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1639),
.B(n_1627),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1639),
.B(n_1628),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1662),
.B(n_1628),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1639),
.B(n_1652),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1662),
.B(n_1628),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1641),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1643),
.B(n_1631),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1643),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1639),
.B(n_1615),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1652),
.B(n_1615),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1652),
.B(n_1615),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1647),
.B(n_1631),
.Y(n_1678)
);

NAND2x1_ASAP7_75t_L g1679 ( 
.A(n_1657),
.B(n_1616),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1655),
.B(n_1625),
.Y(n_1680)
);

INVx3_ASAP7_75t_L g1681 ( 
.A(n_1652),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1645),
.B(n_1616),
.Y(n_1682)
);

OR2x2_ASAP7_75t_L g1683 ( 
.A(n_1655),
.B(n_1636),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1647),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1650),
.B(n_1631),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1650),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_SL g1687 ( 
.A(n_1651),
.B(n_1632),
.Y(n_1687)
);

AND2x4_ASAP7_75t_L g1688 ( 
.A(n_1645),
.B(n_1613),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1645),
.B(n_1616),
.Y(n_1689)
);

INVx3_ASAP7_75t_L g1690 ( 
.A(n_1645),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1656),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1658),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1658),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1634),
.B(n_1619),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1658),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1634),
.B(n_1619),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1674),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1674),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1670),
.B(n_1657),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1674),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1684),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1669),
.B(n_1654),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1684),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1670),
.B(n_1657),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1670),
.B(n_1657),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1667),
.B(n_1665),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1669),
.B(n_1666),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1683),
.B(n_1648),
.Y(n_1708)
);

HB1xp67_ASAP7_75t_L g1709 ( 
.A(n_1683),
.Y(n_1709)
);

INVxp67_ASAP7_75t_L g1710 ( 
.A(n_1687),
.Y(n_1710)
);

NAND2x1p5_ASAP7_75t_L g1711 ( 
.A(n_1687),
.B(n_1638),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1667),
.B(n_1665),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1667),
.B(n_1665),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1672),
.B(n_1660),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1668),
.B(n_1665),
.Y(n_1715)
);

NOR2xp33_ASAP7_75t_L g1716 ( 
.A(n_1683),
.B(n_1596),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1668),
.B(n_1634),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1672),
.B(n_1636),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1692),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1684),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1679),
.B(n_1576),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1668),
.B(n_1649),
.Y(n_1722)
);

INVxp67_ASAP7_75t_L g1723 ( 
.A(n_1675),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1669),
.B(n_1663),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1692),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1686),
.B(n_1633),
.Y(n_1726)
);

INVx1_ASAP7_75t_SL g1727 ( 
.A(n_1675),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1691),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1692),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1671),
.B(n_1663),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1686),
.B(n_1635),
.Y(n_1731)
);

AOI21xp5_ASAP7_75t_L g1732 ( 
.A1(n_1679),
.A2(n_1646),
.B(n_1642),
.Y(n_1732)
);

OAI21xp33_ASAP7_75t_L g1733 ( 
.A1(n_1676),
.A2(n_1642),
.B(n_1651),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1692),
.Y(n_1734)
);

OAI22xp5_ASAP7_75t_L g1735 ( 
.A1(n_1679),
.A2(n_1632),
.B1(n_1661),
.B2(n_1623),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1691),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1675),
.B(n_1649),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1676),
.B(n_1640),
.Y(n_1738)
);

AND2x2_ASAP7_75t_SL g1739 ( 
.A(n_1676),
.B(n_1619),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_1709),
.B(n_1671),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1710),
.B(n_1677),
.Y(n_1741)
);

OAI21xp33_ASAP7_75t_L g1742 ( 
.A1(n_1733),
.A2(n_1677),
.B(n_1682),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1697),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1711),
.B(n_1677),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1697),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1732),
.B(n_1673),
.Y(n_1746)
);

OR2x2_ASAP7_75t_L g1747 ( 
.A(n_1724),
.B(n_1680),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1739),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1698),
.Y(n_1749)
);

AND2x4_ASAP7_75t_SL g1750 ( 
.A(n_1716),
.B(n_1573),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1708),
.B(n_1673),
.Y(n_1751)
);

AOI211x1_ASAP7_75t_L g1752 ( 
.A1(n_1733),
.A2(n_1653),
.B(n_1664),
.C(n_1689),
.Y(n_1752)
);

OR2x2_ASAP7_75t_L g1753 ( 
.A(n_1724),
.B(n_1730),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1714),
.B(n_1678),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1711),
.B(n_1682),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1714),
.B(n_1678),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1730),
.B(n_1680),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1698),
.Y(n_1758)
);

OAI21xp33_ASAP7_75t_L g1759 ( 
.A1(n_1711),
.A2(n_1689),
.B(n_1682),
.Y(n_1759)
);

NOR2xp33_ASAP7_75t_SL g1760 ( 
.A(n_1721),
.B(n_1637),
.Y(n_1760)
);

NOR2xp33_ASAP7_75t_L g1761 ( 
.A(n_1723),
.B(n_1640),
.Y(n_1761)
);

NOR2xp33_ASAP7_75t_L g1762 ( 
.A(n_1727),
.B(n_1638),
.Y(n_1762)
);

INVx1_ASAP7_75t_SL g1763 ( 
.A(n_1727),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1700),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1700),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1702),
.B(n_1685),
.Y(n_1766)
);

HB1xp67_ASAP7_75t_L g1767 ( 
.A(n_1707),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1739),
.B(n_1689),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1702),
.B(n_1685),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1739),
.B(n_1694),
.Y(n_1770)
);

INVx1_ASAP7_75t_SL g1771 ( 
.A(n_1722),
.Y(n_1771)
);

INVx1_ASAP7_75t_SL g1772 ( 
.A(n_1722),
.Y(n_1772)
);

HB1xp67_ASAP7_75t_L g1773 ( 
.A(n_1707),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1719),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1718),
.B(n_1680),
.Y(n_1775)
);

AOI22x1_ASAP7_75t_L g1776 ( 
.A1(n_1748),
.A2(n_1705),
.B1(n_1704),
.B2(n_1699),
.Y(n_1776)
);

AOI22xp33_ASAP7_75t_L g1777 ( 
.A1(n_1746),
.A2(n_1693),
.B1(n_1695),
.B2(n_1625),
.Y(n_1777)
);

INVxp67_ASAP7_75t_L g1778 ( 
.A(n_1767),
.Y(n_1778)
);

HB1xp67_ASAP7_75t_L g1779 ( 
.A(n_1773),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1744),
.B(n_1737),
.Y(n_1780)
);

NAND3xp33_ASAP7_75t_L g1781 ( 
.A(n_1752),
.B(n_1735),
.C(n_1703),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1747),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1745),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1745),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1749),
.Y(n_1785)
);

OR2x2_ASAP7_75t_L g1786 ( 
.A(n_1753),
.B(n_1718),
.Y(n_1786)
);

NAND2xp5_ASAP7_75t_SL g1787 ( 
.A(n_1760),
.B(n_1742),
.Y(n_1787)
);

AOI21xp33_ASAP7_75t_SL g1788 ( 
.A1(n_1762),
.A2(n_1735),
.B(n_1737),
.Y(n_1788)
);

AOI21xp5_ASAP7_75t_L g1789 ( 
.A1(n_1754),
.A2(n_1644),
.B(n_1693),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1749),
.Y(n_1790)
);

NOR2x1_ASAP7_75t_L g1791 ( 
.A(n_1763),
.B(n_1681),
.Y(n_1791)
);

AOI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1756),
.A2(n_1625),
.B1(n_1626),
.B2(n_1659),
.Y(n_1792)
);

AOI22xp33_ASAP7_75t_L g1793 ( 
.A1(n_1751),
.A2(n_1695),
.B1(n_1693),
.B2(n_1625),
.Y(n_1793)
);

INVx3_ASAP7_75t_L g1794 ( 
.A(n_1768),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1747),
.Y(n_1795)
);

OAI22xp5_ASAP7_75t_SL g1796 ( 
.A1(n_1748),
.A2(n_1577),
.B1(n_1575),
.B2(n_1688),
.Y(n_1796)
);

NAND2x1_ASAP7_75t_L g1797 ( 
.A(n_1744),
.B(n_1699),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1771),
.B(n_1738),
.Y(n_1798)
);

BUFx2_ASAP7_75t_L g1799 ( 
.A(n_1753),
.Y(n_1799)
);

OR2x2_ASAP7_75t_L g1800 ( 
.A(n_1740),
.B(n_1701),
.Y(n_1800)
);

INVxp67_ASAP7_75t_L g1801 ( 
.A(n_1741),
.Y(n_1801)
);

OAI221xp5_ASAP7_75t_L g1802 ( 
.A1(n_1781),
.A2(n_1759),
.B1(n_1769),
.B2(n_1766),
.C(n_1770),
.Y(n_1802)
);

OR2x2_ASAP7_75t_L g1803 ( 
.A(n_1799),
.B(n_1772),
.Y(n_1803)
);

OAI32xp33_ASAP7_75t_L g1804 ( 
.A1(n_1787),
.A2(n_1768),
.A3(n_1755),
.B1(n_1770),
.B2(n_1740),
.Y(n_1804)
);

INVx1_ASAP7_75t_SL g1805 ( 
.A(n_1799),
.Y(n_1805)
);

NAND3xp33_ASAP7_75t_SL g1806 ( 
.A(n_1788),
.B(n_1755),
.C(n_1757),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1780),
.B(n_1750),
.Y(n_1807)
);

O2A1O1Ixp33_ASAP7_75t_L g1808 ( 
.A1(n_1787),
.A2(n_1775),
.B(n_1764),
.C(n_1774),
.Y(n_1808)
);

OAI22xp33_ASAP7_75t_L g1809 ( 
.A1(n_1792),
.A2(n_1626),
.B1(n_1757),
.B2(n_1775),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_L g1810 ( 
.A1(n_1777),
.A2(n_1693),
.B1(n_1695),
.B2(n_1774),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1779),
.Y(n_1811)
);

O2A1O1Ixp33_ASAP7_75t_R g1812 ( 
.A1(n_1786),
.A2(n_1695),
.B(n_1626),
.C(n_1726),
.Y(n_1812)
);

AOI211xp5_ASAP7_75t_L g1813 ( 
.A1(n_1789),
.A2(n_1764),
.B(n_1765),
.C(n_1758),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1780),
.B(n_1750),
.Y(n_1814)
);

OAI211xp5_ASAP7_75t_SL g1815 ( 
.A1(n_1801),
.A2(n_1743),
.B(n_1761),
.C(n_1681),
.Y(n_1815)
);

NAND2x1_ASAP7_75t_L g1816 ( 
.A(n_1791),
.B(n_1706),
.Y(n_1816)
);

NOR2xp33_ASAP7_75t_L g1817 ( 
.A(n_1778),
.B(n_1706),
.Y(n_1817)
);

OAI22xp5_ASAP7_75t_L g1818 ( 
.A1(n_1776),
.A2(n_1738),
.B1(n_1694),
.B2(n_1696),
.Y(n_1818)
);

NOR3xp33_ASAP7_75t_L g1819 ( 
.A(n_1794),
.B(n_1725),
.C(n_1719),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1794),
.B(n_1704),
.Y(n_1820)
);

NAND3xp33_ASAP7_75t_L g1821 ( 
.A(n_1794),
.B(n_1703),
.C(n_1701),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1803),
.Y(n_1822)
);

INVx3_ASAP7_75t_L g1823 ( 
.A(n_1816),
.Y(n_1823)
);

INVxp33_ASAP7_75t_L g1824 ( 
.A(n_1811),
.Y(n_1824)
);

AOI22xp33_ASAP7_75t_L g1825 ( 
.A1(n_1806),
.A2(n_1795),
.B1(n_1782),
.B2(n_1793),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1805),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1821),
.Y(n_1827)
);

AOI21xp5_ASAP7_75t_L g1828 ( 
.A1(n_1808),
.A2(n_1797),
.B(n_1795),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1820),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1817),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1813),
.B(n_1782),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1819),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1807),
.Y(n_1833)
);

NOR2x1_ASAP7_75t_L g1834 ( 
.A(n_1826),
.B(n_1797),
.Y(n_1834)
);

NOR2xp33_ASAP7_75t_L g1835 ( 
.A(n_1824),
.B(n_1814),
.Y(n_1835)
);

AOI22xp33_ASAP7_75t_L g1836 ( 
.A1(n_1825),
.A2(n_1809),
.B1(n_1810),
.B2(n_1802),
.Y(n_1836)
);

NOR4xp25_ASAP7_75t_L g1837 ( 
.A(n_1831),
.B(n_1802),
.C(n_1815),
.D(n_1783),
.Y(n_1837)
);

OR2x2_ASAP7_75t_L g1838 ( 
.A(n_1822),
.B(n_1786),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1829),
.B(n_1798),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1833),
.B(n_1804),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1830),
.B(n_1800),
.Y(n_1841)
);

INVxp67_ASAP7_75t_L g1842 ( 
.A(n_1823),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1823),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1832),
.Y(n_1844)
);

NAND2xp5_ASAP7_75t_L g1845 ( 
.A(n_1835),
.B(n_1828),
.Y(n_1845)
);

OAI211xp5_ASAP7_75t_L g1846 ( 
.A1(n_1837),
.A2(n_1825),
.B(n_1827),
.C(n_1785),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1843),
.B(n_1824),
.Y(n_1847)
);

OAI222xp33_ASAP7_75t_L g1848 ( 
.A1(n_1836),
.A2(n_1812),
.B1(n_1800),
.B2(n_1784),
.C1(n_1790),
.C2(n_1818),
.Y(n_1848)
);

AOI211xp5_ASAP7_75t_L g1849 ( 
.A1(n_1840),
.A2(n_1796),
.B(n_1818),
.C(n_1712),
.Y(n_1849)
);

AOI221xp5_ASAP7_75t_L g1850 ( 
.A1(n_1844),
.A2(n_1725),
.B1(n_1734),
.B2(n_1729),
.C(n_1719),
.Y(n_1850)
);

NOR3xp33_ASAP7_75t_L g1851 ( 
.A(n_1846),
.B(n_1842),
.C(n_1841),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1845),
.B(n_1834),
.Y(n_1852)
);

OAI21xp33_ASAP7_75t_SL g1853 ( 
.A1(n_1847),
.A2(n_1838),
.B(n_1839),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1849),
.B(n_1712),
.Y(n_1854)
);

AOI221xp5_ASAP7_75t_L g1855 ( 
.A1(n_1848),
.A2(n_1725),
.B1(n_1734),
.B2(n_1729),
.C(n_1626),
.Y(n_1855)
);

AOI221xp5_ASAP7_75t_L g1856 ( 
.A1(n_1850),
.A2(n_1734),
.B1(n_1729),
.B2(n_1736),
.C(n_1728),
.Y(n_1856)
);

XNOR2xp5_ASAP7_75t_L g1857 ( 
.A(n_1851),
.B(n_1713),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1853),
.Y(n_1858)
);

INVxp67_ASAP7_75t_SL g1859 ( 
.A(n_1852),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1854),
.Y(n_1860)
);

AND2x4_ASAP7_75t_L g1861 ( 
.A(n_1855),
.B(n_1713),
.Y(n_1861)
);

OR2x2_ASAP7_75t_L g1862 ( 
.A(n_1858),
.B(n_1859),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1859),
.B(n_1856),
.Y(n_1863)
);

NAND2x1p5_ASAP7_75t_L g1864 ( 
.A(n_1860),
.B(n_1715),
.Y(n_1864)
);

OAI22xp5_ASAP7_75t_SL g1865 ( 
.A1(n_1862),
.A2(n_1857),
.B1(n_1861),
.B2(n_1736),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1865),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1866),
.B(n_1864),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1866),
.Y(n_1868)
);

AO21x1_ASAP7_75t_L g1869 ( 
.A1(n_1867),
.A2(n_1863),
.B(n_1868),
.Y(n_1869)
);

OAI22xp5_ASAP7_75t_SL g1870 ( 
.A1(n_1867),
.A2(n_1861),
.B1(n_1728),
.B2(n_1720),
.Y(n_1870)
);

AOI21xp5_ASAP7_75t_L g1871 ( 
.A1(n_1869),
.A2(n_1870),
.B(n_1720),
.Y(n_1871)
);

OA21x2_ASAP7_75t_L g1872 ( 
.A1(n_1871),
.A2(n_1715),
.B(n_1717),
.Y(n_1872)
);

OAI211xp5_ASAP7_75t_L g1873 ( 
.A1(n_1872),
.A2(n_1705),
.B(n_1717),
.C(n_1681),
.Y(n_1873)
);

OAI22xp33_ASAP7_75t_L g1874 ( 
.A1(n_1873),
.A2(n_1731),
.B1(n_1726),
.B2(n_1690),
.Y(n_1874)
);

OAI221xp5_ASAP7_75t_R g1875 ( 
.A1(n_1874),
.A2(n_1681),
.B1(n_1690),
.B2(n_1688),
.C(n_1731),
.Y(n_1875)
);

AOI211xp5_ASAP7_75t_L g1876 ( 
.A1(n_1875),
.A2(n_1575),
.B(n_1694),
.C(n_1696),
.Y(n_1876)
);


endmodule