module fake_jpeg_22308_n_139 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_139);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_139;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_96;

BUFx12_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx11_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_11),
.B(n_10),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_4),
.B(n_6),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_7),
.B(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_30),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_23),
.B(n_1),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_31),
.B(n_32),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_1),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_37),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_21),
.B(n_2),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_25),
.Y(n_38)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_38),
.Y(n_43)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_39),
.A2(n_22),
.B1(n_15),
.B2(n_28),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_2),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_2),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_33),
.A2(n_22),
.B1(n_15),
.B2(n_26),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_46),
.A2(n_51),
.B1(n_39),
.B2(n_36),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_32),
.B(n_27),
.Y(n_47)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

FAx1_ASAP7_75t_SL g48 ( 
.A(n_30),
.B(n_27),
.CI(n_26),
.CON(n_48),
.SN(n_48)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_48),
.B(n_19),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_37),
.B(n_29),
.Y(n_50)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_33),
.A2(n_22),
.B1(n_24),
.B2(n_19),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_34),
.B(n_21),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_54),
.B(n_29),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_55),
.B(n_56),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_52),
.B(n_17),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_62),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_54),
.B(n_14),
.Y(n_59)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_61),
.A2(n_67),
.B1(n_71),
.B2(n_72),
.Y(n_76)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_63),
.B(n_65),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_52),
.B(n_48),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_44),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_70),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_14),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_68),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_44),
.Y(n_69)
);

INVx4_ASAP7_75t_SL g80 ( 
.A(n_69),
.Y(n_80)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_62),
.A2(n_64),
.B1(n_57),
.B2(n_60),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_73),
.A2(n_83),
.B1(n_38),
.B2(n_45),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_49),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_47),
.C(n_50),
.Y(n_92)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_79),
.Y(n_93)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_82),
.B(n_85),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_64),
.A2(n_36),
.B1(n_39),
.B2(n_53),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_R g85 ( 
.A1(n_57),
.A2(n_49),
.B1(n_41),
.B2(n_30),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

OAI21xp33_ASAP7_75t_L g89 ( 
.A1(n_81),
.A2(n_84),
.B(n_88),
.Y(n_89)
);

NAND3xp33_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_99),
.C(n_101),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_76),
.A2(n_53),
.B1(n_60),
.B2(n_34),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_76),
.A2(n_53),
.B1(n_35),
.B2(n_43),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_91),
.B(n_94),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_92),
.B(n_41),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_73),
.A2(n_35),
.B1(n_43),
.B2(n_72),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_45),
.C(n_30),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_99),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_101),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_67),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_74),
.A2(n_30),
.B(n_38),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_92),
.Y(n_113)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

AO21x1_ASAP7_75t_L g117 ( 
.A1(n_105),
.A2(n_106),
.B(n_109),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_93),
.Y(n_106)
);

NOR3xp33_ASAP7_75t_SL g107 ( 
.A(n_96),
.B(n_78),
.C(n_87),
.Y(n_107)
);

NAND3xp33_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_110),
.C(n_112),
.Y(n_114)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_115),
.Y(n_121)
);

OAI32xp33_ASAP7_75t_L g115 ( 
.A1(n_108),
.A2(n_90),
.A3(n_91),
.B1(n_98),
.B2(n_83),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_102),
.A2(n_111),
.B(n_103),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_116),
.A2(n_119),
.B1(n_80),
.B2(n_104),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_118),
.B(n_120),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_102),
.A2(n_95),
.B(n_100),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_107),
.A2(n_16),
.B(n_24),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_117),
.A2(n_79),
.B1(n_80),
.B2(n_86),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_125),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_124),
.B(n_126),
.Y(n_127)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

NOR3xp33_ASAP7_75t_SL g126 ( 
.A(n_120),
.B(n_16),
.C(n_82),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_77),
.C(n_44),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_128),
.B(n_126),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_122),
.B(n_3),
.Y(n_130)
);

AOI31xp67_ASAP7_75t_L g134 ( 
.A1(n_130),
.A2(n_8),
.A3(n_12),
.B(n_13),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_129),
.B(n_123),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_132),
.Y(n_136)
);

NOR2xp67_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_3),
.Y(n_133)
);

AOI322xp5_ASAP7_75t_L g135 ( 
.A1(n_133),
.A2(n_134),
.A3(n_130),
.B1(n_13),
.B2(n_12),
.C1(n_25),
.C2(n_18),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_135),
.B(n_25),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_137),
.B(n_138),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_136),
.B(n_18),
.C(n_35),
.Y(n_138)
);


endmodule