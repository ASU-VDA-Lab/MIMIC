module fake_netlist_6_3462_n_15 (n_4, n_2, n_3, n_5, n_1, n_0, n_15);

input n_4;
input n_2;
input n_3;
input n_5;
input n_1;
input n_0;

output n_15;

wire n_7;
wire n_6;
wire n_12;
wire n_14;
wire n_13;
wire n_9;
wire n_11;
wire n_8;
wire n_10;

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_4),
.Y(n_6)
);

CKINVDCx5p33_ASAP7_75t_R g7 ( 
.A(n_5),
.Y(n_7)
);

NOR2xp33_ASAP7_75t_L g8 ( 
.A(n_2),
.B(n_0),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

HB1xp67_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_12),
.B(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

AO221x2_ASAP7_75t_L g15 ( 
.A1(n_14),
.A2(n_11),
.B1(n_9),
.B2(n_6),
.C(n_3),
.Y(n_15)
);


endmodule