module fake_jpeg_26615_n_134 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_134);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_134;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_9),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_7),
.B(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_5),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_29),
.Y(n_37)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_32),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_12),
.Y(n_32)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_21),
.Y(n_33)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_34),
.A2(n_18),
.B1(n_19),
.B2(n_17),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_18),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_35),
.B(n_39),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_27),
.B(n_25),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_36),
.B(n_13),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_18),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_0),
.B(n_1),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_34),
.A2(n_18),
.B1(n_20),
.B2(n_17),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_43),
.A2(n_32),
.B1(n_28),
.B2(n_31),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_18),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_20),
.Y(n_58)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_30),
.B(n_19),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_46),
.A2(n_15),
.B(n_13),
.Y(n_51)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_34),
.B1(n_28),
.B2(n_31),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_48),
.A2(n_57),
.B1(n_46),
.B2(n_40),
.Y(n_76)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_51),
.A2(n_59),
.B(n_46),
.Y(n_65)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_58),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_53),
.A2(n_56),
.B1(n_38),
.B2(n_22),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_55),
.B(n_60),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_22),
.B1(n_26),
.B2(n_16),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_37),
.A2(n_30),
.B1(n_14),
.B2(n_24),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_35),
.B(n_37),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_41),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_62),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_59),
.A2(n_46),
.B(n_44),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_63),
.A2(n_14),
.B(n_16),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_65),
.A2(n_69),
.B(n_51),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_52),
.A2(n_58),
.B1(n_59),
.B2(n_54),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_66),
.A2(n_67),
.B1(n_72),
.B2(n_77),
.Y(n_85)
);

NAND3xp33_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_36),
.C(n_44),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_47),
.A2(n_15),
.B1(n_26),
.B2(n_23),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_54),
.B(n_58),
.Y(n_73)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_76),
.A2(n_50),
.B1(n_48),
.B2(n_56),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_48),
.A2(n_40),
.B1(n_45),
.B2(n_23),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_80),
.A2(n_86),
.B1(n_83),
.B2(n_84),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_67),
.Y(n_96)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_88),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_60),
.C(n_57),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_86),
.C(n_90),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_57),
.C(n_45),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_65),
.A2(n_51),
.B(n_24),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_89),
.A2(n_91),
.B(n_70),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_53),
.C(n_61),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_90),
.B(n_66),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_92),
.A2(n_0),
.B(n_40),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_87),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_94),
.B(n_99),
.Y(n_111)
);

A2O1A1O1Ixp25_ASAP7_75t_L g95 ( 
.A1(n_81),
.A2(n_63),
.B(n_70),
.C(n_76),
.D(n_71),
.Y(n_95)
);

AOI221xp5_ASAP7_75t_L g105 ( 
.A1(n_95),
.A2(n_97),
.B1(n_20),
.B2(n_47),
.C(n_49),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_98),
.Y(n_108)
);

OAI322xp33_ASAP7_75t_L g98 ( 
.A1(n_89),
.A2(n_71),
.A3(n_33),
.B1(n_77),
.B2(n_78),
.C1(n_64),
.C2(n_49),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_78),
.Y(n_100)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_100),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_93),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_103),
.B(n_104),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_100),
.A2(n_85),
.B1(n_91),
.B2(n_82),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_109),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_101),
.Y(n_107)
);

AOI21x1_ASAP7_75t_L g113 ( 
.A1(n_107),
.A2(n_88),
.B(n_47),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_49),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_92),
.C(n_102),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_114),
.Y(n_120)
);

AOI321xp33_ASAP7_75t_L g114 ( 
.A1(n_108),
.A2(n_97),
.A3(n_95),
.B1(n_102),
.B2(n_92),
.C(n_96),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_115),
.B(n_111),
.C(n_109),
.Y(n_119)
);

AOI321xp33_ASAP7_75t_L g117 ( 
.A1(n_108),
.A2(n_7),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C(n_6),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_118),
.Y(n_123)
);

AOI321xp33_ASAP7_75t_L g118 ( 
.A1(n_104),
.A2(n_7),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C(n_6),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_119),
.B(n_8),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_112),
.A2(n_106),
.B(n_107),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g126 ( 
.A1(n_121),
.A2(n_4),
.B(n_8),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_106),
.C(n_41),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_122),
.B(n_116),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_124),
.B(n_125),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_120),
.A2(n_62),
.B1(n_41),
.B2(n_0),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_126),
.A2(n_127),
.B(n_123),
.Y(n_128)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_128),
.Y(n_131)
);

AOI31xp67_ASAP7_75t_SL g129 ( 
.A1(n_125),
.A2(n_8),
.A3(n_10),
.B(n_11),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_129),
.A2(n_0),
.B(n_62),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_132),
.B(n_130),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_133),
.B(n_131),
.Y(n_134)
);


endmodule