module fake_jpeg_30977_n_542 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_542);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_542;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx4f_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_30),
.B(n_9),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_54),
.B(n_82),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

HAxp5_ASAP7_75t_SL g58 ( 
.A(n_34),
.B(n_17),
.CON(n_58),
.SN(n_58)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_58),
.B(n_50),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_61),
.Y(n_121)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_62),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_63),
.Y(n_149)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_64),
.Y(n_137)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_25),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_65),
.B(n_77),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx3_ASAP7_75t_SL g134 ( 
.A(n_66),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_67),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_68),
.Y(n_163)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_72),
.Y(n_144)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_73),
.Y(n_120)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_74),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_76),
.Y(n_168)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_78),
.Y(n_133)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_79),
.Y(n_122)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_80),
.Y(n_147)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_81),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_30),
.B(n_8),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_83),
.Y(n_141)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_25),
.Y(n_84)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_84),
.Y(n_169)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_85),
.Y(n_159)
);

BUFx10_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_86),
.Y(n_117)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_87),
.Y(n_132)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_88),
.Y(n_162)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_90),
.Y(n_127)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_44),
.Y(n_92)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_92),
.Y(n_135)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_93),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_94),
.B(n_103),
.Y(n_139)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_95),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_96),
.Y(n_143)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_97),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g164 ( 
.A(n_98),
.Y(n_164)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_99),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_23),
.Y(n_100)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_100),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_23),
.Y(n_101)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_101),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_29),
.Y(n_102)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_102),
.Y(n_148)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_34),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_26),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_104),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_23),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_106),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_23),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_98),
.A2(n_35),
.B1(n_51),
.B2(n_43),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_115),
.A2(n_138),
.B1(n_157),
.B2(n_39),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_65),
.B(n_35),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_118),
.B(n_123),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_69),
.B(n_51),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_102),
.A2(n_20),
.B1(n_49),
.B2(n_34),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_125),
.A2(n_31),
.B1(n_1),
.B2(n_2),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_43),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_130),
.B(n_140),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_55),
.A2(n_59),
.B1(n_90),
.B2(n_71),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_42),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_105),
.B(n_42),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_142),
.B(n_150),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_58),
.A2(n_38),
.B1(n_32),
.B2(n_40),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_145),
.B(n_167),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_106),
.B(n_53),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_76),
.B(n_21),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_166),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_63),
.A2(n_32),
.B1(n_21),
.B2(n_40),
.Y(n_157)
);

BUFx12_ASAP7_75t_L g165 ( 
.A(n_61),
.Y(n_165)
);

BUFx16f_ASAP7_75t_L g207 ( 
.A(n_165),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_61),
.B(n_53),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_164),
.A2(n_26),
.B1(n_27),
.B2(n_20),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_170),
.Y(n_228)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_121),
.Y(n_171)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_171),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_113),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_172),
.B(n_200),
.Y(n_247)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_144),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_173),
.Y(n_235)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_131),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_174),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_114),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_175),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_114),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_176),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_164),
.A2(n_27),
.B1(n_20),
.B2(n_94),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_177),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_141),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_179),
.B(n_185),
.Y(n_253)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_112),
.Y(n_180)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_180),
.Y(n_241)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_107),
.Y(n_181)
);

INVx5_ASAP7_75t_L g259 ( 
.A(n_181),
.Y(n_259)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_148),
.Y(n_182)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_182),
.Y(n_246)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_124),
.Y(n_183)
);

INVx13_ASAP7_75t_L g249 ( 
.A(n_183),
.Y(n_249)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_116),
.Y(n_184)
);

INVx8_ASAP7_75t_L g238 ( 
.A(n_184),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_167),
.A2(n_96),
.B1(n_68),
.B2(n_67),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_186),
.A2(n_203),
.B1(n_108),
.B2(n_127),
.Y(n_236)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_116),
.Y(n_187)
);

INVx8_ASAP7_75t_L g245 ( 
.A(n_187),
.Y(n_245)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_131),
.Y(n_188)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_188),
.Y(n_254)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_120),
.Y(n_189)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_189),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_153),
.A2(n_20),
.B1(n_94),
.B2(n_77),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_191),
.A2(n_206),
.B1(n_217),
.B2(n_218),
.Y(n_240)
);

AND2x2_ASAP7_75t_SL g192 ( 
.A(n_109),
.B(n_0),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_192),
.B(n_195),
.C(n_202),
.Y(n_230)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_159),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_194),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_162),
.B(n_103),
.C(n_34),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_149),
.Y(n_197)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_197),
.Y(n_251)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_124),
.Y(n_198)
);

INVx13_ASAP7_75t_L g266 ( 
.A(n_198),
.Y(n_266)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_119),
.Y(n_199)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_199),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_158),
.B(n_39),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_158),
.B(n_24),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_201),
.B(n_212),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_139),
.B(n_129),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_155),
.A2(n_49),
.B1(n_24),
.B2(n_19),
.Y(n_203)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_168),
.Y(n_204)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_204),
.Y(n_233)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_168),
.Y(n_205)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_205),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_132),
.A2(n_77),
.B1(n_49),
.B2(n_50),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_155),
.A2(n_49),
.B1(n_19),
.B2(n_37),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_208),
.A2(n_216),
.B1(n_219),
.B2(n_134),
.Y(n_239)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_151),
.Y(n_209)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_209),
.Y(n_267)
);

OAI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_128),
.A2(n_49),
.B1(n_19),
.B2(n_86),
.Y(n_210)
);

OAI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_210),
.A2(n_161),
.B1(n_160),
.B2(n_152),
.Y(n_260)
);

NAND2x1_ASAP7_75t_L g211 ( 
.A(n_125),
.B(n_31),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_211),
.B(n_214),
.Y(n_234)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_169),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_122),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_213),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_137),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_139),
.B(n_50),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_222),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_111),
.A2(n_31),
.B1(n_37),
.B2(n_86),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_147),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_128),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_110),
.A2(n_31),
.B1(n_37),
.B2(n_11),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_129),
.B(n_11),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_220),
.B(n_146),
.Y(n_226)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_135),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_221),
.A2(n_165),
.B1(n_31),
.B2(n_12),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_136),
.B(n_31),
.Y(n_222)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_126),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_223),
.A2(n_134),
.B1(n_132),
.B2(n_161),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_225),
.A2(n_163),
.B1(n_149),
.B2(n_117),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_226),
.B(n_265),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_193),
.B(n_135),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_232),
.B(n_237),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_236),
.A2(n_243),
.B1(n_244),
.B2(n_260),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_192),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_239),
.B(n_215),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_185),
.A2(n_136),
.B1(n_143),
.B2(n_108),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_196),
.A2(n_143),
.B1(n_127),
.B2(n_152),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_192),
.B(n_160),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_202),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g299 ( 
.A1(n_258),
.A2(n_268),
.B1(n_269),
.B2(n_181),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_261),
.A2(n_186),
.B1(n_203),
.B2(n_216),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_178),
.B(n_156),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_211),
.A2(n_133),
.B1(n_117),
.B2(n_163),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_263),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_271),
.B(n_288),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_272),
.A2(n_296),
.B1(n_250),
.B2(n_275),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_273),
.B(n_277),
.Y(n_312)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_238),
.Y(n_274)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_274),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_275),
.A2(n_276),
.B1(n_284),
.B2(n_287),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_253),
.A2(n_195),
.B1(n_196),
.B2(n_219),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_237),
.B(n_202),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_227),
.Y(n_278)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_278),
.Y(n_317)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_227),
.Y(n_281)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_281),
.Y(n_328)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_267),
.Y(n_282)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_282),
.Y(n_335)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_267),
.Y(n_283)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_283),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_253),
.A2(n_196),
.B1(n_189),
.B2(n_217),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_230),
.B(n_215),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_285),
.B(n_290),
.C(n_292),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_232),
.B(n_190),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_286),
.B(n_301),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_253),
.A2(n_213),
.B1(n_183),
.B2(n_221),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_235),
.Y(n_288)
);

OAI32xp33_ASAP7_75t_L g289 ( 
.A1(n_252),
.A2(n_222),
.A3(n_218),
.B1(n_198),
.B2(n_174),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_289),
.B(n_297),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_230),
.B(n_222),
.C(n_188),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_248),
.Y(n_291)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_291),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_231),
.B(n_207),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_L g293 ( 
.A1(n_236),
.A2(n_205),
.B1(n_204),
.B2(n_179),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_293),
.A2(n_295),
.B1(n_304),
.B2(n_306),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_231),
.B(n_234),
.C(n_247),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_294),
.B(n_303),
.C(n_246),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_243),
.A2(n_187),
.B1(n_184),
.B2(n_197),
.Y(n_295)
);

OAI21xp33_ASAP7_75t_SL g296 ( 
.A1(n_228),
.A2(n_250),
.B(n_239),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_235),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_248),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_298),
.B(n_300),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_299),
.A2(n_251),
.B1(n_255),
.B2(n_257),
.Y(n_324)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_233),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_265),
.B(n_223),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_226),
.B(n_182),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_302),
.B(n_305),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_244),
.B(n_233),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_228),
.A2(n_176),
.B1(n_175),
.B2(n_171),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_262),
.B(n_0),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_L g306 ( 
.A1(n_256),
.A2(n_207),
.B1(n_11),
.B2(n_12),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_305),
.Y(n_307)
);

OR2x2_ASAP7_75t_L g344 ( 
.A(n_307),
.B(n_318),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_309),
.A2(n_324),
.B1(n_297),
.B2(n_274),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_275),
.A2(n_264),
.B(n_254),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_310),
.A2(n_321),
.B(n_325),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_280),
.A2(n_240),
.B1(n_264),
.B2(n_256),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_311),
.A2(n_322),
.B1(n_332),
.B2(n_337),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_303),
.A2(n_229),
.B1(n_254),
.B2(n_262),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_314),
.A2(n_249),
.B1(n_1),
.B2(n_3),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_302),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_279),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_319),
.B(n_338),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_273),
.A2(n_229),
.B(n_259),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_280),
.A2(n_229),
.B1(n_245),
.B2(n_238),
.Y(n_322)
);

CKINVDCx14_ASAP7_75t_R g323 ( 
.A(n_277),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_323),
.B(n_271),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_270),
.A2(n_259),
.B(n_207),
.Y(n_325)
);

AND2x2_ASAP7_75t_SL g327 ( 
.A(n_270),
.B(n_246),
.Y(n_327)
);

FAx1_ASAP7_75t_SL g371 ( 
.A(n_327),
.B(n_0),
.CI(n_4),
.CON(n_371),
.SN(n_371)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_290),
.A2(n_300),
.B(n_304),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_329),
.A2(n_278),
.B(n_283),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_286),
.A2(n_245),
.B1(n_251),
.B2(n_255),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_333),
.B(n_313),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_295),
.A2(n_257),
.B1(n_255),
.B2(n_241),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_288),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_287),
.B(n_242),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_339),
.B(n_4),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_276),
.A2(n_257),
.B1(n_241),
.B2(n_242),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_341),
.A2(n_272),
.B1(n_281),
.B2(n_282),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_342),
.B(n_353),
.C(n_354),
.Y(n_375)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_320),
.Y(n_343)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_343),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_345),
.A2(n_367),
.B1(n_308),
.B2(n_323),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_334),
.A2(n_294),
.B(n_289),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_348),
.A2(n_359),
.B(n_374),
.Y(n_391)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_317),
.Y(n_349)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_349),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_313),
.B(n_285),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_350),
.B(n_352),
.Y(n_393)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_320),
.Y(n_351)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_351),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_313),
.B(n_333),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_333),
.B(n_292),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_312),
.B(n_284),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g388 ( 
.A1(n_355),
.A2(n_310),
.B(n_325),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_357),
.A2(n_362),
.B1(n_365),
.B2(n_324),
.Y(n_392)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_358),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g359 ( 
.A1(n_334),
.A2(n_298),
.B(n_291),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_318),
.B(n_0),
.Y(n_360)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_360),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_312),
.B(n_266),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_361),
.B(n_369),
.C(n_371),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_311),
.A2(n_266),
.B1(n_249),
.B2(n_3),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_317),
.Y(n_363)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_363),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_307),
.B(n_0),
.Y(n_364)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_364),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_322),
.A2(n_266),
.B1(n_249),
.B2(n_3),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_315),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_366),
.B(n_370),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_319),
.A2(n_12),
.B1(n_16),
.B2(n_15),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_368),
.B(n_371),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_326),
.B(n_12),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_315),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_330),
.B(n_4),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_372),
.B(n_371),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g373 ( 
.A(n_328),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_373),
.B(n_338),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_SL g435 ( 
.A(n_376),
.B(n_14),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_356),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_378),
.B(n_382),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_381),
.A2(n_383),
.B1(n_396),
.B2(n_400),
.Y(n_411)
);

CKINVDCx14_ASAP7_75t_R g382 ( 
.A(n_358),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_354),
.A2(n_341),
.B1(n_339),
.B2(n_327),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_347),
.A2(n_331),
.B1(n_309),
.B2(n_327),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_384),
.A2(n_387),
.B1(n_392),
.B2(n_401),
.Y(n_408)
);

INVxp33_ASAP7_75t_L g386 ( 
.A(n_360),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_386),
.B(n_399),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_347),
.A2(n_331),
.B1(n_327),
.B2(n_329),
.Y(n_387)
);

AO21x1_ASAP7_75t_L g421 ( 
.A1(n_388),
.A2(n_389),
.B(n_404),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_346),
.A2(n_321),
.B(n_310),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_367),
.A2(n_339),
.B1(n_308),
.B2(n_332),
.Y(n_396)
);

BUFx2_ASAP7_75t_L g398 ( 
.A(n_365),
.Y(n_398)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_398),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g399 ( 
.A(n_349),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_359),
.A2(n_339),
.B1(n_331),
.B2(n_337),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_357),
.A2(n_329),
.B1(n_314),
.B2(n_321),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_344),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_403),
.B(n_378),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_344),
.A2(n_326),
.B(n_325),
.Y(n_404)
);

CKINVDCx14_ASAP7_75t_R g428 ( 
.A(n_405),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_406),
.B(n_372),
.Y(n_414)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_394),
.Y(n_410)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_410),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_391),
.A2(n_346),
.B(n_348),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_413),
.A2(n_417),
.B(n_420),
.Y(n_436)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_414),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_400),
.A2(n_355),
.B1(n_362),
.B2(n_364),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_415),
.A2(n_425),
.B1(n_398),
.B2(n_395),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_416),
.Y(n_439)
);

A2O1A1Ixp33_ASAP7_75t_L g417 ( 
.A1(n_404),
.A2(n_330),
.B(n_363),
.C(n_374),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_393),
.B(n_352),
.C(n_342),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_418),
.B(n_375),
.C(n_376),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_387),
.A2(n_361),
.B1(n_374),
.B2(n_353),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_419),
.A2(n_422),
.B1(n_429),
.B2(n_432),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_391),
.A2(n_316),
.B(n_350),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_384),
.A2(n_316),
.B1(n_336),
.B2(n_335),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_403),
.B(n_336),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_423),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_377),
.A2(n_340),
.B(n_368),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_SL g454 ( 
.A(n_424),
.B(n_380),
.C(n_388),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_394),
.A2(n_335),
.B1(n_328),
.B2(n_340),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_379),
.B(n_369),
.Y(n_426)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_426),
.Y(n_447)
);

OAI21xp33_ASAP7_75t_L g427 ( 
.A1(n_379),
.A2(n_13),
.B(n_15),
.Y(n_427)
);

NAND2xp33_ASAP7_75t_SL g441 ( 
.A(n_427),
.B(n_397),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_401),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_429)
);

NOR3xp33_ASAP7_75t_L g430 ( 
.A(n_390),
.B(n_17),
.C(n_7),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_430),
.Y(n_456)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_385),
.Y(n_431)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_431),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_SL g432 ( 
.A1(n_398),
.A2(n_8),
.B1(n_13),
.B2(n_14),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_390),
.B(n_5),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_433),
.B(n_434),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_392),
.A2(n_5),
.B1(n_8),
.B2(n_14),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_435),
.B(n_380),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_424),
.Y(n_437)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_437),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_407),
.Y(n_438)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_438),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_441),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g443 ( 
.A(n_407),
.Y(n_443)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_443),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_SL g466 ( 
.A(n_444),
.B(n_454),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_423),
.B(n_395),
.Y(n_445)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_445),
.Y(n_470)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_409),
.Y(n_446)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_446),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_418),
.B(n_393),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_449),
.B(n_458),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_451),
.A2(n_455),
.B1(n_408),
.B2(n_383),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_453),
.B(n_420),
.C(n_419),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_415),
.A2(n_402),
.B1(n_380),
.B2(n_381),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_413),
.B(n_375),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_459),
.B(n_463),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_448),
.A2(n_411),
.B1(n_409),
.B2(n_410),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_462),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_464),
.B(n_469),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_436),
.A2(n_421),
.B(n_416),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_468),
.A2(n_442),
.B(n_389),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_458),
.B(n_411),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_449),
.B(n_408),
.C(n_422),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_471),
.B(n_447),
.C(n_454),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_452),
.A2(n_425),
.B1(n_402),
.B2(n_412),
.Y(n_473)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_473),
.Y(n_483)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_450),
.Y(n_474)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_474),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_453),
.B(n_421),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_475),
.B(n_476),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_455),
.B(n_436),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_450),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_477),
.B(n_439),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_SL g478 ( 
.A1(n_468),
.A2(n_438),
.B(n_443),
.Y(n_478)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_478),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_469),
.B(n_451),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_480),
.B(n_486),
.Y(n_497)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_482),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_484),
.B(n_485),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_475),
.B(n_444),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_471),
.B(n_421),
.Y(n_486)
);

XNOR2x1_ASAP7_75t_L g506 ( 
.A(n_487),
.B(n_485),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_463),
.B(n_447),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_488),
.B(n_428),
.C(n_414),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_459),
.B(n_435),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_SL g505 ( 
.A(n_490),
.B(n_491),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_466),
.B(n_445),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_476),
.B(n_456),
.Y(n_492)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_492),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_494),
.A2(n_495),
.B(n_412),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_465),
.B(n_428),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_493),
.A2(n_462),
.B1(n_461),
.B2(n_470),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_496),
.A2(n_499),
.B1(n_503),
.B2(n_504),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_481),
.B(n_464),
.C(n_466),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_498),
.B(n_502),
.C(n_486),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_493),
.A2(n_483),
.B1(n_484),
.B2(n_473),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_481),
.B(n_467),
.C(n_460),
.Y(n_502)
);

NOR2x1_ASAP7_75t_L g504 ( 
.A(n_488),
.B(n_457),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_506),
.B(n_507),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_489),
.A2(n_446),
.B1(n_472),
.B2(n_396),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_509),
.B(n_433),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_511),
.B(n_514),
.Y(n_529)
);

NOR2xp67_ASAP7_75t_SL g512 ( 
.A(n_506),
.B(n_479),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_L g526 ( 
.A1(n_512),
.A2(n_504),
.B(n_509),
.Y(n_526)
);

A2O1A1Ixp33_ASAP7_75t_L g513 ( 
.A1(n_510),
.A2(n_417),
.B(n_406),
.C(n_431),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_513),
.B(n_516),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_508),
.A2(n_440),
.B1(n_429),
.B2(n_434),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_497),
.B(n_480),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_515),
.B(n_498),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_500),
.B(n_479),
.C(n_440),
.Y(n_516)
);

CKINVDCx16_ASAP7_75t_R g517 ( 
.A(n_508),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_517),
.B(n_501),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_500),
.B(n_399),
.C(n_426),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_519),
.B(n_521),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_502),
.B(n_417),
.C(n_385),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_522),
.B(n_505),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_523),
.B(n_524),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_526),
.B(n_527),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_529),
.B(n_501),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g534 ( 
.A1(n_531),
.A2(n_532),
.B(n_524),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_525),
.A2(n_520),
.B1(n_511),
.B2(n_521),
.Y(n_532)
);

OAI311xp33_ASAP7_75t_L g537 ( 
.A1(n_534),
.A2(n_535),
.A3(n_536),
.B1(n_532),
.C1(n_518),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_L g535 ( 
.A1(n_530),
.A2(n_515),
.B(n_503),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_533),
.A2(n_528),
.B(n_518),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g538 ( 
.A(n_537),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_538),
.B(n_499),
.C(n_496),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_SL g540 ( 
.A1(n_539),
.A2(n_513),
.B(n_397),
.Y(n_540)
);

BUFx24_ASAP7_75t_SL g541 ( 
.A(n_540),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_541),
.B(n_507),
.C(n_15),
.Y(n_542)
);


endmodule