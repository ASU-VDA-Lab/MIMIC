module fake_jpeg_12129_n_435 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_435);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_435;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_13),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_7),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g140 ( 
.A(n_47),
.Y(n_140)
);

BUFx24_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_48),
.Y(n_119)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_49),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_37),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_51),
.B(n_60),
.Y(n_103)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_52),
.Y(n_125)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_53),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_55),
.Y(n_124)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_56),
.Y(n_129)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_57),
.Y(n_128)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_58),
.Y(n_130)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_59),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_16),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_19),
.B(n_1),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_62),
.B(n_69),
.Y(n_99)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_29),
.Y(n_63)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_63),
.Y(n_115)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_65),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_16),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_66),
.B(n_68),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_1),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_67),
.B(n_75),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_40),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_38),
.B(n_43),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_20),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_74),
.B(n_77),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_38),
.B(n_2),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_76),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_20),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_45),
.B(n_2),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_78),
.B(n_82),
.Y(n_141)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_79),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_45),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_81),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_23),
.B(n_2),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_83),
.Y(n_133)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_25),
.Y(n_84)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_17),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_86),
.B(n_3),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_87),
.B(n_88),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_21),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_21),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_89),
.B(n_91),
.Y(n_134)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_90),
.B(n_31),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_24),
.B(n_3),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_53),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_92),
.A2(n_96),
.B1(n_97),
.B2(n_104),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_60),
.A2(n_17),
.B1(n_46),
.B2(n_32),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_93),
.A2(n_98),
.B1(n_137),
.B2(n_51),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_76),
.A2(n_41),
.B1(n_25),
.B2(n_44),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_61),
.A2(n_44),
.B1(n_42),
.B2(n_25),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_66),
.A2(n_17),
.B1(n_46),
.B2(n_30),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_62),
.B(n_27),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_101),
.B(n_120),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_52),
.A2(n_44),
.B1(n_42),
.B2(n_25),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_74),
.B(n_24),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_105),
.B(n_135),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_58),
.A2(n_25),
.B1(n_44),
.B2(n_42),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_111),
.A2(n_113),
.B1(n_114),
.B2(n_121),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_79),
.A2(n_42),
.B1(n_45),
.B2(n_33),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_82),
.A2(n_42),
.B1(n_33),
.B2(n_31),
.Y(n_114)
);

NAND2xp33_ASAP7_75t_SL g179 ( 
.A(n_116),
.B(n_56),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_69),
.B(n_35),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_84),
.A2(n_35),
.B1(n_34),
.B2(n_32),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_57),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_49),
.A2(n_30),
.B1(n_34),
.B2(n_5),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_71),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g229 ( 
.A(n_143),
.Y(n_229)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_109),
.Y(n_144)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_144),
.Y(n_194)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_145),
.B(n_149),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_99),
.B(n_81),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_146),
.B(n_153),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_99),
.B(n_101),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_147),
.B(n_180),
.C(n_138),
.Y(n_230)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_95),
.Y(n_148)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_148),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_103),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_150),
.B(n_151),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_131),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_125),
.Y(n_152)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_152),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_89),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_154),
.Y(n_198)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_109),
.Y(n_155)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_155),
.Y(n_200)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_130),
.Y(n_156)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_156),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_137),
.A2(n_47),
.B1(n_54),
.B2(n_72),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_157),
.A2(n_168),
.B1(n_178),
.B2(n_187),
.Y(n_196)
);

NOR2xp67_ASAP7_75t_L g158 ( 
.A(n_105),
.B(n_88),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_158),
.B(n_167),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_106),
.B(n_77),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_160),
.B(n_184),
.Y(n_192)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_161),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_95),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_162),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_127),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_163),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_123),
.Y(n_164)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_164),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_129),
.Y(n_165)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_165),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_108),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_142),
.A2(n_86),
.B1(n_63),
.B2(n_65),
.Y(n_168)
);

OR2x4_ASAP7_75t_L g169 ( 
.A(n_116),
.B(n_48),
.Y(n_169)
);

NOR2x1_ASAP7_75t_R g204 ( 
.A(n_169),
.B(n_176),
.Y(n_204)
);

BUFx5_ASAP7_75t_L g171 ( 
.A(n_132),
.Y(n_171)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_171),
.Y(n_217)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_119),
.Y(n_172)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_172),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_4),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_174),
.B(n_170),
.Y(n_202)
);

INVx13_ASAP7_75t_L g175 ( 
.A(n_129),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_175),
.Y(n_220)
);

OR2x4_ASAP7_75t_L g176 ( 
.A(n_112),
.B(n_48),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_134),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_177),
.B(n_181),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_115),
.A2(n_85),
.B1(n_83),
.B2(n_73),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g215 ( 
.A(n_179),
.B(n_183),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_115),
.B(n_59),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_119),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_126),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_182),
.A2(n_186),
.B1(n_188),
.B2(n_189),
.Y(n_207)
);

INVx13_ASAP7_75t_L g183 ( 
.A(n_129),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_127),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_185),
.A2(n_102),
.B1(n_94),
.B2(n_57),
.Y(n_233)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_124),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_126),
.A2(n_90),
.B1(n_64),
.B2(n_55),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_119),
.Y(n_188)
);

BUFx12f_ASAP7_75t_L g189 ( 
.A(n_128),
.Y(n_189)
);

INVx3_ASAP7_75t_SL g190 ( 
.A(n_132),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_190),
.A2(n_191),
.B1(n_140),
.B2(n_123),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_123),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_153),
.A2(n_107),
.B1(n_133),
.B2(n_140),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_199),
.A2(n_210),
.B1(n_224),
.B2(n_233),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_202),
.B(n_208),
.Y(n_255)
);

A2O1A1Ixp33_ASAP7_75t_L g205 ( 
.A1(n_146),
.A2(n_118),
.B(n_119),
.C(n_135),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_205),
.B(n_214),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_147),
.B(n_100),
.Y(n_208)
);

AO22x1_ASAP7_75t_L g209 ( 
.A1(n_169),
.A2(n_110),
.B1(n_136),
.B2(n_122),
.Y(n_209)
);

AND2x4_ASAP7_75t_SL g260 ( 
.A(n_209),
.B(n_215),
.Y(n_260)
);

OAI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_185),
.A2(n_140),
.B1(n_122),
.B2(n_110),
.Y(n_210)
);

MAJx2_ASAP7_75t_L g212 ( 
.A(n_174),
.B(n_149),
.C(n_173),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_221),
.C(n_230),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_149),
.B(n_107),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_179),
.B(n_133),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_219),
.B(n_227),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_159),
.B(n_117),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_222),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_176),
.B(n_138),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_223),
.B(n_11),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_159),
.A2(n_136),
.B1(n_100),
.B2(n_124),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_144),
.B(n_117),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_166),
.A2(n_180),
.B1(n_182),
.B2(n_155),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_228),
.A2(n_190),
.B1(n_102),
.B2(n_94),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_224),
.A2(n_180),
.B1(n_186),
.B2(n_148),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_235),
.A2(n_241),
.B1(n_244),
.B2(n_248),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_208),
.B(n_184),
.C(n_187),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_237),
.B(n_247),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_192),
.B(n_193),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_238),
.B(n_256),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_239),
.A2(n_249),
.B1(n_254),
.B2(n_217),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_221),
.A2(n_162),
.B1(n_164),
.B2(n_191),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_195),
.Y(n_242)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_242),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_223),
.A2(n_188),
.B(n_165),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_243),
.A2(n_207),
.B(n_229),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_196),
.A2(n_171),
.B1(n_50),
.B2(n_70),
.Y(n_244)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_232),
.Y(n_245)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_245),
.Y(n_279)
);

BUFx4f_ASAP7_75t_L g246 ( 
.A(n_203),
.Y(n_246)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_246),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_189),
.C(n_143),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_196),
.A2(n_172),
.B1(n_87),
.B2(n_70),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_197),
.A2(n_87),
.B1(n_50),
.B2(n_143),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_232),
.Y(n_250)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_250),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_219),
.A2(n_189),
.B1(n_183),
.B2(n_175),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_251),
.A2(n_269),
.B1(n_225),
.B2(n_220),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_197),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_192),
.B(n_4),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_216),
.Y(n_257)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_257),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_215),
.B(n_4),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_258),
.A2(n_215),
.B(n_209),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_226),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_259),
.B(n_262),
.Y(n_287)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_260),
.Y(n_273)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_195),
.Y(n_261)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_261),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_202),
.B(n_6),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_199),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_263),
.A2(n_266),
.B1(n_206),
.B2(n_213),
.Y(n_277)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_198),
.Y(n_264)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_264),
.Y(n_298)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_198),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_265),
.B(n_270),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_214),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_229),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_268),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_220),
.B(n_11),
.Y(n_268)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_194),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_271),
.A2(n_296),
.B(n_234),
.Y(n_323)
);

NAND3xp33_ASAP7_75t_L g305 ( 
.A(n_272),
.B(n_286),
.C(n_269),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_277),
.B(n_240),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_278),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_236),
.B(n_212),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_280),
.B(n_303),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_242),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_281),
.B(n_282),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_260),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_252),
.A2(n_228),
.B1(n_211),
.B2(n_205),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_283),
.A2(n_291),
.B1(n_280),
.B2(n_293),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_255),
.B(n_218),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_261),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_265),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_252),
.A2(n_211),
.B1(n_204),
.B2(n_212),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_237),
.A2(n_204),
.B1(n_206),
.B2(n_209),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_292),
.A2(n_297),
.B1(n_241),
.B2(n_240),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_236),
.B(n_227),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_293),
.B(n_299),
.C(n_302),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_294),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_258),
.A2(n_217),
.B1(n_218),
.B2(n_225),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_253),
.A2(n_201),
.B1(n_216),
.B2(n_213),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_247),
.B(n_194),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_253),
.B(n_200),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_258),
.B(n_200),
.Y(n_303)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_304),
.Y(n_345)
);

OA21x2_ASAP7_75t_SL g340 ( 
.A1(n_305),
.A2(n_324),
.B(n_284),
.Y(n_340)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_301),
.Y(n_307)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_307),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_273),
.A2(n_243),
.B(n_260),
.Y(n_308)
);

AO21x1_ASAP7_75t_L g344 ( 
.A1(n_308),
.A2(n_327),
.B(n_331),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_287),
.B(n_267),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_309),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_276),
.B(n_254),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_310),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_302),
.B(n_264),
.Y(n_311)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_311),
.Y(n_336)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_301),
.Y(n_313)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_313),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_315),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_316),
.A2(n_326),
.B1(n_330),
.B2(n_319),
.Y(n_335)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_275),
.Y(n_317)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_317),
.Y(n_351)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_275),
.Y(n_320)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_320),
.Y(n_353)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_295),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_321),
.Y(n_334)
);

XOR2x1_ASAP7_75t_L g322 ( 
.A(n_291),
.B(n_260),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_322),
.B(n_329),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_323),
.A2(n_325),
.B(n_328),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_285),
.B(n_270),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_292),
.A2(n_248),
.B(n_249),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_295),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_272),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_294),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_271),
.A2(n_239),
.B(n_246),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_278),
.A2(n_263),
.B1(n_266),
.B2(n_257),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_314),
.B(n_274),
.C(n_299),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_332),
.B(n_339),
.C(n_308),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_335),
.A2(n_338),
.B1(n_346),
.B2(n_307),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_319),
.A2(n_283),
.B1(n_300),
.B2(n_277),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_314),
.B(n_274),
.C(n_303),
.Y(n_339)
);

OR2x2_ASAP7_75t_L g360 ( 
.A(n_340),
.B(n_327),
.Y(n_360)
);

MAJx2_ASAP7_75t_L g342 ( 
.A(n_306),
.B(n_298),
.C(n_296),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_342),
.B(n_322),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_316),
.A2(n_298),
.B1(n_284),
.B2(n_288),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_315),
.A2(n_297),
.B1(n_290),
.B2(n_288),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_347),
.A2(n_350),
.B1(n_317),
.B2(n_320),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_318),
.A2(n_290),
.B1(n_279),
.B2(n_257),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_331),
.B(n_279),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_354),
.B(n_355),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_306),
.B(n_246),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_343),
.A2(n_318),
.B1(n_328),
.B2(n_330),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_356),
.B(n_370),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g357 ( 
.A1(n_333),
.A2(n_337),
.B(n_345),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_357),
.B(n_358),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_348),
.B(n_312),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_SL g390 ( 
.A(n_359),
.B(n_362),
.Y(n_390)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_360),
.Y(n_378)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_351),
.Y(n_361)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_361),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_SL g362 ( 
.A(n_354),
.B(n_311),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_351),
.Y(n_363)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_363),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_332),
.B(n_339),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_364),
.B(n_365),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_336),
.B(n_250),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_366),
.B(n_368),
.C(n_373),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_367),
.A2(n_347),
.B1(n_350),
.B2(n_335),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_355),
.B(n_313),
.C(n_323),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_344),
.B(n_329),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_371),
.B(n_372),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_344),
.B(n_325),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_342),
.B(n_321),
.C(n_326),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_352),
.B(n_245),
.C(n_201),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_374),
.B(n_375),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_352),
.B(n_12),
.Y(n_375)
);

OAI322xp33_ASAP7_75t_L g377 ( 
.A1(n_360),
.A2(n_336),
.A3(n_349),
.B1(n_341),
.B2(n_337),
.C1(n_353),
.C2(n_343),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_377),
.B(n_375),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_356),
.Y(n_381)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_381),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_372),
.B(n_334),
.Y(n_382)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_382),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_SL g385 ( 
.A(n_368),
.B(n_341),
.C(n_338),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_385),
.B(n_373),
.C(n_374),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_386),
.A2(n_366),
.B1(n_359),
.B2(n_362),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_371),
.A2(n_346),
.B(n_353),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_389),
.B(n_14),
.Y(n_399)
);

MAJx2_ASAP7_75t_L g412 ( 
.A(n_392),
.B(n_379),
.C(n_384),
.Y(n_412)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_393),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_376),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_394),
.B(n_397),
.Y(n_408)
);

OAI211xp5_ASAP7_75t_L g404 ( 
.A1(n_396),
.A2(n_403),
.B(n_383),
.C(n_387),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_378),
.B(n_369),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_381),
.A2(n_369),
.B1(n_13),
.B2(n_14),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_398),
.B(n_401),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_399),
.B(n_389),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_391),
.B(n_12),
.C(n_13),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_388),
.B(n_14),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_402),
.B(n_13),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_380),
.B(n_12),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_404),
.B(n_405),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_392),
.B(n_391),
.C(n_385),
.Y(n_405)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_407),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_400),
.A2(n_382),
.B(n_380),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_409),
.B(n_413),
.Y(n_418)
);

INVx11_ASAP7_75t_L g411 ( 
.A(n_400),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_411),
.B(n_395),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_412),
.B(n_408),
.C(n_410),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_415),
.B(n_417),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_405),
.B(n_401),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_419),
.B(n_420),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_409),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_406),
.B(n_411),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_421),
.B(n_407),
.Y(n_422)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_422),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_414),
.A2(n_386),
.B1(n_398),
.B2(n_403),
.Y(n_425)
);

OR2x2_ASAP7_75t_L g428 ( 
.A(n_425),
.B(n_416),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_418),
.B(n_399),
.Y(n_426)
);

INVxp33_ASAP7_75t_L g427 ( 
.A(n_426),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_428),
.B(n_423),
.Y(n_431)
);

A2O1A1O1Ixp25_ASAP7_75t_L g430 ( 
.A1(n_429),
.A2(n_424),
.B(n_420),
.C(n_423),
.D(n_412),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_430),
.A2(n_431),
.B(n_427),
.Y(n_432)
);

MAJx2_ASAP7_75t_L g433 ( 
.A(n_432),
.B(n_379),
.C(n_384),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_433),
.B(n_390),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_434),
.B(n_390),
.Y(n_435)
);


endmodule