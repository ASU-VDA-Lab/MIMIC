module fake_jpeg_23678_n_326 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_326);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_326;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g13 ( 
.A(n_12),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

INVx11_ASAP7_75t_SL g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx8_ASAP7_75t_SL g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_18),
.B(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_31),
.Y(n_42)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_30),
.B(n_36),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_18),
.B(n_27),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_32),
.B(n_34),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_37),
.Y(n_41)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_40),
.B(n_45),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_32),
.B(n_17),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_25),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_29),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

BUFx2_ASAP7_75t_R g49 ( 
.A(n_33),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_49),
.A2(n_30),
.B1(n_36),
.B2(n_13),
.Y(n_55)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_52),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_32),
.B(n_17),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_54),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_17),
.Y(n_54)
);

OAI21xp33_ASAP7_75t_L g85 ( 
.A1(n_55),
.A2(n_20),
.B(n_24),
.Y(n_85)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_61),
.Y(n_77)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_59),
.A2(n_44),
.B1(n_36),
.B2(n_30),
.Y(n_84)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_63),
.B(n_65),
.Y(n_89)
);

INVx6_ASAP7_75t_SL g64 ( 
.A(n_49),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_70),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_37),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

BUFx4f_ASAP7_75t_SL g82 ( 
.A(n_67),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_41),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_42),
.A2(n_31),
.B1(n_13),
.B2(n_23),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_71),
.A2(n_73),
.B1(n_23),
.B2(n_20),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_31),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_53),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_40),
.A2(n_31),
.B(n_20),
.C(n_30),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_74),
.B(n_75),
.Y(n_94)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_61),
.A2(n_13),
.B1(n_50),
.B2(n_44),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_76),
.A2(n_81),
.B1(n_92),
.B2(n_96),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_97),
.Y(n_102)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_79),
.B(n_93),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_70),
.A2(n_13),
.B1(n_50),
.B2(n_44),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_84),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_85),
.A2(n_98),
.B1(n_24),
.B2(n_64),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_33),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_73),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_69),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_91),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_90),
.Y(n_117)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_58),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_68),
.A2(n_16),
.B1(n_23),
.B2(n_21),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_39),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_63),
.A2(n_41),
.B1(n_39),
.B2(n_20),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_101),
.A2(n_89),
.B(n_28),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_82),
.Y(n_103)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_103),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_65),
.Y(n_104)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_57),
.Y(n_105)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_109),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_90),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_107),
.Y(n_127)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_80),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_108),
.B(n_111),
.Y(n_138)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_82),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_113),
.Y(n_141)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_116),
.Y(n_129)
);

FAx1_ASAP7_75t_SL g118 ( 
.A(n_92),
.B(n_73),
.CI(n_57),
.CON(n_118),
.SN(n_118)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_118),
.B(n_87),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_80),
.B(n_60),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_119),
.B(n_60),
.Y(n_131)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_120),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_121),
.A2(n_68),
.B1(n_24),
.B2(n_75),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_123),
.A2(n_140),
.B(n_143),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_98),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_126),
.B(n_117),
.C(n_111),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_101),
.A2(n_104),
.B(n_112),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_130),
.A2(n_142),
.B(n_52),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_131),
.B(n_134),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_L g132 ( 
.A1(n_115),
.A2(n_95),
.B1(n_86),
.B2(n_79),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_132),
.A2(n_133),
.B1(n_136),
.B2(n_147),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_101),
.A2(n_84),
.B1(n_86),
.B2(n_93),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_99),
.B(n_77),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_110),
.A2(n_87),
.B1(n_68),
.B2(n_24),
.Y(n_136)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_99),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_146),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_87),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_102),
.A2(n_89),
.B(n_25),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_110),
.A2(n_106),
.B(n_109),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_144),
.A2(n_145),
.B(n_103),
.Y(n_159)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_114),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_118),
.A2(n_74),
.B1(n_59),
.B2(n_80),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_149),
.B(n_150),
.Y(n_179)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_128),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_141),
.Y(n_151)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_120),
.Y(n_152)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_152),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_118),
.Y(n_154)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_154),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_137),
.B(n_108),
.Y(n_155)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_155),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_107),
.Y(n_156)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_156),
.Y(n_195)
);

AO22x1_ASAP7_75t_SL g157 ( 
.A1(n_123),
.A2(n_43),
.B1(n_47),
.B2(n_48),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_157),
.A2(n_135),
.B1(n_138),
.B2(n_43),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_143),
.A2(n_60),
.B1(n_56),
.B2(n_117),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_158),
.A2(n_157),
.B1(n_166),
.B2(n_145),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_159),
.A2(n_164),
.B1(n_173),
.B2(n_16),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_126),
.C(n_142),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_45),
.Y(n_161)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_161),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_131),
.Y(n_185)
);

OAI21x1_ASAP7_75t_L g163 ( 
.A1(n_133),
.A2(n_111),
.B(n_100),
.Y(n_163)
);

A2O1A1Ixp33_ASAP7_75t_SL g194 ( 
.A1(n_163),
.A2(n_167),
.B(n_170),
.C(n_15),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_144),
.A2(n_111),
.B(n_91),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_90),
.Y(n_165)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_165),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_0),
.Y(n_167)
);

NAND3xp33_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_12),
.C(n_11),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_169),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_122),
.A2(n_54),
.B(n_37),
.Y(n_170)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_124),
.Y(n_171)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_171),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_124),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_172),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_147),
.A2(n_146),
.B1(n_129),
.B2(n_134),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_127),
.B(n_83),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_174),
.Y(n_200)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_129),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_113),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_SL g217 ( 
.A(n_176),
.B(n_183),
.C(n_185),
.Y(n_217)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_177),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_181),
.C(n_201),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_160),
.B(n_140),
.C(n_135),
.Y(n_181)
);

MAJx2_ASAP7_75t_L g183 ( 
.A(n_153),
.B(n_140),
.C(n_127),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_186),
.A2(n_188),
.B1(n_158),
.B2(n_175),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_157),
.Y(n_187)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_187),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_153),
.A2(n_113),
.B1(n_25),
.B2(n_15),
.Y(n_188)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_190),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_SL g222 ( 
.A(n_193),
.B(n_194),
.C(n_188),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_173),
.A2(n_19),
.B1(n_22),
.B2(n_35),
.Y(n_196)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_196),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_156),
.B(n_33),
.C(n_48),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_177),
.B(n_172),
.Y(n_202)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_202),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_198),
.B(n_149),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_203),
.B(n_205),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_179),
.B(n_161),
.Y(n_204)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_204),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_184),
.B(n_150),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_179),
.B(n_168),
.Y(n_206)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_206),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_197),
.B(n_154),
.Y(n_207)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_207),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_200),
.B(n_171),
.Y(n_209)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_209),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_190),
.Y(n_211)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_211),
.Y(n_243)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_186),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_212),
.A2(n_220),
.B(n_221),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_213),
.A2(n_194),
.B(n_167),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_191),
.B(n_148),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_214),
.A2(n_224),
.B(n_19),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_180),
.B(n_164),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_215),
.B(n_185),
.Y(n_225)
);

BUFx5_ASAP7_75t_L g216 ( 
.A(n_181),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_216),
.Y(n_241)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_192),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_178),
.B(n_170),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_222),
.A2(n_212),
.B1(n_223),
.B2(n_207),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_182),
.B(n_162),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_225),
.B(n_231),
.Y(n_257)
);

A2O1A1Ixp33_ASAP7_75t_SL g226 ( 
.A1(n_208),
.A2(n_183),
.B(n_187),
.C(n_195),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_226),
.A2(n_22),
.B(n_19),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_217),
.A2(n_189),
.B1(n_176),
.B2(n_201),
.Y(n_227)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_227),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_217),
.A2(n_189),
.B1(n_199),
.B2(n_159),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_228),
.A2(n_229),
.B1(n_244),
.B2(n_213),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_208),
.A2(n_194),
.B1(n_167),
.B2(n_66),
.Y(n_229)
);

HB1xp67_ASAP7_75t_L g230 ( 
.A(n_216),
.Y(n_230)
);

INVxp67_ASAP7_75t_SL g262 ( 
.A(n_230),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_194),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_232),
.B(n_0),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_66),
.C(n_48),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_233),
.B(n_234),
.C(n_218),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_66),
.C(n_47),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_229),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_33),
.C(n_28),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_241),
.B(n_219),
.C(n_206),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_251),
.C(n_225),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_244),
.B(n_220),
.Y(n_248)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_248),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_253),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_258),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_204),
.C(n_222),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_252),
.A2(n_259),
.B(n_261),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_18),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_47),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_255),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_18),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_239),
.A2(n_226),
.B1(n_236),
.B2(n_238),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_258),
.A2(n_34),
.B(n_3),
.Y(n_280)
);

OAI21xp33_ASAP7_75t_L g260 ( 
.A1(n_237),
.A2(n_11),
.B(n_12),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_SL g267 ( 
.A(n_260),
.B(n_264),
.C(n_226),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_245),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_234),
.B(n_18),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_231),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_226),
.A2(n_22),
.B(n_35),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_250),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_266),
.B(n_269),
.C(n_271),
.Y(n_294)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_267),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_268),
.B(n_275),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_232),
.C(n_21),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_21),
.C(n_28),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_272),
.A2(n_278),
.B(n_279),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_37),
.C(n_34),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_33),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_27),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_0),
.C(n_1),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_256),
.A2(n_34),
.B(n_10),
.Y(n_279)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_280),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_292),
.C(n_5),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_270),
.A2(n_261),
.B1(n_254),
.B2(n_257),
.Y(n_282)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_282),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_269),
.A2(n_259),
.B1(n_264),
.B2(n_4),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_285),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_274),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_2),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_27),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_287),
.B(n_288),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_273),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_289)
);

AOI22x1_ASAP7_75t_L g300 ( 
.A1(n_289),
.A2(n_278),
.B1(n_3),
.B2(n_4),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_265),
.B(n_271),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_2),
.Y(n_293)
);

OR2x2_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_290),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_294),
.Y(n_297)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_297),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_281),
.Y(n_299)
);

OA22x2_ASAP7_75t_L g311 ( 
.A1(n_299),
.A2(n_300),
.B1(n_305),
.B2(n_6),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_283),
.A2(n_2),
.B(n_5),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_301),
.B(n_291),
.C(n_292),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_302),
.B(n_304),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_6),
.C(n_7),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_293),
.B(n_284),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_308),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_286),
.C(n_7),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_297),
.A2(n_6),
.B(n_7),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_310),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_6),
.C(n_7),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_313),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_306),
.A2(n_305),
.B1(n_300),
.B2(n_296),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_314),
.B(n_8),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_315),
.A2(n_311),
.B1(n_312),
.B2(n_8),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_318),
.A2(n_319),
.B(n_317),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_320),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_321),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_322),
.A2(n_314),
.B(n_316),
.Y(n_323)
);

AOI21xp33_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_8),
.B(n_9),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_27),
.Y(n_325)
);

FAx1_ASAP7_75t_SL g326 ( 
.A(n_325),
.B(n_27),
.CI(n_82),
.CON(n_326),
.SN(n_326)
);


endmodule