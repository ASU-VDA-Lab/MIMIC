module real_jpeg_4033_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_507;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_0),
.A2(n_37),
.B1(n_42),
.B2(n_47),
.Y(n_36)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_0),
.A2(n_47),
.B1(n_109),
.B2(n_111),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_0),
.A2(n_47),
.B1(n_157),
.B2(n_159),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_0),
.A2(n_47),
.B1(n_233),
.B2(n_235),
.Y(n_232)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_2),
.A2(n_51),
.B1(n_52),
.B2(n_56),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_2),
.A2(n_51),
.B1(n_149),
.B2(n_151),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_2),
.A2(n_51),
.B1(n_239),
.B2(n_240),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_2),
.A2(n_38),
.B1(n_51),
.B2(n_277),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_3),
.A2(n_251),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_3),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_3),
.A2(n_296),
.B1(n_307),
.B2(n_308),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_3),
.A2(n_296),
.B1(n_392),
.B2(n_393),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_L g409 ( 
.A1(n_3),
.A2(n_296),
.B1(n_404),
.B2(n_410),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_4),
.B(n_261),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_4),
.A2(n_260),
.B(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_4),
.B(n_191),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_4),
.B(n_370),
.C(n_372),
.Y(n_369)
);

OAI22xp33_ASAP7_75t_L g374 ( 
.A1(n_4),
.A2(n_375),
.B1(n_376),
.B2(n_378),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_4),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_4),
.B(n_147),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_4),
.A2(n_26),
.B1(n_315),
.B2(n_421),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_5),
.A2(n_289),
.B1(n_291),
.B2(n_292),
.Y(n_288)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_5),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_5),
.A2(n_281),
.B1(n_291),
.B2(n_307),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_5),
.A2(n_291),
.B1(n_378),
.B2(n_382),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_5),
.A2(n_291),
.B1(n_410),
.B2(n_422),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g171 ( 
.A(n_6),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_7),
.A2(n_123),
.B1(n_126),
.B2(n_127),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_7),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_7),
.A2(n_62),
.B1(n_126),
.B2(n_183),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_7),
.A2(n_126),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_7),
.A2(n_126),
.B1(n_266),
.B2(n_269),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_8),
.A2(n_110),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_8),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_8),
.A2(n_188),
.B1(n_281),
.B2(n_283),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g397 ( 
.A1(n_8),
.A2(n_188),
.B1(n_398),
.B2(n_401),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_8),
.A2(n_188),
.B1(n_378),
.B2(n_461),
.Y(n_460)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_9),
.Y(n_135)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_10),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_10),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_10),
.Y(n_316)
);

BUFx5_ASAP7_75t_L g338 ( 
.A(n_10),
.Y(n_338)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_11),
.Y(n_94)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_11),
.Y(n_98)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_11),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_11),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g258 ( 
.A(n_11),
.Y(n_258)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_12),
.Y(n_102)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_13),
.Y(n_508)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_14),
.Y(n_92)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_14),
.Y(n_95)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_14),
.Y(n_110)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_14),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_14),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_14),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_14),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_14),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_14),
.Y(n_262)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_14),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_15),
.Y(n_511)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_16),
.A2(n_80),
.B1(n_82),
.B2(n_83),
.Y(n_79)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_16),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_16),
.A2(n_82),
.B1(n_110),
.B2(n_116),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_16),
.A2(n_82),
.B1(n_169),
.B2(n_172),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_16),
.A2(n_82),
.B1(n_196),
.B2(n_197),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_17),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_507),
.B(n_509),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_495),
.Y(n_19)
);

OAI31xp33_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_220),
.A3(n_241),
.B(n_492),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_200),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_22),
.B(n_200),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_119),
.C(n_163),
.Y(n_22)
);

FAx1_ASAP7_75t_SL g360 ( 
.A(n_23),
.B(n_119),
.CI(n_163),
.CON(n_360),
.SN(n_360)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_86),
.Y(n_23)
);

AOI21xp33_ASAP7_75t_L g219 ( 
.A1(n_24),
.A2(n_25),
.B(n_88),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_48),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_25),
.A2(n_87),
.B1(n_88),
.B2(n_118),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_25),
.A2(n_48),
.B1(n_87),
.B2(n_352),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_34),
.B(n_36),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_26),
.B(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_26),
.A2(n_264),
.B1(n_272),
.B2(n_276),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_26),
.A2(n_276),
.B(n_313),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_26),
.A2(n_175),
.B(n_397),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_26),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_26),
.A2(n_315),
.B1(n_409),
.B2(n_421),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_26),
.A2(n_36),
.B(n_313),
.Y(n_455)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_29),
.Y(n_271)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_29),
.Y(n_404)
);

BUFx5_ASAP7_75t_L g410 ( 
.A(n_29),
.Y(n_410)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_33),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_33),
.Y(n_430)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_36),
.Y(n_176)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_39),
.A2(n_72),
.B1(n_73),
.B2(n_75),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_45),
.Y(n_423)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_46),
.Y(n_400)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_46),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_48),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_59),
.B(n_77),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_50),
.A2(n_60),
.B1(n_78),
.B2(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

OA22x2_ASAP7_75t_L g132 ( 
.A1(n_53),
.A2(n_85),
.B1(n_133),
.B2(n_136),
.Y(n_132)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_54),
.Y(n_159)
);

INVx5_ASAP7_75t_L g380 ( 
.A(n_54),
.Y(n_380)
);

INVx6_ASAP7_75t_L g385 ( 
.A(n_54),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_54),
.Y(n_445)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_55),
.Y(n_158)
);

BUFx5_ASAP7_75t_L g377 ( 
.A(n_55),
.Y(n_377)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_59),
.B(n_161),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_59),
.A2(n_155),
.B(n_156),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_59),
.A2(n_77),
.B(n_156),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_59),
.A2(n_155),
.B1(n_161),
.B2(n_182),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g475 ( 
.A1(n_59),
.A2(n_476),
.B(n_477),
.Y(n_475)
);

INVx1_ASAP7_75t_SL g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_60),
.A2(n_78),
.B1(n_374),
.B2(n_381),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_60),
.A2(n_78),
.B1(n_381),
.B2(n_391),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_60),
.A2(n_78),
.B1(n_391),
.B2(n_460),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_71),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_63),
.B1(n_66),
.B2(n_70),
.Y(n_61)
);

INVx5_ASAP7_75t_L g368 ( 
.A(n_62),
.Y(n_368)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_69),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_70),
.Y(n_392)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx8_ASAP7_75t_L g268 ( 
.A(n_74),
.Y(n_268)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_78),
.Y(n_155)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_79),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_85),
.Y(n_184)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_88),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_108),
.B(n_114),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_89),
.B(n_217),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_89),
.A2(n_191),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_89),
.A2(n_191),
.B1(n_288),
.B2(n_294),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_90),
.A2(n_187),
.B(n_190),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_90),
.A2(n_117),
.B1(n_302),
.B2(n_304),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_90),
.A2(n_117),
.B1(n_187),
.B2(n_295),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g501 ( 
.A1(n_90),
.A2(n_502),
.B(n_503),
.Y(n_501)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_99),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_93),
.B1(n_95),
.B2(n_96),
.Y(n_91)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_103),
.B1(n_104),
.B2(n_106),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_100),
.Y(n_307)
);

INVx6_ASAP7_75t_SL g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_102),
.Y(n_105)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g130 ( 
.A(n_102),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_102),
.Y(n_140)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_104),
.Y(n_144)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_107),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_108),
.B(n_191),
.Y(n_190)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_110),
.Y(n_293)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_113),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g503 ( 
.A(n_114),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_117),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_115),
.Y(n_217)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_116),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g191 ( 
.A(n_117),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_117),
.A2(n_211),
.B(n_216),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_153),
.B(n_162),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_120),
.B(n_153),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_131),
.B1(n_147),
.B2(n_148),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_122),
.A2(n_132),
.B(n_194),
.Y(n_193)
);

OAI32xp33_ASAP7_75t_L g442 ( 
.A1(n_123),
.A2(n_443),
.A3(n_446),
.B1(n_449),
.B2(n_450),
.Y(n_442)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI21xp33_ASAP7_75t_SL g458 ( 
.A1(n_124),
.A2(n_375),
.B(n_449),
.Y(n_458)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_125),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_125),
.Y(n_286)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx5_ASAP7_75t_L g235 ( 
.A(n_130),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_131),
.B(n_195),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_131),
.A2(n_148),
.B(n_206),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_131),
.A2(n_231),
.B(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_131),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_131),
.A2(n_147),
.B1(n_343),
.B2(n_458),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_131),
.A2(n_147),
.B(n_500),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_137),
.Y(n_131)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_132),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_132),
.B(n_232),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_132),
.A2(n_306),
.B1(n_309),
.B2(n_310),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_132),
.A2(n_306),
.B1(n_309),
.B2(n_342),
.Y(n_341)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_134),
.Y(n_452)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_135),
.Y(n_136)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_135),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_141),
.B1(n_144),
.B2(n_145),
.Y(n_137)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_138),
.Y(n_196)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_140),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_140),
.Y(n_256)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_140),
.Y(n_308)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx6_ASAP7_75t_L g448 ( 
.A(n_142),
.Y(n_448)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_143),
.Y(n_146)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_147),
.B(n_195),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_150),
.Y(n_199)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_160),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_154),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_155),
.B(n_375),
.Y(n_419)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_158),
.Y(n_454)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_159),
.Y(n_464)
);

FAx1_ASAP7_75t_SL g200 ( 
.A(n_162),
.B(n_201),
.CI(n_219),
.CON(n_200),
.SN(n_200)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_185),
.C(n_192),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_164),
.B(n_354),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_179),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_165),
.A2(n_179),
.B1(n_180),
.B2(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_165),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_175),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_167),
.A2(n_265),
.B(n_338),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_168),
.Y(n_317)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_170),
.Y(n_277)
);

BUFx5_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_171),
.Y(n_174)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_185),
.A2(n_186),
.B1(n_192),
.B2(n_193),
.Y(n_354)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_194),
.B(n_230),
.Y(n_229)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_198),
.B(n_375),
.Y(n_449)
);

INVx6_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_222),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_200),
.B(n_222),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_210),
.B2(n_218),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_208),
.B2(n_209),
.Y(n_203)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_204),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_204),
.A2(n_209),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_204),
.B(n_228),
.C(n_236),
.Y(n_504)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_205),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_205),
.B(n_209),
.C(n_210),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_207),
.A2(n_232),
.B(n_309),
.Y(n_327)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_210),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_210),
.A2(n_218),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_210),
.B(n_223),
.C(n_226),
.Y(n_497)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_211),
.Y(n_237)
);

INVx8_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx8_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_215),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_221),
.A2(n_493),
.B(n_494),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_236),
.Y(n_226)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_232),
.Y(n_500)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_235),
.Y(n_282)
);

CKINVDCx14_ASAP7_75t_R g502 ( 
.A(n_238),
.Y(n_502)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

OA21x2_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_361),
.B(n_486),
.Y(n_241)
);

NAND3xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_346),
.C(n_358),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_331),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_244),
.A2(n_488),
.B(n_489),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_319),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_245),
.B(n_319),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_299),
.C(n_311),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_246),
.B(n_345),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_278),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_247),
.B(n_279),
.C(n_287),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_263),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_248),
.B(n_263),
.Y(n_334)
);

OAI32xp33_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_251),
.A3(n_253),
.B1(n_255),
.B2(n_259),
.Y(n_248)
);

BUFx12f_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

INVx6_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVxp33_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_273),
.Y(n_272)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g372 ( 
.A(n_277),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_287),
.Y(n_278)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_280),
.Y(n_310)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx4_ASAP7_75t_SL g284 ( 
.A(n_285),
.Y(n_284)
);

INVx5_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_288),
.Y(n_304)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_289),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_299),
.B(n_311),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.C(n_305),
.Y(n_299)
);

FAx1_ASAP7_75t_SL g333 ( 
.A(n_300),
.B(n_301),
.CI(n_305),
.CON(n_333),
.SN(n_333)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_318),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_312),
.B(n_318),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_317),
.Y(n_313)
);

INVx3_ASAP7_75t_SL g314 ( 
.A(n_315),
.Y(n_314)
);

INVx4_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_320),
.B(n_322),
.C(n_324),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_324),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_330),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_326),
.A2(n_327),
.B1(n_328),
.B2(n_329),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_326),
.B(n_329),
.C(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_328),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_330),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_344),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_332),
.B(n_344),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.C(n_335),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_333),
.B(n_484),
.Y(n_483)
);

BUFx24_ASAP7_75t_SL g512 ( 
.A(n_333),
.Y(n_512)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_334),
.B(n_335),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_339),
.C(n_341),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_336),
.A2(n_337),
.B1(n_339),
.B2(n_340),
.Y(n_471)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_SL g470 ( 
.A(n_341),
.B(n_471),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

A2O1A1O1Ixp25_ASAP7_75t_L g486 ( 
.A1(n_346),
.A2(n_358),
.B(n_487),
.C(n_490),
.D(n_491),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_347),
.B(n_357),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_347),
.B(n_357),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_350),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_348),
.B(n_351),
.C(n_356),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_351),
.A2(n_353),
.B1(n_355),
.B2(n_356),
.Y(n_350)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_351),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_353),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_360),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_359),
.B(n_360),
.Y(n_491)
);

BUFx24_ASAP7_75t_SL g515 ( 
.A(n_360),
.Y(n_515)
);

AOI21xp5_ASAP7_75t_L g361 ( 
.A1(n_362),
.A2(n_481),
.B(n_485),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_363),
.A2(n_466),
.B(n_480),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_364),
.A2(n_438),
.B(n_465),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_365),
.A2(n_405),
.B(n_437),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_386),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_366),
.B(n_386),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_373),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_367),
.B(n_373),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_369),
.Y(n_367)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_375),
.B(n_428),
.Y(n_427)
);

INVx3_ASAP7_75t_SL g376 ( 
.A(n_377),
.Y(n_376)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx4_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_385),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_396),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_388),
.A2(n_389),
.B1(n_390),
.B2(n_395),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_388),
.B(n_395),
.C(n_396),
.Y(n_439)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_SL g395 ( 
.A(n_390),
.Y(n_395)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_397),
.Y(n_412)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx6_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx6_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_406),
.A2(n_417),
.B(n_436),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_416),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_407),
.B(n_416),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_408),
.A2(n_411),
.B1(n_412),
.B2(n_413),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_418),
.A2(n_424),
.B(n_435),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_420),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_419),
.B(n_420),
.Y(n_435)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_425),
.B(n_426),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_427),
.B(n_431),
.Y(n_426)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx8_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx4_ASAP7_75t_SL g432 ( 
.A(n_433),
.Y(n_432)
);

INVx4_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_440),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_439),
.B(n_440),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_456),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_441),
.B(n_457),
.C(n_459),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_SL g441 ( 
.A(n_442),
.B(n_455),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_442),
.B(n_455),
.Y(n_474)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx11_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_453),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_459),
.Y(n_456)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_460),
.Y(n_476)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_468),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_467),
.B(n_468),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_469),
.A2(n_470),
.B1(n_472),
.B2(n_473),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_469),
.B(n_475),
.C(n_478),
.Y(n_482)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_474),
.A2(n_475),
.B1(n_478),
.B2(n_479),
.Y(n_473)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_474),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_475),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_483),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_482),
.B(n_483),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_496),
.B(n_505),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_497),
.B(n_498),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_497),
.B(n_498),
.Y(n_506)
);

BUFx24_ASAP7_75t_SL g514 ( 
.A(n_498),
.Y(n_514)
);

FAx1_ASAP7_75t_SL g498 ( 
.A(n_499),
.B(n_501),
.CI(n_504),
.CON(n_498),
.SN(n_498)
);

INVxp67_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx6_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx6_ASAP7_75t_L g510 ( 
.A(n_508),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_510),
.B(n_511),
.Y(n_509)
);


endmodule