module fake_netlist_6_1524_n_760 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_77, n_149, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_760);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_77;
input n_149;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_760;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_226;
wire n_161;
wire n_208;
wire n_462;
wire n_671;
wire n_607;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_725;
wire n_358;
wire n_160;
wire n_751;
wire n_449;
wire n_749;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_742;
wire n_532;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_746;
wire n_609;
wire n_432;
wire n_641;
wire n_693;
wire n_167;
wire n_631;
wire n_174;
wire n_516;
wire n_153;
wire n_720;
wire n_525;
wire n_758;
wire n_611;
wire n_156;
wire n_491;
wire n_656;
wire n_666;
wire n_371;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_163;
wire n_717;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_279;
wire n_686;
wire n_252;
wire n_757;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_411;
wire n_503;
wire n_716;
wire n_152;
wire n_623;
wire n_599;
wire n_513;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_731;
wire n_570;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_683;
wire n_620;
wire n_420;
wire n_608;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_164;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_635;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_728;
wire n_681;
wire n_729;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_688;
wire n_722;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_171;
wire n_678;
wire n_192;
wire n_169;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_SL g152 ( 
.A(n_110),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_94),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_15),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_98),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_115),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_99),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_57),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_136),
.Y(n_159)
);

BUFx10_ASAP7_75t_L g160 ( 
.A(n_131),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_87),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_124),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_60),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_44),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_129),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_123),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_77),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_76),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_14),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_71),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_113),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_101),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_32),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_4),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_25),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_58),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_67),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_81),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_28),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_137),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_64),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_51),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_117),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_141),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_97),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_2),
.Y(n_186)
);

INVx2_ASAP7_75t_SL g187 ( 
.A(n_108),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_83),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_10),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_59),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_73),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_56),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_61),
.Y(n_193)
);

INVxp33_ASAP7_75t_SL g194 ( 
.A(n_96),
.Y(n_194)
);

NOR2xp67_ASAP7_75t_L g195 ( 
.A(n_68),
.B(n_79),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_15),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_145),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_33),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_4),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_78),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_92),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_120),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_150),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_50),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_16),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_41),
.Y(n_206)
);

BUFx10_ASAP7_75t_L g207 ( 
.A(n_62),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_161),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_161),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_161),
.Y(n_210)
);

BUFx8_ASAP7_75t_SL g211 ( 
.A(n_155),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_169),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_196),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_185),
.B(n_200),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_161),
.Y(n_215)
);

AND2x2_ASAP7_75t_SL g216 ( 
.A(n_203),
.B(n_188),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_181),
.Y(n_217)
);

AND2x4_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_22),
.Y(n_218)
);

BUFx12f_ASAP7_75t_L g219 ( 
.A(n_160),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_156),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_160),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_179),
.Y(n_222)
);

NOR2x1_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_0),
.Y(n_223)
);

AND2x4_ASAP7_75t_L g224 ( 
.A(n_179),
.B(n_23),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_160),
.B(n_1),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_3),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_207),
.B(n_3),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_199),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_181),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_181),
.Y(n_230)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_181),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_187),
.B(n_5),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_182),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_182),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_159),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_153),
.Y(n_236)
);

AND2x4_ASAP7_75t_L g237 ( 
.A(n_157),
.B(n_151),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_158),
.B(n_163),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_199),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_166),
.Y(n_240)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_170),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_171),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_207),
.B(n_5),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_172),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_176),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_189),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_177),
.Y(n_247)
);

BUFx12f_ASAP7_75t_L g248 ( 
.A(n_154),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_174),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_162),
.Y(n_250)
);

AND2x6_ASAP7_75t_L g251 ( 
.A(n_224),
.B(n_178),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_215),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_215),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_208),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_220),
.B(n_180),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_208),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_208),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_210),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_210),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_210),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_230),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_230),
.Y(n_262)
);

CKINVDCx6p67_ASAP7_75t_R g263 ( 
.A(n_219),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_230),
.Y(n_264)
);

OAI22xp33_ASAP7_75t_L g265 ( 
.A1(n_227),
.A2(n_205),
.B1(n_186),
.B2(n_173),
.Y(n_265)
);

INVx2_ASAP7_75t_SL g266 ( 
.A(n_249),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_221),
.B(n_194),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_218),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_230),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_231),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_231),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_211),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_214),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_235),
.B(n_184),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_231),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_250),
.B(n_190),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_231),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_234),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_233),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_233),
.Y(n_280)
);

NAND3xp33_ASAP7_75t_L g281 ( 
.A(n_238),
.B(n_192),
.C(n_167),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_L g282 ( 
.A1(n_216),
.A2(n_225),
.B1(n_226),
.B2(n_214),
.Y(n_282)
);

BUFx10_ASAP7_75t_L g283 ( 
.A(n_216),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_234),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_234),
.Y(n_285)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_209),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_234),
.Y(n_287)
);

NAND2xp33_ASAP7_75t_L g288 ( 
.A(n_225),
.B(n_152),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_218),
.B(n_191),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_221),
.B(n_194),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_216),
.B(n_155),
.Y(n_291)
);

INVx2_ASAP7_75t_SL g292 ( 
.A(n_228),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_234),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_234),
.Y(n_294)
);

INVx2_ASAP7_75t_SL g295 ( 
.A(n_239),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_226),
.B(n_173),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_218),
.B(n_198),
.Y(n_297)
);

AOI21x1_ASAP7_75t_L g298 ( 
.A1(n_233),
.A2(n_204),
.B(n_206),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_219),
.B(n_201),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_268),
.B(n_261),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_261),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_268),
.B(n_241),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_278),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_278),
.Y(n_304)
);

AND2x4_ASAP7_75t_L g305 ( 
.A(n_273),
.B(n_218),
.Y(n_305)
);

INVx2_ASAP7_75t_SL g306 ( 
.A(n_266),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_255),
.B(n_248),
.Y(n_307)
);

OR2x2_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_232),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_262),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_274),
.B(n_237),
.Y(n_310)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_286),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_282),
.B(n_248),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_262),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_276),
.B(n_281),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_L g315 ( 
.A1(n_251),
.A2(n_224),
.B1(n_237),
.B2(n_223),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_264),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_264),
.B(n_241),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_289),
.B(n_237),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_271),
.B(n_241),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_275),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_275),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_296),
.A2(n_243),
.B1(n_223),
.B2(n_224),
.Y(n_322)
);

AOI221xp5_ASAP7_75t_L g323 ( 
.A1(n_265),
.A2(n_213),
.B1(n_246),
.B2(n_212),
.C(n_244),
.Y(n_323)
);

NAND2xp33_ASAP7_75t_L g324 ( 
.A(n_251),
.B(n_164),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_288),
.A2(n_237),
.B1(n_224),
.B2(n_165),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_284),
.B(n_241),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_266),
.B(n_168),
.Y(n_327)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_286),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_281),
.B(n_175),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_292),
.B(n_183),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_295),
.B(n_193),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_288),
.B(n_240),
.Y(n_332)
);

AND2x2_ASAP7_75t_SL g333 ( 
.A(n_291),
.B(n_240),
.Y(n_333)
);

INVx4_ASAP7_75t_L g334 ( 
.A(n_251),
.Y(n_334)
);

BUFx4_ASAP7_75t_L g335 ( 
.A(n_272),
.Y(n_335)
);

INVx8_ASAP7_75t_L g336 ( 
.A(n_251),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_295),
.B(n_267),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_284),
.B(n_236),
.Y(n_338)
);

NOR2xp67_ASAP7_75t_SL g339 ( 
.A(n_297),
.B(n_209),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_269),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_L g341 ( 
.A1(n_251),
.A2(n_244),
.B1(n_242),
.B2(n_247),
.Y(n_341)
);

INVxp67_ASAP7_75t_SL g342 ( 
.A(n_286),
.Y(n_342)
);

AND2x4_ASAP7_75t_L g343 ( 
.A(n_298),
.B(n_212),
.Y(n_343)
);

INVx8_ASAP7_75t_L g344 ( 
.A(n_251),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_269),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_251),
.A2(n_242),
.B1(n_245),
.B2(n_247),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_285),
.B(n_236),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_285),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_287),
.A2(n_245),
.B(n_222),
.Y(n_349)
);

NAND3xp33_ASAP7_75t_L g350 ( 
.A(n_290),
.B(n_202),
.C(n_197),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_287),
.B(n_222),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_293),
.Y(n_352)
);

INVxp67_ASAP7_75t_SL g353 ( 
.A(n_293),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_294),
.B(n_209),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_299),
.B(n_209),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_283),
.B(n_209),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_294),
.B(n_209),
.Y(n_357)
);

O2A1O1Ixp33_ASAP7_75t_L g358 ( 
.A1(n_279),
.A2(n_229),
.B(n_217),
.C(n_8),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_270),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_283),
.B(n_217),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_270),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_283),
.B(n_217),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_283),
.A2(n_229),
.B1(n_217),
.B2(n_9),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_314),
.B(n_298),
.Y(n_364)
);

NOR2xp67_ASAP7_75t_L g365 ( 
.A(n_306),
.B(n_252),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_310),
.B(n_277),
.Y(n_366)
);

AOI21xp33_ASAP7_75t_L g367 ( 
.A1(n_322),
.A2(n_6),
.B(n_7),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_333),
.A2(n_263),
.B1(n_280),
.B2(n_259),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_315),
.B(n_252),
.Y(n_369)
);

NOR2xp67_ASAP7_75t_L g370 ( 
.A(n_350),
.B(n_253),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_305),
.B(n_263),
.Y(n_371)
);

NOR2x1p5_ASAP7_75t_SL g372 ( 
.A(n_303),
.B(n_256),
.Y(n_372)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_302),
.A2(n_280),
.B(n_253),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_305),
.B(n_318),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_343),
.B(n_256),
.Y(n_375)
);

AO22x1_ASAP7_75t_L g376 ( 
.A1(n_337),
.A2(n_259),
.B1(n_254),
.B2(n_258),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_308),
.B(n_9),
.Y(n_377)
);

A2O1A1Ixp33_ASAP7_75t_L g378 ( 
.A1(n_332),
.A2(n_254),
.B(n_257),
.C(n_260),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_307),
.B(n_217),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_329),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_356),
.A2(n_217),
.B1(n_229),
.B2(n_85),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_300),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_311),
.Y(n_383)
);

NAND3xp33_ASAP7_75t_L g384 ( 
.A(n_323),
.B(n_229),
.C(n_11),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_330),
.B(n_10),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_353),
.A2(n_229),
.B(n_86),
.Y(n_386)
);

AOI21x1_ASAP7_75t_L g387 ( 
.A1(n_339),
.A2(n_229),
.B(n_84),
.Y(n_387)
);

NAND3xp33_ASAP7_75t_SL g388 ( 
.A(n_325),
.B(n_11),
.C(n_12),
.Y(n_388)
);

NOR2x1p5_ASAP7_75t_L g389 ( 
.A(n_335),
.B(n_12),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_311),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_363),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_355),
.B(n_13),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_360),
.B(n_24),
.Y(n_393)
);

AOI21xp33_ASAP7_75t_L g394 ( 
.A1(n_312),
.A2(n_327),
.B(n_331),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g395 ( 
.A(n_362),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_301),
.B(n_26),
.Y(n_396)
);

OAI21x1_ASAP7_75t_L g397 ( 
.A1(n_346),
.A2(n_90),
.B(n_148),
.Y(n_397)
);

OA22x2_ASAP7_75t_L g398 ( 
.A1(n_309),
.A2(n_321),
.B1(n_313),
.B2(n_316),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_320),
.B(n_17),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_338),
.B(n_18),
.Y(n_400)
);

INVx4_ASAP7_75t_L g401 ( 
.A(n_336),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_341),
.A2(n_91),
.B(n_147),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_324),
.A2(n_328),
.B1(n_342),
.B2(n_334),
.Y(n_403)
);

CKINVDCx6p67_ASAP7_75t_R g404 ( 
.A(n_338),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_334),
.A2(n_89),
.B1(n_146),
.B2(n_144),
.Y(n_405)
);

CKINVDCx10_ASAP7_75t_R g406 ( 
.A(n_349),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_304),
.B(n_19),
.Y(n_407)
);

NOR3xp33_ASAP7_75t_L g408 ( 
.A(n_358),
.B(n_20),
.C(n_21),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_326),
.A2(n_88),
.B(n_143),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_348),
.B(n_27),
.Y(n_410)
);

INVxp67_ASAP7_75t_SL g411 ( 
.A(n_347),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_352),
.B(n_29),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_344),
.A2(n_93),
.B(n_142),
.Y(n_413)
);

NAND3xp33_ASAP7_75t_L g414 ( 
.A(n_347),
.B(n_317),
.C(n_319),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_340),
.A2(n_82),
.B1(n_140),
.B2(n_30),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_351),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_344),
.B(n_20),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_326),
.A2(n_95),
.B(n_31),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_317),
.A2(n_21),
.B1(n_34),
.B2(n_35),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_361),
.B(n_36),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_345),
.B(n_37),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_357),
.A2(n_38),
.B(n_39),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_319),
.A2(n_40),
.B(n_42),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_357),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_354),
.A2(n_43),
.B(n_45),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_359),
.Y(n_426)
);

OAI21x1_ASAP7_75t_L g427 ( 
.A1(n_398),
.A2(n_149),
.B(n_47),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_382),
.B(n_46),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_374),
.A2(n_411),
.B(n_366),
.Y(n_429)
);

NAND3xp33_ASAP7_75t_L g430 ( 
.A(n_384),
.B(n_48),
.C(n_49),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_416),
.B(n_52),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g432 ( 
.A1(n_364),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_398),
.Y(n_433)
);

NAND3xp33_ASAP7_75t_SL g434 ( 
.A(n_385),
.B(n_63),
.C(n_65),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_395),
.A2(n_66),
.B1(n_69),
.B2(n_70),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_377),
.A2(n_72),
.B1(n_74),
.B2(n_75),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_424),
.B(n_379),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_380),
.A2(n_80),
.B1(n_100),
.B2(n_102),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_375),
.A2(n_103),
.B(n_104),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_414),
.A2(n_105),
.B(n_106),
.Y(n_440)
);

OAI21x1_ASAP7_75t_L g441 ( 
.A1(n_373),
.A2(n_139),
.B(n_109),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_426),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_369),
.A2(n_107),
.B(n_111),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_403),
.A2(n_112),
.B1(n_114),
.B2(n_116),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_401),
.A2(n_118),
.B(n_119),
.Y(n_445)
);

NOR4xp25_ASAP7_75t_L g446 ( 
.A(n_367),
.B(n_121),
.C(n_122),
.D(n_125),
.Y(n_446)
);

OAI21x1_ASAP7_75t_L g447 ( 
.A1(n_383),
.A2(n_138),
.B(n_127),
.Y(n_447)
);

NOR4xp25_ASAP7_75t_L g448 ( 
.A(n_391),
.B(n_126),
.C(n_128),
.D(n_130),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_383),
.Y(n_449)
);

INVx4_ASAP7_75t_L g450 ( 
.A(n_401),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_404),
.B(n_132),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_390),
.Y(n_452)
);

INVx1_ASAP7_75t_SL g453 ( 
.A(n_371),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_393),
.A2(n_133),
.B(n_134),
.Y(n_454)
);

OAI21x1_ASAP7_75t_L g455 ( 
.A1(n_390),
.A2(n_135),
.B(n_397),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_402),
.A2(n_396),
.B(n_420),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_400),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_402),
.A2(n_417),
.B(n_423),
.Y(n_458)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_421),
.A2(n_394),
.B(n_410),
.Y(n_459)
);

OAI21x1_ASAP7_75t_L g460 ( 
.A1(n_412),
.A2(n_387),
.B(n_386),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_399),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_372),
.Y(n_462)
);

OAI21x1_ASAP7_75t_L g463 ( 
.A1(n_413),
.A2(n_418),
.B(n_422),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_423),
.A2(n_370),
.B(n_409),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_378),
.A2(n_409),
.B(n_392),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_376),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_368),
.A2(n_381),
.B1(n_405),
.B2(n_391),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_365),
.B(n_407),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_388),
.Y(n_469)
);

OAI21x1_ASAP7_75t_L g470 ( 
.A1(n_425),
.A2(n_415),
.B(n_419),
.Y(n_470)
);

NOR2xp67_ASAP7_75t_SL g471 ( 
.A(n_419),
.B(n_406),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_408),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_389),
.B(n_382),
.Y(n_473)
);

NAND2x1_ASAP7_75t_L g474 ( 
.A(n_401),
.B(n_383),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_398),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_374),
.A2(n_411),
.B(n_344),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_398),
.Y(n_477)
);

OAI21xp33_ASAP7_75t_L g478 ( 
.A1(n_377),
.A2(n_337),
.B(n_296),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_371),
.B(n_273),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_374),
.A2(n_411),
.B(n_344),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_374),
.A2(n_411),
.B(n_344),
.Y(n_481)
);

AOI22xp33_ASAP7_75t_L g482 ( 
.A1(n_467),
.A2(n_477),
.B1(n_475),
.B2(n_433),
.Y(n_482)
);

OR2x6_ASAP7_75t_L g483 ( 
.A(n_472),
.B(n_479),
.Y(n_483)
);

A2O1A1Ixp33_ASAP7_75t_L g484 ( 
.A1(n_464),
.A2(n_478),
.B(n_456),
.C(n_443),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_457),
.B(n_437),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_442),
.B(n_472),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_453),
.B(n_461),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_453),
.B(n_473),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_449),
.Y(n_489)
);

OR2x6_ASAP7_75t_L g490 ( 
.A(n_472),
.B(n_458),
.Y(n_490)
);

AO21x2_ASAP7_75t_L g491 ( 
.A1(n_465),
.A2(n_429),
.B(n_459),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_462),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_466),
.B(n_468),
.Y(n_493)
);

OR2x6_ASAP7_75t_L g494 ( 
.A(n_451),
.B(n_450),
.Y(n_494)
);

OAI211xp5_ASAP7_75t_L g495 ( 
.A1(n_448),
.A2(n_446),
.B(n_443),
.C(n_440),
.Y(n_495)
);

AND2x4_ASAP7_75t_L g496 ( 
.A(n_450),
.B(n_452),
.Y(n_496)
);

AOI21x1_ASAP7_75t_L g497 ( 
.A1(n_476),
.A2(n_481),
.B(n_480),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_462),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_474),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_428),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_427),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_431),
.Y(n_502)
);

NOR2xp67_ASAP7_75t_L g503 ( 
.A(n_434),
.B(n_430),
.Y(n_503)
);

OA21x2_ASAP7_75t_L g504 ( 
.A1(n_465),
.A2(n_470),
.B(n_440),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_441),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_469),
.Y(n_506)
);

OAI21x1_ASAP7_75t_L g507 ( 
.A1(n_447),
.A2(n_445),
.B(n_439),
.Y(n_507)
);

NAND2x1p5_ASAP7_75t_L g508 ( 
.A(n_438),
.B(n_471),
.Y(n_508)
);

AOI222xp33_ASAP7_75t_L g509 ( 
.A1(n_436),
.A2(n_430),
.B1(n_435),
.B2(n_432),
.C1(n_444),
.C2(n_448),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_446),
.B(n_436),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_454),
.Y(n_511)
);

OAI21x1_ASAP7_75t_L g512 ( 
.A1(n_455),
.A2(n_460),
.B(n_463),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_450),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_469),
.Y(n_514)
);

INVxp67_ASAP7_75t_L g515 ( 
.A(n_479),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_450),
.Y(n_516)
);

OR2x2_ASAP7_75t_L g517 ( 
.A(n_479),
.B(n_273),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_457),
.B(n_382),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_433),
.Y(n_519)
);

OR2x2_ASAP7_75t_L g520 ( 
.A(n_479),
.B(n_273),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_457),
.B(n_382),
.Y(n_521)
);

AO21x2_ASAP7_75t_L g522 ( 
.A1(n_464),
.A2(n_465),
.B(n_456),
.Y(n_522)
);

CKINVDCx8_ASAP7_75t_R g523 ( 
.A(n_469),
.Y(n_523)
);

OAI21x1_ASAP7_75t_SL g524 ( 
.A1(n_440),
.A2(n_443),
.B(n_431),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_519),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g526 ( 
.A(n_482),
.B(n_490),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_492),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_498),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_492),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_485),
.B(n_518),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_498),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_492),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_483),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_482),
.Y(n_534)
);

OR2x2_ASAP7_75t_L g535 ( 
.A(n_490),
.B(n_483),
.Y(n_535)
);

NOR2x1_ASAP7_75t_L g536 ( 
.A(n_490),
.B(n_493),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_521),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_513),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_489),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_513),
.Y(n_540)
);

NAND3xp33_ASAP7_75t_L g541 ( 
.A(n_509),
.B(n_484),
.C(n_495),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_501),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_486),
.B(n_488),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_486),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_486),
.B(n_515),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_487),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_513),
.Y(n_547)
);

HB1xp67_ASAP7_75t_L g548 ( 
.A(n_483),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_500),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_522),
.Y(n_550)
);

INVx1_ASAP7_75t_SL g551 ( 
.A(n_517),
.Y(n_551)
);

OA21x2_ASAP7_75t_L g552 ( 
.A1(n_484),
.A2(n_510),
.B(n_512),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_502),
.B(n_520),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_522),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_506),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_511),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_504),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_504),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_508),
.B(n_504),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_542),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_526),
.B(n_508),
.Y(n_561)
);

INVx1_ASAP7_75t_SL g562 ( 
.A(n_551),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_526),
.B(n_503),
.Y(n_563)
);

AND2x4_ASAP7_75t_SL g564 ( 
.A(n_544),
.B(n_494),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_534),
.B(n_506),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_530),
.B(n_514),
.Y(n_566)
);

OR2x2_ASAP7_75t_L g567 ( 
.A(n_541),
.B(n_491),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_534),
.B(n_491),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_542),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_538),
.Y(n_570)
);

INVx1_ASAP7_75t_SL g571 ( 
.A(n_546),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_L g572 ( 
.A1(n_536),
.A2(n_524),
.B1(n_514),
.B2(n_494),
.Y(n_572)
);

AND2x4_ASAP7_75t_L g573 ( 
.A(n_544),
.B(n_494),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_556),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_L g575 ( 
.A1(n_537),
.A2(n_523),
.B1(n_496),
.B2(n_513),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_543),
.B(n_496),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_553),
.B(n_537),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_543),
.B(n_549),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_549),
.B(n_496),
.Y(n_579)
);

HB1xp67_ASAP7_75t_L g580 ( 
.A(n_555),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_553),
.B(n_523),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_556),
.Y(n_582)
);

OR2x2_ASAP7_75t_L g583 ( 
.A(n_559),
.B(n_505),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_525),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_545),
.B(n_516),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_525),
.B(n_507),
.Y(n_586)
);

INVx3_ASAP7_75t_SL g587 ( 
.A(n_538),
.Y(n_587)
);

BUFx2_ASAP7_75t_L g588 ( 
.A(n_535),
.Y(n_588)
);

INVxp67_ASAP7_75t_L g589 ( 
.A(n_548),
.Y(n_589)
);

BUFx2_ASAP7_75t_L g590 ( 
.A(n_535),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_528),
.B(n_507),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_557),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_558),
.Y(n_593)
);

AND2x4_ASAP7_75t_L g594 ( 
.A(n_533),
.B(n_499),
.Y(n_594)
);

AND2x2_ASAP7_75t_L g595 ( 
.A(n_528),
.B(n_516),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_550),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_550),
.Y(n_597)
);

BUFx3_ASAP7_75t_L g598 ( 
.A(n_533),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_531),
.Y(n_599)
);

BUFx2_ASAP7_75t_L g600 ( 
.A(n_536),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_554),
.Y(n_601)
);

INVx1_ASAP7_75t_SL g602 ( 
.A(n_533),
.Y(n_602)
);

HB1xp67_ASAP7_75t_L g603 ( 
.A(n_580),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_592),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_592),
.Y(n_605)
);

AND2x4_ASAP7_75t_L g606 ( 
.A(n_573),
.B(n_559),
.Y(n_606)
);

OR2x2_ASAP7_75t_L g607 ( 
.A(n_567),
.B(n_554),
.Y(n_607)
);

AND2x4_ASAP7_75t_L g608 ( 
.A(n_598),
.B(n_540),
.Y(n_608)
);

INVx3_ASAP7_75t_R g609 ( 
.A(n_594),
.Y(n_609)
);

OR2x2_ASAP7_75t_L g610 ( 
.A(n_567),
.B(n_568),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_593),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_593),
.Y(n_612)
);

INVxp67_ASAP7_75t_SL g613 ( 
.A(n_577),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_578),
.B(n_539),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_563),
.B(n_552),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_578),
.B(n_539),
.Y(n_616)
);

OR2x2_ASAP7_75t_L g617 ( 
.A(n_568),
.B(n_552),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_560),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_563),
.B(n_552),
.Y(n_619)
);

OR2x2_ASAP7_75t_L g620 ( 
.A(n_588),
.B(n_552),
.Y(n_620)
);

NAND2x1p5_ASAP7_75t_L g621 ( 
.A(n_600),
.B(n_512),
.Y(n_621)
);

HB1xp67_ASAP7_75t_L g622 ( 
.A(n_571),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_598),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_565),
.B(n_529),
.Y(n_624)
);

HB1xp67_ASAP7_75t_L g625 ( 
.A(n_588),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_565),
.B(n_529),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_561),
.B(n_529),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_560),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_561),
.B(n_527),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_596),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_569),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_590),
.B(n_527),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_569),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_566),
.B(n_540),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_596),
.Y(n_635)
);

OR2x2_ASAP7_75t_L g636 ( 
.A(n_610),
.B(n_583),
.Y(n_636)
);

HB1xp67_ASAP7_75t_L g637 ( 
.A(n_625),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_634),
.B(n_572),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_623),
.Y(n_639)
);

BUFx2_ASAP7_75t_L g640 ( 
.A(n_621),
.Y(n_640)
);

AND2x2_ASAP7_75t_SL g641 ( 
.A(n_606),
.B(n_600),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_613),
.B(n_562),
.Y(n_642)
);

NOR2x1_ASAP7_75t_L g643 ( 
.A(n_623),
.B(n_574),
.Y(n_643)
);

OR2x2_ASAP7_75t_L g644 ( 
.A(n_610),
.B(n_597),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_615),
.B(n_586),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_604),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_604),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_605),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_619),
.B(n_597),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_603),
.B(n_589),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_605),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_622),
.B(n_624),
.Y(n_652)
);

OR2x2_ASAP7_75t_L g653 ( 
.A(n_620),
.B(n_601),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_624),
.B(n_581),
.Y(n_654)
);

BUFx2_ASAP7_75t_L g655 ( 
.A(n_621),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_611),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_626),
.B(n_602),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_611),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_612),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_606),
.B(n_591),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_612),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_630),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_626),
.B(n_584),
.Y(n_663)
);

NAND2x1p5_ASAP7_75t_L g664 ( 
.A(n_643),
.B(n_641),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_646),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_640),
.B(n_606),
.Y(n_666)
);

HB1xp67_ASAP7_75t_L g667 ( 
.A(n_637),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_646),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_647),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_641),
.B(n_606),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_638),
.B(n_614),
.Y(n_671)
);

AND2x4_ASAP7_75t_L g672 ( 
.A(n_640),
.B(n_655),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_642),
.B(n_632),
.Y(n_673)
);

OR2x2_ASAP7_75t_L g674 ( 
.A(n_636),
.B(n_620),
.Y(n_674)
);

BUFx2_ASAP7_75t_L g675 ( 
.A(n_639),
.Y(n_675)
);

AOI22xp5_ASAP7_75t_L g676 ( 
.A1(n_641),
.A2(n_575),
.B1(n_573),
.B2(n_594),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_647),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_652),
.B(n_654),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_648),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_648),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_660),
.B(n_627),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_656),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_651),
.Y(n_683)
);

OAI211xp5_ASAP7_75t_SL g684 ( 
.A1(n_671),
.A2(n_650),
.B(n_657),
.C(n_643),
.Y(n_684)
);

OAI221xp5_ASAP7_75t_L g685 ( 
.A1(n_671),
.A2(n_585),
.B1(n_616),
.B2(n_655),
.C(n_639),
.Y(n_685)
);

OR2x2_ASAP7_75t_L g686 ( 
.A(n_674),
.B(n_636),
.Y(n_686)
);

AOI22xp5_ASAP7_75t_L g687 ( 
.A1(n_676),
.A2(n_664),
.B1(n_666),
.B2(n_670),
.Y(n_687)
);

AOI31xp33_ASAP7_75t_L g688 ( 
.A1(n_664),
.A2(n_644),
.A3(n_609),
.B(n_663),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_669),
.Y(n_689)
);

A2O1A1Ixp33_ASAP7_75t_L g690 ( 
.A1(n_666),
.A2(n_598),
.B(n_573),
.C(n_564),
.Y(n_690)
);

INVx2_ASAP7_75t_SL g691 ( 
.A(n_667),
.Y(n_691)
);

OAI21xp5_ASAP7_75t_SL g692 ( 
.A1(n_678),
.A2(n_660),
.B(n_573),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_665),
.Y(n_693)
);

HB1xp67_ASAP7_75t_L g694 ( 
.A(n_667),
.Y(n_694)
);

OAI22xp33_ASAP7_75t_L g695 ( 
.A1(n_673),
.A2(n_607),
.B1(n_644),
.B2(n_617),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_665),
.Y(n_696)
);

BUFx3_ASAP7_75t_L g697 ( 
.A(n_691),
.Y(n_697)
);

AOI221xp5_ASAP7_75t_L g698 ( 
.A1(n_684),
.A2(n_683),
.B1(n_680),
.B2(n_679),
.C(n_677),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_687),
.B(n_675),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_689),
.Y(n_700)
);

INVx1_ASAP7_75t_SL g701 ( 
.A(n_694),
.Y(n_701)
);

OAI32xp33_ASAP7_75t_L g702 ( 
.A1(n_685),
.A2(n_682),
.A3(n_668),
.B1(n_653),
.B2(n_658),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_701),
.B(n_692),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_698),
.B(n_681),
.Y(n_704)
);

AOI211xp5_ASAP7_75t_L g705 ( 
.A1(n_702),
.A2(n_685),
.B(n_695),
.C(n_690),
.Y(n_705)
);

NOR3xp33_ASAP7_75t_L g706 ( 
.A(n_699),
.B(n_688),
.C(n_540),
.Y(n_706)
);

OAI21xp33_ASAP7_75t_SL g707 ( 
.A1(n_699),
.A2(n_688),
.B(n_686),
.Y(n_707)
);

AOI21xp5_ASAP7_75t_L g708 ( 
.A1(n_700),
.A2(n_672),
.B(n_666),
.Y(n_708)
);

AOI21xp33_ASAP7_75t_SL g709 ( 
.A1(n_707),
.A2(n_672),
.B(n_696),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_706),
.B(n_697),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_704),
.Y(n_711)
);

NAND4xp75_ASAP7_75t_L g712 ( 
.A(n_708),
.B(n_595),
.C(n_579),
.D(n_662),
.Y(n_712)
);

BUFx8_ASAP7_75t_SL g713 ( 
.A(n_710),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_711),
.B(n_705),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_714),
.B(n_710),
.Y(n_715)
);

CKINVDCx14_ASAP7_75t_R g716 ( 
.A(n_713),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_714),
.B(n_709),
.Y(n_717)
);

NOR2x1_ASAP7_75t_L g718 ( 
.A(n_715),
.B(n_717),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_716),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_717),
.Y(n_720)
);

XOR2xp5_ASAP7_75t_L g721 ( 
.A(n_716),
.B(n_712),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_716),
.B(n_703),
.Y(n_722)
);

NOR2x2_ASAP7_75t_L g723 ( 
.A(n_716),
.B(n_693),
.Y(n_723)
);

OAI22x1_ASAP7_75t_L g724 ( 
.A1(n_721),
.A2(n_672),
.B1(n_587),
.B2(n_697),
.Y(n_724)
);

BUFx2_ASAP7_75t_L g725 ( 
.A(n_719),
.Y(n_725)
);

AOI22xp5_ASAP7_75t_L g726 ( 
.A1(n_722),
.A2(n_608),
.B1(n_662),
.B2(n_668),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_718),
.B(n_682),
.Y(n_727)
);

AND3x4_ASAP7_75t_L g728 ( 
.A(n_720),
.B(n_608),
.C(n_594),
.Y(n_728)
);

AND2x4_ASAP7_75t_L g729 ( 
.A(n_723),
.B(n_645),
.Y(n_729)
);

OAI22xp5_ASAP7_75t_L g730 ( 
.A1(n_718),
.A2(n_651),
.B1(n_658),
.B2(n_653),
.Y(n_730)
);

OR4x1_ASAP7_75t_L g731 ( 
.A(n_725),
.B(n_635),
.C(n_630),
.D(n_574),
.Y(n_731)
);

AOI31xp33_ASAP7_75t_L g732 ( 
.A1(n_727),
.A2(n_579),
.A3(n_576),
.B(n_595),
.Y(n_732)
);

OAI22xp5_ASAP7_75t_L g733 ( 
.A1(n_729),
.A2(n_661),
.B1(n_659),
.B2(n_656),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_726),
.B(n_576),
.Y(n_734)
);

OAI221xp5_ASAP7_75t_L g735 ( 
.A1(n_730),
.A2(n_621),
.B1(n_587),
.B2(n_540),
.C(n_659),
.Y(n_735)
);

OAI22xp5_ASAP7_75t_L g736 ( 
.A1(n_728),
.A2(n_661),
.B1(n_617),
.B2(n_608),
.Y(n_736)
);

OA22x2_ASAP7_75t_L g737 ( 
.A1(n_724),
.A2(n_587),
.B1(n_564),
.B2(n_594),
.Y(n_737)
);

OA21x2_ASAP7_75t_L g738 ( 
.A1(n_732),
.A2(n_635),
.B(n_497),
.Y(n_738)
);

OAI22x1_ASAP7_75t_L g739 ( 
.A1(n_734),
.A2(n_609),
.B1(n_633),
.B2(n_631),
.Y(n_739)
);

AOI21xp5_ASAP7_75t_L g740 ( 
.A1(n_737),
.A2(n_564),
.B(n_516),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_735),
.A2(n_632),
.B1(n_627),
.B2(n_629),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_731),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_733),
.Y(n_743)
);

OA22x2_ASAP7_75t_L g744 ( 
.A1(n_736),
.A2(n_633),
.B1(n_631),
.B2(n_628),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_732),
.B(n_547),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_742),
.B(n_649),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_744),
.Y(n_747)
);

OAI22xp5_ASAP7_75t_L g748 ( 
.A1(n_743),
.A2(n_607),
.B1(n_628),
.B2(n_618),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_738),
.Y(n_749)
);

AOI22xp5_ASAP7_75t_L g750 ( 
.A1(n_745),
.A2(n_739),
.B1(n_740),
.B2(n_741),
.Y(n_750)
);

OAI21xp5_ASAP7_75t_L g751 ( 
.A1(n_742),
.A2(n_531),
.B(n_591),
.Y(n_751)
);

AOI221xp5_ASAP7_75t_L g752 ( 
.A1(n_743),
.A2(n_570),
.B1(n_538),
.B2(n_547),
.C(n_618),
.Y(n_752)
);

AOI21x1_ASAP7_75t_L g753 ( 
.A1(n_749),
.A2(n_516),
.B(n_599),
.Y(n_753)
);

AOI21xp5_ASAP7_75t_L g754 ( 
.A1(n_746),
.A2(n_538),
.B(n_547),
.Y(n_754)
);

AOI21xp5_ASAP7_75t_L g755 ( 
.A1(n_751),
.A2(n_538),
.B(n_547),
.Y(n_755)
);

AOI21xp5_ASAP7_75t_L g756 ( 
.A1(n_747),
.A2(n_750),
.B(n_752),
.Y(n_756)
);

AND3x1_ASAP7_75t_L g757 ( 
.A(n_756),
.B(n_748),
.C(n_499),
.Y(n_757)
);

AO21x2_ASAP7_75t_L g758 ( 
.A1(n_753),
.A2(n_532),
.B(n_582),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_757),
.B(n_754),
.Y(n_759)
);

AOI21xp33_ASAP7_75t_L g760 ( 
.A1(n_759),
.A2(n_758),
.B(n_755),
.Y(n_760)
);


endmodule