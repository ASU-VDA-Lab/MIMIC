module real_aes_10469_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_673;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_364;
wire n_319;
wire n_112;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_94;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_455;
wire n_310;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_89;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_87;
wire n_676;
wire n_658;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_88;
wire n_159;
wire n_108;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
wire n_91;
INVxp33_ASAP7_75t_L g516 ( .A(n_0), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_0), .A2(n_76), .B1(n_620), .B2(n_625), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_1), .B(n_152), .Y(n_151) );
AOI22xp5_ASAP7_75t_L g202 ( .A1(n_2), .A2(n_62), .B1(n_150), .B2(n_203), .Y(n_202) );
HB1xp67_ASAP7_75t_L g709 ( .A(n_2), .Y(n_709) );
AND2x2_ASAP7_75t_L g503 ( .A(n_3), .B(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_3), .B(n_58), .Y(n_532) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_3), .Y(n_542) );
INVx1_ASAP7_75t_L g587 ( .A(n_3), .Y(n_587) );
INVxp67_ASAP7_75t_L g552 ( .A(n_4), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g651 ( .A1(n_4), .A2(n_21), .B1(n_625), .B2(n_652), .Y(n_651) );
HB1xp67_ASAP7_75t_L g680 ( .A(n_5), .Y(n_680) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_6), .Y(n_156) );
INVx2_ASAP7_75t_L g600 ( .A(n_7), .Y(n_600) );
OR2x2_ASAP7_75t_L g631 ( .A(n_7), .B(n_598), .Y(n_631) );
INVx1_ASAP7_75t_L g502 ( .A(n_8), .Y(n_502) );
OR2x2_ASAP7_75t_L g531 ( .A(n_8), .B(n_532), .Y(n_531) );
BUFx2_ASAP7_75t_L g544 ( .A(n_8), .Y(n_544) );
BUFx2_ASAP7_75t_L g594 ( .A(n_8), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g170 ( .A1(n_9), .A2(n_29), .B1(n_171), .B2(n_172), .Y(n_170) );
AOI22xp5_ASAP7_75t_L g216 ( .A1(n_10), .A2(n_44), .B1(n_172), .B2(n_174), .Y(n_216) );
NAND3xp33_ASAP7_75t_L g196 ( .A(n_11), .B(n_139), .C(n_172), .Y(n_196) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_12), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_13), .B(n_117), .Y(n_136) );
NAND2xp5_ASAP7_75t_SL g135 ( .A(n_14), .B(n_92), .Y(n_135) );
NAND3xp33_ASAP7_75t_L g191 ( .A(n_15), .B(n_89), .C(n_142), .Y(n_191) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_15), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g201 ( .A1(n_16), .A2(n_20), .B1(n_142), .B2(n_171), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_17), .B(n_117), .Y(n_116) );
BUFx6f_ASAP7_75t_L g89 ( .A(n_18), .Y(n_89) );
INVxp67_ASAP7_75t_L g546 ( .A(n_19), .Y(n_546) );
AOI221xp5_ASAP7_75t_L g643 ( .A1(n_19), .A2(n_46), .B1(n_644), .B2(n_645), .C(n_648), .Y(n_643) );
INVxp67_ASAP7_75t_L g560 ( .A(n_21), .Y(n_560) );
BUFx6f_ASAP7_75t_L g93 ( .A(n_22), .Y(n_93) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_23), .B(n_233), .Y(n_232) );
INVx1_ASAP7_75t_L g598 ( .A(n_24), .Y(n_598) );
INVx1_ASAP7_75t_L g618 ( .A(n_24), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g173 ( .A1(n_25), .A2(n_37), .B1(n_174), .B2(n_177), .Y(n_173) );
OAI221xp5_ASAP7_75t_L g523 ( .A1(n_26), .A2(n_33), .B1(n_524), .B2(n_533), .C(n_537), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g632 ( .A1(n_26), .A2(n_33), .B1(n_633), .B2(n_638), .Y(n_632) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_27), .B(n_89), .Y(n_189) );
OAI21x1_ASAP7_75t_L g109 ( .A1(n_28), .A2(n_48), .B(n_110), .Y(n_109) );
AND2x2_ASAP7_75t_L g218 ( .A(n_30), .B(n_128), .Y(n_218) );
AND2x6_ASAP7_75t_L g83 ( .A(n_31), .B(n_84), .Y(n_83) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_31), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g721 ( .A(n_31), .B(n_673), .Y(n_721) );
NAND2x1p5_ASAP7_75t_L g197 ( .A(n_32), .B(n_128), .Y(n_197) );
INVx1_ASAP7_75t_L g569 ( .A(n_34), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g121 ( .A(n_35), .B(n_92), .Y(n_121) );
INVx1_ASAP7_75t_L g84 ( .A(n_36), .Y(n_84) );
HB1xp67_ASAP7_75t_L g673 ( .A(n_36), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_38), .B(n_128), .Y(n_143) );
NAND2xp5_ASAP7_75t_SL g141 ( .A(n_39), .B(n_142), .Y(n_141) );
INVx1_ASAP7_75t_L g580 ( .A(n_40), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_41), .B(n_142), .Y(n_231) );
NAND2x1_ASAP7_75t_L g127 ( .A(n_42), .B(n_128), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_43), .B(n_139), .Y(n_149) );
INVx2_ASAP7_75t_L g499 ( .A(n_45), .Y(n_499) );
INVxp33_ASAP7_75t_L g567 ( .A(n_46), .Y(n_567) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_47), .B(n_225), .Y(n_224) );
CKINVDCx5p33_ASAP7_75t_R g228 ( .A(n_49), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_50), .B(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g572 ( .A(n_51), .Y(n_572) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_52), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g215 ( .A1(n_53), .A2(n_56), .B1(n_142), .B2(n_171), .Y(n_215) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_54), .Y(n_160) );
BUFx10_ASAP7_75t_L g706 ( .A(n_55), .Y(n_706) );
INVx1_ASAP7_75t_SL g206 ( .A(n_57), .Y(n_206) );
INVx2_ASAP7_75t_L g504 ( .A(n_58), .Y(n_504) );
CKINVDCx5p33_ASAP7_75t_R g180 ( .A(n_59), .Y(n_180) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_60), .Y(n_125) );
INVxp33_ASAP7_75t_L g511 ( .A(n_61), .Y(n_511) );
AOI221xp5_ASAP7_75t_L g609 ( .A1(n_61), .A2(n_63), .B1(n_610), .B2(n_613), .C(n_616), .Y(n_609) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_62), .Y(n_717) );
INVxp33_ASAP7_75t_L g505 ( .A(n_63), .Y(n_505) );
INVx1_ASAP7_75t_L g689 ( .A(n_64), .Y(n_689) );
INVx2_ASAP7_75t_L g110 ( .A(n_65), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_66), .B(n_139), .Y(n_193) );
INVx1_ASAP7_75t_L g576 ( .A(n_67), .Y(n_576) );
CKINVDCx5p33_ASAP7_75t_R g687 ( .A(n_68), .Y(n_687) );
NAND2xp5_ASAP7_75t_SL g113 ( .A(n_69), .B(n_114), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g606 ( .A(n_70), .Y(n_606) );
INVx2_ASAP7_75t_L g500 ( .A(n_71), .Y(n_500) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_72), .B(n_118), .Y(n_229) );
BUFx3_ASAP7_75t_L g603 ( .A(n_73), .Y(n_603) );
INVx1_ASAP7_75t_L g628 ( .A(n_73), .Y(n_628) );
BUFx3_ASAP7_75t_L g605 ( .A(n_74), .Y(n_605) );
INVx1_ASAP7_75t_L g624 ( .A(n_74), .Y(n_624) );
XNOR2xp5_ASAP7_75t_L g488 ( .A(n_75), .B(n_489), .Y(n_488) );
INVxp33_ASAP7_75t_L g493 ( .A(n_76), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_94), .B(n_487), .Y(n_77) );
BUFx2_ASAP7_75t_L g78 ( .A(n_79), .Y(n_78) );
AND2x2_ASAP7_75t_L g79 ( .A(n_80), .B(n_85), .Y(n_79) );
HB1xp67_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_81), .B(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
OAI21xp5_ASAP7_75t_L g161 ( .A1(n_82), .A2(n_151), .B(n_162), .Y(n_161) );
INVx8_ASAP7_75t_L g166 ( .A(n_82), .Y(n_166) );
INVx8_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
BUFx2_ASAP7_75t_L g126 ( .A(n_83), .Y(n_126) );
OAI21x1_ASAP7_75t_L g133 ( .A1(n_83), .A2(n_134), .B(n_137), .Y(n_133) );
OAI21x1_ASAP7_75t_L g187 ( .A1(n_83), .A2(n_188), .B(n_192), .Y(n_187) );
INVx1_ASAP7_75t_L g235 ( .A(n_83), .Y(n_235) );
INVxp67_ASAP7_75t_SL g85 ( .A(n_86), .Y(n_85) );
AO21x1_ASAP7_75t_L g719 ( .A1(n_86), .A2(n_720), .B(n_721), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g86 ( .A(n_87), .B(n_90), .Y(n_86) );
BUFx2_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
AOI21x1_ASAP7_75t_L g120 ( .A1(n_88), .A2(n_121), .B(n_122), .Y(n_120) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_88), .Y(n_169) );
INVx3_ASAP7_75t_L g204 ( .A(n_88), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_88), .A2(n_231), .B(n_232), .Y(n_230) );
BUFx12f_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
INVx5_ASAP7_75t_L g119 ( .A(n_89), .Y(n_119) );
OAI22xp5_ASAP7_75t_L g137 ( .A1(n_89), .A2(n_138), .B1(n_140), .B2(n_141), .Y(n_137) );
INVx5_ASAP7_75t_L g139 ( .A(n_89), .Y(n_139) );
OAI321xp33_ASAP7_75t_L g147 ( .A1(n_89), .A2(n_142), .A3(n_148), .B1(n_149), .B2(n_150), .C(n_151), .Y(n_147) );
HB1xp67_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_92), .Y(n_91) );
INVx1_ASAP7_75t_L g123 ( .A(n_92), .Y(n_123) );
INVx2_ASAP7_75t_L g150 ( .A(n_92), .Y(n_150) );
INVx2_ASAP7_75t_L g158 ( .A(n_92), .Y(n_158) );
OR2x2_ASAP7_75t_L g159 ( .A(n_92), .B(n_160), .Y(n_159) );
BUFx6f_ASAP7_75t_L g92 ( .A(n_93), .Y(n_92) );
INVx2_ASAP7_75t_L g115 ( .A(n_93), .Y(n_115) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_93), .Y(n_118) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_93), .Y(n_142) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_93), .Y(n_172) );
INVx1_ASAP7_75t_L g176 ( .A(n_93), .Y(n_176) );
INVx1_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
NOR3x2_ASAP7_75t_L g95 ( .A(n_96), .B(n_364), .C(n_459), .Y(n_95) );
OR2x2_ASAP7_75t_L g96 ( .A(n_97), .B(n_307), .Y(n_96) );
NAND3xp33_ASAP7_75t_L g97 ( .A(n_98), .B(n_253), .C(n_286), .Y(n_97) );
AOI221xp5_ASAP7_75t_L g98 ( .A1(n_99), .A2(n_182), .B1(n_207), .B2(n_236), .C(n_240), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
OR2x2_ASAP7_75t_L g100 ( .A(n_101), .B(n_144), .Y(n_100) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_101), .B(n_363), .Y(n_420) );
INVx2_ASAP7_75t_SL g431 ( .A(n_101), .Y(n_431) );
OR2x2_ASAP7_75t_L g101 ( .A(n_102), .B(n_130), .Y(n_101) );
INVx1_ASAP7_75t_L g289 ( .A(n_102), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_102), .B(n_130), .Y(n_339) );
AND2x2_ASAP7_75t_L g433 ( .A(n_102), .B(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
OR2x2_ASAP7_75t_L g336 ( .A(n_103), .B(n_163), .Y(n_336) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_103), .Y(n_359) );
INVx2_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g257 ( .A(n_104), .Y(n_257) );
OAI21x1_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_111), .B(n_127), .Y(n_104) );
OAI21x1_ASAP7_75t_L g132 ( .A1(n_105), .A2(n_133), .B(n_143), .Y(n_132) );
OAI21x1_ASAP7_75t_L g247 ( .A1(n_105), .A2(n_111), .B(n_127), .Y(n_247) );
OAI21x1_ASAP7_75t_L g270 ( .A1(n_105), .A2(n_133), .B(n_143), .Y(n_270) );
INVx3_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
AO31x2_ASAP7_75t_L g199 ( .A1(n_106), .A2(n_166), .A3(n_200), .B(n_205), .Y(n_199) );
INVx4_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx3_ASAP7_75t_L g167 ( .A(n_107), .Y(n_167) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_107), .Y(n_276) );
BUFx6f_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx2_ASAP7_75t_L g129 ( .A(n_108), .Y(n_129) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_108), .B(n_235), .Y(n_234) );
INVx2_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g152 ( .A(n_109), .Y(n_152) );
OAI21x1_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_120), .B(n_126), .Y(n_111) );
AOI21x1_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_116), .B(n_119), .Y(n_112) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx2_ASAP7_75t_L g177 ( .A(n_115), .Y(n_177) );
INVxp67_ASAP7_75t_L g190 ( .A(n_117), .Y(n_190) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g171 ( .A(n_118), .Y(n_171) );
INVx2_ASAP7_75t_L g233 ( .A(n_118), .Y(n_233) );
AOI21x1_ASAP7_75t_L g134 ( .A1(n_119), .A2(n_135), .B(n_136), .Y(n_134) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_119), .A2(n_154), .B(n_159), .Y(n_153) );
CKINVDCx6p67_ASAP7_75t_R g178 ( .A(n_119), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g122 ( .A(n_123), .B(n_124), .Y(n_122) );
INVx1_ASAP7_75t_L g140 ( .A(n_123), .Y(n_140) );
INVx4_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx3_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx2_ASAP7_75t_SL g325 ( .A(n_131), .Y(n_325) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g321 ( .A(n_132), .Y(n_321) );
O2A1O1Ixp33_ASAP7_75t_L g227 ( .A1(n_139), .A2(n_142), .B(n_228), .C(n_229), .Y(n_227) );
INVx2_ASAP7_75t_SL g195 ( .A(n_142), .Y(n_195) );
INVx1_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x2_ASAP7_75t_L g284 ( .A(n_145), .B(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g305 ( .A(n_145), .B(n_306), .Y(n_305) );
BUFx3_ASAP7_75t_L g328 ( .A(n_145), .Y(n_328) );
AND2x2_ASAP7_75t_L g145 ( .A(n_146), .B(n_163), .Y(n_145) );
INVx2_ASAP7_75t_L g239 ( .A(n_146), .Y(n_239) );
INVx1_ASAP7_75t_L g249 ( .A(n_146), .Y(n_249) );
OAI21x1_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_153), .B(n_161), .Y(n_146) );
HB1xp67_ASAP7_75t_L g162 ( .A(n_152), .Y(n_162) );
INVx1_ASAP7_75t_L g181 ( .A(n_152), .Y(n_181) );
BUFx5_ASAP7_75t_L g213 ( .A(n_152), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_155), .B(n_157), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g259 ( .A(n_163), .Y(n_259) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g238 ( .A(n_164), .Y(n_238) );
AOI21x1_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_168), .B(n_179), .Y(n_164) );
AND2x2_ASAP7_75t_L g165 ( .A(n_166), .B(n_167), .Y(n_165) );
INVx2_ASAP7_75t_L g186 ( .A(n_167), .Y(n_186) );
OAI22xp5_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_170), .B1(n_173), .B2(n_178), .Y(n_168) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g203 ( .A(n_176), .Y(n_203) );
OAI22xp5_ASAP7_75t_L g200 ( .A1(n_178), .A2(n_201), .B1(n_202), .B2(n_204), .Y(n_200) );
OA22x2_ASAP7_75t_L g214 ( .A1(n_178), .A2(n_204), .B1(n_215), .B2(n_216), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_180), .B(n_181), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_181), .B(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g225 ( .A(n_181), .Y(n_225) );
INVxp67_ASAP7_75t_SL g182 ( .A(n_183), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_184), .B(n_198), .Y(n_183) );
INVx2_ASAP7_75t_L g302 ( .A(n_184), .Y(n_302) );
NOR2xp67_ASAP7_75t_L g410 ( .A(n_184), .B(n_411), .Y(n_410) );
NAND2xp33_ASAP7_75t_SL g453 ( .A(n_184), .B(n_377), .Y(n_453) );
BUFx3_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AND2x2_ASAP7_75t_L g221 ( .A(n_185), .B(n_222), .Y(n_221) );
AND2x2_ASAP7_75t_L g296 ( .A(n_185), .B(n_223), .Y(n_296) );
OAI21x1_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_187), .B(n_197), .Y(n_185) );
OAI21x1_ASAP7_75t_L g264 ( .A1(n_186), .A2(n_187), .B(n_197), .Y(n_264) );
OAI21xp5_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_190), .B(n_191), .Y(n_188) );
OAI21xp5_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_196), .Y(n_192) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NOR2x1_ASAP7_75t_L g219 ( .A(n_198), .B(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g443 ( .A(n_198), .Y(n_443) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_198), .Y(n_467) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g265 ( .A(n_199), .Y(n_265) );
INVx1_ASAP7_75t_L g293 ( .A(n_199), .Y(n_293) );
AND2x2_ASAP7_75t_L g301 ( .A(n_199), .B(n_275), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_199), .B(n_210), .Y(n_378) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_199), .Y(n_457) );
OAI22xp33_ASAP7_75t_SL g461 ( .A1(n_207), .A2(n_462), .B1(n_463), .B2(n_464), .Y(n_461) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_219), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_208), .B(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g330 ( .A(n_208), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g441 ( .A(n_208), .Y(n_441) );
AND2x2_ASAP7_75t_L g486 ( .A(n_208), .B(n_340), .Y(n_486) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g349 ( .A(n_209), .B(n_340), .Y(n_349) );
AND2x2_ASAP7_75t_L g421 ( .A(n_209), .B(n_422), .Y(n_421) );
NOR2x1_ASAP7_75t_L g435 ( .A(n_209), .B(n_292), .Y(n_435) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g252 ( .A(n_210), .Y(n_252) );
INVx1_ASAP7_75t_L g283 ( .A(n_210), .Y(n_283) );
INVxp67_ASAP7_75t_SL g298 ( .A(n_210), .Y(n_298) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_210), .Y(n_485) );
OAI21x1_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_214), .B(n_217), .Y(n_210) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
OA21x2_ASAP7_75t_L g275 ( .A1(n_214), .A2(n_276), .B(n_277), .Y(n_275) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVxp67_ASAP7_75t_L g277 ( .A(n_218), .Y(n_277) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_L g251 ( .A(n_221), .B(n_252), .Y(n_251) );
INVx1_ASAP7_75t_L g342 ( .A(n_221), .Y(n_342) );
INVx2_ASAP7_75t_L g274 ( .A(n_222), .Y(n_274) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g282 ( .A(n_223), .Y(n_282) );
NAND2x1p5_ASAP7_75t_L g223 ( .A(n_224), .B(n_226), .Y(n_223) );
OAI21x1_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_230), .B(n_234), .Y(n_226) );
NAND3xp33_ASAP7_75t_L g440 ( .A(n_236), .B(n_441), .C(n_442), .Y(n_440) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
OR2x2_ASAP7_75t_L g288 ( .A(n_237), .B(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g318 ( .A(n_237), .B(n_319), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_237), .B(n_339), .Y(n_338) );
OR2x2_ASAP7_75t_L g413 ( .A(n_237), .B(n_245), .Y(n_413) );
OR2x2_ASAP7_75t_L g439 ( .A(n_237), .B(n_339), .Y(n_439) );
NOR2xp67_ASAP7_75t_L g458 ( .A(n_237), .B(n_306), .Y(n_458) );
OR2x2_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
AND2x2_ASAP7_75t_L g248 ( .A(n_238), .B(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_238), .B(n_285), .Y(n_346) );
AND2x2_ASAP7_75t_L g268 ( .A(n_239), .B(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g385 ( .A(n_239), .B(n_270), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_241), .B(n_250), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
AND2x4_ASAP7_75t_L g242 ( .A(n_243), .B(n_248), .Y(n_242) );
OR2x2_ASAP7_75t_L g452 ( .A(n_243), .B(n_346), .Y(n_452) );
INVx2_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g389 ( .A(n_244), .B(n_325), .Y(n_389) );
AND2x2_ASAP7_75t_L g425 ( .A(n_244), .B(n_268), .Y(n_425) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g271 ( .A(n_245), .B(n_258), .Y(n_271) );
AND2x2_ASAP7_75t_L g397 ( .A(n_245), .B(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g405 ( .A(n_245), .B(n_332), .Y(n_405) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_245), .Y(n_418) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g324 ( .A(n_246), .B(n_259), .Y(n_324) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g371 ( .A(n_247), .B(n_249), .Y(n_371) );
AND2x2_ASAP7_75t_L g334 ( .A(n_248), .B(n_320), .Y(n_334) );
INVx2_ASAP7_75t_L g363 ( .A(n_248), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_248), .B(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g403 ( .A(n_249), .Y(n_403) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx2_ASAP7_75t_L g313 ( .A(n_252), .Y(n_313) );
AND2x2_ASAP7_75t_L g476 ( .A(n_252), .B(n_281), .Y(n_476) );
AOI322xp5_ASAP7_75t_L g253 ( .A1(n_254), .A2(n_260), .A3(n_266), .B1(n_271), .B2(n_272), .C1(n_278), .C2(n_284), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
A2O1A1Ixp33_ASAP7_75t_L g479 ( .A1(n_255), .A2(n_480), .B(n_482), .C(n_486), .Y(n_479) );
BUFx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AOI32xp33_ASAP7_75t_L g454 ( .A1(n_256), .A2(n_384), .A3(n_422), .B1(n_455), .B2(n_458), .Y(n_454) );
AND2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
BUFx2_ASAP7_75t_L g304 ( .A(n_257), .Y(n_304) );
INVxp67_ASAP7_75t_SL g327 ( .A(n_257), .Y(n_327) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_259), .Y(n_370) );
NOR2x1p5_ASAP7_75t_L g380 ( .A(n_261), .B(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g272 ( .A(n_262), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g262 ( .A(n_263), .B(n_265), .Y(n_262) );
AND2x2_ASAP7_75t_L g332 ( .A(n_263), .B(n_274), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_263), .B(n_282), .Y(n_395) );
INVx1_ASAP7_75t_L g434 ( .A(n_263), .Y(n_434) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g356 ( .A(n_264), .B(n_275), .Y(n_356) );
AND2x4_ASAP7_75t_L g281 ( .A(n_265), .B(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g412 ( .A(n_265), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_266), .B(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_267), .B(n_336), .Y(n_335) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g285 ( .A(n_270), .Y(n_285) );
INVx1_ASAP7_75t_L g386 ( .A(n_271), .Y(n_386) );
AND2x4_ASAP7_75t_L g463 ( .A(n_271), .B(n_325), .Y(n_463) );
INVx2_ASAP7_75t_L g387 ( .A(n_273), .Y(n_387) );
AND2x4_ASAP7_75t_L g409 ( .A(n_273), .B(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
AND2x2_ASAP7_75t_L g340 ( .A(n_274), .B(n_293), .Y(n_340) );
INVx2_ASAP7_75t_L g355 ( .A(n_274), .Y(n_355) );
INVx3_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
OAI22xp33_ASAP7_75t_L g406 ( .A1(n_279), .A2(n_407), .B1(n_408), .B2(n_413), .Y(n_406) );
OR2x6_ASAP7_75t_L g279 ( .A(n_280), .B(n_283), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x4_ASAP7_75t_L g314 ( .A(n_281), .B(n_302), .Y(n_314) );
INVx1_ASAP7_75t_L g390 ( .A(n_281), .Y(n_390) );
AND2x2_ASAP7_75t_L g422 ( .A(n_282), .B(n_412), .Y(n_422) );
AND2x2_ASAP7_75t_L g382 ( .A(n_283), .B(n_355), .Y(n_382) );
AND2x2_ASAP7_75t_L g450 ( .A(n_283), .B(n_296), .Y(n_450) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_284), .Y(n_350) );
INVx2_ASAP7_75t_L g306 ( .A(n_285), .Y(n_306) );
AOI22xp5_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_290), .B1(n_299), .B2(n_303), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_289), .B(n_385), .Y(n_407) );
AOI221xp5_ASAP7_75t_SL g343 ( .A1(n_290), .A2(n_344), .B1(n_347), .B2(n_350), .C(n_351), .Y(n_343) );
AND2x4_ASAP7_75t_L g290 ( .A(n_291), .B(n_294), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NOR2xp67_ASAP7_75t_L g354 ( .A(n_293), .B(n_355), .Y(n_354) );
BUFx2_ASAP7_75t_L g424 ( .A(n_294), .Y(n_424) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NAND3xp33_ASAP7_75t_L g347 ( .A(n_295), .B(n_330), .C(n_348), .Y(n_347) );
NAND2x1p5_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
INVx2_ASAP7_75t_L g376 ( .A(n_296), .Y(n_376) );
AND2x2_ASAP7_75t_L g455 ( .A(n_296), .B(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
AND2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_305), .Y(n_303) );
AND2x4_ASAP7_75t_L g402 ( .A(n_306), .B(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_343), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_315), .B(n_329), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND2x1p5_ASAP7_75t_L g310 ( .A(n_311), .B(n_314), .Y(n_310) );
AOI21xp5_ASAP7_75t_L g391 ( .A1(n_311), .A2(n_392), .B(n_406), .Y(n_391) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g361 ( .A(n_313), .B(n_332), .Y(n_361) );
NAND3xp33_ASAP7_75t_L g315 ( .A(n_316), .B(n_322), .C(n_326), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_319), .Y(n_481) );
INVx2_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g419 ( .A(n_321), .B(n_403), .Y(n_419) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
INVx2_ASAP7_75t_L g464 ( .A(n_323), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx2_ASAP7_75t_L g449 ( .A(n_324), .Y(n_449) );
AND2x2_ASAP7_75t_L g366 ( .A(n_325), .B(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g472 ( .A(n_325), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
OAI21xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_333), .B(n_337), .Y(n_329) );
INVx2_ASAP7_75t_L g446 ( .A(n_331), .Y(n_446) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NOR2x1_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
AOI22xp5_ASAP7_75t_L g337 ( .A1(n_334), .A2(n_338), .B1(n_340), .B2(n_341), .Y(n_337) );
INVx2_ASAP7_75t_L g367 ( .A(n_336), .Y(n_367) );
OAI221xp5_ASAP7_75t_L g468 ( .A1(n_336), .A2(n_469), .B1(n_474), .B2(n_477), .C(n_479), .Y(n_468) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_SL g398 ( .A(n_346), .Y(n_398) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_357), .B1(n_360), .B2(n_362), .Y(n_351) );
INVx1_ASAP7_75t_L g462 ( .A(n_352), .Y(n_462) );
INVx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_354), .B(n_356), .Y(n_353) );
INVx1_ASAP7_75t_L g430 ( .A(n_355), .Y(n_430) );
AND2x4_ASAP7_75t_L g436 ( .A(n_356), .B(n_422), .Y(n_436) );
OR2x2_ASAP7_75t_L g362 ( .A(n_358), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g368 ( .A(n_360), .Y(n_368) );
INVx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g466 ( .A(n_361), .B(n_467), .Y(n_466) );
NAND4xp75_ASAP7_75t_L g364 ( .A(n_365), .B(n_391), .C(n_414), .D(n_437), .Y(n_364) );
AOI221x1_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_368), .B1(n_369), .B2(n_372), .C(n_383), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_369), .B(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_379), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_377), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_377), .B(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g470 ( .A(n_377), .B(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_378), .B(n_395), .Y(n_473) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
OAI32xp33_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_386), .A3(n_387), .B1(n_388), .B2(n_390), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
A2O1A1Ixp33_ASAP7_75t_L g432 ( .A1(n_385), .A2(n_433), .B(n_435), .C(n_436), .Y(n_432) );
AND2x2_ASAP7_75t_L g447 ( .A(n_385), .B(n_448), .Y(n_447) );
OAI22xp33_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_396), .B1(n_399), .B2(n_404), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx2_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx4_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_402), .Y(n_478) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVxp67_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
A2O1A1Ixp33_ASAP7_75t_L g451 ( .A1(n_413), .A2(n_452), .B(n_453), .C(n_454), .Y(n_451) );
NOR2xp67_ASAP7_75t_L g414 ( .A(n_415), .B(n_426), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_416), .B(n_423), .Y(n_415) );
OAI21xp33_ASAP7_75t_SL g416 ( .A1(n_417), .A2(n_420), .B(n_421), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_424), .B(n_425), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_427), .B(n_432), .Y(n_426) );
NAND2x1_ASAP7_75t_SL g427 ( .A(n_428), .B(n_431), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g471 ( .A(n_430), .Y(n_471) );
AND2x2_ASAP7_75t_L g475 ( .A(n_433), .B(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_434), .B(n_485), .Y(n_484) );
AOI221x1_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_444), .B1(n_447), .B2(n_450), .C(n_451), .Y(n_437) );
NAND2xp5_ASAP7_75t_SL g438 ( .A(n_439), .B(n_440), .Y(n_438) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OR2x2_ASAP7_75t_L g483 ( .A(n_443), .B(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
OR2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_468), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_461), .B(n_465), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_472), .B(n_473), .Y(n_469) );
INVxp67_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVxp67_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
OAI221xp5_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_489), .B1(n_671), .B2(n_676), .C(n_713), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_489), .A2(n_714), .B1(n_717), .B2(n_718), .Y(n_713) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_588), .Y(n_489) );
NOR3xp33_ASAP7_75t_L g490 ( .A(n_491), .B(n_523), .C(n_539), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_492), .B(n_510), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_493), .A2(n_494), .B1(n_505), .B2(n_506), .Y(n_492) );
AND2x4_ASAP7_75t_L g494 ( .A(n_495), .B(n_501), .Y(n_494) );
INVx3_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx3_ASAP7_75t_L g571 ( .A(n_496), .Y(n_571) );
INVx3_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
BUFx6f_ASAP7_75t_L g554 ( .A(n_497), .Y(n_554) );
AND2x4_ASAP7_75t_L g497 ( .A(n_498), .B(n_500), .Y(n_497) );
AND2x4_ASAP7_75t_L g508 ( .A(n_498), .B(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g515 ( .A(n_499), .B(n_500), .Y(n_515) );
INVx1_ASAP7_75t_L g522 ( .A(n_499), .Y(n_522) );
INVx1_ASAP7_75t_L g529 ( .A(n_499), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_499), .B(n_520), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_499), .B(n_500), .Y(n_559) );
INVx1_ASAP7_75t_L g565 ( .A(n_499), .Y(n_565) );
INVx1_ASAP7_75t_L g509 ( .A(n_500), .Y(n_509) );
INVx2_ASAP7_75t_L g520 ( .A(n_500), .Y(n_520) );
INVx1_ASAP7_75t_L g566 ( .A(n_500), .Y(n_566) );
AND2x6_ASAP7_75t_L g506 ( .A(n_501), .B(n_507), .Y(n_506) );
AND2x4_ASAP7_75t_L g512 ( .A(n_501), .B(n_513), .Y(n_512) );
AND2x2_ASAP7_75t_L g517 ( .A(n_501), .B(n_518), .Y(n_517) );
AND2x4_ASAP7_75t_L g501 ( .A(n_502), .B(n_503), .Y(n_501) );
INVx1_ASAP7_75t_L g584 ( .A(n_502), .Y(n_584) );
INVx1_ASAP7_75t_L g543 ( .A(n_504), .Y(n_543) );
INVx1_ASAP7_75t_L g586 ( .A(n_504), .Y(n_586) );
NAND2x1p5_ASAP7_75t_L g538 ( .A(n_507), .B(n_530), .Y(n_538) );
BUFx3_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B1(n_516), .B2(n_517), .Y(n_510) );
INVx2_ASAP7_75t_SL g513 ( .A(n_514), .Y(n_513) );
INVx3_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
BUFx6f_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AND2x4_ASAP7_75t_L g519 ( .A(n_520), .B(n_521), .Y(n_519) );
INVx1_ASAP7_75t_L g536 ( .A(n_520), .Y(n_536) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_SL g524 ( .A(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
NAND2x1_ASAP7_75t_SL g526 ( .A(n_527), .B(n_530), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
NAND2x1p5_ASAP7_75t_L g534 ( .A(n_530), .B(n_535), .Y(n_534) );
INVx3_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
OR2x2_ASAP7_75t_L g591 ( .A(n_531), .B(n_558), .Y(n_591) );
BUFx4f_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
BUFx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
OAI33xp33_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_545), .A3(n_555), .B1(n_568), .B2(n_573), .B3(n_581), .Y(n_539) );
OR2x6_ASAP7_75t_L g540 ( .A(n_541), .B(n_544), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .Y(n_541) );
BUFx2_ASAP7_75t_L g670 ( .A(n_544), .Y(n_670) );
OAI22xp5_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_547), .B1(n_552), .B2(n_553), .Y(n_545) );
OAI22xp5_ASAP7_75t_L g568 ( .A1(n_547), .A2(n_569), .B1(n_570), .B2(n_572), .Y(n_568) );
INVx2_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx4_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
OAI22xp33_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_560), .B1(n_561), .B2(n_567), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx2_ASAP7_75t_SL g557 ( .A(n_558), .Y(n_557) );
INVx2_ASAP7_75t_SL g575 ( .A(n_558), .Y(n_575) );
BUFx6f_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
BUFx6f_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
AND2x2_ASAP7_75t_L g579 ( .A(n_565), .B(n_566), .Y(n_579) );
AOI221xp5_ASAP7_75t_L g608 ( .A1(n_569), .A2(n_609), .B1(n_619), .B2(n_629), .C(n_632), .Y(n_608) );
INVx2_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_572), .A2(n_576), .B1(n_660), .B2(n_665), .Y(n_659) );
OAI22xp33_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_576), .B1(n_577), .B2(n_580), .Y(n_573) );
INVx3_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
BUFx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx3_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AOI221xp5_ASAP7_75t_L g642 ( .A1(n_580), .A2(n_643), .B1(n_651), .B2(n_654), .C(n_656), .Y(n_642) );
CKINVDCx8_ASAP7_75t_R g581 ( .A(n_582), .Y(n_581) );
INVx5_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
OR2x6_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
NAND2x1p5_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
AOI21xp33_ASAP7_75t_SL g588 ( .A1(n_589), .A2(n_606), .B(n_607), .Y(n_588) );
INVx5_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AND2x4_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AND2x4_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
AND2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_601), .Y(n_595) );
AND2x4_ASAP7_75t_L g634 ( .A(n_596), .B(n_635), .Y(n_634) );
AND2x4_ASAP7_75t_L g639 ( .A(n_596), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g658 ( .A(n_596), .Y(n_658) );
AND2x4_ASAP7_75t_L g596 ( .A(n_597), .B(n_599), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x4_ASAP7_75t_L g617 ( .A(n_599), .B(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g650 ( .A(n_600), .B(n_618), .Y(n_650) );
INVx6_ASAP7_75t_L g615 ( .A(n_601), .Y(n_615) );
AND2x4_ASAP7_75t_L g601 ( .A(n_602), .B(n_604), .Y(n_601) );
INVx1_ASAP7_75t_L g641 ( .A(n_602), .Y(n_641) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g612 ( .A(n_603), .B(n_605), .Y(n_612) );
AND2x4_ASAP7_75t_L g623 ( .A(n_603), .B(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g637 ( .A(n_604), .Y(n_637) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
AND2x4_ASAP7_75t_L g627 ( .A(n_605), .B(n_628), .Y(n_627) );
AOI31xp33_ASAP7_75t_L g607 ( .A1(n_608), .A2(n_642), .A3(n_659), .B(n_668), .Y(n_607) );
BUFx4f_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AND2x4_ASAP7_75t_L g655 ( .A(n_611), .B(n_630), .Y(n_655) );
BUFx6f_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
BUFx6f_ASAP7_75t_L g647 ( .A(n_612), .Y(n_647) );
BUFx6f_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
BUFx6f_ASAP7_75t_L g653 ( .A(n_615), .Y(n_653) );
CKINVDCx5p33_ASAP7_75t_R g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx2_ASAP7_75t_SL g621 ( .A(n_622), .Y(n_621) );
AND2x4_ASAP7_75t_L g629 ( .A(n_622), .B(n_630), .Y(n_629) );
BUFx6f_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
BUFx2_ASAP7_75t_L g644 ( .A(n_623), .Y(n_644) );
INVx1_ASAP7_75t_L g664 ( .A(n_624), .Y(n_664) );
BUFx6f_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
BUFx6f_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx2_ASAP7_75t_L g667 ( .A(n_627), .Y(n_667) );
INVx1_ASAP7_75t_L g663 ( .A(n_628), .Y(n_663) );
INVx2_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
OR2x2_ASAP7_75t_L g661 ( .A(n_631), .B(n_662), .Y(n_661) );
OR2x2_ASAP7_75t_L g666 ( .A(n_631), .B(n_667), .Y(n_666) );
INVx2_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
INVx2_ASAP7_75t_SL g708 ( .A(n_634), .Y(n_708) );
INVx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_L g704 ( .A(n_636), .Y(n_704) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx2_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
BUFx3_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
BUFx6f_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AND2x4_ASAP7_75t_L g656 ( .A(n_646), .B(n_657), .Y(n_656) );
BUFx6f_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx3_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
BUFx3_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx2_ASAP7_75t_SL g701 ( .A(n_650), .Y(n_701) );
INVx4_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
BUFx6f_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
INVx6_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
OR2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
INVx4_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
BUFx8_ASAP7_75t_SL g668 ( .A(n_669), .Y(n_668) );
INVx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
BUFx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_673), .B(n_674), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_673), .B(n_675), .Y(n_697) );
INVx1_ASAP7_75t_SL g720 ( .A(n_673), .Y(n_720) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_693), .B1(n_709), .B2(n_710), .Y(n_676) );
OAI22xp5_ASAP7_75t_L g714 ( .A1(n_677), .A2(n_709), .B1(n_715), .B2(n_716), .Y(n_714) );
AOI22xp5_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_682), .B1(n_691), .B2(n_692), .Y(n_677) );
INVx1_ASAP7_75t_L g691 ( .A(n_678), .Y(n_691) );
XNOR2xp5_ASAP7_75t_SL g678 ( .A(n_679), .B(n_681), .Y(n_678) );
CKINVDCx5p33_ASAP7_75t_R g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g692 ( .A(n_682), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_684), .B1(n_685), .B2(n_686), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
OAI22xp5_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_688), .B1(n_689), .B2(n_690), .Y(n_686) );
INVx1_ASAP7_75t_L g690 ( .A(n_687), .Y(n_690) );
CKINVDCx14_ASAP7_75t_R g688 ( .A(n_689), .Y(n_688) );
INVx8_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx8_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
CKINVDCx20_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
BUFx4f_ASAP7_75t_L g715 ( .A(n_696), .Y(n_715) );
OR2x6_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .Y(n_696) );
OR2x4_ASAP7_75t_L g712 ( .A(n_697), .B(n_699), .Y(n_712) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
AOI31xp33_ASAP7_75t_L g699 ( .A1(n_700), .A2(n_702), .A3(n_705), .B(n_707), .Y(n_699) );
BUFx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVxp67_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx6_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVxp67_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
BUFx6f_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx2_ASAP7_75t_L g716 ( .A(n_711), .Y(n_716) );
INVx8_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
BUFx2_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
endmodule