module fake_aes_3013_n_17 (n_1, n_2, n_0, n_17);
input n_1;
input n_2;
input n_0;
output n_17;
wire n_11;
wire n_13;
wire n_16;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_14;
wire n_7;
wire n_15;
wire n_10;
wire n_8;
INVx3_ASAP7_75t_L g3 ( .A(n_2), .Y(n_3) );
NAND2xp5_ASAP7_75t_SL g4 ( .A(n_2), .B(n_0), .Y(n_4) );
NAND2xp5_ASAP7_75t_SL g5 ( .A(n_0), .B(n_2), .Y(n_5) );
AOI211x1_ASAP7_75t_L g6 ( .A1(n_4), .A2(n_0), .B(n_1), .C(n_2), .Y(n_6) );
NAND3xp33_ASAP7_75t_L g7 ( .A(n_5), .B(n_0), .C(n_1), .Y(n_7) );
NAND2xp5_ASAP7_75t_L g8 ( .A(n_7), .B(n_3), .Y(n_8) );
INVx2_ASAP7_75t_L g9 ( .A(n_6), .Y(n_9) );
INVx2_ASAP7_75t_L g10 ( .A(n_8), .Y(n_10) );
NAND2xp5_ASAP7_75t_L g11 ( .A(n_9), .B(n_3), .Y(n_11) );
NOR2xp33_ASAP7_75t_L g12 ( .A(n_10), .B(n_0), .Y(n_12) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_11), .B(n_3), .Y(n_13) );
NOR2x1_ASAP7_75t_L g14 ( .A(n_12), .B(n_0), .Y(n_14) );
NOR2x1_ASAP7_75t_L g15 ( .A(n_13), .B(n_1), .Y(n_15) );
OAI22xp5_ASAP7_75t_SL g16 ( .A1(n_14), .A2(n_1), .B1(n_2), .B2(n_15), .Y(n_16) );
AOI22xp5_ASAP7_75t_SL g17 ( .A1(n_16), .A2(n_1), .B1(n_2), .B2(n_12), .Y(n_17) );
endmodule