module fake_jpeg_7083_n_317 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_33),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_42),
.Y(n_52)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx3_ASAP7_75t_SL g58 ( 
.A(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_17),
.B(n_16),
.Y(n_42)
);

HAxp5_ASAP7_75t_SL g43 ( 
.A(n_22),
.B(n_15),
.CON(n_43),
.SN(n_43)
);

NOR2xp67_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_17),
.Y(n_64)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_25),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_36),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_46),
.Y(n_75)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_48),
.B(n_54),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_28),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_SL g73 ( 
.A(n_49),
.B(n_40),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_43),
.A2(n_31),
.B1(n_21),
.B2(n_32),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_50),
.A2(n_60),
.B1(n_34),
.B2(n_26),
.Y(n_70)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_56),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_44),
.A2(n_34),
.B1(n_26),
.B2(n_22),
.Y(n_53)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_53),
.A2(n_64),
.B(n_28),
.C(n_20),
.Y(n_84)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_59),
.B(n_63),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_39),
.A2(n_31),
.B1(n_21),
.B2(n_32),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_44),
.A2(n_18),
.B1(n_32),
.B2(n_21),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_62),
.A2(n_23),
.B1(n_30),
.B2(n_34),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_23),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_35),
.B(n_33),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_65),
.B(n_66),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_35),
.B(n_33),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_35),
.B(n_30),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_67),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_70),
.B(n_79),
.Y(n_115)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_71),
.B(n_76),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_44),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_72),
.B(n_73),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_64),
.A2(n_39),
.B1(n_40),
.B2(n_38),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_74),
.A2(n_81),
.B1(n_91),
.B2(n_62),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g76 ( 
.A(n_68),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_56),
.A2(n_23),
.B1(n_30),
.B2(n_22),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_77),
.A2(n_84),
.B(n_85),
.Y(n_123)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

FAx1_ASAP7_75t_SL g79 ( 
.A(n_50),
.B(n_40),
.CI(n_38),
.CON(n_79),
.SN(n_79)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_49),
.A2(n_40),
.B1(n_38),
.B2(n_18),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_53),
.A2(n_31),
.B1(n_18),
.B2(n_26),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_82),
.A2(n_88),
.B1(n_53),
.B2(n_70),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_56),
.A2(n_28),
.B1(n_11),
.B2(n_14),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_87),
.Y(n_104)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_62),
.A2(n_38),
.B1(n_25),
.B2(n_28),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_55),
.A2(n_25),
.B1(n_28),
.B2(n_27),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_57),
.B(n_28),
.C(n_25),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_47),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_58),
.A2(n_28),
.B1(n_9),
.B2(n_10),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_93),
.Y(n_121)
);

AND2x2_ASAP7_75t_SL g95 ( 
.A(n_58),
.B(n_27),
.Y(n_95)
);

AOI32xp33_ASAP7_75t_L g103 ( 
.A1(n_95),
.A2(n_58),
.A3(n_68),
.B1(n_66),
.B2(n_65),
.Y(n_103)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_96),
.B(n_99),
.Y(n_127)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_76),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_100),
.A2(n_110),
.B1(n_118),
.B2(n_88),
.Y(n_124)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_101),
.B(n_106),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_60),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_102),
.B(n_105),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_SL g148 ( 
.A(n_103),
.B(n_119),
.C(n_120),
.Y(n_148)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_95),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_107),
.B(n_108),
.Y(n_152)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_89),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_109),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_86),
.Y(n_112)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_112),
.Y(n_133)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_113),
.Y(n_135)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_114),
.A2(n_90),
.B1(n_80),
.B2(n_75),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_116),
.B(n_73),
.C(n_92),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_84),
.A2(n_55),
.B1(n_59),
.B2(n_68),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_69),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_72),
.B(n_48),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_55),
.Y(n_122)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_122),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_124),
.A2(n_101),
.B1(n_106),
.B2(n_121),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_102),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_125),
.A2(n_141),
.B1(n_144),
.B2(n_145),
.Y(n_154)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_129),
.B(n_132),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_109),
.A2(n_84),
.B(n_77),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_100),
.A2(n_72),
.B1(n_79),
.B2(n_82),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_131),
.A2(n_142),
.B1(n_150),
.B2(n_83),
.Y(n_164)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_134),
.B(n_138),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_123),
.A2(n_79),
.B(n_74),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_136),
.Y(n_179)
);

XNOR2x1_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_73),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_140),
.C(n_108),
.Y(n_160)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_113),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_139),
.A2(n_146),
.B1(n_112),
.B2(n_107),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_115),
.A2(n_74),
.B1(n_70),
.B2(n_79),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_92),
.B1(n_75),
.B2(n_80),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_97),
.A2(n_81),
.B1(n_91),
.B2(n_55),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_117),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_97),
.A2(n_81),
.B1(n_59),
.B2(n_85),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_149),
.A2(n_67),
.B1(n_63),
.B2(n_51),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_110),
.A2(n_94),
.B1(n_83),
.B2(n_45),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_152),
.B(n_114),
.Y(n_153)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_153),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_125),
.B(n_105),
.Y(n_156)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_156),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_127),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_157),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_158),
.A2(n_161),
.B1(n_164),
.B2(n_167),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_160),
.B(n_163),
.C(n_171),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_124),
.A2(n_123),
.B1(n_117),
.B2(n_121),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_147),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_162),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_119),
.C(n_103),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_125),
.B(n_94),
.Y(n_165)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_165),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_46),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_166),
.A2(n_170),
.B(n_173),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_136),
.A2(n_51),
.B1(n_93),
.B2(n_54),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_150),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_168),
.B(n_169),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_144),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_46),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_69),
.C(n_54),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_141),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_172),
.B(n_180),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_58),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_151),
.B(n_104),
.C(n_98),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_178),
.C(n_149),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_133),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_175),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_176),
.A2(n_52),
.B1(n_45),
.B2(n_99),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_131),
.B(n_52),
.Y(n_178)
);

INVx13_ASAP7_75t_L g180 ( 
.A(n_132),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_145),
.B(n_48),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_181),
.A2(n_133),
.B1(n_138),
.B2(n_135),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_182),
.A2(n_183),
.B1(n_129),
.B2(n_146),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_128),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_148),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_195),
.C(n_198),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_154),
.B(n_130),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_207),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_190),
.B(n_173),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_155),
.A2(n_179),
.B(n_170),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_196),
.A2(n_197),
.B(n_199),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_155),
.A2(n_179),
.B(n_165),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_160),
.B(n_148),
.C(n_126),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_168),
.A2(n_126),
.B1(n_45),
.B2(n_96),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_200),
.A2(n_156),
.B1(n_161),
.B2(n_174),
.Y(n_226)
);

AOI21x1_ASAP7_75t_L g202 ( 
.A1(n_181),
.A2(n_133),
.B(n_24),
.Y(n_202)
);

OAI21xp33_ASAP7_75t_L g216 ( 
.A1(n_202),
.A2(n_204),
.B(n_157),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_172),
.A2(n_139),
.B1(n_135),
.B2(n_128),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_205),
.A2(n_206),
.B1(n_175),
.B2(n_159),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_158),
.A2(n_61),
.B1(n_27),
.B2(n_24),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_154),
.B(n_24),
.Y(n_207)
);

A2O1A1O1Ixp25_ASAP7_75t_L g209 ( 
.A1(n_164),
.A2(n_19),
.B(n_15),
.C(n_13),
.D(n_12),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_209),
.B(n_12),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_163),
.B(n_61),
.C(n_19),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_210),
.B(n_171),
.C(n_167),
.Y(n_222)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_204),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_211),
.B(n_212),
.Y(n_243)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_194),
.Y(n_212)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_205),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_214),
.B(n_221),
.Y(n_244)
);

INVx13_ASAP7_75t_L g215 ( 
.A(n_186),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_215),
.B(n_216),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_193),
.B(n_162),
.Y(n_219)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_219),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_220),
.A2(n_232),
.B(n_233),
.Y(n_239)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_199),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_227),
.C(n_231),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_223),
.A2(n_228),
.B1(n_202),
.B2(n_203),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_187),
.B(n_177),
.Y(n_224)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_224),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_188),
.B(n_180),
.Y(n_225)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_225),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_229),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_192),
.B(n_166),
.C(n_176),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_203),
.A2(n_173),
.B1(n_183),
.B2(n_61),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_183),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_201),
.B(n_13),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_230),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_192),
.B(n_61),
.C(n_19),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_200),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_191),
.B(n_0),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_190),
.B(n_13),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_234),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_235),
.A2(n_209),
.B1(n_206),
.B2(n_12),
.Y(n_255)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_237),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_189),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_240),
.B(n_241),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_217),
.B(n_185),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_198),
.C(n_195),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_242),
.B(n_250),
.C(n_253),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_211),
.A2(n_184),
.B1(n_197),
.B2(n_196),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_248),
.A2(n_249),
.B1(n_231),
.B2(n_233),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_214),
.A2(n_232),
.B1(n_213),
.B2(n_223),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_217),
.B(n_184),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_210),
.C(n_207),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_255),
.B(n_235),
.Y(n_260)
);

MAJx2_ASAP7_75t_L g256 ( 
.A(n_240),
.B(n_213),
.C(n_226),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_256),
.A2(n_265),
.B(n_253),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_243),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_266),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_252),
.B(n_219),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_258),
.A2(n_263),
.B(n_269),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_222),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_242),
.C(n_238),
.Y(n_273)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_260),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_244),
.A2(n_247),
.B(n_245),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_261),
.A2(n_270),
.B(n_215),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g262 ( 
.A(n_237),
.Y(n_262)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_262),
.Y(n_277)
);

INVxp33_ASAP7_75t_L g263 ( 
.A(n_239),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_248),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_264),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_236),
.A2(n_221),
.B1(n_212),
.B2(n_228),
.Y(n_265)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_239),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_249),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_276),
.C(n_279),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_254),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_238),
.C(n_250),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_261),
.A2(n_268),
.B(n_267),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_278),
.A2(n_281),
.B(n_283),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_251),
.C(n_255),
.Y(n_279)
);

NOR3xp33_ASAP7_75t_SL g280 ( 
.A(n_256),
.B(n_246),
.C(n_254),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_280),
.B(n_263),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_259),
.C(n_265),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_285),
.B(n_289),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_288),
.C(n_294),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_246),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_274),
.B(n_0),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_282),
.A2(n_11),
.B(n_10),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_290),
.B(n_291),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_0),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_272),
.B(n_9),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_292),
.B(n_293),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_1),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_276),
.B(n_1),
.Y(n_294)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_288),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_298),
.A2(n_301),
.B(n_303),
.Y(n_307)
);

AOI322xp5_ASAP7_75t_L g300 ( 
.A1(n_286),
.A2(n_280),
.A3(n_282),
.B1(n_279),
.B2(n_273),
.C1(n_5),
.C2(n_6),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_300),
.B(n_302),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_287),
.B(n_1),
.Y(n_301)
);

AOI322xp5_ASAP7_75t_L g302 ( 
.A1(n_294),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_5),
.C1(n_6),
.C2(n_7),
.Y(n_302)
);

AOI31xp67_ASAP7_75t_SL g303 ( 
.A1(n_295),
.A2(n_2),
.A3(n_3),
.B(n_4),
.Y(n_303)
);

A2O1A1Ixp33_ASAP7_75t_SL g306 ( 
.A1(n_298),
.A2(n_295),
.B(n_3),
.C(n_7),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_306),
.A2(n_7),
.B(n_8),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_296),
.B(n_2),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_308),
.A2(n_309),
.B(n_310),
.Y(n_311)
);

NAND2x1_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_2),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_299),
.B(n_3),
.Y(n_310)
);

OA21x2_ASAP7_75t_L g312 ( 
.A1(n_305),
.A2(n_297),
.B(n_304),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_312),
.B(n_313),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_307),
.C(n_306),
.Y(n_315)
);

OAI21xp33_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_311),
.B(n_7),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_8),
.Y(n_317)
);


endmodule