module fake_jpeg_30369_n_382 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_382);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_382;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_10),
.B(n_6),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_2),
.B(n_12),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx5p33_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

INVx6_ASAP7_75t_SL g41 ( 
.A(n_4),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_47),
.Y(n_94)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_21),
.B(n_9),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_52),
.Y(n_81)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_21),
.B(n_15),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_57),
.Y(n_84)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_56),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_31),
.B(n_14),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_31),
.B(n_13),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_58),
.B(n_68),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx5_ASAP7_75t_SL g97 ( 
.A(n_62),
.Y(n_97)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_17),
.B(n_13),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_64),
.B(n_69),
.Y(n_101)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_65),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_67),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_17),
.B(n_12),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_37),
.B(n_11),
.Y(n_69)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_70),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_72),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_74),
.Y(n_86)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_75),
.B(n_77),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_76),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_18),
.Y(n_77)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_78),
.B(n_26),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_79),
.B(n_26),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_60),
.A2(n_43),
.B1(n_28),
.B2(n_29),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_80),
.A2(n_112),
.B1(n_0),
.B2(n_1),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_56),
.A2(n_59),
.B1(n_44),
.B2(n_47),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_82),
.A2(n_45),
.B1(n_40),
.B2(n_35),
.Y(n_142)
);

NOR2x1_ASAP7_75t_L g90 ( 
.A(n_52),
.B(n_37),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_90),
.B(n_127),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_49),
.B(n_42),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_91),
.B(n_105),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_79),
.B(n_29),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_92),
.B(n_103),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_55),
.A2(n_41),
.B1(n_27),
.B2(n_33),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_99),
.A2(n_111),
.B1(n_114),
.B2(n_123),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_79),
.B(n_34),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_67),
.B(n_42),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_65),
.B(n_19),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_107),
.B(n_116),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_53),
.A2(n_33),
.B1(n_27),
.B2(n_35),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_78),
.A2(n_33),
.B1(n_27),
.B2(n_24),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_63),
.A2(n_33),
.B1(n_27),
.B2(n_35),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_66),
.B(n_19),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_119),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_52),
.B(n_28),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_61),
.B(n_34),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_120),
.B(n_0),
.Y(n_168)
);

BUFx12_ASAP7_75t_L g121 ( 
.A(n_70),
.Y(n_121)
);

INVx13_ASAP7_75t_L g165 ( 
.A(n_121),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_72),
.A2(n_33),
.B1(n_27),
.B2(n_35),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g172 ( 
.A(n_129),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_97),
.A2(n_48),
.B1(n_46),
.B2(n_51),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_130),
.A2(n_148),
.B1(n_93),
.B2(n_94),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_115),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_132),
.B(n_133),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_116),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_90),
.A2(n_39),
.B1(n_24),
.B2(n_25),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_134),
.A2(n_161),
.B(n_5),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_126),
.A2(n_77),
.B1(n_76),
.B2(n_74),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_136),
.A2(n_151),
.B1(n_157),
.B2(n_162),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_91),
.B(n_73),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_137),
.Y(n_183)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_83),
.Y(n_138)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_138),
.Y(n_178)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_83),
.Y(n_140)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_140),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_105),
.A2(n_39),
.B(n_25),
.C(n_10),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_141),
.B(n_145),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_142),
.A2(n_146),
.B1(n_150),
.B2(n_163),
.Y(n_176)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_143),
.Y(n_177)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_87),
.Y(n_144)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

O2A1O1Ixp33_ASAP7_75t_L g145 ( 
.A1(n_107),
.A2(n_100),
.B(n_127),
.C(n_110),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_108),
.A2(n_71),
.B1(n_62),
.B2(n_45),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_97),
.A2(n_40),
.B1(n_35),
.B2(n_26),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_89),
.Y(n_149)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_149),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_109),
.A2(n_40),
.B1(n_26),
.B2(n_4),
.Y(n_150)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_89),
.Y(n_153)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_153),
.Y(n_189)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_124),
.Y(n_154)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_154),
.Y(n_194)
);

BUFx12_ASAP7_75t_L g155 ( 
.A(n_121),
.Y(n_155)
);

INVx4_ASAP7_75t_SL g174 ( 
.A(n_155),
.Y(n_174)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_113),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_158),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_126),
.A2(n_40),
.B1(n_26),
.B2(n_4),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_117),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_81),
.B(n_40),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_159),
.B(n_167),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_112),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_164),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_86),
.A2(n_0),
.B(n_1),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_108),
.A2(n_8),
.B1(n_1),
.B2(n_4),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_162),
.A2(n_151),
.B1(n_133),
.B2(n_170),
.Y(n_192)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_85),
.A2(n_122),
.B1(n_113),
.B2(n_106),
.Y(n_163)
);

INVx4_ASAP7_75t_SL g164 ( 
.A(n_85),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_101),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_168),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_84),
.B(n_0),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_117),
.B(n_1),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_169),
.B(n_5),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_122),
.B(n_5),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_170),
.B(n_102),
.Y(n_202)
);

OAI21xp33_ASAP7_75t_SL g175 ( 
.A1(n_161),
.A2(n_104),
.B(n_106),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_175),
.A2(n_209),
.B(n_128),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_160),
.A2(n_94),
.B1(n_93),
.B2(n_86),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_182),
.A2(n_205),
.B1(n_164),
.B2(n_149),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_152),
.B(n_95),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_184),
.B(n_203),
.Y(n_239)
);

NAND3xp33_ASAP7_75t_L g186 ( 
.A(n_147),
.B(n_104),
.C(n_125),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_193),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_188),
.A2(n_192),
.B1(n_150),
.B2(n_144),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_139),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_190),
.B(n_191),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_134),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_195),
.A2(n_206),
.B(n_193),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_131),
.B(n_98),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_202),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_145),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_198),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_135),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_135),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_199),
.B(n_200),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_135),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_152),
.B(n_95),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_143),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_204),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_142),
.A2(n_102),
.B1(n_131),
.B2(n_137),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_147),
.B(n_125),
.C(n_98),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_208),
.B(n_121),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_137),
.A2(n_88),
.B(n_6),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_181),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_212),
.B(n_214),
.Y(n_245)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_178),
.Y(n_213)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_213),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_196),
.B(n_159),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_208),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_215),
.B(n_216),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_132),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_181),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_217),
.B(n_221),
.Y(n_264)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_178),
.Y(n_219)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_219),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_220),
.A2(n_224),
.B1(n_228),
.B2(n_232),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_173),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_201),
.B(n_167),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_222),
.B(n_230),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_223),
.A2(n_225),
.B(n_238),
.Y(n_250)
);

OAI22x1_ASAP7_75t_L g225 ( 
.A1(n_175),
.A2(n_141),
.B1(n_165),
.B2(n_96),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_173),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_226),
.B(n_229),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_205),
.A2(n_140),
.B1(n_153),
.B2(n_138),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_192),
.B(n_156),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_201),
.B(n_166),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_172),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_231),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_185),
.A2(n_154),
.B1(n_144),
.B2(n_164),
.Y(n_232)
);

AO22x1_ASAP7_75t_L g233 ( 
.A1(n_185),
.A2(n_186),
.B1(n_171),
.B2(n_183),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_236),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_242),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_158),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_234),
.C(n_215),
.Y(n_257)
);

NAND2x1p5_ASAP7_75t_L g236 ( 
.A(n_171),
.B(n_88),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_176),
.A2(n_129),
.B1(n_96),
.B2(n_165),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_237),
.A2(n_188),
.B1(n_172),
.B2(n_180),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_206),
.B(n_129),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_179),
.Y(n_243)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_243),
.Y(n_247)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_179),
.Y(n_244)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_244),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_221),
.Y(n_252)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_252),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_223),
.A2(n_195),
.B(n_203),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_253),
.Y(n_297)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_213),
.Y(n_256)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_256),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_271),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_233),
.A2(n_191),
.B(n_184),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_262),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_239),
.B(n_187),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_241),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_233),
.A2(n_176),
.B(n_187),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_219),
.Y(n_263)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_263),
.Y(n_292)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_243),
.Y(n_265)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_265),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_266),
.A2(n_172),
.B1(n_177),
.B2(n_194),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_216),
.B(n_182),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_235),
.C(n_214),
.Y(n_285)
);

INVx2_ASAP7_75t_SL g268 ( 
.A(n_231),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_268),
.B(n_272),
.Y(n_277)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_244),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_270),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_242),
.A2(n_207),
.B(n_189),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_228),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_237),
.A2(n_207),
.B1(n_189),
.B2(n_180),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_274),
.A2(n_232),
.B1(n_217),
.B2(n_224),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_272),
.A2(n_226),
.B1(n_225),
.B2(n_220),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_278),
.A2(n_279),
.B1(n_296),
.B2(n_274),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_267),
.A2(n_218),
.B1(n_241),
.B2(n_212),
.Y(n_279)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_280),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_262),
.A2(n_249),
.B1(n_229),
.B2(n_251),
.Y(n_283)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_283),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_284),
.B(n_269),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_285),
.B(n_271),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_264),
.B(n_240),
.Y(n_286)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_286),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_257),
.B(n_210),
.C(n_230),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_255),
.C(n_258),
.Y(n_299)
);

AOI221xp5_ASAP7_75t_L g288 ( 
.A1(n_259),
.A2(n_238),
.B1(n_227),
.B2(n_236),
.C(n_210),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_249),
.Y(n_309)
);

AOI322xp5_ASAP7_75t_L g289 ( 
.A1(n_250),
.A2(n_236),
.A3(n_222),
.B1(n_211),
.B2(n_165),
.C1(n_177),
.C2(n_194),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_250),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_211),
.Y(n_290)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_290),
.Y(n_307)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_291),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_245),
.B(n_174),
.Y(n_293)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_293),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_261),
.A2(n_174),
.B1(n_6),
.B2(n_7),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_255),
.B(n_174),
.Y(n_298)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_298),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_299),
.B(n_300),
.C(n_304),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_258),
.C(n_261),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_301),
.B(n_305),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_302),
.A2(n_279),
.B1(n_278),
.B2(n_297),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_276),
.B(n_261),
.C(n_253),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_248),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_314),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_310),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_285),
.B(n_266),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_311),
.A2(n_294),
.B1(n_295),
.B2(n_292),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_282),
.B(n_247),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_313),
.Y(n_331)
);

XOR2x2_ASAP7_75t_L g314 ( 
.A(n_275),
.B(n_247),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_298),
.B(n_254),
.C(n_265),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_318),
.B(n_293),
.C(n_283),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_299),
.B(n_275),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_321),
.B(n_334),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_323),
.B(n_310),
.C(n_308),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_324),
.B(n_335),
.C(n_318),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_303),
.A2(n_290),
.B1(n_296),
.B2(n_277),
.Y(n_325)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_325),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_303),
.A2(n_277),
.B1(n_297),
.B2(n_294),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_326),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g327 ( 
.A1(n_309),
.A2(n_307),
.B(n_315),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_327),
.A2(n_306),
.B(n_312),
.Y(n_346)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_307),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_329),
.B(n_330),
.Y(n_340)
);

O2A1O1Ixp33_ASAP7_75t_L g330 ( 
.A1(n_315),
.A2(n_280),
.B(n_292),
.C(n_281),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_306),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_332),
.B(n_333),
.Y(n_343)
);

NOR3xp33_ASAP7_75t_SL g334 ( 
.A(n_301),
.B(n_295),
.C(n_281),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_300),
.B(n_246),
.C(n_263),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_337),
.B(n_344),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_338),
.B(n_339),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_321),
.B(n_304),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_322),
.B(n_335),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_322),
.B(n_317),
.C(n_314),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_345),
.B(n_347),
.C(n_319),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_346),
.B(n_348),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_319),
.B(n_316),
.C(n_312),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_SL g348 ( 
.A(n_320),
.B(n_316),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_342),
.A2(n_329),
.B1(n_333),
.B2(n_324),
.Y(n_349)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_349),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_342),
.A2(n_330),
.B1(n_327),
.B2(n_334),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_350),
.B(n_353),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_351),
.B(n_155),
.C(n_6),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_336),
.A2(n_331),
.B1(n_328),
.B2(n_254),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_338),
.B(n_320),
.C(n_331),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_354),
.B(n_356),
.C(n_352),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_340),
.A2(n_343),
.B(n_347),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_355),
.B(n_357),
.Y(n_366)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_341),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_354),
.B(n_339),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_360),
.B(n_361),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_356),
.B(n_348),
.C(n_268),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_362),
.A2(n_358),
.B(n_7),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_355),
.A2(n_270),
.B1(n_256),
.B2(n_246),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_363),
.B(n_364),
.Y(n_374)
);

O2A1O1Ixp33_ASAP7_75t_L g364 ( 
.A1(n_350),
.A2(n_268),
.B(n_155),
.C(n_7),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_365),
.B(n_351),
.C(n_349),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_369),
.B(n_372),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_370),
.B(n_373),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g371 ( 
.A1(n_361),
.A2(n_366),
.B(n_359),
.Y(n_371)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_371),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_367),
.B(n_358),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_362),
.B(n_155),
.C(n_5),
.Y(n_373)
);

AOI21x1_ASAP7_75t_L g375 ( 
.A1(n_368),
.A2(n_364),
.B(n_8),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_375),
.A2(n_374),
.B(n_377),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_379),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_376),
.A2(n_378),
.B(n_374),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_381),
.B(n_380),
.Y(n_382)
);


endmodule