module fake_jpeg_7075_n_339 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_36),
.Y(n_51)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_37),
.B(n_39),
.Y(n_54)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_38),
.B(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_23),
.B(n_7),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_44),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_43),
.B(n_23),
.Y(n_56)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_26),
.Y(n_64)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_46),
.B(n_49),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_27),
.B1(n_32),
.B2(n_19),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_47),
.A2(n_50),
.B1(n_72),
.B2(n_30),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_38),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_60),
.Y(n_74)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_38),
.A2(n_27),
.B1(n_23),
.B2(n_30),
.Y(n_50)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_52),
.B(n_55),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_56),
.B(n_59),
.Y(n_87)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_28),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_64),
.B(n_67),
.Y(n_95)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_35),
.B(n_32),
.C(n_20),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_70),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_43),
.B(n_30),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_69),
.A2(n_33),
.B(n_29),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_38),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_69),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_34),
.A2(n_27),
.B1(n_20),
.B2(n_18),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_35),
.B(n_18),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_19),
.Y(n_93)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_56),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_77),
.Y(n_128)
);

NAND2xp33_ASAP7_75t_SL g78 ( 
.A(n_73),
.B(n_28),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_78),
.A2(n_84),
.B(n_92),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_80),
.A2(n_49),
.B1(n_14),
.B2(n_9),
.Y(n_116)
);

BUFx12_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_81),
.Y(n_102)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_66),
.B(n_35),
.Y(n_84)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_88),
.Y(n_113)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_91),
.Y(n_127)
);

AND2x2_ASAP7_75t_SL g92 ( 
.A(n_73),
.B(n_41),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_54),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_62),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_94),
.B(n_96),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_60),
.A2(n_44),
.B(n_33),
.C(n_16),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_97),
.B(n_93),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_54),
.B(n_16),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_57),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_92),
.A2(n_44),
.B1(n_55),
.B2(n_59),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_100),
.A2(n_115),
.B1(n_121),
.B2(n_84),
.Y(n_130)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_104),
.B(n_107),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_106),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_98),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_110),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_51),
.C(n_68),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_109),
.B(n_97),
.C(n_94),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_71),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_96),
.A2(n_65),
.B1(n_58),
.B2(n_52),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_111),
.A2(n_116),
.B1(n_125),
.B2(n_93),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_112),
.B(n_122),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_76),
.A2(n_61),
.B1(n_67),
.B2(n_70),
.Y(n_115)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_118),
.B(n_119),
.Y(n_150)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_95),
.B(n_16),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_74),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_92),
.A2(n_41),
.B1(n_26),
.B2(n_21),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_123),
.A2(n_95),
.B(n_78),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_92),
.A2(n_48),
.B1(n_13),
.B2(n_8),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_124),
.A2(n_84),
.B(n_83),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_77),
.A2(n_41),
.B1(n_31),
.B2(n_22),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_81),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_126),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_129),
.B(n_139),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_130),
.A2(n_149),
.B1(n_151),
.B2(n_126),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_128),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_131),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_132),
.B(n_133),
.C(n_155),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_108),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_101),
.A2(n_84),
.B1(n_74),
.B2(n_76),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_134),
.Y(n_170)
);

BUFx24_ASAP7_75t_SL g137 ( 
.A(n_103),
.Y(n_137)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_137),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_138),
.A2(n_147),
.B1(n_146),
.B2(n_152),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_74),
.Y(n_140)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_140),
.Y(n_169)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_142),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_103),
.B(n_76),
.Y(n_143)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_143),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_128),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_144),
.Y(n_165)
);

A2O1A1Ixp33_ASAP7_75t_SL g146 ( 
.A1(n_111),
.A2(n_31),
.B(n_22),
.C(n_16),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_146),
.A2(n_156),
.B(n_29),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_118),
.A2(n_119),
.B1(n_117),
.B2(n_115),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_148),
.A2(n_153),
.B(n_141),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_109),
.A2(n_79),
.B1(n_90),
.B2(n_88),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_120),
.A2(n_79),
.B1(n_90),
.B2(n_86),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_112),
.Y(n_152)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_112),
.Y(n_153)
);

BUFx24_ASAP7_75t_L g178 ( 
.A(n_153),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_102),
.B(n_91),
.C(n_81),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_91),
.C(n_81),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_147),
.A2(n_106),
.B1(n_107),
.B2(n_86),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_158),
.B(n_162),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_129),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_160),
.A2(n_175),
.B(n_180),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_142),
.A2(n_89),
.B1(n_105),
.B2(n_104),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_163),
.A2(n_168),
.B1(n_171),
.B2(n_174),
.Y(n_185)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_164),
.B(n_179),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_133),
.B(n_16),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_166),
.A2(n_167),
.B(n_146),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_130),
.A2(n_105),
.B1(n_113),
.B2(n_63),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_149),
.A2(n_143),
.B1(n_132),
.B2(n_140),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_135),
.A2(n_113),
.B1(n_31),
.B2(n_22),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_138),
.A2(n_91),
.B(n_29),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_135),
.A2(n_22),
.B1(n_31),
.B2(n_26),
.Y(n_176)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_176),
.Y(n_187)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_136),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_148),
.A2(n_0),
.B(n_1),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_145),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_181),
.B(n_150),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_139),
.A2(n_26),
.B1(n_24),
.B2(n_114),
.Y(n_184)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_184),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_161),
.B(n_151),
.Y(n_186)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_186),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_134),
.Y(n_188)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_188),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_SL g224 ( 
.A(n_189),
.B(n_209),
.C(n_176),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_165),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_192),
.B(n_193),
.Y(n_233)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_164),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_162),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_194),
.B(n_199),
.Y(n_218)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_195),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_173),
.Y(n_196)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_196),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_155),
.C(n_156),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_197),
.B(n_202),
.C(n_203),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_198),
.A2(n_208),
.B(n_167),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_177),
.B(n_154),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_174),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_200),
.B(n_201),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_168),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_183),
.B(n_146),
.C(n_154),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_171),
.B(n_146),
.C(n_127),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_179),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_204),
.B(n_182),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_173),
.B(n_0),
.Y(n_206)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_206),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_158),
.B(n_24),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_157),
.B(n_1),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_160),
.B(n_127),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_210),
.B(n_175),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_178),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_211),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_194),
.A2(n_163),
.B1(n_170),
.B2(n_172),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_212),
.A2(n_215),
.B1(n_208),
.B2(n_231),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_189),
.B(n_166),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_216),
.Y(n_243)
);

OAI22xp33_ASAP7_75t_L g217 ( 
.A1(n_201),
.A2(n_172),
.B1(n_170),
.B2(n_180),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_217),
.A2(n_226),
.B1(n_191),
.B2(n_208),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_207),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_220),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_166),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_234),
.C(n_236),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_224),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_193),
.Y(n_227)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_227),
.Y(n_238)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_228),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_198),
.A2(n_182),
.B(n_178),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_205),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_185),
.A2(n_178),
.B1(n_184),
.B2(n_114),
.Y(n_230)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_230),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_210),
.B(n_24),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_192),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_235),
.B(n_196),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_202),
.B(n_188),
.C(n_203),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_205),
.B(n_24),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_237),
.B(n_236),
.C(n_225),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_255),
.C(n_256),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_241),
.A2(n_244),
.B(n_254),
.Y(n_264)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_233),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_245),
.B(n_247),
.Y(n_278)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_218),
.Y(n_247)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_213),
.B(n_206),
.Y(n_250)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_250),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_219),
.B(n_211),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_251),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_209),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_253),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_223),
.B(n_200),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_221),
.C(n_216),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_234),
.B(n_190),
.C(n_191),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_222),
.B(n_187),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_260),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_230),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_259),
.B(n_229),
.Y(n_263)
);

BUFx24_ASAP7_75t_SL g260 ( 
.A(n_237),
.Y(n_260)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_263),
.Y(n_280)
);

XNOR2x1_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_214),
.Y(n_266)
);

XNOR2x1_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_239),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_253),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_269),
.A2(n_270),
.B(n_271),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_212),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_241),
.A2(n_226),
.B(n_217),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_259),
.A2(n_248),
.B1(n_256),
.B2(n_240),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_272),
.A2(n_275),
.B1(n_265),
.B2(n_262),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_243),
.B(n_224),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_279),
.C(n_2),
.Y(n_292)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_238),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_261),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_242),
.B(n_187),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_277),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_252),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_243),
.B(n_255),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_285),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_263),
.A2(n_248),
.B1(n_246),
.B2(n_238),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_283),
.A2(n_291),
.B1(n_264),
.B2(n_2),
.Y(n_303)
);

CKINVDCx14_ASAP7_75t_R g299 ( 
.A(n_284),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_239),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_246),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_286),
.B(n_287),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_227),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_268),
.B(n_8),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_288),
.B(n_294),
.Y(n_297)
);

OR2x2_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_269),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_262),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_272),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_295),
.C(n_271),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_266),
.B(n_9),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_278),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_265),
.B(n_2),
.C(n_3),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_300),
.B(n_293),
.Y(n_315)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_301),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_302),
.A2(n_303),
.B(n_10),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_280),
.B(n_264),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_304),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_279),
.C(n_5),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_307),
.C(n_309),
.Y(n_318)
);

INVx11_ASAP7_75t_L g306 ( 
.A(n_289),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_306),
.B(n_308),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_281),
.B(n_4),
.C(n_5),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_285),
.B(n_4),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_282),
.B(n_5),
.C(n_6),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_290),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_312),
.A2(n_313),
.B(n_314),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_299),
.B(n_283),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_297),
.B(n_295),
.Y(n_314)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_315),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_296),
.B(n_307),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_317),
.B(n_305),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_296),
.B(n_6),
.C(n_7),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g324 ( 
.A1(n_319),
.A2(n_320),
.B(n_309),
.Y(n_324)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_311),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_322),
.A2(n_325),
.B(n_326),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_323),
.B(n_327),
.C(n_302),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_324),
.Y(n_331)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_319),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_316),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_318),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_330),
.B(n_332),
.C(n_333),
.Y(n_335)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_321),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_323),
.B(n_318),
.C(n_310),
.Y(n_333)
);

O2A1O1Ixp33_ASAP7_75t_SL g334 ( 
.A1(n_331),
.A2(n_306),
.B(n_317),
.C(n_328),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_334),
.A2(n_329),
.B(n_11),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_336),
.A2(n_10),
.B(n_11),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_337),
.A2(n_335),
.B(n_13),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_15),
.B1(n_11),
.B2(n_14),
.Y(n_339)
);


endmodule