module fake_jpeg_9233_n_249 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_249);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_249;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_37),
.Y(n_58)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_38),
.B(n_44),
.Y(n_50)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

CKINVDCx6p67_ASAP7_75t_R g60 ( 
.A(n_40),
.Y(n_60)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_19),
.B(n_1),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_41),
.A2(n_34),
.B1(n_23),
.B2(n_32),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_45),
.A2(n_53),
.B1(n_54),
.B2(n_64),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_44),
.A2(n_26),
.B1(n_28),
.B2(n_24),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_42),
.Y(n_68)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_65),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_26),
.B1(n_34),
.B2(n_32),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_34),
.B1(n_23),
.B2(n_24),
.Y(n_54)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_44),
.B(n_22),
.Y(n_57)
);

OAI21xp33_ASAP7_75t_L g84 ( 
.A1(n_57),
.A2(n_37),
.B(n_35),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_44),
.B(n_27),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_62),
.Y(n_67)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_27),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_44),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_36),
.A2(n_20),
.B1(n_19),
.B2(n_22),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_60),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_66),
.B(n_70),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_68),
.B(n_83),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_38),
.C(n_43),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_69),
.B(n_71),
.C(n_86),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_50),
.C(n_57),
.Y(n_71)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_72),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_52),
.A2(n_36),
.B1(n_39),
.B2(n_20),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_52),
.A2(n_39),
.B1(n_36),
.B2(n_38),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_49),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_79),
.B(n_89),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

O2A1O1Ixp33_ASAP7_75t_L g111 ( 
.A1(n_82),
.A2(n_29),
.B(n_40),
.C(n_46),
.Y(n_111)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_84),
.A2(n_85),
.B1(n_31),
.B2(n_18),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_62),
.A2(n_39),
.B1(n_38),
.B2(n_43),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_88),
.Y(n_100)
);

AO22x2_ASAP7_75t_L g93 ( 
.A1(n_82),
.A2(n_49),
.B1(n_56),
.B2(n_51),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_93),
.A2(n_111),
.B1(n_40),
.B2(n_73),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_86),
.A2(n_58),
.B(n_55),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_94),
.A2(n_96),
.B(n_104),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_67),
.A2(n_58),
.B(n_55),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_103),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_75),
.A2(n_39),
.B1(n_65),
.B2(n_33),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_101),
.A2(n_93),
.B1(n_109),
.B2(n_110),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_67),
.B(n_37),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_69),
.A2(n_35),
.B(n_29),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_27),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_108),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_27),
.Y(n_108)
);

AO22x1_ASAP7_75t_L g112 ( 
.A1(n_87),
.A2(n_40),
.B1(n_33),
.B2(n_31),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_115),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_113),
.A2(n_92),
.B(n_95),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_68),
.B(n_1),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_93),
.A2(n_90),
.B1(n_79),
.B2(n_72),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_116),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_95),
.A2(n_92),
.B(n_97),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_117),
.A2(n_120),
.B(n_134),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_93),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_119),
.B(n_121),
.Y(n_145)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_81),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_123),
.B(n_126),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_90),
.C(n_77),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_138),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_25),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_129),
.B(n_130),
.Y(n_152)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_101),
.Y(n_130)
);

OAI21xp33_ASAP7_75t_L g131 ( 
.A1(n_108),
.A2(n_1),
.B(n_2),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_131),
.B(n_2),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_93),
.A2(n_80),
.B1(n_70),
.B2(n_88),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_132),
.A2(n_139),
.B1(n_110),
.B2(n_109),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_96),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_133),
.B(n_112),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_94),
.B(n_78),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_136),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_78),
.Y(n_136)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_137),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_31),
.C(n_18),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_111),
.A2(n_18),
.B1(n_25),
.B2(n_5),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_99),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_151),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_123),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_144),
.B(n_148),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_146),
.A2(n_130),
.B1(n_119),
.B2(n_121),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_118),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_118),
.B(n_104),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_139),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_99),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_150),
.A2(n_158),
.B(n_160),
.Y(n_169)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_122),
.B(n_99),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_154),
.B(n_157),
.Y(n_178)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_132),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_126),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_161),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_127),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_137),
.Y(n_162)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_162),
.Y(n_168)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_134),
.Y(n_163)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_163),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_164),
.A2(n_167),
.B1(n_170),
.B2(n_180),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_165),
.A2(n_157),
.B(n_163),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_162),
.A2(n_119),
.B1(n_120),
.B2(n_136),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_155),
.A2(n_125),
.B1(n_124),
.B2(n_117),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_152),
.Y(n_171)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_171),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_142),
.Y(n_172)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_172),
.Y(n_187)
);

AOI322xp5_ASAP7_75t_SL g174 ( 
.A1(n_158),
.A2(n_128),
.A3(n_124),
.B1(n_138),
.B2(n_15),
.C1(n_16),
.C2(n_14),
.Y(n_174)
);

AOI322xp5_ASAP7_75t_L g189 ( 
.A1(n_174),
.A2(n_148),
.A3(n_150),
.B1(n_144),
.B2(n_15),
.C1(n_14),
.C2(n_10),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_147),
.B(n_128),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_183),
.C(n_156),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_142),
.Y(n_177)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_177),
.Y(n_190)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_145),
.Y(n_179)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_179),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_153),
.A2(n_112),
.B1(n_100),
.B2(n_102),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_140),
.Y(n_181)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_181),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_153),
.A2(n_105),
.B1(n_25),
.B2(n_6),
.Y(n_182)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_182),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_147),
.B(n_105),
.C(n_25),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_176),
.B(n_156),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_185),
.B(n_192),
.C(n_193),
.Y(n_213)
);

NAND4xp25_ASAP7_75t_SL g188 ( 
.A(n_175),
.B(n_141),
.C(n_161),
.D(n_159),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_173),
.Y(n_208)
);

NOR3xp33_ASAP7_75t_L g209 ( 
.A(n_189),
.B(n_201),
.C(n_196),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_168),
.A2(n_178),
.B1(n_177),
.B2(n_172),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_191),
.A2(n_180),
.B1(n_169),
.B2(n_166),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_167),
.B(n_154),
.Y(n_193)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_195),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_151),
.C(n_143),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_196),
.B(n_201),
.Y(n_202)
);

OAI31xp33_ASAP7_75t_L g200 ( 
.A1(n_178),
.A2(n_150),
.A3(n_146),
.B(n_149),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_200),
.A2(n_166),
.B1(n_164),
.B2(n_169),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_140),
.C(n_141),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_181),
.Y(n_203)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_203),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_186),
.B(n_171),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_206),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_197),
.B(n_184),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_207),
.A2(n_214),
.B(n_193),
.Y(n_221)
);

OR2x2_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_209),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_210),
.A2(n_211),
.B1(n_199),
.B2(n_194),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_198),
.A2(n_165),
.B1(n_5),
.B2(n_6),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_3),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_212),
.B(n_211),
.Y(n_218)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_188),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_205),
.A2(n_190),
.B1(n_187),
.B2(n_200),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_215),
.A2(n_213),
.B1(n_11),
.B2(n_12),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_203),
.A2(n_195),
.B(n_192),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_217),
.A2(n_210),
.B(n_213),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_218),
.B(n_223),
.Y(n_231)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_219),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_221),
.B(n_224),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_3),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_202),
.B(n_7),
.C(n_8),
.Y(n_224)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_225),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_212),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_227),
.B(n_223),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_229),
.Y(n_234)
);

OAI21x1_ASAP7_75t_L g229 ( 
.A1(n_220),
.A2(n_218),
.B(n_224),
.Y(n_229)
);

INVx11_ASAP7_75t_L g232 ( 
.A(n_216),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_232),
.B(n_222),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_225),
.B(n_217),
.C(n_231),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_235),
.B(n_231),
.C(n_226),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_236),
.A2(n_237),
.B(n_230),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_215),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_238),
.B(n_228),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_239),
.B(n_241),
.C(n_242),
.Y(n_245)
);

INVx13_ASAP7_75t_L g240 ( 
.A(n_234),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_240),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_239),
.A2(n_233),
.B(n_235),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_244),
.B(n_13),
.C(n_7),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_243),
.A2(n_240),
.B1(n_241),
.B2(n_13),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_246),
.A2(n_247),
.B1(n_245),
.B2(n_7),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_248),
.B(n_12),
.Y(n_249)
);


endmodule