module fake_jpeg_5386_n_44 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_44);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_44;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx12f_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_6),
.Y(n_9)
);

AND2x2_ASAP7_75t_SL g10 ( 
.A(n_3),
.B(n_6),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_2),
.B(n_4),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_9),
.B(n_0),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_16),
.B(n_21),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_19),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_15),
.A2(n_0),
.B1(n_1),
.B2(n_14),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_18),
.A2(n_12),
.B1(n_13),
.B2(n_20),
.Y(n_25)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

O2A1O1Ixp33_ASAP7_75t_L g20 ( 
.A1(n_10),
.A2(n_0),
.B(n_1),
.C(n_14),
.Y(n_20)
);

XNOR2x1_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_24),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_15),
.B(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_17),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_7),
.B(n_12),
.C(n_8),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_13),
.C(n_22),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_12),
.B(n_8),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_25),
.A2(n_27),
.B1(n_32),
.B2(n_26),
.Y(n_39)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_30),
.C(n_26),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_17),
.B(n_23),
.C(n_24),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_32),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_30),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_35),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_26),
.A2(n_25),
.B1(n_31),
.B2(n_29),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_34),
.Y(n_42)
);

AOI31xp67_ASAP7_75t_L g40 ( 
.A1(n_39),
.A2(n_28),
.A3(n_35),
.B(n_37),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_40),
.A2(n_42),
.B1(n_36),
.B2(n_38),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_41),
.Y(n_44)
);


endmodule