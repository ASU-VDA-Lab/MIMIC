module fake_jpeg_26961_n_251 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_251);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_251;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_14),
.B(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx1_ASAP7_75t_SL g45 ( 
.A(n_33),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_41),
.Y(n_47)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_35),
.B(n_38),
.Y(n_44)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_21),
.B(n_9),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_42),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_40),
.A2(n_32),
.B1(n_21),
.B2(n_31),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_46),
.A2(n_58),
.B1(n_30),
.B2(n_19),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_32),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_53),
.Y(n_65)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_30),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_56),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_35),
.B(n_19),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_57),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_35),
.A2(n_31),
.B1(n_24),
.B2(n_28),
.Y(n_58)
);

NAND2xp33_ASAP7_75t_SL g59 ( 
.A(n_54),
.B(n_39),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_59),
.B(n_74),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_47),
.B(n_34),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_60),
.B(n_61),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_38),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_55),
.B(n_34),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_66),
.Y(n_92)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_63),
.Y(n_98)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_64),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_49),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_43),
.A2(n_31),
.B1(n_16),
.B2(n_28),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_52),
.A2(n_39),
.B(n_1),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_18),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_56),
.A2(n_33),
.B1(n_40),
.B2(n_36),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_71),
.A2(n_78),
.B1(n_57),
.B2(n_43),
.Y(n_86)
);

CKINVDCx9p33_ASAP7_75t_R g73 ( 
.A(n_45),
.Y(n_73)
);

INVx6_ASAP7_75t_SL g101 ( 
.A(n_73),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_38),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_83),
.Y(n_96)
);

AO22x2_ASAP7_75t_L g78 ( 
.A1(n_51),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_42),
.Y(n_80)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_53),
.A2(n_38),
.B(n_35),
.C(n_34),
.Y(n_81)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_22),
.Y(n_95)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

OR2x2_ASAP7_75t_SL g83 ( 
.A(n_50),
.B(n_27),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g84 ( 
.A(n_54),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_49),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_86),
.A2(n_70),
.B(n_66),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_88),
.B(n_95),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_65),
.A2(n_57),
.B1(n_43),
.B2(n_33),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_89),
.A2(n_93),
.B1(n_78),
.B2(n_75),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_71),
.A2(n_33),
.B1(n_36),
.B2(n_37),
.Y(n_93)
);

AND2x6_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_68),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_97),
.B(n_108),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_65),
.B(n_48),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_102),
.B(n_109),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_78),
.A2(n_36),
.B1(n_25),
.B2(n_24),
.Y(n_103)
);

OAI21xp33_ASAP7_75t_L g128 ( 
.A1(n_103),
.A2(n_107),
.B(n_0),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_78),
.A2(n_25),
.B1(n_27),
.B2(n_18),
.Y(n_107)
);

AND2x6_ASAP7_75t_L g108 ( 
.A(n_78),
.B(n_11),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_77),
.B(n_48),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_111),
.B(n_112),
.Y(n_160)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_83),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_113),
.B(n_125),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_110),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_117),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_69),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_116),
.B(n_129),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_110),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_118),
.A2(n_86),
.B1(n_93),
.B2(n_94),
.Y(n_140)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_104),
.Y(n_119)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_63),
.C(n_77),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_120),
.B(n_90),
.C(n_23),
.Y(n_146)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_122),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_91),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_131),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_64),
.Y(n_125)
);

OAI32xp33_ASAP7_75t_L g126 ( 
.A1(n_97),
.A2(n_59),
.A3(n_22),
.B1(n_73),
.B2(n_75),
.Y(n_126)
);

OAI32xp33_ASAP7_75t_L g148 ( 
.A1(n_126),
.A2(n_131),
.A3(n_115),
.B1(n_117),
.B2(n_111),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_84),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_127),
.B(n_134),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_128),
.A2(n_133),
.B1(n_100),
.B2(n_101),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_98),
.B(n_26),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_88),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_96),
.B(n_70),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_105),
.A2(n_85),
.B(n_1),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_135),
.A2(n_87),
.B(n_90),
.Y(n_149)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g145 ( 
.A(n_136),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_114),
.A2(n_105),
.B(n_94),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_137),
.A2(n_141),
.B(n_143),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_140),
.A2(n_154),
.B1(n_155),
.B2(n_23),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_133),
.A2(n_100),
.B(n_108),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_98),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_142),
.B(n_144),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_100),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_146),
.B(n_48),
.C(n_132),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_135),
.A2(n_104),
.B(n_1),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_147),
.A2(n_148),
.B(n_0),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_149),
.A2(n_159),
.B(n_23),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_112),
.A2(n_79),
.B1(n_101),
.B2(n_72),
.Y(n_151)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_151),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_72),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_157),
.Y(n_163)
);

AO22x1_ASAP7_75t_L g153 ( 
.A1(n_118),
.A2(n_79),
.B1(n_80),
.B2(n_72),
.Y(n_153)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_130),
.A2(n_126),
.B1(n_121),
.B2(n_129),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_121),
.A2(n_124),
.B1(n_123),
.B2(n_136),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_124),
.B(n_80),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_132),
.A2(n_26),
.B(n_20),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_173),
.C(n_146),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_162),
.B(n_26),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_165),
.B(n_177),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_149),
.A2(n_119),
.B(n_122),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_169),
.A2(n_170),
.B(n_183),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_145),
.Y(n_171)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_171),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_161),
.B(n_20),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_172),
.B(n_144),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_23),
.C(n_20),
.Y(n_173)
);

INVx13_ASAP7_75t_L g174 ( 
.A(n_145),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_174),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_176),
.A2(n_184),
.B1(n_143),
.B2(n_151),
.Y(n_188)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_138),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_150),
.B(n_9),
.Y(n_178)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_178),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_138),
.Y(n_179)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_179),
.Y(n_191)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_180),
.Y(n_195)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_155),
.Y(n_181)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_181),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_160),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_182),
.A2(n_159),
.B1(n_158),
.B2(n_156),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_147),
.A2(n_0),
.B(n_2),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_186),
.B(n_164),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_187),
.B(n_192),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_182),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_168),
.B(n_142),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_168),
.B(n_154),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_187),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_181),
.A2(n_140),
.B1(n_148),
.B2(n_153),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_194),
.A2(n_175),
.B1(n_170),
.B2(n_167),
.Y(n_206)
);

OAI222xp33_ASAP7_75t_L g198 ( 
.A1(n_183),
.A2(n_141),
.B1(n_137),
.B2(n_157),
.C1(n_139),
.C2(n_153),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_198),
.A2(n_176),
.B1(n_199),
.B2(n_194),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_200),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_172),
.B(n_158),
.C(n_3),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_201),
.B(n_184),
.C(n_173),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_202),
.B(n_212),
.C(n_193),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_203),
.B(n_163),
.Y(n_221)
);

OR2x2_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_207),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_206),
.A2(n_208),
.B1(n_211),
.B2(n_197),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_196),
.A2(n_175),
.B1(n_167),
.B2(n_174),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_209),
.B(n_201),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_174),
.Y(n_210)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_210),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_198),
.A2(n_179),
.B1(n_177),
.B2(n_180),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_186),
.B(n_163),
.C(n_166),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_199),
.A2(n_166),
.B(n_169),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_213),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_216),
.C(n_214),
.Y(n_229)
);

NOR2x1_ASAP7_75t_SL g218 ( 
.A(n_212),
.B(n_189),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_218),
.A2(n_205),
.B(n_206),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_191),
.C(n_192),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_219),
.B(n_214),
.C(n_171),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_221),
.B(n_203),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_195),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_222),
.B(n_223),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_213),
.B(n_185),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_225),
.B(n_205),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_229),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_197),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_227),
.B(n_228),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_231),
.A2(n_232),
.B(n_233),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_171),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_230),
.A2(n_224),
.B1(n_221),
.B2(n_217),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_237),
.Y(n_243)
);

A2O1A1O1Ixp25_ASAP7_75t_L g237 ( 
.A1(n_233),
.A2(n_219),
.B(n_216),
.C(n_226),
.D(n_7),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_231),
.A2(n_11),
.B(n_5),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_239),
.B(n_12),
.C(n_5),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_235),
.A2(n_11),
.B1(n_5),
.B2(n_6),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_240),
.B(n_241),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_238),
.B(n_15),
.C(n_7),
.Y(n_242)
);

O2A1O1Ixp33_ASAP7_75t_SL g244 ( 
.A1(n_242),
.A2(n_10),
.B(n_12),
.C(n_13),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g247 ( 
.A1(n_244),
.A2(n_245),
.B(n_10),
.Y(n_247)
);

AOI221xp5_ASAP7_75t_L g246 ( 
.A1(n_243),
.A2(n_236),
.B1(n_10),
.B2(n_13),
.C(n_14),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_246),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_247),
.B(n_15),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_248),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_13),
.C(n_15),
.Y(n_251)
);


endmodule