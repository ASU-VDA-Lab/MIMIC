module real_jpeg_5707_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_0),
.B(n_126),
.Y(n_125)
);

AND2x2_ASAP7_75t_SL g159 ( 
.A(n_0),
.B(n_160),
.Y(n_159)
);

AND2x2_ASAP7_75t_SL g170 ( 
.A(n_0),
.B(n_171),
.Y(n_170)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_2),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_2),
.B(n_111),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_2),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_2),
.B(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_2),
.B(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_2),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_2),
.B(n_261),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_3),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_4),
.B(n_38),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_4),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_4),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_4),
.B(n_28),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_5),
.B(n_60),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_5),
.B(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_5),
.Y(n_116)
);

AND2x2_ASAP7_75t_SL g146 ( 
.A(n_5),
.B(n_147),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_5),
.B(n_113),
.Y(n_173)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_7),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_7),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_8),
.B(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_8),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_8),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_9),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_9),
.B(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_9),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_9),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_9),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_9),
.B(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_9),
.B(n_286),
.Y(n_285)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_11),
.Y(n_66)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_11),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_11),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_12),
.Y(n_82)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_12),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g165 ( 
.A(n_12),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_13),
.B(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_13),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_13),
.B(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_13),
.B(n_111),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_13),
.B(n_269),
.Y(n_268)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_14),
.Y(n_118)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_14),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_14),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_15),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_15),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_15),
.B(n_134),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_15),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_15),
.B(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_15),
.B(n_280),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_187),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_185),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_152),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_19),
.B(n_152),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_102),
.C(n_136),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_20),
.B(n_191),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_67),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_21),
.B(n_68),
.C(n_83),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_43),
.C(n_57),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_22),
.B(n_216),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_37),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_31),
.B2(n_36),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_25),
.B(n_31),
.C(n_37),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_27),
.Y(n_25)
);

OR2x2_ASAP7_75t_SL g44 ( 
.A(n_26),
.B(n_45),
.Y(n_44)
);

OR2x2_ASAP7_75t_SL g70 ( 
.A(n_26),
.B(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_29),
.B(n_98),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_30),
.Y(n_238)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_30),
.Y(n_273)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_34),
.Y(n_160)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_35),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g207 ( 
.A(n_35),
.Y(n_207)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx8_ASAP7_75t_L g229 ( 
.A(n_42),
.Y(n_229)
);

BUFx5_ASAP7_75t_L g292 ( 
.A(n_42),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_43),
.A2(n_57),
.B1(n_58),
.B2(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_43),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_48),
.C(n_51),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_44),
.A2(n_51),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_44),
.Y(n_200)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_48),
.B(n_199),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_50),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_51),
.Y(n_201)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_55),
.Y(n_213)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_63),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_59),
.A2(n_169),
.B1(n_170),
.B2(n_172),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_59),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_59),
.A2(n_63),
.B1(n_64),
.B2(n_172),
.Y(n_214)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_62),
.Y(n_144)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_62),
.Y(n_283)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_83),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_74),
.B2(n_75),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_70),
.B(n_76),
.C(n_81),
.Y(n_184)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_80),
.B2(n_81),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_77),
.B(n_125),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_77),
.B(n_125),
.Y(n_233)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_79),
.Y(n_91)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_79),
.Y(n_171)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_79),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_79),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_92),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_84),
.A2(n_85),
.B(n_88),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_84),
.B(n_93),
.C(n_97),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_88),
.Y(n_84)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_87),
.Y(n_182)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_90),
.Y(n_131)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_97),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_102),
.B(n_136),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_120),
.C(n_122),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_103),
.A2(n_120),
.B1(n_121),
.B2(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_103),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_109),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_104),
.B(n_110),
.C(n_115),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_105),
.B(n_291),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_105),
.B(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_107),
.Y(n_106)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_114),
.B1(n_115),
.B2(n_119),
.Y(n_109)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_117),
.Y(n_163)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_117),
.Y(n_232)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_118),
.Y(n_275)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_122),
.B(n_195),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_129),
.C(n_132),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_123),
.A2(n_124),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_128),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_129),
.A2(n_130),
.B1(n_132),
.B2(n_133),
.Y(n_321)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_135),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_151),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_138),
.B(n_139),
.C(n_151),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_145),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_146),
.C(n_149),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_149),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_175),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_166),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_161),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_173),
.B2(n_174),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_169),
.A2(n_170),
.B1(n_225),
.B2(n_226),
.Y(n_262)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_170),
.B(n_225),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_173),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_184),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_218),
.B(n_329),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_192),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_190),
.B(n_192),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_197),
.C(n_215),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_193),
.A2(n_194),
.B1(n_325),
.B2(n_326),
.Y(n_324)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_197),
.B(n_215),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_202),
.C(n_214),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_198),
.B(n_315),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_202),
.B(n_214),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_208),
.C(n_209),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_203),
.A2(n_204),
.B1(n_209),
.B2(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_208),
.B(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_209),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_237),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_210),
.B(n_294),
.Y(n_293)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx8_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_323),
.B(n_328),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_310),
.B(n_322),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_263),
.B(n_309),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_249),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_222),
.B(n_249),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_234),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_223),
.B(n_235),
.C(n_246),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_230),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_224),
.B(n_231),
.C(n_233),
.Y(n_318)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx8_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_246),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_239),
.C(n_241),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_236),
.B(n_251),
.Y(n_250)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_239),
.A2(n_240),
.B1(n_241),
.B2(n_242),
.Y(n_251)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx8_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

BUFx5_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_252),
.C(n_262),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_250),
.B(n_306),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_252),
.A2(n_253),
.B1(n_262),
.B2(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_259),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_254),
.A2(n_255),
.B1(n_259),
.B2(n_260),
.Y(n_276)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx5_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_262),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_303),
.B(n_308),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_288),
.B(n_302),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_266),
.B(n_277),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_266),
.B(n_277),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_276),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_274),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_268),
.B(n_274),
.C(n_276),
.Y(n_304)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx5_ASAP7_75t_SL g270 ( 
.A(n_271),
.Y(n_270)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_284),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_278),
.A2(n_279),
.B1(n_284),
.B2(n_285),
.Y(n_300)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx6_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx8_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_296),
.B(n_301),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_293),
.Y(n_289)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_300),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_297),
.B(n_300),
.Y(n_301)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_305),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_312),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_313),
.A2(n_314),
.B1(n_316),
.B2(n_317),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_313),
.B(n_318),
.C(n_319),
.Y(n_327)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_324),
.B(n_327),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_327),
.Y(n_328)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_325),
.Y(n_326)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);


endmodule