module real_aes_2356_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_504;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_754;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_288;
wire n_147;
wire n_756;
wire n_150;
wire n_404;
wire n_598;
wire n_735;
wire n_728;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_0), .B(n_147), .Y(n_461) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_1), .A2(n_155), .B(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_2), .B(n_766), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_3), .B(n_147), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_4), .B(n_174), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_5), .B(n_174), .Y(n_472) );
INVx1_ASAP7_75t_L g143 ( .A(n_6), .Y(n_143) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_7), .A2(n_106), .B1(n_726), .B2(n_731), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_8), .B(n_174), .Y(n_501) );
CKINVDCx16_ASAP7_75t_R g766 ( .A(n_9), .Y(n_766) );
NAND2xp33_ASAP7_75t_L g542 ( .A(n_10), .B(n_172), .Y(n_542) );
AND2x2_ASAP7_75t_L g177 ( .A(n_11), .B(n_178), .Y(n_177) );
AND2x2_ASAP7_75t_L g188 ( .A(n_12), .B(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g134 ( .A(n_13), .Y(n_134) );
AOI221x1_ASAP7_75t_L g447 ( .A1(n_14), .A2(n_26), .B1(n_147), .B2(n_155), .C(n_448), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_15), .B(n_174), .Y(n_243) );
CKINVDCx16_ASAP7_75t_R g116 ( .A(n_16), .Y(n_116) );
NOR3xp33_ASAP7_75t_L g764 ( .A(n_16), .B(n_765), .C(n_767), .Y(n_764) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_17), .B(n_147), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g107 ( .A1(n_18), .A2(n_88), .B1(n_108), .B2(n_109), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_18), .Y(n_108) );
AO21x2_ASAP7_75t_L g536 ( .A1(n_19), .A2(n_189), .B(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_20), .B(n_132), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_21), .B(n_174), .Y(n_525) );
AO21x1_ASAP7_75t_L g467 ( .A1(n_22), .A2(n_147), .B(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_23), .B(n_147), .Y(n_228) );
INVx1_ASAP7_75t_L g119 ( .A(n_24), .Y(n_119) );
AOI22xp33_ASAP7_75t_L g137 ( .A1(n_25), .A2(n_92), .B1(n_138), .B2(n_147), .Y(n_137) );
NAND2x1_ASAP7_75t_L g459 ( .A(n_27), .B(n_174), .Y(n_459) );
NAND2x1_ASAP7_75t_L g500 ( .A(n_28), .B(n_172), .Y(n_500) );
OR2x2_ASAP7_75t_L g135 ( .A(n_29), .B(n_89), .Y(n_135) );
OA21x2_ASAP7_75t_L g167 ( .A1(n_29), .A2(n_89), .B(n_134), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_30), .B(n_172), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_31), .B(n_174), .Y(n_541) );
AO21x2_ASAP7_75t_L g238 ( .A1(n_32), .A2(n_178), .B(n_239), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_33), .B(n_172), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_34), .A2(n_155), .B(n_184), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_35), .B(n_174), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_36), .A2(n_155), .B(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g145 ( .A(n_37), .B(n_146), .Y(n_145) );
AND2x2_ASAP7_75t_L g153 ( .A(n_37), .B(n_143), .Y(n_153) );
INVx1_ASAP7_75t_L g159 ( .A(n_37), .Y(n_159) );
OR2x6_ASAP7_75t_L g117 ( .A(n_38), .B(n_118), .Y(n_117) );
INVxp67_ASAP7_75t_L g767 ( .A(n_38), .Y(n_767) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_39), .B(n_147), .Y(n_482) );
OAI22xp5_ASAP7_75t_SL g750 ( .A1(n_40), .A2(n_751), .B1(n_752), .B2(n_755), .Y(n_750) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_40), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_41), .B(n_147), .Y(n_187) );
XNOR2xp5_ASAP7_75t_L g106 ( .A(n_42), .B(n_107), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_43), .B(n_174), .Y(n_213) );
CKINVDCx20_ASAP7_75t_R g529 ( .A(n_44), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_45), .B(n_172), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_46), .B(n_147), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_47), .A2(n_155), .B(n_170), .Y(n_169) );
AOI22xp5_ASAP7_75t_L g752 ( .A1(n_48), .A2(n_63), .B1(n_753), .B2(n_754), .Y(n_752) );
CKINVDCx20_ASAP7_75t_R g754 ( .A(n_48), .Y(n_754) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_49), .A2(n_155), .B(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_50), .B(n_172), .Y(n_200) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_51), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_52), .B(n_172), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_53), .B(n_147), .Y(n_240) );
CKINVDCx20_ASAP7_75t_R g742 ( .A(n_54), .Y(n_742) );
INVx1_ASAP7_75t_L g141 ( .A(n_55), .Y(n_141) );
INVx1_ASAP7_75t_L g150 ( .A(n_55), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_56), .B(n_174), .Y(n_173) );
AND2x2_ASAP7_75t_L g208 ( .A(n_57), .B(n_132), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_58), .B(n_172), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_59), .B(n_174), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_60), .B(n_172), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_61), .A2(n_155), .B(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_62), .B(n_147), .Y(n_176) );
CKINVDCx20_ASAP7_75t_R g753 ( .A(n_63), .Y(n_753) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_64), .B(n_147), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_65), .A2(n_155), .B(n_221), .Y(n_220) );
AND2x2_ASAP7_75t_L g234 ( .A(n_66), .B(n_133), .Y(n_234) );
AO21x1_ASAP7_75t_L g469 ( .A1(n_67), .A2(n_155), .B(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_68), .B(n_147), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_69), .B(n_172), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_70), .B(n_147), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_71), .B(n_172), .Y(n_244) );
AOI22xp5_ASAP7_75t_L g154 ( .A1(n_72), .A2(n_96), .B1(n_155), .B2(n_157), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_73), .B(n_174), .Y(n_231) );
AND2x2_ASAP7_75t_L g483 ( .A(n_74), .B(n_133), .Y(n_483) );
INVx1_ASAP7_75t_L g146 ( .A(n_75), .Y(n_146) );
INVx1_ASAP7_75t_L g152 ( .A(n_75), .Y(n_152) );
AND2x2_ASAP7_75t_L g503 ( .A(n_76), .B(n_178), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_77), .B(n_172), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_78), .A2(n_155), .B(n_212), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g197 ( .A1(n_79), .A2(n_155), .B(n_198), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_80), .A2(n_155), .B(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g225 ( .A(n_81), .B(n_133), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g131 ( .A(n_82), .B(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g120 ( .A(n_83), .Y(n_120) );
AND2x2_ASAP7_75t_L g488 ( .A(n_84), .B(n_178), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g527 ( .A(n_85), .B(n_147), .Y(n_527) );
AND2x2_ASAP7_75t_L g201 ( .A(n_86), .B(n_189), .Y(n_201) );
AND2x2_ASAP7_75t_L g468 ( .A(n_87), .B(n_215), .Y(n_468) );
INVx1_ASAP7_75t_L g109 ( .A(n_88), .Y(n_109) );
AND2x2_ASAP7_75t_L g462 ( .A(n_90), .B(n_178), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_91), .B(n_172), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_93), .B(n_174), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_94), .B(n_172), .Y(n_449) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_95), .A2(n_155), .B(n_524), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_97), .A2(n_155), .B(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_98), .B(n_174), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_99), .B(n_174), .Y(n_493) );
BUFx2_ASAP7_75t_L g233 ( .A(n_100), .Y(n_233) );
BUFx2_ASAP7_75t_L g738 ( .A(n_101), .Y(n_738) );
BUFx2_ASAP7_75t_SL g746 ( .A(n_101), .Y(n_746) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_102), .A2(n_155), .B(n_540), .Y(n_539) );
AOI21xp33_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_760), .B(n_768), .Y(n_103) );
OA21x2_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_735), .B(n_743), .Y(n_104) );
OAI21xp5_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_110), .B(n_725), .Y(n_105) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OAI22xp5_ASAP7_75t_L g111 ( .A1(n_112), .A2(n_121), .B1(n_440), .B2(n_720), .Y(n_111) );
CKINVDCx6p67_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
CKINVDCx11_ASAP7_75t_R g727 ( .A(n_113), .Y(n_727) );
INVx3_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_115), .Y(n_114) );
AND2x6_ASAP7_75t_SL g115 ( .A(n_116), .B(n_117), .Y(n_115) );
OR2x6_ASAP7_75t_SL g723 ( .A(n_116), .B(n_724), .Y(n_723) );
OR2x2_ASAP7_75t_L g734 ( .A(n_116), .B(n_117), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_116), .B(n_724), .Y(n_741) );
CKINVDCx5p33_ASAP7_75t_R g724 ( .A(n_117), .Y(n_724) );
INVx1_ASAP7_75t_L g763 ( .A(n_118), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_120), .Y(n_118) );
INVx4_ASAP7_75t_L g728 ( .A(n_121), .Y(n_728) );
AOI22x1_ASAP7_75t_L g749 ( .A1(n_121), .A2(n_728), .B1(n_750), .B2(n_756), .Y(n_749) );
OR2x6_ASAP7_75t_L g121 ( .A(n_122), .B(n_377), .Y(n_121) );
NAND3xp33_ASAP7_75t_L g122 ( .A(n_123), .B(n_293), .C(n_330), .Y(n_122) );
NOR3xp33_ASAP7_75t_L g123 ( .A(n_124), .B(n_261), .C(n_276), .Y(n_123) );
OAI221xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_205), .B1(n_235), .B2(n_247), .C(n_248), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
NAND2xp5_ASAP7_75t_SL g126 ( .A(n_127), .B(n_190), .Y(n_126) );
OAI22xp33_ASAP7_75t_SL g321 ( .A1(n_127), .A2(n_285), .B1(n_322), .B2(n_325), .Y(n_321) );
OR2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_162), .Y(n_127) );
OAI21xp33_ASAP7_75t_SL g331 ( .A1(n_128), .A2(n_332), .B(n_338), .Y(n_331) );
OR2x2_ASAP7_75t_L g360 ( .A(n_128), .B(n_192), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_128), .B(n_280), .Y(n_361) );
INVx2_ASAP7_75t_L g392 ( .A(n_128), .Y(n_392) );
INVx2_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_129), .B(n_252), .Y(n_373) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
OR2x2_ASAP7_75t_L g247 ( .A(n_130), .B(n_165), .Y(n_247) );
BUFx3_ASAP7_75t_L g273 ( .A(n_130), .Y(n_273) );
AND2x2_ASAP7_75t_L g409 ( .A(n_130), .B(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g432 ( .A(n_130), .B(n_193), .Y(n_432) );
AND2x4_ASAP7_75t_L g130 ( .A(n_131), .B(n_136), .Y(n_130) );
AND2x4_ASAP7_75t_L g204 ( .A(n_131), .B(n_136), .Y(n_204) );
AO21x2_ASAP7_75t_L g136 ( .A1(n_132), .A2(n_137), .B(n_154), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g181 ( .A(n_132), .Y(n_181) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_132), .A2(n_196), .B(n_197), .Y(n_195) );
OA21x2_ASAP7_75t_L g446 ( .A1(n_132), .A2(n_447), .B(n_451), .Y(n_446) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_132), .A2(n_490), .B(n_491), .Y(n_489) );
OA21x2_ASAP7_75t_L g590 ( .A1(n_132), .A2(n_447), .B(n_451), .Y(n_590) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x2_ASAP7_75t_SL g133 ( .A(n_134), .B(n_135), .Y(n_133) );
AND2x4_ASAP7_75t_L g215 ( .A(n_134), .B(n_135), .Y(n_215) );
AND2x4_ASAP7_75t_L g138 ( .A(n_139), .B(n_144), .Y(n_138) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_142), .Y(n_139) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
AND2x2_ASAP7_75t_L g156 ( .A(n_141), .B(n_143), .Y(n_156) );
AND2x4_ASAP7_75t_L g174 ( .A(n_141), .B(n_151), .Y(n_174) );
HB1xp67_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
BUFx3_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
AND2x6_ASAP7_75t_L g155 ( .A(n_145), .B(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g161 ( .A(n_146), .Y(n_161) );
AND2x6_ASAP7_75t_L g172 ( .A(n_146), .B(n_149), .Y(n_172) );
AND2x4_ASAP7_75t_L g147 ( .A(n_148), .B(n_153), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_149), .B(n_151), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx5_ASAP7_75t_L g175 ( .A(n_153), .Y(n_175) );
AND2x4_ASAP7_75t_L g157 ( .A(n_156), .B(n_158), .Y(n_157) );
NOR2x1p5_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
INVx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_SL g162 ( .A(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_163), .B(n_193), .Y(n_352) );
INVx1_ASAP7_75t_L g389 ( .A(n_163), .Y(n_389) );
AND2x2_ASAP7_75t_L g163 ( .A(n_164), .B(n_179), .Y(n_163) );
AND2x2_ASAP7_75t_L g203 ( .A(n_164), .B(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g410 ( .A(n_164), .Y(n_410) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g253 ( .A(n_165), .Y(n_253) );
AND2x2_ASAP7_75t_L g254 ( .A(n_165), .B(n_179), .Y(n_254) );
AND2x2_ASAP7_75t_L g275 ( .A(n_165), .B(n_194), .Y(n_275) );
AND2x2_ASAP7_75t_L g357 ( .A(n_165), .B(n_180), .Y(n_357) );
AO21x2_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_168), .B(n_177), .Y(n_165) );
INVx4_ASAP7_75t_L g178 ( .A(n_166), .Y(n_178) );
INVx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
BUFx4f_ASAP7_75t_L g189 ( .A(n_167), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_169), .B(n_176), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_173), .B(n_175), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_172), .B(n_233), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_175), .A2(n_185), .B(n_186), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_175), .A2(n_199), .B(n_200), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_175), .A2(n_213), .B(n_214), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g221 ( .A1(n_175), .A2(n_222), .B(n_223), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_175), .A2(n_231), .B(n_232), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_175), .A2(n_243), .B(n_244), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g448 ( .A1(n_175), .A2(n_449), .B(n_450), .Y(n_448) );
AOI21xp5_ASAP7_75t_L g458 ( .A1(n_175), .A2(n_459), .B(n_460), .Y(n_458) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_175), .A2(n_471), .B(n_472), .Y(n_470) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_175), .A2(n_480), .B(n_481), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_175), .A2(n_493), .B(n_494), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_175), .A2(n_500), .B(n_501), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_175), .A2(n_525), .B(n_526), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_175), .A2(n_541), .B(n_542), .Y(n_540) );
INVx3_ASAP7_75t_L g218 ( .A(n_178), .Y(n_218) );
AND2x4_ASAP7_75t_SL g250 ( .A(n_179), .B(n_194), .Y(n_250) );
INVx1_ASAP7_75t_L g281 ( .A(n_179), .Y(n_281) );
INVx2_ASAP7_75t_L g289 ( .A(n_179), .Y(n_289) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_179), .Y(n_313) );
INVx3_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
HB1xp67_ASAP7_75t_L g202 ( .A(n_180), .Y(n_202) );
AOI21x1_ASAP7_75t_L g180 ( .A1(n_181), .A2(n_182), .B(n_188), .Y(n_180) );
AO21x2_ASAP7_75t_L g496 ( .A1(n_181), .A2(n_497), .B(n_503), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_183), .B(n_187), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_189), .A2(n_228), .B(n_229), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_191), .B(n_203), .Y(n_190) );
AND2x2_ASAP7_75t_L g428 ( .A(n_191), .B(n_291), .Y(n_428) );
INVx1_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_193), .B(n_202), .Y(n_192) );
NAND2x1p5_ASAP7_75t_L g287 ( .A(n_193), .B(n_288), .Y(n_287) );
AND2x2_ASAP7_75t_L g339 ( .A(n_193), .B(n_254), .Y(n_339) );
AND2x2_ASAP7_75t_L g356 ( .A(n_193), .B(n_357), .Y(n_356) );
INVx4_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
AND2x4_ASAP7_75t_L g280 ( .A(n_194), .B(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g296 ( .A(n_194), .Y(n_296) );
AND2x2_ASAP7_75t_L g340 ( .A(n_194), .B(n_341), .Y(n_340) );
OR2x2_ASAP7_75t_L g347 ( .A(n_194), .B(n_348), .Y(n_347) );
NOR2x1_ASAP7_75t_L g362 ( .A(n_194), .B(n_253), .Y(n_362) );
BUFx2_ASAP7_75t_L g372 ( .A(n_194), .Y(n_372) );
AND2x2_ASAP7_75t_L g397 ( .A(n_194), .B(n_357), .Y(n_397) );
AND2x2_ASAP7_75t_L g418 ( .A(n_194), .B(n_419), .Y(n_418) );
OR2x6_ASAP7_75t_L g194 ( .A(n_195), .B(n_201), .Y(n_194) );
INVx1_ASAP7_75t_L g349 ( .A(n_202), .Y(n_349) );
NAND2xp5_ASAP7_75t_SL g295 ( .A(n_203), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g379 ( .A(n_203), .B(n_250), .Y(n_379) );
INVx3_ASAP7_75t_L g286 ( .A(n_204), .Y(n_286) );
AND2x2_ASAP7_75t_L g419 ( .A(n_204), .B(n_341), .Y(n_419) );
INVx1_ASAP7_75t_SL g205 ( .A(n_206), .Y(n_205) );
AOI22xp5_ASAP7_75t_L g248 ( .A1(n_206), .A2(n_249), .B1(n_254), .B2(n_255), .Y(n_248) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_216), .Y(n_206) );
INVx4_ASAP7_75t_L g246 ( .A(n_207), .Y(n_246) );
INVx2_ASAP7_75t_L g283 ( .A(n_207), .Y(n_283) );
NAND2x1_ASAP7_75t_L g309 ( .A(n_207), .B(n_226), .Y(n_309) );
OR2x2_ASAP7_75t_L g324 ( .A(n_207), .B(n_259), .Y(n_324) );
OR2x2_ASAP7_75t_SL g351 ( .A(n_207), .B(n_323), .Y(n_351) );
AND2x2_ASAP7_75t_L g364 ( .A(n_207), .B(n_238), .Y(n_364) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_207), .Y(n_385) );
OR2x6_ASAP7_75t_L g207 ( .A(n_208), .B(n_209), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_210), .A2(n_211), .B(n_215), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_215), .A2(n_240), .B(n_241), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_215), .B(n_474), .Y(n_473) );
INVx1_ASAP7_75t_SL g521 ( .A(n_215), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_215), .A2(n_538), .B(n_539), .Y(n_537) );
INVx2_ASAP7_75t_L g264 ( .A(n_216), .Y(n_264) );
AND2x2_ASAP7_75t_L g396 ( .A(n_216), .B(n_370), .Y(n_396) );
NOR2x1_ASAP7_75t_SL g216 ( .A(n_217), .B(n_226), .Y(n_216) );
AND2x2_ASAP7_75t_L g237 ( .A(n_217), .B(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g413 ( .A(n_217), .B(n_336), .Y(n_413) );
AO21x1_ASAP7_75t_SL g217 ( .A1(n_218), .A2(n_219), .B(n_225), .Y(n_217) );
AO21x2_ASAP7_75t_L g260 ( .A1(n_218), .A2(n_219), .B(n_225), .Y(n_260) );
AO21x2_ASAP7_75t_L g455 ( .A1(n_218), .A2(n_456), .B(n_462), .Y(n_455) );
AO21x2_ASAP7_75t_L g476 ( .A1(n_218), .A2(n_477), .B(n_483), .Y(n_476) );
AO21x2_ASAP7_75t_L g510 ( .A1(n_218), .A2(n_477), .B(n_483), .Y(n_510) );
AO21x2_ASAP7_75t_L g514 ( .A1(n_218), .A2(n_456), .B(n_462), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_220), .B(n_224), .Y(n_219) );
OR2x2_ASAP7_75t_L g245 ( .A(n_226), .B(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g256 ( .A(n_226), .B(n_246), .Y(n_256) );
AND2x2_ASAP7_75t_L g302 ( .A(n_226), .B(n_259), .Y(n_302) );
OR2x2_ASAP7_75t_L g323 ( .A(n_226), .B(n_238), .Y(n_323) );
INVx2_ASAP7_75t_SL g329 ( .A(n_226), .Y(n_329) );
AND2x2_ASAP7_75t_L g335 ( .A(n_226), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g345 ( .A(n_226), .B(n_328), .Y(n_345) );
BUFx2_ASAP7_75t_L g367 ( .A(n_226), .Y(n_367) );
OR2x6_ASAP7_75t_L g226 ( .A(n_227), .B(n_234), .Y(n_226) );
INVx2_ASAP7_75t_L g414 ( .A(n_235), .Y(n_414) );
OR2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_245), .Y(n_235) );
OR2x2_ASAP7_75t_L g439 ( .A(n_236), .B(n_283), .Y(n_439) );
INVx2_ASAP7_75t_SL g236 ( .A(n_237), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_237), .B(n_246), .Y(n_305) );
AND2x2_ASAP7_75t_L g376 ( .A(n_237), .B(n_256), .Y(n_376) );
INVx1_ASAP7_75t_L g258 ( .A(n_238), .Y(n_258) );
HB1xp67_ASAP7_75t_L g267 ( .A(n_238), .Y(n_267) );
INVx1_ASAP7_75t_L g300 ( .A(n_238), .Y(n_300) );
INVx2_ASAP7_75t_L g336 ( .A(n_238), .Y(n_336) );
NOR2xp67_ASAP7_75t_L g266 ( .A(n_246), .B(n_267), .Y(n_266) );
BUFx2_ASAP7_75t_L g326 ( .A(n_246), .Y(n_326) );
INVx2_ASAP7_75t_SL g402 ( .A(n_247), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g303 ( .A1(n_249), .A2(n_304), .B1(n_306), .B2(n_310), .Y(n_303) );
AND2x2_ASAP7_75t_SL g249 ( .A(n_250), .B(n_251), .Y(n_249) );
AND2x2_ASAP7_75t_L g430 ( .A(n_250), .B(n_286), .Y(n_430) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_252), .B(n_296), .Y(n_375) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g341 ( .A(n_253), .B(n_289), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_254), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g284 ( .A(n_255), .Y(n_284) );
AOI221xp5_ASAP7_75t_L g398 ( .A1(n_255), .A2(n_399), .B1(n_403), .B2(n_405), .C(n_407), .Y(n_398) );
AND2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
AND2x2_ASAP7_75t_L g268 ( .A(n_256), .B(n_269), .Y(n_268) );
INVxp67_ASAP7_75t_SL g292 ( .A(n_256), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_256), .B(n_299), .Y(n_354) );
INVx1_ASAP7_75t_SL g350 ( .A(n_257), .Y(n_350) );
AOI221xp5_ASAP7_75t_SL g378 ( .A1(n_257), .A2(n_268), .B1(n_379), .B2(n_380), .C(n_383), .Y(n_378) );
AOI322xp5_ASAP7_75t_L g411 ( .A1(n_257), .A2(n_329), .A3(n_356), .B1(n_412), .B2(n_414), .C1(n_415), .C2(n_418), .Y(n_411) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
BUFx2_ASAP7_75t_L g278 ( .A(n_258), .Y(n_278) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_259), .Y(n_270) );
INVx2_ASAP7_75t_L g328 ( .A(n_259), .Y(n_328) );
AND2x2_ASAP7_75t_L g369 ( .A(n_259), .B(n_370), .Y(n_369) );
INVx3_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
OA21x2_ASAP7_75t_SL g261 ( .A1(n_262), .A2(n_268), .B(n_271), .Y(n_261) );
AOI211xp5_ASAP7_75t_L g431 ( .A1(n_262), .A2(n_432), .B(n_433), .C(n_437), .Y(n_431) );
INVx1_ASAP7_75t_SL g262 ( .A(n_263), .Y(n_262) );
OR2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
OR2x2_ASAP7_75t_L g320 ( .A(n_264), .B(n_282), .Y(n_320) );
OR2x2_ASAP7_75t_L g404 ( .A(n_264), .B(n_299), .Y(n_404) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g344 ( .A(n_266), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g422 ( .A(n_269), .Y(n_422) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g308 ( .A(n_270), .Y(n_308) );
INVx1_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
OR2x2_ASAP7_75t_L g277 ( .A(n_273), .B(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
AND2x2_ASAP7_75t_L g312 ( .A(n_275), .B(n_313), .Y(n_312) );
OAI322xp33_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_279), .A3(n_282), .B1(n_284), .B2(n_285), .C1(n_290), .C2(n_292), .Y(n_276) );
INVx1_ASAP7_75t_L g318 ( .A(n_277), .Y(n_318) );
OR2x2_ASAP7_75t_L g290 ( .A(n_279), .B(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_279), .B(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g301 ( .A(n_283), .B(n_302), .Y(n_301) );
OAI32xp33_ASAP7_75t_L g346 ( .A1(n_283), .A2(n_347), .A3(n_350), .B1(n_351), .B2(n_352), .Y(n_346) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_287), .Y(n_285) );
INVx2_ASAP7_75t_L g291 ( .A(n_286), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_286), .B(n_349), .Y(n_348) );
NOR2x1_ASAP7_75t_L g388 ( .A(n_286), .B(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g412 ( .A(n_286), .B(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g333 ( .A(n_287), .Y(n_333) );
INVx1_ASAP7_75t_SL g288 ( .A(n_289), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_291), .B(n_357), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g293 ( .A(n_294), .B(n_314), .Y(n_293) );
OAI21xp33_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_297), .B(n_303), .Y(n_294) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
AND2x4_ASAP7_75t_SL g298 ( .A(n_299), .B(n_301), .Y(n_298) );
INVx3_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g363 ( .A(n_302), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_305), .A2(n_325), .B1(n_427), .B2(n_429), .Y(n_426) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
A2O1A1Ixp33_ASAP7_75t_L g353 ( .A1(n_307), .A2(n_354), .B(n_355), .C(n_358), .Y(n_353) );
OR2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_309), .Y(n_307) );
INVx3_ASAP7_75t_L g435 ( .A(n_309), .Y(n_435) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx2_ASAP7_75t_L g316 ( .A(n_313), .Y(n_316) );
AO21x1_ASAP7_75t_L g314 ( .A1(n_315), .A2(n_317), .B(n_321), .Y(n_314) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g381 ( .A(n_316), .Y(n_381) );
AND2x2_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_322), .B(n_408), .Y(n_407) );
OR2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx1_ASAP7_75t_L g337 ( .A(n_324), .Y(n_337) );
OR2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
INVx1_ASAP7_75t_L g394 ( .A(n_327), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
NOR3xp33_ASAP7_75t_L g330 ( .A(n_331), .B(n_353), .C(n_365), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
OAI21xp5_ASAP7_75t_SL g395 ( .A1(n_334), .A2(n_396), .B(n_397), .Y(n_395) );
AND2x4_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
INVx1_ASAP7_75t_L g370 ( .A(n_336), .Y(n_370) );
O2A1O1Ixp5_ASAP7_75t_SL g338 ( .A1(n_339), .A2(n_340), .B(n_342), .C(n_346), .Y(n_338) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_348), .Y(n_438) );
INVx2_ASAP7_75t_L g423 ( .A(n_351), .Y(n_423) );
AOI21xp33_ASAP7_75t_L g437 ( .A1(n_352), .A2(n_438), .B(n_439), .Y(n_437) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g417 ( .A(n_357), .Y(n_417) );
OAI31xp33_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_361), .A3(n_362), .B(n_363), .Y(n_358) );
INVx1_ASAP7_75t_SL g359 ( .A(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g436 ( .A(n_364), .Y(n_436) );
OAI21xp5_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_371), .B(n_374), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
BUFx2_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g386 ( .A(n_369), .Y(n_386) );
AOI21xp33_ASAP7_75t_SL g433 ( .A1(n_371), .A2(n_434), .B(n_436), .Y(n_433) );
OR2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
INVx2_ASAP7_75t_L g401 ( .A(n_372), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_372), .B(n_392), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_372), .B(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g382 ( .A(n_373), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
NAND5xp2_ASAP7_75t_L g377 ( .A(n_378), .B(n_398), .C(n_411), .D(n_420), .E(n_431), .Y(n_377) );
AND2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
OAI221xp5_ASAP7_75t_L g383 ( .A1(n_384), .A2(n_387), .B1(n_390), .B2(n_393), .C(n_395), .Y(n_383) );
OR2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVxp67_ASAP7_75t_SL g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVxp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_401), .B(n_402), .Y(n_400) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
AOI21xp5_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_424), .B(n_426), .Y(n_420) );
AND2x4_ASAP7_75t_L g421 ( .A(n_422), .B(n_423), .Y(n_421) );
INVx1_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
INVxp67_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx3_ASAP7_75t_L g730 ( .A(n_440), .Y(n_730) );
NAND4xp75_ASAP7_75t_L g440 ( .A(n_441), .B(n_630), .C(n_670), .D(n_699), .Y(n_440) );
NOR2x1_ASAP7_75t_L g441 ( .A(n_442), .B(n_592), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_443), .B(n_549), .Y(n_442) );
AOI21xp5_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_484), .B(n_504), .Y(n_443) );
AND2x2_ASAP7_75t_SL g444 ( .A(n_445), .B(n_452), .Y(n_444) );
AND2x4_ASAP7_75t_L g548 ( .A(n_445), .B(n_509), .Y(n_548) );
INVx1_ASAP7_75t_SL g601 ( .A(n_445), .Y(n_601) );
AOI21xp33_ASAP7_75t_L g636 ( .A1(n_445), .A2(n_637), .B(n_640), .Y(n_636) );
A2O1A1Ixp33_ASAP7_75t_SL g640 ( .A1(n_445), .A2(n_641), .B(n_642), .C(n_643), .Y(n_640) );
NAND2x1_ASAP7_75t_L g681 ( .A(n_445), .B(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_445), .B(n_642), .Y(n_703) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g507 ( .A(n_446), .Y(n_507) );
HB1xp67_ASAP7_75t_L g580 ( .A(n_446), .Y(n_580) );
AND2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_463), .Y(n_452) );
AND2x2_ASAP7_75t_L g572 ( .A(n_453), .B(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g653 ( .A(n_453), .B(n_509), .Y(n_653) );
INVx1_ASAP7_75t_L g713 ( .A(n_453), .Y(n_713) );
BUFx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AND2x2_ASAP7_75t_L g557 ( .A(n_454), .B(n_475), .Y(n_557) );
AND2x2_ASAP7_75t_L g682 ( .A(n_454), .B(n_476), .Y(n_682) );
AND2x2_ASAP7_75t_L g687 ( .A(n_454), .B(n_647), .Y(n_687) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVxp67_ASAP7_75t_L g563 ( .A(n_455), .Y(n_563) );
BUFx3_ASAP7_75t_L g596 ( .A(n_455), .Y(n_596) );
AND2x2_ASAP7_75t_L g642 ( .A(n_455), .B(n_476), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_457), .B(n_461), .Y(n_456) );
AND2x2_ASAP7_75t_L g627 ( .A(n_463), .B(n_506), .Y(n_627) );
AND2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_475), .Y(n_463) );
AND2x4_ASAP7_75t_L g509 ( .A(n_464), .B(n_510), .Y(n_509) );
OR2x2_ASAP7_75t_L g619 ( .A(n_464), .B(n_603), .Y(n_619) );
AND2x2_ASAP7_75t_SL g662 ( .A(n_464), .B(n_590), .Y(n_662) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
BUFx2_ASAP7_75t_L g598 ( .A(n_465), .Y(n_598) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g559 ( .A(n_466), .Y(n_559) );
OAI21x1_ASAP7_75t_SL g466 ( .A1(n_467), .A2(n_469), .B(n_473), .Y(n_466) );
INVx1_ASAP7_75t_L g474 ( .A(n_468), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_475), .B(n_559), .Y(n_562) );
AND2x2_ASAP7_75t_L g647 ( .A(n_475), .B(n_590), .Y(n_647) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AND2x2_ASAP7_75t_L g644 ( .A(n_476), .B(n_507), .Y(n_644) );
AND2x2_ASAP7_75t_L g664 ( .A(n_476), .B(n_590), .Y(n_664) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_478), .B(n_482), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_484), .B(n_553), .Y(n_582) );
AOI221xp5_ASAP7_75t_L g675 ( .A1(n_484), .A2(n_676), .B1(n_677), .B2(n_678), .C(n_680), .Y(n_675) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
OAI332xp33_ASAP7_75t_L g709 ( .A1(n_485), .A2(n_569), .A3(n_576), .B1(n_635), .B2(n_710), .B3(n_711), .C1(n_712), .C2(n_714), .Y(n_709) );
NAND2x1p5_ASAP7_75t_L g485 ( .A(n_486), .B(n_495), .Y(n_485) );
AND2x2_ASAP7_75t_L g515 ( .A(n_486), .B(n_496), .Y(n_515) );
AND2x2_ASAP7_75t_L g532 ( .A(n_486), .B(n_533), .Y(n_532) );
INVx4_ASAP7_75t_L g544 ( .A(n_486), .Y(n_544) );
AND2x2_ASAP7_75t_SL g604 ( .A(n_486), .B(n_545), .Y(n_604) );
INVx5_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NOR2x1_ASAP7_75t_SL g566 ( .A(n_487), .B(n_533), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_487), .B(n_495), .Y(n_570) );
AND2x2_ASAP7_75t_L g577 ( .A(n_487), .B(n_496), .Y(n_577) );
BUFx2_ASAP7_75t_L g612 ( .A(n_487), .Y(n_612) );
AND2x2_ASAP7_75t_L g667 ( .A(n_487), .B(n_536), .Y(n_667) );
OR2x6_ASAP7_75t_L g487 ( .A(n_488), .B(n_489), .Y(n_487) );
OR2x2_ASAP7_75t_L g535 ( .A(n_495), .B(n_536), .Y(n_535) );
AND2x4_ASAP7_75t_L g545 ( .A(n_495), .B(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g585 ( .A(n_495), .Y(n_585) );
AND2x2_ASAP7_75t_L g655 ( .A(n_495), .B(n_554), .Y(n_655) );
AND2x2_ASAP7_75t_L g668 ( .A(n_495), .B(n_669), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_495), .B(n_669), .Y(n_686) );
INVx4_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_496), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_498), .B(n_502), .Y(n_497) );
OAI32xp33_ASAP7_75t_L g504 ( .A1(n_505), .A2(n_511), .A3(n_516), .B1(n_530), .B2(n_547), .Y(n_504) );
INVx2_ASAP7_75t_L g613 ( .A(n_505), .Y(n_613) );
OR2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_508), .Y(n_505) );
INVx1_ASAP7_75t_L g624 ( .A(n_506), .Y(n_624) );
BUFx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
AND2x4_ASAP7_75t_L g558 ( .A(n_507), .B(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g691 ( .A(n_507), .B(n_596), .Y(n_691) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g603 ( .A(n_510), .Y(n_603) );
INVx1_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_515), .Y(n_512) );
INVx2_ASAP7_75t_L g591 ( .A(n_513), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_513), .B(n_634), .Y(n_633) );
BUFx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AND2x4_ASAP7_75t_SL g602 ( .A(n_514), .B(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g679 ( .A(n_514), .Y(n_679) );
AND2x2_ASAP7_75t_L g697 ( .A(n_514), .B(n_559), .Y(n_697) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
NOR2xp67_ASAP7_75t_SL g641 ( .A(n_517), .B(n_570), .Y(n_641) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_518), .B(n_552), .Y(n_639) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_L g715 ( .A(n_519), .B(n_585), .Y(n_715) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g546 ( .A(n_520), .Y(n_546) );
INVx2_ASAP7_75t_L g587 ( .A(n_520), .Y(n_587) );
AO21x2_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_522), .B(n_528), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g528 ( .A(n_521), .B(n_529), .Y(n_528) );
AO21x2_ASAP7_75t_L g533 ( .A1(n_521), .A2(n_522), .B(n_528), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_523), .B(n_527), .Y(n_522) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_531), .B(n_543), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_531), .B(n_589), .Y(n_674) );
AND2x4_ASAP7_75t_L g531 ( .A(n_532), .B(n_534), .Y(n_531) );
AND3x2_ASAP7_75t_L g629 ( .A(n_532), .B(n_576), .C(n_585), .Y(n_629) );
AND2x2_ASAP7_75t_L g553 ( .A(n_533), .B(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_533), .B(n_536), .Y(n_610) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
OR2x2_ASAP7_75t_L g564 ( .A(n_535), .B(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g554 ( .A(n_536), .Y(n_554) );
INVx1_ASAP7_75t_L g569 ( .A(n_536), .Y(n_569) );
BUFx3_ASAP7_75t_L g576 ( .A(n_536), .Y(n_576) );
AND2x2_ASAP7_75t_L g586 ( .A(n_536), .B(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
AND2x4_ASAP7_75t_L g595 ( .A(n_544), .B(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_544), .B(n_554), .Y(n_638) );
AND2x2_ASAP7_75t_L g594 ( .A(n_545), .B(n_569), .Y(n_594) );
INVx2_ASAP7_75t_L g621 ( .A(n_545), .Y(n_621) );
INVx1_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
AOI211xp5_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_555), .B(n_560), .C(n_581), .Y(n_549) );
OAI21xp5_ASAP7_75t_L g701 ( .A1(n_550), .A2(n_677), .B(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_553), .B(n_612), .Y(n_611) );
AOI211xp5_ASAP7_75t_SL g631 ( .A1(n_553), .A2(n_632), .B(n_636), .C(n_645), .Y(n_631) );
AND2x2_ASAP7_75t_L g617 ( .A(n_554), .B(n_577), .Y(n_617) );
OR2x2_ASAP7_75t_L g620 ( .A(n_554), .B(n_621), .Y(n_620) );
INVx1_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_557), .B(n_558), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g707 ( .A(n_557), .B(n_662), .Y(n_707) );
NAND2xp5_ASAP7_75t_SL g616 ( .A(n_558), .B(n_603), .Y(n_616) );
AOI221xp5_ASAP7_75t_L g672 ( .A1(n_558), .A2(n_584), .B1(n_664), .B2(n_667), .C(n_673), .Y(n_672) );
AND2x4_ASAP7_75t_L g589 ( .A(n_559), .B(n_590), .Y(n_589) );
OR2x2_ASAP7_75t_L g635 ( .A(n_559), .B(n_590), .Y(n_635) );
OAI221xp5_ASAP7_75t_SL g560 ( .A1(n_561), .A2(n_564), .B1(n_567), .B2(n_571), .C(n_574), .Y(n_560) );
AND2x2_ASAP7_75t_L g706 ( .A(n_561), .B(n_707), .Y(n_706) );
OR2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
INVx1_ASAP7_75t_L g573 ( .A(n_562), .Y(n_573) );
INVx1_ASAP7_75t_L g659 ( .A(n_563), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g680 ( .A(n_564), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g578 ( .A(n_566), .B(n_569), .Y(n_578) );
AND2x2_ASAP7_75t_L g654 ( .A(n_566), .B(n_655), .Y(n_654) );
OR2x2_ASAP7_75t_L g567 ( .A(n_568), .B(n_570), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_SL g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g579 ( .A(n_573), .B(n_580), .Y(n_579) );
OAI21xp5_ASAP7_75t_SL g574 ( .A1(n_575), .A2(n_578), .B(n_579), .Y(n_574) );
INVx1_ASAP7_75t_L g698 ( .A(n_575), .Y(n_698) );
AND2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
AND2x2_ASAP7_75t_L g677 ( .A(n_576), .B(n_604), .Y(n_677) );
AND2x2_ASAP7_75t_SL g650 ( .A(n_577), .B(n_586), .Y(n_650) );
AOI21xp33_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_583), .B(n_588), .Y(n_581) );
OAI22xp33_ASAP7_75t_L g618 ( .A1(n_582), .A2(n_616), .B1(n_619), .B2(n_620), .Y(n_618) );
INVx1_ASAP7_75t_L g688 ( .A(n_582), .Y(n_688) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
INVx1_ASAP7_75t_L g608 ( .A(n_585), .Y(n_608) );
INVx1_ASAP7_75t_L g669 ( .A(n_587), .Y(n_669) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_589), .B(n_591), .Y(n_588) );
NAND2xp5_ASAP7_75t_SL g710 ( .A(n_589), .B(n_659), .Y(n_710) );
AND2x2_ASAP7_75t_L g678 ( .A(n_590), .B(n_679), .Y(n_678) );
OAI211xp5_ASAP7_75t_L g671 ( .A1(n_591), .A2(n_672), .B(n_675), .C(n_683), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_593), .B(n_614), .Y(n_592) );
AOI322xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_595), .A3(n_597), .B1(n_599), .B2(n_604), .C1(n_605), .C2(n_613), .Y(n_593) );
CKINVDCx16_ASAP7_75t_R g711 ( .A(n_595), .Y(n_711) );
AND2x2_ASAP7_75t_L g661 ( .A(n_596), .B(n_662), .Y(n_661) );
INVx1_ASAP7_75t_SL g695 ( .A(n_596), .Y(n_695) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NOR2xp33_ASAP7_75t_SL g646 ( .A(n_598), .B(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_SL g652 ( .A(n_598), .B(n_644), .Y(n_652) );
AND2x2_ASAP7_75t_L g676 ( .A(n_598), .B(n_642), .Y(n_676) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
INVx1_ASAP7_75t_L g648 ( .A(n_602), .Y(n_648) );
NAND2xp33_ASAP7_75t_SL g605 ( .A(n_606), .B(n_611), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
AOI221xp5_ASAP7_75t_SL g651 ( .A1(n_607), .A2(n_652), .B1(n_653), .B2(n_654), .C(n_656), .Y(n_651) );
AND2x2_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
INVxp67_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g718 ( .A(n_610), .Y(n_718) );
AOI211xp5_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_617), .B(n_618), .C(n_622), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_SL g693 ( .A(n_617), .Y(n_693) );
INVx1_ASAP7_75t_L g625 ( .A(n_619), .Y(n_625) );
OR2x2_ASAP7_75t_L g712 ( .A(n_619), .B(n_713), .Y(n_712) );
INVx2_ASAP7_75t_SL g708 ( .A(n_620), .Y(n_708) );
AOI21xp33_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_626), .B(n_628), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_624), .B(n_642), .Y(n_719) );
INVx1_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_651), .Y(n_630) );
INVx1_ASAP7_75t_SL g632 ( .A(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_634), .B(n_658), .Y(n_657) );
INVx1_ASAP7_75t_SL g634 ( .A(n_635), .Y(n_634) );
OR2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_639), .Y(n_637) );
OR2x2_ASAP7_75t_L g685 ( .A(n_638), .B(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AOI21xp33_ASAP7_75t_SL g645 ( .A1(n_646), .A2(n_648), .B(n_649), .Y(n_645) );
INVx2_ASAP7_75t_SL g649 ( .A(n_650), .Y(n_649) );
AOI31xp33_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_660), .A3(n_663), .B(n_665), .Y(n_656) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_662), .B(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_SL g665 ( .A(n_666), .Y(n_665) );
AND2x4_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
AOI221xp5_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_687), .B1(n_688), .B2(n_689), .C(n_692), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVxp67_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
OAI22xp5_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_694), .B1(n_696), .B2(n_698), .Y(n_692) );
CKINVDCx16_ASAP7_75t_R g696 ( .A(n_697), .Y(n_696) );
NOR3xp33_ASAP7_75t_L g699 ( .A(n_700), .B(n_709), .C(n_716), .Y(n_699) );
NAND2xp5_ASAP7_75t_SL g700 ( .A(n_701), .B(n_704), .Y(n_700) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_705), .B(n_708), .Y(n_704) );
INVxp67_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_717), .B(n_719), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
BUFx4f_ASAP7_75t_SL g720 ( .A(n_721), .Y(n_720) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_SL g729 ( .A(n_722), .Y(n_729) );
CKINVDCx11_ASAP7_75t_R g722 ( .A(n_723), .Y(n_722) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_728), .B1(n_729), .B2(n_730), .Y(n_726) );
CKINVDCx5p33_ASAP7_75t_R g731 ( .A(n_732), .Y(n_731) );
CKINVDCx5p33_ASAP7_75t_R g732 ( .A(n_733), .Y(n_732) );
INVx3_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_736), .B(n_739), .Y(n_735) );
HB1xp67_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
HB1xp67_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVxp67_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
AOI21xp5_ASAP7_75t_L g747 ( .A1(n_740), .A2(n_748), .B(n_757), .Y(n_747) );
NOR2xp33_ASAP7_75t_SL g740 ( .A(n_741), .B(n_742), .Y(n_740) );
BUFx2_ASAP7_75t_R g759 ( .A(n_741), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_744), .B(n_747), .Y(n_743) );
HB1xp67_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
CKINVDCx5p33_ASAP7_75t_R g745 ( .A(n_746), .Y(n_745) );
INVx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g756 ( .A(n_750), .Y(n_756) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_SL g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_SL g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
CKINVDCx20_ASAP7_75t_R g770 ( .A(n_761), .Y(n_770) );
INVx2_ASAP7_75t_SL g761 ( .A(n_762), .Y(n_761) );
AND2x2_ASAP7_75t_SL g762 ( .A(n_763), .B(n_764), .Y(n_762) );
NOR2xp33_ASAP7_75t_L g768 ( .A(n_769), .B(n_770), .Y(n_768) );
endmodule