module real_jpeg_31266_n_15 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_328;
wire n_149;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_0),
.Y(n_146)
);

BUFx12f_ASAP7_75t_L g277 ( 
.A(n_0),
.Y(n_277)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

OAI21xp33_ASAP7_75t_L g125 ( 
.A1(n_1),
.A2(n_126),
.B(n_127),
.Y(n_125)
);

OAI32xp33_ASAP7_75t_L g205 ( 
.A1(n_1),
.A2(n_206),
.A3(n_210),
.B1(n_213),
.B2(n_220),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_1),
.A2(n_58),
.B1(n_237),
.B2(n_242),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_1),
.B(n_282),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_1),
.B(n_352),
.Y(n_351)
);

AO22x1_ASAP7_75t_L g198 ( 
.A1(n_2),
.A2(n_199),
.B1(n_200),
.B2(n_204),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_2),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_2),
.A2(n_199),
.B1(n_391),
.B2(n_395),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_3),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_3),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_3),
.Y(n_380)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_4),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_4),
.Y(n_177)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_5),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_6),
.Y(n_82)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_6),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_6),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_7),
.A2(n_86),
.B1(n_89),
.B2(n_90),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_7),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_7),
.A2(n_89),
.B1(n_134),
.B2(n_138),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_7),
.A2(n_89),
.B1(n_260),
.B2(n_263),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_7),
.A2(n_89),
.B1(n_365),
.B2(n_369),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_8),
.Y(n_289)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_8),
.Y(n_360)
);

OAI22x1_ASAP7_75t_L g295 ( 
.A1(n_9),
.A2(n_296),
.B1(n_301),
.B2(n_302),
.Y(n_295)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_9),
.Y(n_301)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_10),
.Y(n_71)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_10),
.Y(n_96)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_10),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_11),
.A2(n_42),
.B1(n_47),
.B2(n_53),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_11),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_11),
.A2(n_53),
.B1(n_231),
.B2(n_233),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_11),
.A2(n_53),
.B1(n_400),
.B2(n_403),
.Y(n_399)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_12),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_12),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_12),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_12),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_13),
.A2(n_332),
.B1(n_334),
.B2(n_335),
.Y(n_331)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_13),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_14),
.A2(n_31),
.B1(n_34),
.B2(n_38),
.Y(n_30)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_14),
.A2(n_38),
.B1(n_180),
.B2(n_183),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_14),
.A2(n_38),
.B1(n_308),
.B2(n_311),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_317),
.Y(n_15)
);

HB1xp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_266),
.B(n_316),
.Y(n_17)
);

O2A1O1Ixp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_159),
.B(n_188),
.C(n_189),
.Y(n_18)
);

AOI21x1_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_123),
.B(n_158),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_54),
.Y(n_20)
);

NOR2xp67_ASAP7_75t_L g158 ( 
.A(n_21),
.B(n_54),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_29),
.B1(n_39),
.B2(n_40),
.Y(n_21)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_22),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_22),
.B(n_133),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_22),
.A2(n_295),
.B1(n_328),
.B2(n_331),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_26),
.Y(n_22)
);

INVx3_ASAP7_75t_SL g39 ( 
.A(n_23),
.Y(n_39)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_25),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_25),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_25),
.Y(n_197)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_28),
.Y(n_149)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_28),
.Y(n_203)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_28),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

OAI21xp33_ASAP7_75t_SL g153 ( 
.A1(n_30),
.A2(n_154),
.B(n_156),
.Y(n_153)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_33),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_37),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_39),
.B(n_295),
.Y(n_294)
);

INVxp33_ASAP7_75t_SL g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_41),
.A2(n_126),
.B(n_127),
.Y(n_162)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22x1_ASAP7_75t_L g93 ( 
.A1(n_45),
.A2(n_94),
.B1(n_97),
.B2(n_100),
.Y(n_93)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_52),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_83),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_55),
.B(n_83),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_62),
.B1(n_72),
.B2(n_78),
.Y(n_55)
);

INVxp67_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

OAI21xp33_ASAP7_75t_L g103 ( 
.A1(n_57),
.A2(n_58),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_58),
.B(n_142),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_58),
.B(n_152),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_58),
.B(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_58),
.B(n_221),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_58),
.A2(n_385),
.B(n_386),
.Y(n_384)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_59),
.Y(n_212)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_61),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_61),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_65),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_79),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_82),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_102),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_84),
.A2(n_111),
.B(n_230),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_92),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_85),
.B(n_110),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_85),
.A2(n_92),
.B1(n_110),
.B2(n_389),
.Y(n_388)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g152 ( 
.A(n_92),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_93),
.Y(n_228)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_99),
.Y(n_304)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_99),
.Y(n_333)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_110),
.Y(n_102)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_108),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g174 ( 
.A(n_109),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_110),
.A2(n_226),
.B1(n_227),
.B2(n_229),
.Y(n_225)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_116),
.B1(n_118),
.B2(n_121),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_SL g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_115),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_115),
.Y(n_234)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_115),
.Y(n_394)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

OAI21xp33_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_150),
.B(n_157),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_140),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_126),
.A2(n_198),
.B(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_133),
.Y(n_127)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_147),
.Y(n_140)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_146),
.Y(n_330)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_153),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_151),
.B(n_153),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_152),
.A2(n_179),
.B(n_187),
.Y(n_178)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_156),
.A2(n_196),
.B(n_198),
.Y(n_195)
);

INVxp67_ASAP7_75t_SL g278 ( 
.A(n_156),
.Y(n_278)
);

NOR2xp67_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_160),
.B(n_161),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_191),
.C(n_192),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_178),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_164),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_165),
.A2(n_306),
.B(n_312),
.Y(n_305)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_165),
.Y(n_408)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_166),
.B(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_167),
.B(n_249),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_170),
.B1(n_173),
.B2(n_175),
.Y(n_167)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_169),
.Y(n_223)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_172),
.Y(n_255)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_174),
.Y(n_232)
);

INVx5_ASAP7_75t_SL g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_177),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_179),
.Y(n_226)
);

INVx1_ASAP7_75t_SL g180 ( 
.A(n_181),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_184),
.Y(n_183)
);

INVx4_ASAP7_75t_SL g184 ( 
.A(n_185),
.Y(n_184)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_193),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g315 ( 
.A(n_190),
.B(n_193),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_224),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_194),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_205),
.Y(n_194)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_R g274 ( 
.A(n_198),
.B(n_275),
.Y(n_274)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_201),
.Y(n_200)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_202),
.Y(n_204)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_205),
.A2(n_274),
.B(n_278),
.Y(n_273)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_208),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_209),
.Y(n_402)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_216),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_219),
.Y(n_252)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_235),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_225),
.B(n_235),
.C(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

OA21x2_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_247),
.B(n_258),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_241),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_241),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_241),
.Y(n_342)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_241),
.Y(n_407)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_SL g250 ( 
.A(n_246),
.Y(n_250)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_246),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_246),
.Y(n_310)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

NAND2xp33_ASAP7_75t_SL g312 ( 
.A(n_248),
.B(n_259),
.Y(n_312)
);

AOI22x1_ASAP7_75t_L g397 ( 
.A1(n_248),
.A2(n_307),
.B1(n_398),
.B2(n_408),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_253),
.B2(n_256),
.Y(n_249)
);

INVx2_ASAP7_75t_SL g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_254),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx8_ASAP7_75t_L g292 ( 
.A(n_257),
.Y(n_292)
);

INVxp67_ASAP7_75t_SL g260 ( 
.A(n_261),
.Y(n_260)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_315),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_313),
.Y(n_267)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_268),
.B(n_313),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_279),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_272),
.B2(n_273),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_270),
.B(n_273),
.C(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx8_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_279),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_305),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_293),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_281),
.B(n_305),
.C(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_282),
.B(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_283),
.B(n_373),
.Y(n_372)
);

AOI22x1_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_288),
.B1(n_290),
.B2(n_291),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx8_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_288),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_289),
.Y(n_345)
);

INVx5_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx5_ASAP7_75t_L g356 ( 
.A(n_292),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_293),
.Y(n_324)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_310),
.Y(n_311)
);

NAND2xp33_ASAP7_75t_SL g317 ( 
.A(n_318),
.B(n_412),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_320),
.B(n_409),
.Y(n_319)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_320),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_361),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_322),
.A2(n_323),
.B1(n_325),
.B2(n_326),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_338),
.Y(n_326)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_SL g329 ( 
.A(n_330),
.Y(n_329)
);

BUFx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

AOI32xp33_ASAP7_75t_L g338 ( 
.A1(n_339),
.A2(n_343),
.A3(n_346),
.B1(n_351),
.B2(n_355),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_345),
.Y(n_376)
);

INVx4_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx11_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

BUFx12f_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx6_ASAP7_75t_L g354 ( 
.A(n_350),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g370 ( 
.A(n_350),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_350),
.Y(n_375)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_351),
.Y(n_386)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

NAND2xp33_ASAP7_75t_R g355 ( 
.A(n_356),
.B(n_357),
.Y(n_355)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_360),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_387),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_371),
.Y(n_362)
);

INVx3_ASAP7_75t_SL g365 ( 
.A(n_366),
.Y(n_365)
);

INVx4_ASAP7_75t_SL g366 ( 
.A(n_367),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_369),
.Y(n_385)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_372),
.B(n_384),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_374),
.A2(n_376),
.B1(n_377),
.B2(n_381),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx6_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_382),
.Y(n_381)
);

INVx4_ASAP7_75t_SL g382 ( 
.A(n_383),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_397),
.Y(n_387)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

BUFx4f_ASAP7_75t_SL g392 ( 
.A(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

BUFx2_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_410),
.B(n_413),
.Y(n_412)
);


endmodule