module fake_netlist_5_1162_n_324 (n_91, n_82, n_10, n_24, n_86, n_83, n_61, n_90, n_75, n_65, n_78, n_74, n_57, n_96, n_37, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_0, n_58, n_9, n_69, n_18, n_42, n_22, n_1, n_45, n_46, n_21, n_94, n_38, n_80, n_4, n_35, n_73, n_17, n_92, n_19, n_30, n_5, n_33, n_14, n_84, n_23, n_29, n_79, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_71, n_85, n_95, n_59, n_26, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_36, n_76, n_87, n_27, n_64, n_77, n_81, n_28, n_89, n_70, n_68, n_93, n_72, n_32, n_41, n_56, n_51, n_63, n_97, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_324);

input n_91;
input n_82;
input n_10;
input n_24;
input n_86;
input n_83;
input n_61;
input n_90;
input n_75;
input n_65;
input n_78;
input n_74;
input n_57;
input n_96;
input n_37;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_42;
input n_22;
input n_1;
input n_45;
input n_46;
input n_21;
input n_94;
input n_38;
input n_80;
input n_4;
input n_35;
input n_73;
input n_17;
input n_92;
input n_19;
input n_30;
input n_5;
input n_33;
input n_14;
input n_84;
input n_23;
input n_29;
input n_79;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_71;
input n_85;
input n_95;
input n_59;
input n_26;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_81;
input n_28;
input n_89;
input n_70;
input n_68;
input n_93;
input n_72;
input n_32;
input n_41;
input n_56;
input n_51;
input n_63;
input n_97;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;

output n_324;

wire n_137;
wire n_294;
wire n_318;
wire n_194;
wire n_316;
wire n_248;
wire n_136;
wire n_124;
wire n_146;
wire n_315;
wire n_268;
wire n_127;
wire n_235;
wire n_226;
wire n_111;
wire n_155;
wire n_116;
wire n_284;
wire n_245;
wire n_139;
wire n_105;
wire n_280;
wire n_254;
wire n_302;
wire n_265;
wire n_293;
wire n_244;
wire n_173;
wire n_198;
wire n_247;
wire n_314;
wire n_321;
wire n_292;
wire n_212;
wire n_119;
wire n_275;
wire n_252;
wire n_295;
wire n_133;
wire n_147;
wire n_307;
wire n_150;
wire n_106;
wire n_209;
wire n_259;
wire n_301;
wire n_186;
wire n_134;
wire n_191;
wire n_171;
wire n_153;
wire n_204;
wire n_250;
wire n_260;
wire n_298;
wire n_320;
wire n_286;
wire n_122;
wire n_282;
wire n_132;
wire n_101;
wire n_281;
wire n_240;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_152;
wire n_317;
wire n_323;
wire n_195;
wire n_227;
wire n_271;
wire n_123;
wire n_167;
wire n_234;
wire n_308;
wire n_267;
wire n_297;
wire n_156;
wire n_225;
wire n_219;
wire n_157;
wire n_131;
wire n_192;
wire n_223;
wire n_158;
wire n_138;
wire n_264;
wire n_109;
wire n_163;
wire n_276;
wire n_183;
wire n_185;
wire n_243;
wire n_169;
wire n_255;
wire n_215;
wire n_196;
wire n_211;
wire n_218;
wire n_181;
wire n_290;
wire n_221;
wire n_178;
wire n_287;
wire n_104;
wire n_141;
wire n_145;
wire n_313;
wire n_216;
wire n_168;
wire n_164;
wire n_311;
wire n_208;
wire n_142;
wire n_214;
wire n_140;
wire n_299;
wire n_303;
wire n_296;
wire n_241;
wire n_184;
wire n_144;
wire n_114;
wire n_165;
wire n_213;
wire n_129;
wire n_197;
wire n_107;
wire n_236;
wire n_249;
wire n_304;
wire n_203;
wire n_274;
wire n_277;
wire n_149;
wire n_309;
wire n_130;
wire n_322;
wire n_258;
wire n_151;
wire n_306;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_224;
wire n_228;
wire n_283;
wire n_112;
wire n_239;
wire n_310;
wire n_170;
wire n_102;
wire n_161;
wire n_273;
wire n_270;
wire n_230;
wire n_118;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_172;
wire n_206;
wire n_217;
wire n_312;
wire n_210;
wire n_176;
wire n_182;
wire n_143;
wire n_237;
wire n_180;
wire n_207;
wire n_229;
wire n_108;
wire n_177;
wire n_117;
wire n_233;
wire n_205;
wire n_113;
wire n_246;
wire n_179;
wire n_125;
wire n_269;
wire n_128;
wire n_285;
wire n_120;
wire n_232;
wire n_135;
wire n_126;
wire n_202;
wire n_266;
wire n_272;
wire n_193;
wire n_251;
wire n_160;
wire n_154;
wire n_148;
wire n_300;
wire n_159;
wire n_175;
wire n_262;
wire n_238;
wire n_319;
wire n_121;
wire n_242;
wire n_200;
wire n_162;
wire n_222;
wire n_115;
wire n_199;
wire n_187;
wire n_103;
wire n_166;
wire n_256;
wire n_305;
wire n_278;
wire n_110;

INVxp67_ASAP7_75t_SL g101 ( 
.A(n_7),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_0),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_33),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_23),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_35),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_66),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_46),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_64),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_70),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_41),
.Y(n_114)
);

CKINVDCx5p33_ASAP7_75t_R g115 ( 
.A(n_52),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_50),
.Y(n_116)
);

INVxp33_ASAP7_75t_SL g117 ( 
.A(n_19),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_62),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_94),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_84),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_14),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_5),
.Y(n_122)
);

INVxp33_ASAP7_75t_L g123 ( 
.A(n_43),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_8),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_18),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_29),
.Y(n_129)
);

INVxp67_ASAP7_75t_SL g130 ( 
.A(n_63),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_77),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_36),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_6),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_11),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_85),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_44),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_15),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_81),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_56),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_73),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_96),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_49),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_79),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_42),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_48),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_93),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_90),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g149 ( 
.A(n_92),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_100),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_10),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_30),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_67),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_68),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_91),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_1),
.Y(n_156)
);

OAI21x1_ASAP7_75t_L g157 ( 
.A1(n_107),
.A2(n_54),
.B(n_98),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_149),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_115),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_109),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_110),
.A2(n_126),
.B1(n_117),
.B2(n_101),
.Y(n_161)
);

AND2x4_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_1),
.Y(n_162)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_122),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_104),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_134),
.Y(n_165)
);

OA21x2_ASAP7_75t_L g166 ( 
.A1(n_102),
.A2(n_2),
.B(n_3),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_131),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_103),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_105),
.Y(n_169)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_131),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_106),
.Y(n_171)
);

AND2x6_ASAP7_75t_L g172 ( 
.A(n_131),
.B(n_9),
.Y(n_172)
);

NAND2xp33_ASAP7_75t_L g173 ( 
.A(n_149),
.B(n_3),
.Y(n_173)
);

AND2x4_ASAP7_75t_L g174 ( 
.A(n_128),
.B(n_4),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_148),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_108),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_133),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_111),
.Y(n_178)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_140),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_149),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_159),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_179),
.B(n_119),
.Y(n_182)
);

AND2x6_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_112),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_163),
.B(n_143),
.Y(n_184)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_172),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_170),
.Y(n_186)
);

INVx3_ASAP7_75t_R g187 ( 
.A(n_162),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_160),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_161),
.B(n_150),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_168),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_113),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_114),
.Y(n_192)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_172),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_170),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_156),
.B(n_174),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_167),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_172),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_176),
.B(n_116),
.Y(n_199)
);

AOI21x1_ASAP7_75t_L g200 ( 
.A1(n_158),
.A2(n_155),
.B(n_154),
.Y(n_200)
);

OR2x6_ASAP7_75t_L g201 ( 
.A(n_164),
.B(n_118),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_178),
.Y(n_202)
);

AND2x4_ASAP7_75t_L g203 ( 
.A(n_165),
.B(n_130),
.Y(n_203)
);

NAND2xp33_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_149),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_173),
.A2(n_137),
.B1(n_152),
.B2(n_151),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_177),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_181),
.B(n_175),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_184),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_186),
.Y(n_209)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_201),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_120),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_188),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_183),
.B(n_180),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_197),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_183),
.B(n_121),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_124),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_200),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_196),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_191),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_194),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_190),
.Y(n_221)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_185),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_192),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_202),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_125),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_189),
.B(n_127),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_199),
.Y(n_227)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_193),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_193),
.B(n_129),
.Y(n_230)
);

A2O1A1Ixp33_ASAP7_75t_L g231 ( 
.A1(n_204),
.A2(n_157),
.B(n_141),
.C(n_153),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_226),
.A2(n_198),
.B1(n_139),
.B2(n_147),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_212),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_208),
.A2(n_198),
.B1(n_138),
.B2(n_146),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_214),
.Y(n_235)
);

NAND2x1p5_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_166),
.Y(n_236)
);

AO22x1_ASAP7_75t_L g237 ( 
.A1(n_219),
.A2(n_145),
.B1(n_144),
.B2(n_142),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_209),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_220),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_132),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_135),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_218),
.Y(n_242)
);

BUFx8_ASAP7_75t_SL g243 ( 
.A(n_221),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_224),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_216),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_229),
.A2(n_57),
.B(n_97),
.Y(n_246)
);

AND2x2_ASAP7_75t_SL g247 ( 
.A(n_207),
.B(n_225),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_223),
.Y(n_248)
);

AO32x1_ASAP7_75t_L g249 ( 
.A1(n_230),
.A2(n_12),
.A3(n_13),
.B1(n_16),
.B2(n_17),
.Y(n_249)
);

O2A1O1Ixp33_ASAP7_75t_SL g250 ( 
.A1(n_231),
.A2(n_20),
.B(n_21),
.C(n_22),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_227),
.B(n_24),
.Y(n_251)
);

O2A1O1Ixp5_ASAP7_75t_L g252 ( 
.A1(n_215),
.A2(n_25),
.B(n_26),
.C(n_27),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g253 ( 
.A(n_206),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_213),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_244),
.Y(n_255)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_238),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_235),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_248),
.B(n_210),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_235),
.Y(n_259)
);

AO31x2_ASAP7_75t_L g260 ( 
.A1(n_241),
.A2(n_211),
.A3(n_217),
.B(n_222),
.Y(n_260)
);

AO21x2_ASAP7_75t_L g261 ( 
.A1(n_251),
.A2(n_217),
.B(n_228),
.Y(n_261)
);

OAI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_253),
.A2(n_228),
.B1(n_222),
.B2(n_32),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_240),
.A2(n_228),
.B1(n_222),
.B2(n_34),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_28),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_242),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_245),
.A2(n_31),
.B1(n_37),
.B2(n_38),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_233),
.B(n_39),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g268 ( 
.A1(n_254),
.A2(n_95),
.B1(n_40),
.B2(n_45),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_247),
.B(n_47),
.Y(n_269)
);

INVx5_ASAP7_75t_L g270 ( 
.A(n_254),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_239),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_259),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_259),
.Y(n_273)
);

NAND3xp33_ASAP7_75t_L g274 ( 
.A(n_269),
.B(n_237),
.C(n_234),
.Y(n_274)
);

OAI221xp5_ASAP7_75t_L g275 ( 
.A1(n_267),
.A2(n_232),
.B1(n_238),
.B2(n_236),
.C(n_252),
.Y(n_275)
);

AO21x2_ASAP7_75t_L g276 ( 
.A1(n_264),
.A2(n_250),
.B(n_246),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_257),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_265),
.Y(n_278)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_270),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_255),
.Y(n_280)
);

AOI21xp33_ASAP7_75t_SL g281 ( 
.A1(n_266),
.A2(n_243),
.B(n_51),
.Y(n_281)
);

AOI222xp33_ASAP7_75t_L g282 ( 
.A1(n_266),
.A2(n_268),
.B1(n_271),
.B2(n_258),
.C1(n_256),
.C2(n_263),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_268),
.A2(n_249),
.B1(n_53),
.B2(n_55),
.Y(n_283)
);

INVx6_ASAP7_75t_L g284 ( 
.A(n_256),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_272),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_273),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_278),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_277),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_280),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_279),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_284),
.Y(n_291)
);

NAND3xp33_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_263),
.C(n_270),
.Y(n_292)
);

BUFx4f_ASAP7_75t_SL g293 ( 
.A(n_281),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_293),
.A2(n_282),
.B1(n_283),
.B2(n_275),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_287),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_288),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_285),
.Y(n_297)
);

NOR3xp33_ASAP7_75t_L g298 ( 
.A(n_292),
.B(n_283),
.C(n_262),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_286),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_290),
.Y(n_300)
);

AOI221xp5_ASAP7_75t_L g301 ( 
.A1(n_294),
.A2(n_276),
.B1(n_261),
.B2(n_58),
.C(n_59),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_300),
.B(n_260),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_295),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_296),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_297),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_299),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_303),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_305),
.B(n_298),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_306),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_304),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_307),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_308),
.A2(n_301),
.B(n_298),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_311),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_312),
.A2(n_302),
.B1(n_309),
.B2(n_310),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_313),
.B(n_314),
.Y(n_315)
);

INVx2_ASAP7_75t_SL g316 ( 
.A(n_315),
.Y(n_316)
);

OR2x6_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_60),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_317),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_318),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_319),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_320),
.A2(n_65),
.B1(n_71),
.B2(n_72),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_321),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_322),
.A2(n_75),
.B1(n_76),
.B2(n_78),
.Y(n_323)
);

OAI22xp33_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_83),
.B1(n_87),
.B2(n_88),
.Y(n_324)
);


endmodule