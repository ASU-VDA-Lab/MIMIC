module fake_aes_3782_n_539 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_539);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_539;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g77 ( .A(n_35), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_31), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_27), .Y(n_79) );
INVxp67_ASAP7_75t_L g80 ( .A(n_68), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_23), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_16), .Y(n_82) );
BUFx3_ASAP7_75t_L g83 ( .A(n_7), .Y(n_83) );
CKINVDCx16_ASAP7_75t_R g84 ( .A(n_28), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_63), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_19), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_46), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_71), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_14), .Y(n_89) );
INVxp67_ASAP7_75t_L g90 ( .A(n_22), .Y(n_90) );
INVx1_ASAP7_75t_SL g91 ( .A(n_69), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_20), .Y(n_92) );
INVxp67_ASAP7_75t_SL g93 ( .A(n_48), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_59), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_60), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_36), .Y(n_96) );
BUFx8_ASAP7_75t_SL g97 ( .A(n_16), .Y(n_97) );
CKINVDCx20_ASAP7_75t_R g98 ( .A(n_34), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_17), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_76), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_55), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_49), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_8), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_67), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_57), .Y(n_105) );
INVxp67_ASAP7_75t_L g106 ( .A(n_6), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_18), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_7), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_24), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_25), .Y(n_110) );
INVxp33_ASAP7_75t_SL g111 ( .A(n_15), .Y(n_111) );
INVx3_ASAP7_75t_L g112 ( .A(n_83), .Y(n_112) );
HB1xp67_ASAP7_75t_L g113 ( .A(n_83), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_106), .B(n_0), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_77), .Y(n_115) );
BUFx6f_ASAP7_75t_L g116 ( .A(n_100), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_100), .Y(n_117) );
AND2x2_ASAP7_75t_L g118 ( .A(n_84), .B(n_0), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_77), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_81), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_82), .B(n_1), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_81), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_85), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_85), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_86), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_86), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_89), .B(n_1), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_87), .Y(n_128) );
OA21x2_ASAP7_75t_L g129 ( .A1(n_87), .A2(n_41), .B(n_74), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_78), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_79), .Y(n_131) );
INVx2_ASAP7_75t_L g132 ( .A(n_88), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g133 ( .A(n_103), .B(n_2), .Y(n_133) );
BUFx3_ASAP7_75t_L g134 ( .A(n_92), .Y(n_134) );
INVx6_ASAP7_75t_L g135 ( .A(n_130), .Y(n_135) );
OR2x2_ASAP7_75t_L g136 ( .A(n_113), .B(n_108), .Y(n_136) );
BUFx2_ASAP7_75t_L g137 ( .A(n_118), .Y(n_137) );
CKINVDCx16_ASAP7_75t_R g138 ( .A(n_118), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_115), .B(n_95), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_116), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_126), .Y(n_141) );
INVx4_ASAP7_75t_L g142 ( .A(n_112), .Y(n_142) );
AND2x4_ASAP7_75t_L g143 ( .A(n_115), .B(n_109), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_131), .B(n_101), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_116), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_131), .B(n_101), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g147 ( .A(n_119), .B(n_80), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_119), .B(n_104), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_116), .Y(n_149) );
OAI21xp33_ASAP7_75t_L g150 ( .A1(n_122), .A2(n_110), .B(n_107), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_116), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_126), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_126), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_126), .Y(n_154) );
AND2x2_ASAP7_75t_L g155 ( .A(n_122), .B(n_90), .Y(n_155) );
INVx2_ASAP7_75t_SL g156 ( .A(n_134), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_124), .B(n_111), .Y(n_157) );
AND2x2_ASAP7_75t_L g158 ( .A(n_124), .B(n_93), .Y(n_158) );
AND2x2_ASAP7_75t_L g159 ( .A(n_128), .B(n_98), .Y(n_159) );
AND2x4_ASAP7_75t_L g160 ( .A(n_128), .B(n_94), .Y(n_160) );
INVx1_ASAP7_75t_SL g161 ( .A(n_159), .Y(n_161) );
INVx3_ASAP7_75t_SL g162 ( .A(n_138), .Y(n_162) );
BUFx3_ASAP7_75t_L g163 ( .A(n_156), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_140), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_142), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_142), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_142), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_142), .Y(n_168) );
INVx2_ASAP7_75t_SL g169 ( .A(n_136), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_155), .B(n_134), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_140), .Y(n_171) );
AND2x4_ASAP7_75t_L g172 ( .A(n_158), .B(n_127), .Y(n_172) );
BUFx3_ASAP7_75t_L g173 ( .A(n_156), .Y(n_173) );
OR2x4_ASAP7_75t_L g174 ( .A(n_136), .B(n_157), .Y(n_174) );
AND2x4_ASAP7_75t_L g175 ( .A(n_158), .B(n_127), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_155), .B(n_134), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_143), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_143), .Y(n_178) );
HB1xp67_ASAP7_75t_L g179 ( .A(n_159), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_143), .B(n_114), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_143), .B(n_121), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_145), .Y(n_182) );
NAND2x1p5_ASAP7_75t_L g183 ( .A(n_160), .B(n_123), .Y(n_183) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_140), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_144), .B(n_132), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_160), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_146), .B(n_132), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_160), .B(n_112), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_145), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_160), .B(n_112), .Y(n_190) );
INVx4_ASAP7_75t_L g191 ( .A(n_135), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_139), .Y(n_192) );
AND2x4_ASAP7_75t_L g193 ( .A(n_137), .B(n_133), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_140), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_167), .Y(n_195) );
NAND3xp33_ASAP7_75t_L g196 ( .A(n_192), .B(n_150), .C(n_148), .Y(n_196) );
OAI22xp5_ASAP7_75t_L g197 ( .A1(n_192), .A2(n_138), .B1(n_137), .B2(n_98), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_183), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_183), .Y(n_199) );
INVx5_ASAP7_75t_L g200 ( .A(n_191), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_169), .B(n_139), .Y(n_201) );
BUFx6f_ASAP7_75t_L g202 ( .A(n_183), .Y(n_202) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_163), .Y(n_203) );
INVx5_ASAP7_75t_L g204 ( .A(n_191), .Y(n_204) );
BUFx8_ASAP7_75t_SL g205 ( .A(n_193), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_181), .A2(n_147), .B(n_148), .Y(n_206) );
BUFx6f_ASAP7_75t_L g207 ( .A(n_163), .Y(n_207) );
AOI22xp5_ASAP7_75t_L g208 ( .A1(n_161), .A2(n_150), .B1(n_105), .B2(n_102), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_167), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_177), .Y(n_210) );
OAI21x1_ASAP7_75t_L g211 ( .A1(n_164), .A2(n_129), .B(n_145), .Y(n_211) );
OAI21xp5_ASAP7_75t_L g212 ( .A1(n_177), .A2(n_129), .B(n_153), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_193), .B(n_111), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_178), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_178), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_165), .Y(n_216) );
INVx3_ASAP7_75t_L g217 ( .A(n_163), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_186), .Y(n_218) );
AND2x4_ASAP7_75t_L g219 ( .A(n_169), .B(n_102), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_174), .B(n_193), .Y(n_220) );
BUFx3_ASAP7_75t_L g221 ( .A(n_173), .Y(n_221) );
CKINVDCx5p33_ASAP7_75t_R g222 ( .A(n_162), .Y(n_222) );
INVx3_ASAP7_75t_L g223 ( .A(n_173), .Y(n_223) );
AND2x2_ASAP7_75t_L g224 ( .A(n_193), .B(n_120), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_186), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_165), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_166), .Y(n_227) );
AO21x2_ASAP7_75t_L g228 ( .A1(n_212), .A2(n_123), .B(n_125), .Y(n_228) );
AOI22xp33_ASAP7_75t_L g229 ( .A1(n_219), .A2(n_179), .B1(n_162), .B2(n_175), .Y(n_229) );
AND2x4_ASAP7_75t_L g230 ( .A(n_198), .B(n_172), .Y(n_230) );
OAI22xp5_ASAP7_75t_L g231 ( .A1(n_208), .A2(n_174), .B1(n_170), .B2(n_176), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_210), .Y(n_232) );
AND2x4_ASAP7_75t_L g233 ( .A(n_198), .B(n_172), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_216), .Y(n_234) );
OAI21xp5_ASAP7_75t_L g235 ( .A1(n_196), .A2(n_168), .B(n_166), .Y(n_235) );
AOI22xp5_ASAP7_75t_L g236 ( .A1(n_219), .A2(n_162), .B1(n_174), .B2(n_172), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_201), .B(n_224), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_224), .Y(n_238) );
BUFx2_ASAP7_75t_L g239 ( .A(n_202), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_219), .B(n_172), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_201), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_216), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_210), .Y(n_243) );
OAI22xp5_ASAP7_75t_L g244 ( .A1(n_208), .A2(n_188), .B1(n_190), .B2(n_175), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_214), .Y(n_245) );
CKINVDCx5p33_ASAP7_75t_R g246 ( .A(n_205), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_220), .B(n_175), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_214), .Y(n_248) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_219), .B(n_175), .Y(n_249) );
AND2x4_ASAP7_75t_L g250 ( .A(n_199), .B(n_180), .Y(n_250) );
AOI22xp33_ASAP7_75t_SL g251 ( .A1(n_197), .A2(n_105), .B1(n_97), .B2(n_185), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_215), .Y(n_252) );
CKINVDCx16_ASAP7_75t_R g253 ( .A(n_202), .Y(n_253) );
OR2x2_ASAP7_75t_L g254 ( .A(n_213), .B(n_187), .Y(n_254) );
BUFx6f_ASAP7_75t_L g255 ( .A(n_239), .Y(n_255) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_240), .A2(n_196), .B(n_249), .C(n_254), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_234), .Y(n_257) );
OR2x6_ASAP7_75t_L g258 ( .A(n_234), .B(n_202), .Y(n_258) );
AOI22xp33_ASAP7_75t_L g259 ( .A1(n_251), .A2(n_199), .B1(n_202), .B2(n_225), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_241), .B(n_202), .Y(n_260) );
HB1xp67_ASAP7_75t_L g261 ( .A(n_253), .Y(n_261) );
AND2x4_ASAP7_75t_L g262 ( .A(n_232), .B(n_202), .Y(n_262) );
AND2x4_ASAP7_75t_L g263 ( .A(n_232), .B(n_215), .Y(n_263) );
AND2x4_ASAP7_75t_L g264 ( .A(n_248), .B(n_218), .Y(n_264) );
OAI22xp5_ASAP7_75t_L g265 ( .A1(n_236), .A2(n_229), .B1(n_244), .B2(n_237), .Y(n_265) );
AND2x2_ASAP7_75t_L g266 ( .A(n_230), .B(n_218), .Y(n_266) );
OAI22xp5_ASAP7_75t_L g267 ( .A1(n_231), .A2(n_221), .B1(n_207), .B2(n_203), .Y(n_267) );
BUFx4f_ASAP7_75t_SL g268 ( .A(n_230), .Y(n_268) );
OAI221xp5_ASAP7_75t_L g269 ( .A1(n_247), .A2(n_222), .B1(n_206), .B2(n_225), .C(n_120), .Y(n_269) );
NAND3xp33_ASAP7_75t_L g270 ( .A(n_235), .B(n_130), .C(n_116), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g271 ( .A1(n_230), .A2(n_97), .B1(n_227), .B2(n_216), .Y(n_271) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_233), .A2(n_227), .B1(n_226), .B2(n_209), .Y(n_272) );
AOI222xp33_ASAP7_75t_L g273 ( .A1(n_238), .A2(n_125), .B1(n_123), .B2(n_120), .C1(n_226), .C2(n_117), .Y(n_273) );
NAND3xp33_ASAP7_75t_L g274 ( .A(n_248), .B(n_130), .C(n_116), .Y(n_274) );
INVx3_ASAP7_75t_L g275 ( .A(n_242), .Y(n_275) );
OA21x2_ASAP7_75t_L g276 ( .A1(n_242), .A2(n_212), .B(n_211), .Y(n_276) );
OAI22xp33_ASAP7_75t_L g277 ( .A1(n_268), .A2(n_246), .B1(n_254), .B2(n_252), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_257), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_257), .Y(n_279) );
INVx1_ASAP7_75t_SL g280 ( .A(n_261), .Y(n_280) );
AO21x2_ASAP7_75t_L g281 ( .A1(n_270), .A2(n_228), .B(n_211), .Y(n_281) );
NOR2x1_ASAP7_75t_R g282 ( .A(n_262), .B(n_246), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_260), .B(n_233), .Y(n_283) );
AOI222xp33_ASAP7_75t_L g284 ( .A1(n_265), .A2(n_233), .B1(n_245), .B2(n_243), .C1(n_250), .C2(n_125), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_257), .Y(n_285) );
OAI22xp5_ASAP7_75t_L g286 ( .A1(n_256), .A2(n_239), .B1(n_250), .B2(n_221), .Y(n_286) );
AOI22xp33_ASAP7_75t_L g287 ( .A1(n_259), .A2(n_250), .B1(n_226), .B2(n_112), .Y(n_287) );
OAI22xp5_ASAP7_75t_L g288 ( .A1(n_272), .A2(n_221), .B1(n_207), .B2(n_203), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_263), .Y(n_289) );
AOI221xp5_ASAP7_75t_L g290 ( .A1(n_271), .A2(n_117), .B1(n_126), .B2(n_130), .C(n_99), .Y(n_290) );
BUFx3_ASAP7_75t_L g291 ( .A(n_255), .Y(n_291) );
INVxp67_ASAP7_75t_L g292 ( .A(n_262), .Y(n_292) );
OAI33xp33_ASAP7_75t_L g293 ( .A1(n_267), .A2(n_96), .A3(n_152), .B1(n_153), .B2(n_154), .B3(n_141), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_263), .Y(n_294) );
BUFx3_ASAP7_75t_L g295 ( .A(n_255), .Y(n_295) );
BUFx2_ASAP7_75t_L g296 ( .A(n_258), .Y(n_296) );
OAI221xp5_ASAP7_75t_L g297 ( .A1(n_269), .A2(n_130), .B1(n_126), .B2(n_195), .C(n_209), .Y(n_297) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_262), .Y(n_298) );
INVx4_ASAP7_75t_L g299 ( .A(n_291), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_280), .B(n_260), .Y(n_300) );
INVx2_ASAP7_75t_SL g301 ( .A(n_291), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_279), .B(n_275), .Y(n_302) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_280), .Y(n_303) );
INVx4_ASAP7_75t_L g304 ( .A(n_291), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_278), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_279), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_278), .Y(n_307) );
AND2x2_ASAP7_75t_SL g308 ( .A(n_296), .B(n_255), .Y(n_308) );
INVx5_ASAP7_75t_SL g309 ( .A(n_282), .Y(n_309) );
OAI33xp33_ASAP7_75t_L g310 ( .A1(n_277), .A2(n_154), .A3(n_152), .B1(n_141), .B2(n_270), .B3(n_274), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_278), .B(n_275), .Y(n_311) );
OAI31xp33_ASAP7_75t_SL g312 ( .A1(n_286), .A2(n_263), .A3(n_264), .B(n_266), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_285), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_285), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_285), .Y(n_315) );
OAI31xp33_ASAP7_75t_L g316 ( .A1(n_286), .A2(n_266), .A3(n_264), .B(n_263), .Y(n_316) );
OAI31xp33_ASAP7_75t_L g317 ( .A1(n_297), .A2(n_264), .A3(n_262), .B(n_275), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_289), .Y(n_318) );
AOI221xp5_ASAP7_75t_L g319 ( .A1(n_290), .A2(n_264), .B1(n_130), .B2(n_91), .C(n_274), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_289), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_294), .Y(n_321) );
OAI31xp33_ASAP7_75t_L g322 ( .A1(n_287), .A2(n_294), .A3(n_288), .B(n_283), .Y(n_322) );
AND2x4_ASAP7_75t_L g323 ( .A(n_295), .B(n_258), .Y(n_323) );
OA211x2_ASAP7_75t_L g324 ( .A1(n_282), .A2(n_258), .B(n_273), .C(n_255), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_283), .B(n_275), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_296), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_298), .Y(n_327) );
OAI33xp33_ASAP7_75t_L g328 ( .A1(n_292), .A2(n_149), .A3(n_151), .B1(n_4), .B2(n_5), .B3(n_6), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_318), .B(n_295), .Y(n_329) );
INVx1_ASAP7_75t_SL g330 ( .A(n_303), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_306), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_318), .B(n_295), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_305), .Y(n_333) );
OR2x2_ASAP7_75t_L g334 ( .A(n_327), .B(n_255), .Y(n_334) );
OR2x2_ASAP7_75t_L g335 ( .A(n_327), .B(n_255), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_320), .B(n_284), .Y(n_336) );
OR2x2_ASAP7_75t_L g337 ( .A(n_320), .B(n_281), .Y(n_337) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_300), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_306), .Y(n_339) );
OR2x2_ASAP7_75t_L g340 ( .A(n_321), .B(n_281), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_321), .B(n_284), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_302), .B(n_273), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_325), .B(n_2), .Y(n_343) );
INVx1_ASAP7_75t_SL g344 ( .A(n_308), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_302), .B(n_258), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_305), .Y(n_346) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_307), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_307), .B(n_281), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_313), .Y(n_349) );
INVxp67_ASAP7_75t_SL g350 ( .A(n_313), .Y(n_350) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_314), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_314), .B(n_258), .Y(n_352) );
NOR2x1p5_ASAP7_75t_L g353 ( .A(n_309), .B(n_3), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_315), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_315), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_326), .B(n_228), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_311), .B(n_281), .Y(n_357) );
INVx6_ASAP7_75t_L g358 ( .A(n_299), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_311), .Y(n_359) );
AND2x2_ASAP7_75t_SL g360 ( .A(n_312), .B(n_308), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_326), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_323), .B(n_276), .Y(n_362) );
INVx2_ASAP7_75t_SL g363 ( .A(n_299), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_316), .B(n_228), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_308), .Y(n_365) );
AOI33xp33_ASAP7_75t_L g366 ( .A1(n_301), .A2(n_149), .A3(n_151), .B1(n_5), .B2(n_8), .B3(n_9), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_299), .B(n_3), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_301), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_323), .Y(n_369) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_304), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_304), .B(n_288), .Y(n_371) );
OR2x2_ASAP7_75t_L g372 ( .A(n_304), .B(n_276), .Y(n_372) );
OAI31xp33_ASAP7_75t_SL g373 ( .A1(n_324), .A2(n_4), .A3(n_9), .B(n_10), .Y(n_373) );
OAI21x1_ASAP7_75t_SL g374 ( .A1(n_363), .A2(n_372), .B(n_368), .Y(n_374) );
OR2x2_ASAP7_75t_L g375 ( .A(n_338), .B(n_323), .Y(n_375) );
O2A1O1Ixp33_ASAP7_75t_L g376 ( .A1(n_367), .A2(n_343), .B(n_353), .C(n_330), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_331), .B(n_322), .Y(n_377) );
NOR2x1_ASAP7_75t_L g378 ( .A(n_368), .B(n_309), .Y(n_378) );
NAND2xp5_ASAP7_75t_SL g379 ( .A(n_360), .B(n_309), .Y(n_379) );
OAI21xp33_ASAP7_75t_L g380 ( .A1(n_373), .A2(n_319), .B(n_309), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_347), .B(n_317), .Y(n_381) );
OR2x2_ASAP7_75t_L g382 ( .A(n_351), .B(n_10), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_331), .Y(n_383) );
INVx1_ASAP7_75t_SL g384 ( .A(n_358), .Y(n_384) );
AND2x4_ASAP7_75t_L g385 ( .A(n_369), .B(n_11), .Y(n_385) );
AND2x4_ASAP7_75t_L g386 ( .A(n_369), .B(n_11), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_370), .B(n_12), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_359), .B(n_12), .Y(n_388) );
AND2x4_ASAP7_75t_L g389 ( .A(n_363), .B(n_13), .Y(n_389) );
NOR2xp67_ASAP7_75t_L g390 ( .A(n_372), .B(n_13), .Y(n_390) );
OR2x2_ASAP7_75t_L g391 ( .A(n_350), .B(n_14), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_339), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_339), .Y(n_393) );
INVxp33_ASAP7_75t_L g394 ( .A(n_334), .Y(n_394) );
OAI21xp5_ASAP7_75t_L g395 ( .A1(n_366), .A2(n_328), .B(n_129), .Y(n_395) );
AND2x4_ASAP7_75t_L g396 ( .A(n_365), .B(n_15), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_361), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_361), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_355), .Y(n_399) );
OR2x2_ASAP7_75t_L g400 ( .A(n_359), .B(n_276), .Y(n_400) );
NOR3xp33_ASAP7_75t_L g401 ( .A(n_364), .B(n_310), .C(n_293), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_336), .B(n_276), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_355), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_349), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_336), .B(n_129), .Y(n_405) );
INVx2_ASAP7_75t_SL g406 ( .A(n_358), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_362), .B(n_21), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_349), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_362), .B(n_26), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_354), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_341), .B(n_151), .Y(n_411) );
OR2x2_ASAP7_75t_L g412 ( .A(n_334), .B(n_335), .Y(n_412) );
OAI21xp33_ASAP7_75t_L g413 ( .A1(n_360), .A2(n_149), .B(n_140), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_329), .B(n_29), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_358), .B(n_30), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_329), .B(n_32), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_354), .Y(n_417) );
HB1xp67_ASAP7_75t_L g418 ( .A(n_358), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_332), .Y(n_419) );
OAI21xp5_ASAP7_75t_L g420 ( .A1(n_341), .A2(n_209), .B(n_195), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_332), .B(n_140), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_365), .B(n_33), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_335), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_333), .Y(n_424) );
OR2x2_ASAP7_75t_L g425 ( .A(n_345), .B(n_195), .Y(n_425) );
INVxp67_ASAP7_75t_L g426 ( .A(n_374), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_397), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_375), .B(n_344), .Y(n_428) );
NAND2x1_ASAP7_75t_L g429 ( .A(n_378), .B(n_371), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_398), .Y(n_430) );
INVxp67_ASAP7_75t_L g431 ( .A(n_418), .Y(n_431) );
AOI21xp5_ASAP7_75t_L g432 ( .A1(n_413), .A2(n_352), .B(n_371), .Y(n_432) );
OR2x2_ASAP7_75t_L g433 ( .A(n_412), .B(n_357), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_394), .B(n_357), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_419), .B(n_348), .Y(n_435) );
AOI21xp5_ASAP7_75t_L g436 ( .A1(n_413), .A2(n_342), .B(n_356), .Y(n_436) );
NOR2x1_ASAP7_75t_L g437 ( .A(n_379), .B(n_346), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g438 ( .A1(n_380), .A2(n_348), .B1(n_346), .B2(n_333), .Y(n_438) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_384), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_383), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_423), .B(n_340), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_402), .B(n_340), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_399), .B(n_337), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_403), .B(n_337), .Y(n_444) );
XOR2xp5_ASAP7_75t_L g445 ( .A(n_406), .B(n_37), .Y(n_445) );
OAI21xp33_ASAP7_75t_L g446 ( .A1(n_380), .A2(n_207), .B(n_203), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_384), .B(n_38), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_392), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_393), .Y(n_449) );
AND2x4_ASAP7_75t_L g450 ( .A(n_400), .B(n_39), .Y(n_450) );
CKINVDCx16_ASAP7_75t_R g451 ( .A(n_389), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_404), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_408), .B(n_40), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_410), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_417), .Y(n_455) );
XNOR2xp5_ASAP7_75t_L g456 ( .A(n_387), .B(n_42), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_424), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_382), .Y(n_458) );
AND2x4_ASAP7_75t_SL g459 ( .A(n_389), .B(n_207), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_377), .B(n_43), .Y(n_460) );
INVx2_ASAP7_75t_SL g461 ( .A(n_385), .Y(n_461) );
O2A1O1Ixp5_ASAP7_75t_L g462 ( .A1(n_377), .A2(n_217), .B(n_223), .C(n_191), .Y(n_462) );
NOR2xp67_ASAP7_75t_SL g463 ( .A(n_391), .B(n_207), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_401), .B(n_44), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_381), .Y(n_465) );
NOR3xp33_ASAP7_75t_L g466 ( .A(n_376), .B(n_223), .C(n_217), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_407), .B(n_45), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_409), .B(n_47), .Y(n_468) );
NAND2xp33_ASAP7_75t_SL g469 ( .A(n_385), .B(n_207), .Y(n_469) );
AOI21xp5_ASAP7_75t_L g470 ( .A1(n_390), .A2(n_204), .B(n_200), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_396), .B(n_203), .Y(n_471) );
OAI22x1_ASAP7_75t_L g472 ( .A1(n_396), .A2(n_204), .B1(n_200), .B2(n_217), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_425), .Y(n_473) );
AOI31xp33_ASAP7_75t_L g474 ( .A1(n_386), .A2(n_50), .A3(n_51), .B(n_52), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_388), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_L g476 ( .A1(n_395), .A2(n_223), .B(n_217), .C(n_173), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_386), .Y(n_477) );
AOI311xp33_ASAP7_75t_L g478 ( .A1(n_420), .A2(n_53), .A3(n_54), .B(n_56), .C(n_58), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_L g479 ( .A1(n_395), .A2(n_223), .B(n_168), .C(n_194), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_411), .Y(n_480) );
AOI221xp5_ASAP7_75t_L g481 ( .A1(n_420), .A2(n_204), .B1(n_200), .B2(n_164), .C(n_194), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_405), .B(n_61), .Y(n_482) );
INVx2_ASAP7_75t_SL g483 ( .A(n_414), .Y(n_483) );
A2O1A1Ixp33_ASAP7_75t_L g484 ( .A1(n_415), .A2(n_204), .B(n_200), .C(n_203), .Y(n_484) );
AOI222xp33_ASAP7_75t_L g485 ( .A1(n_416), .A2(n_135), .B1(n_200), .B2(n_204), .C1(n_203), .C2(n_182), .Y(n_485) );
AOI21xp33_ASAP7_75t_L g486 ( .A1(n_421), .A2(n_62), .B(n_64), .Y(n_486) );
NAND3xp33_ASAP7_75t_L g487 ( .A(n_422), .B(n_204), .C(n_200), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_380), .A2(n_204), .B1(n_200), .B2(n_135), .Y(n_488) );
XNOR2xp5_ASAP7_75t_L g489 ( .A(n_379), .B(n_65), .Y(n_489) );
INVx1_ASAP7_75t_SL g490 ( .A(n_384), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_412), .B(n_66), .Y(n_491) );
OAI221xp5_ASAP7_75t_SL g492 ( .A1(n_376), .A2(n_70), .B1(n_72), .B2(n_73), .C(n_75), .Y(n_492) );
BUFx6f_ASAP7_75t_L g493 ( .A(n_389), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_376), .B(n_135), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_377), .B(n_135), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g496 ( .A1(n_380), .A2(n_191), .B1(n_164), .B2(n_194), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_397), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_377), .B(n_182), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_465), .B(n_426), .Y(n_499) );
AOI221x1_ASAP7_75t_L g500 ( .A1(n_446), .A2(n_466), .B1(n_464), .B2(n_460), .C(n_495), .Y(n_500) );
NAND3xp33_ASAP7_75t_L g501 ( .A(n_488), .B(n_438), .C(n_496), .Y(n_501) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_451), .A2(n_461), .B1(n_477), .B2(n_458), .Y(n_502) );
AOI22xp5_ASAP7_75t_L g503 ( .A1(n_494), .A2(n_483), .B1(n_475), .B2(n_473), .Y(n_503) );
AOI211xp5_ASAP7_75t_SL g504 ( .A1(n_474), .A2(n_492), .B(n_464), .C(n_460), .Y(n_504) );
OA33x2_ASAP7_75t_L g505 ( .A1(n_442), .A2(n_441), .A3(n_498), .B1(n_443), .B2(n_444), .B3(n_453), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_439), .Y(n_506) );
O2A1O1Ixp33_ASAP7_75t_SL g507 ( .A1(n_429), .A2(n_471), .B(n_456), .C(n_489), .Y(n_507) );
NAND4xp25_ASAP7_75t_L g508 ( .A(n_478), .B(n_437), .C(n_479), .D(n_476), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_433), .Y(n_509) );
OAI21x1_ASAP7_75t_L g510 ( .A1(n_432), .A2(n_462), .B(n_436), .Y(n_510) );
OAI22xp33_ASAP7_75t_L g511 ( .A1(n_493), .A2(n_490), .B1(n_487), .B2(n_431), .Y(n_511) );
AOI211xp5_ASAP7_75t_L g512 ( .A1(n_469), .A2(n_493), .B(n_463), .C(n_484), .Y(n_512) );
AOI22xp33_ASAP7_75t_SL g513 ( .A1(n_493), .A2(n_459), .B1(n_428), .B2(n_480), .Y(n_513) );
AOI221xp5_ASAP7_75t_L g514 ( .A1(n_497), .A2(n_449), .B1(n_448), .B2(n_427), .C(n_430), .Y(n_514) );
AOI21xp33_ASAP7_75t_L g515 ( .A1(n_491), .A2(n_472), .B(n_445), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_499), .B(n_440), .Y(n_516) );
XNOR2xp5_ASAP7_75t_L g517 ( .A(n_502), .B(n_434), .Y(n_517) );
OAI22xp5_ASAP7_75t_L g518 ( .A1(n_513), .A2(n_442), .B1(n_441), .B2(n_435), .Y(n_518) );
NOR2x1_ASAP7_75t_SL g519 ( .A(n_506), .B(n_447), .Y(n_519) );
OAI211xp5_ASAP7_75t_SL g520 ( .A1(n_504), .A2(n_485), .B(n_486), .C(n_481), .Y(n_520) );
AOI221xp5_ASAP7_75t_L g521 ( .A1(n_507), .A2(n_444), .B1(n_443), .B2(n_455), .C(n_454), .Y(n_521) );
AOI22xp5_ASAP7_75t_L g522 ( .A1(n_503), .A2(n_452), .B1(n_457), .B2(n_450), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_509), .Y(n_523) );
OAI311xp33_ASAP7_75t_L g524 ( .A1(n_508), .A2(n_453), .A3(n_468), .B1(n_467), .C1(n_482), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_523), .Y(n_525) );
NAND4xp25_ASAP7_75t_L g526 ( .A(n_521), .B(n_512), .C(n_500), .D(n_515), .Y(n_526) );
AOI31xp33_ASAP7_75t_L g527 ( .A1(n_518), .A2(n_512), .A3(n_511), .B(n_501), .Y(n_527) );
NOR3xp33_ASAP7_75t_L g528 ( .A(n_520), .B(n_510), .C(n_514), .Y(n_528) );
INVxp67_ASAP7_75t_L g529 ( .A(n_517), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_525), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_528), .Y(n_531) );
OAI22xp5_ASAP7_75t_L g532 ( .A1(n_527), .A2(n_522), .B1(n_516), .B2(n_524), .Y(n_532) );
INVx3_ASAP7_75t_L g533 ( .A(n_530), .Y(n_533) );
OR3x2_ASAP7_75t_L g534 ( .A(n_531), .B(n_526), .C(n_529), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_533), .Y(n_535) );
OAI22xp5_ASAP7_75t_L g536 ( .A1(n_534), .A2(n_532), .B1(n_519), .B2(n_505), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g537 ( .A1(n_536), .A2(n_533), .B1(n_450), .B2(n_470), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_537), .Y(n_538) );
AOI221xp5_ASAP7_75t_L g539 ( .A1(n_538), .A2(n_535), .B1(n_189), .B2(n_184), .C(n_171), .Y(n_539) );
endmodule