module real_jpeg_28334_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_200;
wire n_164;
wire n_140;
wire n_126;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_216;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_0),
.A2(n_29),
.B1(n_61),
.B2(n_64),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_0),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_0),
.A2(n_30),
.B1(n_64),
.B2(n_74),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_0),
.A2(n_35),
.B1(n_41),
.B2(n_64),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_0),
.A2(n_56),
.B1(n_57),
.B2(n_64),
.Y(n_201)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_2),
.A2(n_35),
.B1(n_41),
.B2(n_42),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_2),
.A2(n_42),
.B1(n_56),
.B2(n_57),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

AOI21xp5_ASAP7_75t_L g28 ( 
.A1(n_3),
.A2(n_27),
.B(n_29),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_3),
.A2(n_25),
.B1(n_30),
.B2(n_74),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_3),
.B(n_57),
.Y(n_157)
);

A2O1A1O1Ixp25_ASAP7_75t_L g159 ( 
.A1(n_3),
.A2(n_57),
.B(n_91),
.C(n_157),
.D(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_3),
.B(n_54),
.Y(n_164)
);

OAI21xp33_ASAP7_75t_L g187 ( 
.A1(n_3),
.A2(n_34),
.B(n_170),
.Y(n_187)
);

A2O1A1O1Ixp25_ASAP7_75t_L g197 ( 
.A1(n_3),
.A2(n_53),
.B(n_61),
.C(n_66),
.D(n_198),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_3),
.B(n_61),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_4),
.A2(n_30),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_4),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_4),
.A2(n_29),
.B1(n_61),
.B2(n_73),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_4),
.A2(n_56),
.B1(n_57),
.B2(n_73),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_4),
.A2(n_35),
.B1(n_41),
.B2(n_73),
.Y(n_177)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_7),
.A2(n_56),
.B1(n_57),
.B2(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_7),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_7),
.A2(n_29),
.B1(n_61),
.B2(n_89),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_7),
.A2(n_35),
.B1(n_41),
.B2(n_89),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_8),
.A2(n_29),
.B1(n_61),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_8),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_8),
.A2(n_30),
.B1(n_68),
.B2(n_74),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g103 ( 
.A1(n_8),
.A2(n_56),
.B1(n_57),
.B2(n_68),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_8),
.A2(n_35),
.B1(n_41),
.B2(n_68),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_10),
.A2(n_35),
.B1(n_41),
.B2(n_128),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_10),
.Y(n_128)
);

O2A1O1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_11),
.A2(n_57),
.B(n_92),
.C(n_95),
.Y(n_91)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_11),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_12),
.A2(n_35),
.B1(n_41),
.B2(n_86),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_12),
.Y(n_86)
);

BUFx24_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_15),
.A2(n_35),
.B1(n_41),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_15),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_15),
.A2(n_48),
.B1(n_56),
.B2(n_57),
.Y(n_130)
);

INVx11_ASAP7_75t_SL g37 ( 
.A(n_16),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_136),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_134),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_111),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_20),
.B(n_111),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_82),
.C(n_98),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_21),
.B(n_149),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_49),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_22),
.B(n_50),
.C(n_81),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_31),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_23),
.A2(n_24),
.B1(n_31),
.B2(n_32),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

A2O1A1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_26),
.B(n_28),
.C(n_30),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_25),
.B(n_75),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_25),
.B(n_97),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_25),
.B(n_46),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_26),
.A2(n_27),
.B1(n_29),
.B2(n_61),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_26),
.A2(n_27),
.B1(n_30),
.B2(n_74),
.Y(n_79)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_29),
.A2(n_58),
.B1(n_59),
.B2(n_61),
.Y(n_60)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

AOI32xp33_ASAP7_75t_L g205 ( 
.A1(n_29),
.A2(n_57),
.A3(n_198),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_30),
.Y(n_74)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_39),
.B1(n_43),
.B2(n_47),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_33),
.A2(n_43),
.B1(n_176),
.B2(n_178),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_34),
.A2(n_46),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_34),
.A2(n_85),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_34),
.A2(n_40),
.B1(n_44),
.B2(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_34),
.A2(n_169),
.B(n_170),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_34),
.B(n_172),
.Y(n_185)
);

NAND2x1_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_38),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_35),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_35),
.A2(n_41),
.B1(n_93),
.B2(n_94),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_35),
.B(n_93),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

AOI32xp33_ASAP7_75t_L g156 ( 
.A1(n_41),
.A2(n_56),
.A3(n_94),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_41),
.B(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_44),
.A2(n_177),
.B(n_184),
.Y(n_183)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx5_ASAP7_75t_SL g126 ( 
.A(n_45),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_45),
.B(n_171),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_45),
.A2(n_185),
.B(n_204),
.Y(n_203)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_47),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_51),
.B1(n_70),
.B2(n_81),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_62),
.B(n_65),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_53),
.A2(n_54),
.B1(n_63),
.B2(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_53),
.B(n_123),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_60),
.Y(n_53)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_56),
.Y(n_57)
);

NAND2xp33_ASAP7_75t_SL g207 ( 
.A(n_56),
.B(n_58),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_57),
.B(n_93),
.Y(n_92)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_58),
.Y(n_206)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_69),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_67),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_69),
.A2(n_121),
.B(n_122),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_69),
.A2(n_110),
.B(n_122),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_70),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_75),
.B(n_77),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_72),
.A2(n_76),
.B1(n_78),
.B2(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_76),
.B(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_76),
.B(n_80),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_80),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_78),
.A2(n_105),
.B(n_106),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_82),
.B(n_98),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_87),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_83),
.B(n_87),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_90),
.B1(n_96),
.B2(n_97),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_88),
.A2(n_97),
.B(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_90),
.A2(n_96),
.B1(n_97),
.B2(n_130),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_90),
.A2(n_216),
.B(n_217),
.Y(n_215)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_91),
.B(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_91),
.A2(n_95),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_95),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_97),
.B(n_103),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_97),
.A2(n_101),
.B(n_167),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_104),
.C(n_108),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_99),
.A2(n_100),
.B1(n_108),
.B2(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_104),
.B(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_111)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_112),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_113),
.B(n_124),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_115),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_119),
.B2(n_120),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_129),
.Y(n_124)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_131),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_150),
.B(n_224),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_148),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_138),
.B(n_148),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_142),
.C(n_143),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_139),
.B(n_222),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_142),
.B(n_143),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_145),
.C(n_147),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_144),
.B(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_145),
.B(n_147),
.Y(n_212)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_146),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_219),
.B(n_223),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_209),
.B(n_218),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_193),
.B(n_208),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_173),
.B(n_192),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_161),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_155),
.B(n_161),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_159),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_160),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_168),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_165),
.B2(n_166),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_166),
.C(n_168),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_167),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_169),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_180),
.B(n_191),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_179),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_175),
.B(n_179),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_186),
.B(n_190),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_182),
.B(n_183),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_194),
.B(n_195),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_196),
.B(n_210),
.Y(n_218)
);

FAx1_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_199),
.CI(n_202),
.CON(n_196),
.SN(n_196)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_201),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_205),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_213),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_214),
.C(n_215),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_220),
.B(n_221),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);


endmodule