module fake_ibex_49_n_985 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_148, n_2, n_76, n_8, n_118, n_183, n_67, n_9, n_164, n_38, n_198, n_124, n_37, n_110, n_193, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_191, n_178, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_180, n_194, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_192, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_179, n_72, n_166, n_195, n_163, n_26, n_188, n_114, n_199, n_34, n_97, n_102, n_197, n_181, n_15, n_131, n_123, n_24, n_52, n_189, n_99, n_135, n_105, n_156, n_126, n_187, n_1, n_154, n_182, n_111, n_196, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_186, n_50, n_11, n_92, n_144, n_170, n_101, n_190, n_113, n_138, n_96, n_185, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_184, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_985);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_183;
input n_67;
input n_9;
input n_164;
input n_38;
input n_198;
input n_124;
input n_37;
input n_110;
input n_193;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_191;
input n_178;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_180;
input n_194;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_192;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_179;
input n_72;
input n_166;
input n_195;
input n_163;
input n_26;
input n_188;
input n_114;
input n_199;
input n_34;
input n_97;
input n_102;
input n_197;
input n_181;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_189;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_187;
input n_1;
input n_154;
input n_182;
input n_111;
input n_196;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_186;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_190;
input n_113;
input n_138;
input n_96;
input n_185;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_184;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_985;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_946;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_926;
wire n_328;
wire n_293;
wire n_341;
wire n_372;
wire n_418;
wire n_256;
wire n_510;
wire n_947;
wire n_845;
wire n_981;
wire n_972;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_956;
wire n_790;
wire n_920;
wire n_452;
wire n_664;
wire n_255;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_873;
wire n_962;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_957;
wire n_678;
wire n_663;
wire n_969;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_961;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_974;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_457;
wire n_412;
wire n_494;
wire n_226;
wire n_930;
wire n_336;
wire n_959;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_727;
wire n_216;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_963;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_498;
wire n_708;
wire n_317;
wire n_375;
wire n_340;
wire n_280;
wire n_698;
wire n_901;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_326;
wire n_327;
wire n_879;
wire n_723;
wire n_270;
wire n_346;
wire n_383;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_948;
wire n_859;
wire n_259;
wire n_339;
wire n_276;
wire n_470;
wire n_770;
wire n_965;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_941;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_936;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_533;
wire n_508;
wire n_939;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_928;
wire n_967;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_982;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_929;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_977;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_923;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_933;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_938;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_720;
wire n_710;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_944;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_524;
wire n_349;
wire n_765;
wire n_857;
wire n_849;
wire n_980;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_917;
wire n_388;
wire n_953;
wire n_625;
wire n_968;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_931;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_858;
wire n_207;
wire n_922;
wire n_438;
wire n_851;
wire n_689;
wire n_960;
wire n_793;
wire n_676;
wire n_937;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_973;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_514;
wire n_488;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_635;
wire n_979;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_966;
wire n_359;
wire n_826;
wire n_299;
wire n_433;
wire n_262;
wire n_439;
wire n_704;
wire n_949;
wire n_924;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_796;
wire n_837;
wire n_797;
wire n_477;
wire n_640;
wire n_954;
wire n_363;
wire n_402;
wire n_725;
wire n_369;
wire n_976;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_935;
wire n_869;
wire n_925;
wire n_718;
wire n_918;
wire n_801;
wire n_672;
wire n_722;
wire n_401;
wire n_554;
wire n_553;
wire n_735;
wire n_305;
wire n_882;
wire n_942;
wire n_713;
wire n_307;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_392;
wire n_206;
wire n_354;
wire n_630;
wire n_567;
wire n_516;
wire n_548;
wire n_943;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_940;
wire n_200;
wire n_506;
wire n_444;
wire n_564;
wire n_562;
wire n_868;
wire n_546;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_975;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_520;
wire n_411;
wire n_784;
wire n_684;
wire n_775;
wire n_934;
wire n_927;
wire n_658;
wire n_512;
wire n_615;
wire n_950;
wire n_685;
wire n_397;
wire n_366;
wire n_283;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_971;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_978;
wire n_818;
wire n_653;
wire n_238;
wire n_214;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_951;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_919;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_320;
wire n_288;
wire n_247;
wire n_379;
wire n_285;
wire n_551;
wire n_612;
wire n_291;
wire n_318;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_955;
wire n_342;
wire n_233;
wire n_385;
wire n_414;
wire n_430;
wire n_741;
wire n_729;
wire n_603;
wire n_378;
wire n_486;
wire n_952;
wire n_422;
wire n_264;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_820;
wire n_670;
wire n_805;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_958;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_250;
wire n_945;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_528;
wire n_683;
wire n_631;
wire n_260;
wire n_620;
wire n_836;
wire n_794;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_970;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_396;
wire n_252;
wire n_697;
wire n_816;
wire n_874;
wire n_912;
wire n_921;
wire n_890;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_964;
wire n_424;
wire n_565;
wire n_916;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_984;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_202;
wire n_298;
wire n_231;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_932;
wire n_657;
wire n_764;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_54),
.Y(n_200)
);

INVxp33_ASAP7_75t_SL g201 ( 
.A(n_117),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_143),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_137),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_11),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_83),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_139),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_96),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_138),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_73),
.Y(n_209)
);

BUFx10_ASAP7_75t_L g210 ( 
.A(n_184),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_155),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_75),
.Y(n_212)
);

BUFx10_ASAP7_75t_L g213 ( 
.A(n_44),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_120),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_32),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_111),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_51),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_156),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_148),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_114),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_21),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_50),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_72),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_141),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_39),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_169),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_60),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_88),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_22),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_79),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_174),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_146),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_159),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_158),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_86),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_8),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_61),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_194),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_53),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_66),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_102),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_109),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_196),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_112),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_90),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_95),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_176),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_166),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_147),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_173),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_6),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_182),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_16),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_31),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_19),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_52),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_24),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_149),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_185),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_142),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_36),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_108),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_177),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_127),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_9),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_18),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_190),
.Y(n_267)
);

INVxp67_ASAP7_75t_SL g268 ( 
.A(n_67),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_57),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_2),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_94),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_38),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_100),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_32),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_84),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_104),
.Y(n_276)
);

BUFx10_ASAP7_75t_L g277 ( 
.A(n_136),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_46),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_107),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_40),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_164),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_195),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_154),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_188),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_165),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_150),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_33),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_179),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_99),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_129),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_24),
.Y(n_291)
);

BUFx8_ASAP7_75t_SL g292 ( 
.A(n_199),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_37),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_140),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_93),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_186),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_192),
.Y(n_297)
);

NOR2xp67_ASAP7_75t_L g298 ( 
.A(n_26),
.B(n_175),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_41),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_13),
.Y(n_300)
);

BUFx10_ASAP7_75t_L g301 ( 
.A(n_193),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_11),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_25),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_78),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_29),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_82),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_76),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_87),
.Y(n_308)
);

BUFx5_ASAP7_75t_L g309 ( 
.A(n_92),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_55),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_122),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_70),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_45),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_116),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_144),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_119),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_20),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_68),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_153),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_35),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_74),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_64),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_20),
.Y(n_323)
);

NOR2xp67_ASAP7_75t_L g324 ( 
.A(n_8),
.B(n_0),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_98),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_1),
.Y(n_326)
);

INVx4_ASAP7_75t_L g327 ( 
.A(n_310),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_211),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_241),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_300),
.B(n_0),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_309),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_309),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_302),
.Y(n_333)
);

INVx5_ASAP7_75t_L g334 ( 
.A(n_211),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_241),
.B(n_1),
.Y(n_335)
);

AND2x4_ASAP7_75t_L g336 ( 
.A(n_266),
.B(n_2),
.Y(n_336)
);

OAI22x1_ASAP7_75t_SL g337 ( 
.A1(n_274),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_292),
.Y(n_338)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_266),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_211),
.Y(n_340)
);

AND2x4_ASAP7_75t_L g341 ( 
.A(n_302),
.B(n_234),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_309),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_221),
.Y(n_343)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_210),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_309),
.Y(n_345)
);

AND2x6_ASAP7_75t_L g346 ( 
.A(n_269),
.B(n_299),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_211),
.Y(n_347)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_210),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_236),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_320),
.B(n_3),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_238),
.B(n_4),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_274),
.A2(n_326),
.B1(n_270),
.B2(n_291),
.Y(n_352)
);

AND2x4_ASAP7_75t_L g353 ( 
.A(n_269),
.B(n_5),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_238),
.B(n_6),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_309),
.B(n_7),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_251),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_303),
.B(n_7),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_309),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_326),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_308),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_255),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_265),
.B(n_10),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_203),
.B(n_205),
.Y(n_363)
);

AND2x4_ASAP7_75t_L g364 ( 
.A(n_299),
.B(n_12),
.Y(n_364)
);

BUFx8_ASAP7_75t_SL g365 ( 
.A(n_292),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_287),
.Y(n_366)
);

INVx3_ASAP7_75t_L g367 ( 
.A(n_213),
.Y(n_367)
);

OA21x2_ASAP7_75t_L g368 ( 
.A1(n_242),
.A2(n_306),
.B(n_284),
.Y(n_368)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_213),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_206),
.B(n_13),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_242),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_247),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_284),
.Y(n_373)
);

AND2x4_ASAP7_75t_L g374 ( 
.A(n_318),
.B(n_14),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_308),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_308),
.Y(n_376)
);

INVx5_ASAP7_75t_L g377 ( 
.A(n_311),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_306),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_264),
.Y(n_379)
);

AND2x4_ASAP7_75t_L g380 ( 
.A(n_318),
.B(n_15),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_325),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_311),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_325),
.Y(n_383)
);

INVx6_ASAP7_75t_L g384 ( 
.A(n_277),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_277),
.B(n_17),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_204),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_311),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_305),
.A2(n_18),
.B1(n_19),
.B2(n_21),
.Y(n_388)
);

OAI21x1_ASAP7_75t_L g389 ( 
.A1(n_208),
.A2(n_115),
.B(n_197),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_209),
.Y(n_390)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_311),
.Y(n_391)
);

AND2x4_ASAP7_75t_L g392 ( 
.A(n_317),
.B(n_22),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_323),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_212),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_301),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_214),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_301),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_216),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_222),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_225),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_226),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_227),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_331),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_336),
.Y(n_404)
);

OAI22xp33_ASAP7_75t_L g405 ( 
.A1(n_333),
.A2(n_253),
.B1(n_215),
.B2(n_229),
.Y(n_405)
);

INVx8_ASAP7_75t_L g406 ( 
.A(n_341),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_331),
.Y(n_407)
);

INVx4_ASAP7_75t_L g408 ( 
.A(n_353),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_327),
.B(n_249),
.Y(n_409)
);

BUFx10_ASAP7_75t_L g410 ( 
.A(n_384),
.Y(n_410)
);

NOR2x1p5_ASAP7_75t_L g411 ( 
.A(n_338),
.B(n_254),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_346),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_332),
.Y(n_413)
);

BUFx2_ASAP7_75t_L g414 ( 
.A(n_333),
.Y(n_414)
);

AOI22xp33_ASAP7_75t_L g415 ( 
.A1(n_392),
.A2(n_201),
.B1(n_322),
.B2(n_297),
.Y(n_415)
);

BUFx2_ASAP7_75t_L g416 ( 
.A(n_386),
.Y(n_416)
);

CKINVDCx6p67_ASAP7_75t_R g417 ( 
.A(n_351),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_332),
.Y(n_418)
);

INVx2_ASAP7_75t_SL g419 ( 
.A(n_384),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_342),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_342),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_327),
.B(n_257),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_327),
.B(n_261),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_392),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_353),
.B(n_233),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_345),
.Y(n_426)
);

INVx2_ASAP7_75t_SL g427 ( 
.A(n_384),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_345),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_329),
.B(n_272),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_339),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_353),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_358),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_341),
.B(n_293),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_358),
.Y(n_434)
);

OR2x2_ASAP7_75t_L g435 ( 
.A(n_349),
.B(n_324),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_341),
.B(n_200),
.Y(n_436)
);

INVx2_ASAP7_75t_SL g437 ( 
.A(n_384),
.Y(n_437)
);

AOI22xp33_ASAP7_75t_SL g438 ( 
.A1(n_359),
.A2(n_264),
.B1(n_288),
.B2(n_240),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_368),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_364),
.Y(n_440)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_351),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_368),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_365),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_364),
.B(n_237),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_364),
.Y(n_445)
);

BUFx4f_ASAP7_75t_L g446 ( 
.A(n_374),
.Y(n_446)
);

INVx4_ASAP7_75t_L g447 ( 
.A(n_374),
.Y(n_447)
);

AOI22xp33_ASAP7_75t_L g448 ( 
.A1(n_368),
.A2(n_267),
.B1(n_271),
.B2(n_273),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_340),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_340),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_344),
.B(n_243),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_374),
.Y(n_452)
);

INVx1_ASAP7_75t_SL g453 ( 
.A(n_338),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_381),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_380),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_380),
.Y(n_456)
);

INVx8_ASAP7_75t_L g457 ( 
.A(n_346),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_380),
.Y(n_458)
);

BUFx6f_ASAP7_75t_SL g459 ( 
.A(n_395),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_401),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_344),
.B(n_202),
.Y(n_461)
);

AND2x6_ASAP7_75t_L g462 ( 
.A(n_354),
.B(n_245),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_360),
.Y(n_463)
);

AOI21x1_ASAP7_75t_L g464 ( 
.A1(n_389),
.A2(n_259),
.B(n_246),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_360),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_365),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_360),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_360),
.Y(n_468)
);

INVx5_ASAP7_75t_L g469 ( 
.A(n_346),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_354),
.A2(n_288),
.B1(n_239),
.B2(n_258),
.Y(n_470)
);

OAI21xp33_ASAP7_75t_SL g471 ( 
.A1(n_363),
.A2(n_298),
.B(n_278),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_375),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_371),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_375),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_348),
.B(n_217),
.Y(n_475)
);

BUFx10_ASAP7_75t_L g476 ( 
.A(n_397),
.Y(n_476)
);

OR2x6_ASAP7_75t_L g477 ( 
.A(n_372),
.B(n_276),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_346),
.Y(n_478)
);

INVx2_ASAP7_75t_SL g479 ( 
.A(n_348),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_371),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_373),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_379),
.Y(n_482)
);

OAI22xp33_ASAP7_75t_L g483 ( 
.A1(n_388),
.A2(n_350),
.B1(n_330),
.B2(n_335),
.Y(n_483)
);

AOI22xp33_ASAP7_75t_SL g484 ( 
.A1(n_385),
.A2(n_268),
.B1(n_282),
.B2(n_296),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_375),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_375),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_373),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_378),
.Y(n_488)
);

NAND2xp33_ASAP7_75t_L g489 ( 
.A(n_346),
.B(n_218),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_376),
.Y(n_490)
);

CKINVDCx14_ASAP7_75t_R g491 ( 
.A(n_379),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g492 ( 
.A(n_399),
.B(n_279),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_367),
.B(n_219),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_376),
.Y(n_494)
);

BUFx10_ASAP7_75t_L g495 ( 
.A(n_398),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_367),
.B(n_281),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_399),
.Y(n_497)
);

INVx2_ASAP7_75t_SL g498 ( 
.A(n_367),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_376),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_376),
.Y(n_500)
);

NAND2xp33_ASAP7_75t_R g501 ( 
.A(n_385),
.B(n_220),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_399),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_390),
.B(n_286),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_352),
.Y(n_504)
);

BUFx10_ASAP7_75t_L g505 ( 
.A(n_370),
.Y(n_505)
);

INVx4_ASAP7_75t_L g506 ( 
.A(n_369),
.Y(n_506)
);

INVx6_ASAP7_75t_L g507 ( 
.A(n_334),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_382),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_369),
.Y(n_509)
);

CKINVDCx6p67_ASAP7_75t_R g510 ( 
.A(n_357),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_381),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_343),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_390),
.B(n_289),
.Y(n_513)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_383),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_382),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_382),
.Y(n_516)
);

NOR3xp33_ASAP7_75t_L g517 ( 
.A(n_405),
.B(n_362),
.C(n_355),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_495),
.B(n_394),
.Y(n_518)
);

BUFx6f_ASAP7_75t_SL g519 ( 
.A(n_476),
.Y(n_519)
);

INVx8_ASAP7_75t_L g520 ( 
.A(n_406),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_484),
.A2(n_355),
.B1(n_366),
.B2(n_393),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_484),
.A2(n_356),
.B1(n_361),
.B2(n_396),
.Y(n_522)
);

INVx8_ASAP7_75t_L g523 ( 
.A(n_406),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_433),
.B(n_394),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_436),
.B(n_396),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_L g526 ( 
.A1(n_415),
.A2(n_402),
.B1(n_400),
.B2(n_383),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_406),
.A2(n_337),
.B1(n_304),
.B2(n_312),
.Y(n_527)
);

AOI22xp33_ASAP7_75t_L g528 ( 
.A1(n_462),
.A2(n_294),
.B1(n_313),
.B2(n_316),
.Y(n_528)
);

INVx2_ASAP7_75t_SL g529 ( 
.A(n_410),
.Y(n_529)
);

INVx4_ASAP7_75t_L g530 ( 
.A(n_457),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_446),
.B(n_223),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_414),
.B(n_207),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_424),
.B(n_228),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_506),
.B(n_230),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_511),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_416),
.B(n_224),
.Y(n_536)
);

NOR2xp67_ASAP7_75t_SL g537 ( 
.A(n_469),
.B(n_231),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_454),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_514),
.Y(n_539)
);

NAND2xp33_ASAP7_75t_L g540 ( 
.A(n_457),
.B(n_232),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_409),
.B(n_235),
.Y(n_541)
);

O2A1O1Ixp5_ASAP7_75t_L g542 ( 
.A1(n_425),
.A2(n_389),
.B(n_283),
.C(n_280),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_409),
.B(n_244),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_441),
.B(n_248),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_441),
.B(n_250),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_462),
.A2(n_295),
.B1(n_256),
.B2(n_260),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_512),
.B(n_262),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_475),
.B(n_263),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_417),
.B(n_252),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_491),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_L g551 ( 
.A1(n_483),
.A2(n_307),
.B1(n_314),
.B2(n_319),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_460),
.Y(n_552)
);

AND2x4_ASAP7_75t_SL g553 ( 
.A(n_410),
.B(n_328),
.Y(n_553)
);

NOR3xp33_ASAP7_75t_L g554 ( 
.A(n_405),
.B(n_275),
.C(n_285),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_422),
.B(n_290),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_423),
.B(n_315),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_SL g557 ( 
.A(n_469),
.B(n_408),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_462),
.A2(n_321),
.B1(n_377),
.B2(n_334),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g559 ( 
.A1(n_483),
.A2(n_377),
.B1(n_334),
.B2(n_391),
.Y(n_559)
);

NOR2xp67_ASAP7_75t_L g560 ( 
.A(n_443),
.B(n_23),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_510),
.B(n_23),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_430),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_473),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_404),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_509),
.B(n_334),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_451),
.B(n_334),
.Y(n_566)
);

BUFx8_ASAP7_75t_L g567 ( 
.A(n_459),
.Y(n_567)
);

BUFx5_ASAP7_75t_L g568 ( 
.A(n_412),
.Y(n_568)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_462),
.A2(n_377),
.B1(n_387),
.B2(n_391),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_480),
.Y(n_570)
);

NOR2xp67_ASAP7_75t_L g571 ( 
.A(n_429),
.B(n_25),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_451),
.B(n_377),
.Y(n_572)
);

AND2x6_ASAP7_75t_SL g573 ( 
.A(n_477),
.B(n_466),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_481),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_496),
.B(n_377),
.Y(n_575)
);

OR2x6_ASAP7_75t_L g576 ( 
.A(n_477),
.B(n_391),
.Y(n_576)
);

A2O1A1Ixp33_ASAP7_75t_L g577 ( 
.A1(n_431),
.A2(n_391),
.B(n_387),
.C(n_347),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_496),
.B(n_328),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_487),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_462),
.B(n_328),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_488),
.Y(n_581)
);

OR2x2_ASAP7_75t_L g582 ( 
.A(n_453),
.B(n_27),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_SL g583 ( 
.A1(n_504),
.A2(n_491),
.B1(n_482),
.B2(n_438),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_479),
.B(n_42),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_498),
.B(n_43),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_440),
.Y(n_586)
);

INVxp67_ASAP7_75t_L g587 ( 
.A(n_501),
.Y(n_587)
);

OAI21xp5_ASAP7_75t_L g588 ( 
.A1(n_439),
.A2(n_391),
.B(n_387),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_445),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_445),
.Y(n_590)
);

A2O1A1Ixp33_ASAP7_75t_L g591 ( 
.A1(n_452),
.A2(n_387),
.B(n_347),
.C(n_328),
.Y(n_591)
);

OAI22xp5_ASAP7_75t_L g592 ( 
.A1(n_438),
.A2(n_470),
.B1(n_477),
.B2(n_458),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_455),
.B(n_347),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_456),
.B(n_387),
.Y(n_594)
);

A2O1A1Ixp33_ASAP7_75t_L g595 ( 
.A1(n_442),
.A2(n_28),
.B(n_30),
.C(n_31),
.Y(n_595)
);

AO221x1_ASAP7_75t_L g596 ( 
.A1(n_501),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.C(n_37),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_419),
.B(n_47),
.Y(n_597)
);

AOI22xp33_ASAP7_75t_L g598 ( 
.A1(n_448),
.A2(n_34),
.B1(n_38),
.B2(n_48),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_408),
.B(n_49),
.Y(n_599)
);

O2A1O1Ixp5_ASAP7_75t_L g600 ( 
.A1(n_425),
.A2(n_56),
.B(n_58),
.C(n_59),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_427),
.B(n_437),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_497),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_447),
.B(n_62),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_447),
.Y(n_604)
);

OAI22xp33_ASAP7_75t_L g605 ( 
.A1(n_435),
.A2(n_444),
.B1(n_461),
.B2(n_493),
.Y(n_605)
);

NOR2xp67_ASAP7_75t_L g606 ( 
.A(n_471),
.B(n_63),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_448),
.A2(n_65),
.B1(n_69),
.B2(n_71),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_442),
.Y(n_608)
);

BUFx3_ASAP7_75t_L g609 ( 
.A(n_513),
.Y(n_609)
);

AOI22xp33_ASAP7_75t_L g610 ( 
.A1(n_513),
.A2(n_77),
.B1(n_80),
.B2(n_81),
.Y(n_610)
);

O2A1O1Ixp5_ASAP7_75t_L g611 ( 
.A1(n_464),
.A2(n_198),
.B(n_85),
.C(n_89),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_520),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_536),
.B(n_505),
.Y(n_613)
);

INVxp67_ASAP7_75t_L g614 ( 
.A(n_519),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_532),
.B(n_505),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_604),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_518),
.Y(n_617)
);

INVx1_ASAP7_75t_SL g618 ( 
.A(n_520),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_518),
.B(n_503),
.Y(n_619)
);

AOI21xp5_ASAP7_75t_L g620 ( 
.A1(n_608),
.A2(n_489),
.B(n_478),
.Y(n_620)
);

AO22x1_ASAP7_75t_L g621 ( 
.A1(n_567),
.A2(n_411),
.B1(n_434),
.B2(n_432),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g622 ( 
.A1(n_588),
.A2(n_492),
.B(n_407),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_L g623 ( 
.A1(n_588),
.A2(n_403),
.B(n_413),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_561),
.B(n_403),
.Y(n_624)
);

CKINVDCx10_ASAP7_75t_R g625 ( 
.A(n_519),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g626 ( 
.A(n_549),
.B(n_413),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_524),
.B(n_418),
.Y(n_627)
);

NOR2xp67_ASAP7_75t_L g628 ( 
.A(n_550),
.B(n_91),
.Y(n_628)
);

OR2x6_ASAP7_75t_L g629 ( 
.A(n_523),
.B(n_420),
.Y(n_629)
);

NAND3xp33_ASAP7_75t_L g630 ( 
.A(n_554),
.B(n_420),
.C(n_421),
.Y(n_630)
);

BUFx8_ASAP7_75t_L g631 ( 
.A(n_582),
.Y(n_631)
);

AOI21xp5_ASAP7_75t_L g632 ( 
.A1(n_566),
.A2(n_421),
.B(n_426),
.Y(n_632)
);

AO21x1_ASAP7_75t_L g633 ( 
.A1(n_559),
.A2(n_578),
.B(n_526),
.Y(n_633)
);

AOI21xp5_ASAP7_75t_L g634 ( 
.A1(n_572),
.A2(n_428),
.B(n_432),
.Y(n_634)
);

A2O1A1Ixp33_ASAP7_75t_L g635 ( 
.A1(n_525),
.A2(n_434),
.B(n_502),
.C(n_516),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_605),
.B(n_507),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_564),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_517),
.B(n_507),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_587),
.B(n_544),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_586),
.Y(n_640)
);

O2A1O1Ixp33_ASAP7_75t_L g641 ( 
.A1(n_551),
.A2(n_515),
.B(n_508),
.C(n_500),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_604),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_SL g643 ( 
.A(n_530),
.B(n_449),
.Y(n_643)
);

CKINVDCx16_ASAP7_75t_R g644 ( 
.A(n_592),
.Y(n_644)
);

A2O1A1Ixp33_ASAP7_75t_L g645 ( 
.A1(n_521),
.A2(n_500),
.B(n_499),
.C(n_494),
.Y(n_645)
);

INVx2_ASAP7_75t_SL g646 ( 
.A(n_567),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_545),
.B(n_97),
.Y(n_647)
);

AOI21xp5_ASAP7_75t_L g648 ( 
.A1(n_575),
.A2(n_533),
.B(n_547),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_535),
.B(n_539),
.Y(n_649)
);

NOR3xp33_ASAP7_75t_L g650 ( 
.A(n_592),
.B(n_490),
.C(n_486),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_SL g651 ( 
.A(n_530),
.B(n_449),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_609),
.B(n_101),
.Y(n_652)
);

A2O1A1Ixp33_ASAP7_75t_L g653 ( 
.A1(n_522),
.A2(n_485),
.B(n_474),
.C(n_472),
.Y(n_653)
);

INVx2_ASAP7_75t_SL g654 ( 
.A(n_529),
.Y(n_654)
);

AOI21x1_ASAP7_75t_L g655 ( 
.A1(n_599),
.A2(n_468),
.B(n_467),
.Y(n_655)
);

AOI22xp33_ASAP7_75t_L g656 ( 
.A1(n_596),
.A2(n_465),
.B1(n_463),
.B2(n_450),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_583),
.B(n_103),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_548),
.B(n_105),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_576),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_528),
.B(n_106),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_541),
.B(n_110),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_562),
.Y(n_662)
);

AOI21xp5_ASAP7_75t_L g663 ( 
.A1(n_593),
.A2(n_113),
.B(n_118),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_551),
.B(n_563),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_534),
.B(n_121),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_546),
.B(n_123),
.Y(n_666)
);

OAI22xp5_ASAP7_75t_L g667 ( 
.A1(n_576),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_555),
.B(n_128),
.Y(n_668)
);

AO22x1_ASAP7_75t_L g669 ( 
.A1(n_573),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_669)
);

BUFx2_ASAP7_75t_L g670 ( 
.A(n_570),
.Y(n_670)
);

OAI21xp5_ASAP7_75t_L g671 ( 
.A1(n_611),
.A2(n_606),
.B(n_526),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g672 ( 
.A1(n_594),
.A2(n_133),
.B(n_134),
.Y(n_672)
);

AOI21xp5_ASAP7_75t_L g673 ( 
.A1(n_594),
.A2(n_135),
.B(n_145),
.Y(n_673)
);

OAI21xp5_ASAP7_75t_L g674 ( 
.A1(n_600),
.A2(n_151),
.B(n_152),
.Y(n_674)
);

A2O1A1Ixp33_ASAP7_75t_L g675 ( 
.A1(n_589),
.A2(n_157),
.B(n_160),
.C(n_161),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g676 ( 
.A1(n_557),
.A2(n_162),
.B(n_163),
.Y(n_676)
);

CKINVDCx10_ASAP7_75t_R g677 ( 
.A(n_527),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_574),
.B(n_579),
.Y(n_678)
);

BUFx2_ASAP7_75t_L g679 ( 
.A(n_581),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_590),
.Y(n_680)
);

OAI21xp5_ASAP7_75t_L g681 ( 
.A1(n_599),
.A2(n_167),
.B(n_168),
.Y(n_681)
);

NOR3xp33_ASAP7_75t_L g682 ( 
.A(n_543),
.B(n_170),
.C(n_171),
.Y(n_682)
);

OAI22xp5_ASAP7_75t_L g683 ( 
.A1(n_598),
.A2(n_172),
.B1(n_178),
.B2(n_180),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_556),
.B(n_181),
.Y(n_684)
);

OAI21xp5_ASAP7_75t_L g685 ( 
.A1(n_603),
.A2(n_607),
.B(n_580),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_538),
.Y(n_686)
);

A2O1A1Ixp33_ASAP7_75t_L g687 ( 
.A1(n_571),
.A2(n_183),
.B(n_187),
.C(n_189),
.Y(n_687)
);

AND2x6_ASAP7_75t_SL g688 ( 
.A(n_601),
.B(n_191),
.Y(n_688)
);

AOI21xp5_ASAP7_75t_L g689 ( 
.A1(n_603),
.A2(n_565),
.B(n_531),
.Y(n_689)
);

INVx1_ASAP7_75t_SL g690 ( 
.A(n_553),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_558),
.B(n_540),
.Y(n_691)
);

O2A1O1Ixp33_ASAP7_75t_L g692 ( 
.A1(n_595),
.A2(n_591),
.B(n_577),
.C(n_585),
.Y(n_692)
);

BUFx6f_ASAP7_75t_L g693 ( 
.A(n_612),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_612),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_617),
.B(n_584),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_613),
.B(n_560),
.Y(n_696)
);

A2O1A1Ixp33_ASAP7_75t_L g697 ( 
.A1(n_648),
.A2(n_597),
.B(n_569),
.C(n_610),
.Y(n_697)
);

AOI21xp5_ASAP7_75t_L g698 ( 
.A1(n_623),
.A2(n_622),
.B(n_671),
.Y(n_698)
);

AO31x2_ASAP7_75t_L g699 ( 
.A1(n_633),
.A2(n_602),
.A3(n_552),
.B(n_568),
.Y(n_699)
);

AOI21xp5_ASAP7_75t_L g700 ( 
.A1(n_685),
.A2(n_568),
.B(n_537),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_649),
.Y(n_701)
);

AO31x2_ASAP7_75t_L g702 ( 
.A1(n_653),
.A2(n_568),
.A3(n_645),
.B(n_635),
.Y(n_702)
);

AOI21xp33_ASAP7_75t_L g703 ( 
.A1(n_615),
.A2(n_568),
.B(n_691),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_670),
.B(n_679),
.Y(n_704)
);

NOR4xp25_ASAP7_75t_L g705 ( 
.A(n_664),
.B(n_641),
.C(n_656),
.D(n_657),
.Y(n_705)
);

OAI21xp5_ASAP7_75t_L g706 ( 
.A1(n_638),
.A2(n_630),
.B(n_619),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_626),
.B(n_644),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_618),
.B(n_624),
.Y(n_708)
);

NOR2xp67_ASAP7_75t_L g709 ( 
.A(n_646),
.B(n_614),
.Y(n_709)
);

BUFx6f_ASAP7_75t_L g710 ( 
.A(n_629),
.Y(n_710)
);

AO31x2_ASAP7_75t_L g711 ( 
.A1(n_683),
.A2(n_675),
.A3(n_687),
.B(n_667),
.Y(n_711)
);

NOR2xp67_ASAP7_75t_L g712 ( 
.A(n_654),
.B(n_625),
.Y(n_712)
);

AOI21xp5_ASAP7_75t_L g713 ( 
.A1(n_685),
.A2(n_620),
.B(n_634),
.Y(n_713)
);

AND2x6_ASAP7_75t_L g714 ( 
.A(n_659),
.B(n_652),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_SL g715 ( 
.A1(n_629),
.A2(n_659),
.B(n_681),
.Y(n_715)
);

OR2x2_ASAP7_75t_SL g716 ( 
.A(n_677),
.B(n_688),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_SL g717 ( 
.A(n_659),
.B(n_690),
.Y(n_717)
);

OAI22xp33_ASAP7_75t_L g718 ( 
.A1(n_627),
.A2(n_678),
.B1(n_662),
.B2(n_637),
.Y(n_718)
);

O2A1O1Ixp5_ASAP7_75t_L g719 ( 
.A1(n_668),
.A2(n_684),
.B(n_665),
.C(n_666),
.Y(n_719)
);

BUFx3_ASAP7_75t_L g720 ( 
.A(n_631),
.Y(n_720)
);

INVx3_ASAP7_75t_L g721 ( 
.A(n_631),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_639),
.B(n_640),
.Y(n_722)
);

A2O1A1Ixp33_ASAP7_75t_L g723 ( 
.A1(n_658),
.A2(n_647),
.B(n_661),
.C(n_636),
.Y(n_723)
);

OAI21xp5_ASAP7_75t_L g724 ( 
.A1(n_692),
.A2(n_632),
.B(n_689),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_616),
.Y(n_725)
);

BUFx3_ASAP7_75t_L g726 ( 
.A(n_686),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_680),
.B(n_621),
.Y(n_727)
);

AOI221x1_ASAP7_75t_L g728 ( 
.A1(n_663),
.A2(n_673),
.B1(n_672),
.B2(n_676),
.C(n_660),
.Y(n_728)
);

AND2x4_ASAP7_75t_L g729 ( 
.A(n_628),
.B(n_642),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_669),
.Y(n_730)
);

OAI21x1_ASAP7_75t_L g731 ( 
.A1(n_643),
.A2(n_651),
.B(n_655),
.Y(n_731)
);

AO32x2_ASAP7_75t_L g732 ( 
.A1(n_667),
.A2(n_559),
.A3(n_526),
.B1(n_551),
.B2(n_592),
.Y(n_732)
);

AOI21xp5_ASAP7_75t_L g733 ( 
.A1(n_648),
.A2(n_623),
.B(n_446),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_649),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_649),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_649),
.Y(n_736)
);

BUFx2_ASAP7_75t_L g737 ( 
.A(n_612),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_649),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_617),
.B(n_649),
.Y(n_739)
);

AOI21xp5_ASAP7_75t_L g740 ( 
.A1(n_648),
.A2(n_623),
.B(n_446),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_L g741 ( 
.A1(n_644),
.A2(n_592),
.B1(n_554),
.B2(n_617),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_617),
.B(n_649),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_612),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_617),
.B(n_649),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_617),
.B(n_649),
.Y(n_745)
);

AOI221x1_ASAP7_75t_L g746 ( 
.A1(n_671),
.A2(n_650),
.B1(n_674),
.B2(n_682),
.C(n_681),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_SL g747 ( 
.A(n_618),
.B(n_519),
.Y(n_747)
);

NAND2x1_ASAP7_75t_L g748 ( 
.A(n_629),
.B(n_612),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_617),
.B(n_649),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_617),
.B(n_649),
.Y(n_750)
);

INVx2_ASAP7_75t_SL g751 ( 
.A(n_612),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_617),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_649),
.Y(n_753)
);

INVx3_ASAP7_75t_L g754 ( 
.A(n_612),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_617),
.B(n_649),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_617),
.B(n_649),
.Y(n_756)
);

OA21x2_ASAP7_75t_L g757 ( 
.A1(n_671),
.A2(n_674),
.B(n_633),
.Y(n_757)
);

OAI21xp5_ASAP7_75t_L g758 ( 
.A1(n_648),
.A2(n_623),
.B(n_542),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_613),
.B(n_615),
.Y(n_759)
);

AOI21xp5_ASAP7_75t_L g760 ( 
.A1(n_648),
.A2(n_623),
.B(n_446),
.Y(n_760)
);

AOI21xp5_ASAP7_75t_L g761 ( 
.A1(n_648),
.A2(n_623),
.B(n_446),
.Y(n_761)
);

AOI21xp5_ASAP7_75t_L g762 ( 
.A1(n_648),
.A2(n_623),
.B(n_446),
.Y(n_762)
);

AOI21xp5_ASAP7_75t_L g763 ( 
.A1(n_648),
.A2(n_623),
.B(n_446),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_617),
.B(n_649),
.Y(n_764)
);

A2O1A1Ixp33_ASAP7_75t_L g765 ( 
.A1(n_648),
.A2(n_639),
.B(n_617),
.C(n_658),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_649),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_648),
.A2(n_623),
.B(n_446),
.Y(n_767)
);

NAND3xp33_ASAP7_75t_L g768 ( 
.A(n_671),
.B(n_656),
.C(n_471),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_617),
.B(n_649),
.Y(n_769)
);

INVx5_ASAP7_75t_L g770 ( 
.A(n_612),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_648),
.A2(n_623),
.B(n_446),
.Y(n_771)
);

INVxp67_ASAP7_75t_L g772 ( 
.A(n_617),
.Y(n_772)
);

HB1xp67_ASAP7_75t_L g773 ( 
.A(n_612),
.Y(n_773)
);

AO32x2_ASAP7_75t_L g774 ( 
.A1(n_667),
.A2(n_559),
.A3(n_526),
.B1(n_551),
.B2(n_592),
.Y(n_774)
);

BUFx6f_ASAP7_75t_L g775 ( 
.A(n_612),
.Y(n_775)
);

BUFx6f_ASAP7_75t_L g776 ( 
.A(n_612),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_648),
.A2(n_623),
.B(n_446),
.Y(n_777)
);

AO31x2_ASAP7_75t_L g778 ( 
.A1(n_633),
.A2(n_653),
.A3(n_645),
.B(n_559),
.Y(n_778)
);

NOR2xp67_ASAP7_75t_SL g779 ( 
.A(n_770),
.B(n_720),
.Y(n_779)
);

AND2x4_ASAP7_75t_L g780 ( 
.A(n_701),
.B(n_734),
.Y(n_780)
);

AND2x4_ASAP7_75t_L g781 ( 
.A(n_735),
.B(n_736),
.Y(n_781)
);

INVx3_ASAP7_75t_SL g782 ( 
.A(n_770),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_738),
.Y(n_783)
);

HB1xp67_ASAP7_75t_L g784 ( 
.A(n_752),
.Y(n_784)
);

OAI21xp5_ASAP7_75t_L g785 ( 
.A1(n_768),
.A2(n_765),
.B(n_706),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_718),
.A2(n_761),
.B(n_760),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_753),
.B(n_766),
.Y(n_787)
);

OAI21xp5_ASAP7_75t_L g788 ( 
.A1(n_724),
.A2(n_705),
.B(n_771),
.Y(n_788)
);

OR2x2_ASAP7_75t_L g789 ( 
.A(n_704),
.B(n_739),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_742),
.Y(n_790)
);

BUFx3_ASAP7_75t_L g791 ( 
.A(n_770),
.Y(n_791)
);

INVx3_ASAP7_75t_L g792 ( 
.A(n_694),
.Y(n_792)
);

OAI22xp5_ASAP7_75t_L g793 ( 
.A1(n_744),
.A2(n_745),
.B1(n_756),
.B2(n_764),
.Y(n_793)
);

OA21x2_ASAP7_75t_L g794 ( 
.A1(n_746),
.A2(n_731),
.B(n_758),
.Y(n_794)
);

AND2x2_ASAP7_75t_SL g795 ( 
.A(n_710),
.B(n_747),
.Y(n_795)
);

OAI21x1_ASAP7_75t_L g796 ( 
.A1(n_700),
.A2(n_767),
.B(n_763),
.Y(n_796)
);

NAND2x1p5_ASAP7_75t_L g797 ( 
.A(n_748),
.B(n_743),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_749),
.Y(n_798)
);

OAI21x1_ASAP7_75t_L g799 ( 
.A1(n_733),
.A2(n_777),
.B(n_762),
.Y(n_799)
);

AO31x2_ASAP7_75t_L g800 ( 
.A1(n_740),
.A2(n_728),
.A3(n_723),
.B(n_697),
.Y(n_800)
);

CKINVDCx11_ASAP7_75t_R g801 ( 
.A(n_743),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_750),
.Y(n_802)
);

OAI21x1_ASAP7_75t_SL g803 ( 
.A1(n_755),
.A2(n_769),
.B(n_727),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_772),
.Y(n_804)
);

CKINVDCx16_ASAP7_75t_R g805 ( 
.A(n_716),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_722),
.Y(n_806)
);

OA21x2_ASAP7_75t_L g807 ( 
.A1(n_719),
.A2(n_703),
.B(n_695),
.Y(n_807)
);

OAI21xp5_ASAP7_75t_L g808 ( 
.A1(n_757),
.A2(n_741),
.B(n_715),
.Y(n_808)
);

OA21x2_ASAP7_75t_L g809 ( 
.A1(n_699),
.A2(n_729),
.B(n_702),
.Y(n_809)
);

OA21x2_ASAP7_75t_L g810 ( 
.A1(n_699),
.A2(n_702),
.B(n_778),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_707),
.A2(n_730),
.B1(n_759),
.B2(n_696),
.Y(n_811)
);

BUFx12f_ASAP7_75t_L g812 ( 
.A(n_775),
.Y(n_812)
);

HB1xp67_ASAP7_75t_L g813 ( 
.A(n_708),
.Y(n_813)
);

CKINVDCx20_ASAP7_75t_R g814 ( 
.A(n_737),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_699),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_773),
.B(n_751),
.Y(n_816)
);

INVx3_ASAP7_75t_L g817 ( 
.A(n_776),
.Y(n_817)
);

AOI21xp33_ASAP7_75t_L g818 ( 
.A1(n_717),
.A2(n_710),
.B(n_725),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_726),
.B(n_754),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_711),
.A2(n_725),
.B(n_732),
.Y(n_820)
);

OAI21xp5_ASAP7_75t_L g821 ( 
.A1(n_714),
.A2(n_732),
.B(n_774),
.Y(n_821)
);

OR2x6_ASAP7_75t_L g822 ( 
.A(n_712),
.B(n_721),
.Y(n_822)
);

AND2x4_ASAP7_75t_L g823 ( 
.A(n_709),
.B(n_714),
.Y(n_823)
);

NAND2x1p5_ASAP7_75t_L g824 ( 
.A(n_714),
.B(n_732),
.Y(n_824)
);

HB1xp67_ASAP7_75t_L g825 ( 
.A(n_752),
.Y(n_825)
);

HB1xp67_ASAP7_75t_L g826 ( 
.A(n_752),
.Y(n_826)
);

AOI22xp5_ASAP7_75t_L g827 ( 
.A1(n_759),
.A2(n_379),
.B1(n_644),
.B2(n_592),
.Y(n_827)
);

NAND2x1p5_ASAP7_75t_L g828 ( 
.A(n_770),
.B(n_612),
.Y(n_828)
);

BUFx3_ASAP7_75t_L g829 ( 
.A(n_770),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_759),
.B(n_644),
.Y(n_830)
);

HB1xp67_ASAP7_75t_L g831 ( 
.A(n_752),
.Y(n_831)
);

AND2x4_ASAP7_75t_L g832 ( 
.A(n_701),
.B(n_736),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_720),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_739),
.B(n_742),
.Y(n_834)
);

INVxp67_ASAP7_75t_L g835 ( 
.A(n_739),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_701),
.Y(n_836)
);

INVx3_ASAP7_75t_L g837 ( 
.A(n_693),
.Y(n_837)
);

BUFx3_ASAP7_75t_L g838 ( 
.A(n_770),
.Y(n_838)
);

AO31x2_ASAP7_75t_L g839 ( 
.A1(n_746),
.A2(n_633),
.A3(n_698),
.B(n_713),
.Y(n_839)
);

HB1xp67_ASAP7_75t_L g840 ( 
.A(n_780),
.Y(n_840)
);

HB1xp67_ASAP7_75t_L g841 ( 
.A(n_780),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_793),
.B(n_835),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_835),
.B(n_834),
.Y(n_843)
);

BUFx4f_ASAP7_75t_SL g844 ( 
.A(n_814),
.Y(n_844)
);

HB1xp67_ASAP7_75t_L g845 ( 
.A(n_781),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_803),
.Y(n_846)
);

BUFx2_ASAP7_75t_L g847 ( 
.A(n_824),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_790),
.B(n_798),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_783),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_802),
.B(n_787),
.Y(n_850)
);

BUFx3_ASAP7_75t_L g851 ( 
.A(n_828),
.Y(n_851)
);

OAI21xp5_ASAP7_75t_L g852 ( 
.A1(n_788),
.A2(n_785),
.B(n_820),
.Y(n_852)
);

CKINVDCx6p67_ASAP7_75t_R g853 ( 
.A(n_782),
.Y(n_853)
);

HB1xp67_ASAP7_75t_L g854 ( 
.A(n_781),
.Y(n_854)
);

HB1xp67_ASAP7_75t_L g855 ( 
.A(n_832),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_836),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_815),
.Y(n_857)
);

INVx2_ASAP7_75t_SL g858 ( 
.A(n_782),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_806),
.B(n_813),
.Y(n_859)
);

OR2x2_ASAP7_75t_L g860 ( 
.A(n_789),
.B(n_813),
.Y(n_860)
);

BUFx2_ASAP7_75t_L g861 ( 
.A(n_784),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_808),
.B(n_821),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_825),
.B(n_826),
.Y(n_863)
);

AND2x4_ASAP7_75t_L g864 ( 
.A(n_808),
.B(n_821),
.Y(n_864)
);

HB1xp67_ASAP7_75t_L g865 ( 
.A(n_832),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_826),
.B(n_831),
.Y(n_866)
);

OA21x2_ASAP7_75t_L g867 ( 
.A1(n_796),
.A2(n_786),
.B(n_799),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_830),
.B(n_827),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_839),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_812),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_863),
.B(n_810),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_843),
.B(n_804),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_861),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_866),
.B(n_810),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_861),
.Y(n_875)
);

OR2x2_ASAP7_75t_L g876 ( 
.A(n_860),
.B(n_809),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_842),
.B(n_843),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_850),
.B(n_811),
.Y(n_878)
);

INVx2_ASAP7_75t_SL g879 ( 
.A(n_851),
.Y(n_879)
);

INVxp67_ASAP7_75t_SL g880 ( 
.A(n_842),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_867),
.Y(n_881)
);

OR2x2_ASAP7_75t_L g882 ( 
.A(n_860),
.B(n_800),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_850),
.B(n_811),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_852),
.B(n_800),
.Y(n_884)
);

AND2x4_ASAP7_75t_L g885 ( 
.A(n_847),
.B(n_800),
.Y(n_885)
);

NOR2x1_ASAP7_75t_SL g886 ( 
.A(n_846),
.B(n_822),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_852),
.B(n_794),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_857),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_862),
.B(n_807),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_848),
.B(n_816),
.Y(n_890)
);

AND2x4_ASAP7_75t_SL g891 ( 
.A(n_840),
.B(n_841),
.Y(n_891)
);

INVx3_ASAP7_75t_L g892 ( 
.A(n_881),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_888),
.Y(n_893)
);

OR2x2_ASAP7_75t_L g894 ( 
.A(n_880),
.B(n_862),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_888),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_877),
.B(n_862),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_877),
.B(n_864),
.Y(n_897)
);

HB1xp67_ASAP7_75t_L g898 ( 
.A(n_873),
.Y(n_898)
);

BUFx3_ASAP7_75t_L g899 ( 
.A(n_891),
.Y(n_899)
);

NAND2x1p5_ASAP7_75t_L g900 ( 
.A(n_879),
.B(n_846),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_871),
.B(n_864),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_871),
.B(n_864),
.Y(n_902)
);

BUFx3_ASAP7_75t_L g903 ( 
.A(n_891),
.Y(n_903)
);

HB1xp67_ASAP7_75t_L g904 ( 
.A(n_875),
.Y(n_904)
);

OR2x2_ASAP7_75t_L g905 ( 
.A(n_876),
.B(n_882),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_885),
.B(n_864),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_874),
.B(n_869),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_901),
.B(n_902),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_893),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_893),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_901),
.B(n_902),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_896),
.B(n_889),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_895),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_896),
.B(n_889),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_897),
.B(n_887),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_897),
.B(n_887),
.Y(n_916)
);

HB1xp67_ASAP7_75t_L g917 ( 
.A(n_898),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_907),
.B(n_884),
.Y(n_918)
);

AND2x2_ASAP7_75t_L g919 ( 
.A(n_907),
.B(n_884),
.Y(n_919)
);

OR2x2_ASAP7_75t_L g920 ( 
.A(n_905),
.B(n_876),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_906),
.B(n_874),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_909),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_917),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_908),
.B(n_906),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_909),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_913),
.Y(n_926)
);

AND2x2_ASAP7_75t_L g927 ( 
.A(n_908),
.B(n_911),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_918),
.B(n_898),
.Y(n_928)
);

INVx1_ASAP7_75t_SL g929 ( 
.A(n_920),
.Y(n_929)
);

HB1xp67_ASAP7_75t_L g930 ( 
.A(n_920),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_911),
.B(n_906),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_912),
.B(n_906),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_918),
.B(n_904),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_919),
.B(n_904),
.Y(n_934)
);

AOI221xp5_ASAP7_75t_L g935 ( 
.A1(n_923),
.A2(n_916),
.B1(n_915),
.B2(n_919),
.C(n_912),
.Y(n_935)
);

HB1xp67_ASAP7_75t_L g936 ( 
.A(n_930),
.Y(n_936)
);

NAND3xp33_ASAP7_75t_SL g937 ( 
.A(n_929),
.B(n_900),
.C(n_833),
.Y(n_937)
);

NOR2x1_ASAP7_75t_L g938 ( 
.A(n_934),
.B(n_899),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_922),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_928),
.B(n_805),
.Y(n_940)
);

A2O1A1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_924),
.A2(n_903),
.B(n_899),
.C(n_891),
.Y(n_941)
);

NOR2x2_ASAP7_75t_L g942 ( 
.A(n_927),
.B(n_822),
.Y(n_942)
);

OAI221xp5_ASAP7_75t_L g943 ( 
.A1(n_933),
.A2(n_822),
.B1(n_868),
.B2(n_878),
.C(n_883),
.Y(n_943)
);

AND2x4_ASAP7_75t_L g944 ( 
.A(n_924),
.B(n_921),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_922),
.Y(n_945)
);

OAI221xp5_ASAP7_75t_L g946 ( 
.A1(n_938),
.A2(n_926),
.B1(n_925),
.B2(n_931),
.C(n_932),
.Y(n_946)
);

A2O1A1Ixp33_ASAP7_75t_L g947 ( 
.A1(n_937),
.A2(n_927),
.B(n_931),
.C(n_932),
.Y(n_947)
);

AOI22xp5_ASAP7_75t_L g948 ( 
.A1(n_943),
.A2(n_921),
.B1(n_915),
.B2(n_916),
.Y(n_948)
);

INVxp67_ASAP7_75t_L g949 ( 
.A(n_940),
.Y(n_949)
);

AOI221xp5_ASAP7_75t_L g950 ( 
.A1(n_935),
.A2(n_936),
.B1(n_939),
.B2(n_945),
.C(n_944),
.Y(n_950)
);

AOI22xp33_ASAP7_75t_L g951 ( 
.A1(n_944),
.A2(n_894),
.B1(n_905),
.B2(n_899),
.Y(n_951)
);

AOI221xp5_ASAP7_75t_L g952 ( 
.A1(n_950),
.A2(n_949),
.B1(n_946),
.B2(n_947),
.C(n_948),
.Y(n_952)
);

OAI32xp33_ASAP7_75t_L g953 ( 
.A1(n_951),
.A2(n_942),
.A3(n_903),
.B1(n_900),
.B2(n_894),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_948),
.Y(n_954)
);

AOI221xp5_ASAP7_75t_L g955 ( 
.A1(n_952),
.A2(n_925),
.B1(n_941),
.B2(n_872),
.C(n_910),
.Y(n_955)
);

NOR2x1_ASAP7_75t_L g956 ( 
.A(n_954),
.B(n_823),
.Y(n_956)
);

NOR3xp33_ASAP7_75t_L g957 ( 
.A(n_955),
.B(n_956),
.C(n_953),
.Y(n_957)
);

CKINVDCx20_ASAP7_75t_R g958 ( 
.A(n_955),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_958),
.B(n_914),
.Y(n_959)
);

OAI311xp33_ASAP7_75t_L g960 ( 
.A1(n_957),
.A2(n_859),
.A3(n_844),
.B1(n_890),
.C1(n_848),
.Y(n_960)
);

INVx1_ASAP7_75t_SL g961 ( 
.A(n_959),
.Y(n_961)
);

OAI22xp33_ASAP7_75t_L g962 ( 
.A1(n_960),
.A2(n_853),
.B1(n_870),
.B2(n_903),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_961),
.Y(n_963)
);

AND2x4_ASAP7_75t_SL g964 ( 
.A(n_962),
.B(n_870),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_961),
.B(n_914),
.Y(n_965)
);

AO22x2_ASAP7_75t_L g966 ( 
.A1(n_963),
.A2(n_858),
.B1(n_823),
.B2(n_829),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_965),
.B(n_858),
.Y(n_967)
);

AOI22xp5_ASAP7_75t_L g968 ( 
.A1(n_964),
.A2(n_853),
.B1(n_795),
.B2(n_779),
.Y(n_968)
);

BUFx2_ASAP7_75t_L g969 ( 
.A(n_963),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_963),
.B(n_886),
.Y(n_970)
);

NAND2x1p5_ASAP7_75t_L g971 ( 
.A(n_969),
.B(n_791),
.Y(n_971)
);

NAND2x1p5_ASAP7_75t_L g972 ( 
.A(n_968),
.B(n_838),
.Y(n_972)
);

AOI22xp33_ASAP7_75t_L g973 ( 
.A1(n_970),
.A2(n_801),
.B1(n_879),
.B2(n_892),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_966),
.A2(n_967),
.B(n_828),
.Y(n_974)
);

XNOR2xp5_ASAP7_75t_L g975 ( 
.A(n_968),
.B(n_845),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_SL g976 ( 
.A1(n_969),
.A2(n_886),
.B(n_819),
.Y(n_976)
);

AOI22x1_ASAP7_75t_SL g977 ( 
.A1(n_969),
.A2(n_837),
.B1(n_817),
.B2(n_792),
.Y(n_977)
);

AO21x2_ASAP7_75t_L g978 ( 
.A1(n_974),
.A2(n_818),
.B(n_859),
.Y(n_978)
);

OAI21xp5_ASAP7_75t_L g979 ( 
.A1(n_971),
.A2(n_818),
.B(n_797),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_973),
.B(n_849),
.Y(n_980)
);

OA22x2_ASAP7_75t_L g981 ( 
.A1(n_975),
.A2(n_854),
.B1(n_855),
.B2(n_865),
.Y(n_981)
);

OAI21xp5_ASAP7_75t_L g982 ( 
.A1(n_981),
.A2(n_972),
.B(n_976),
.Y(n_982)
);

OAI22xp5_ASAP7_75t_L g983 ( 
.A1(n_980),
.A2(n_977),
.B1(n_856),
.B2(n_849),
.Y(n_983)
);

OR2x6_ASAP7_75t_L g984 ( 
.A(n_982),
.B(n_979),
.Y(n_984)
);

AOI22xp33_ASAP7_75t_L g985 ( 
.A1(n_984),
.A2(n_983),
.B1(n_978),
.B2(n_851),
.Y(n_985)
);


endmodule