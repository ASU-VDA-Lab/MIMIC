module fake_jpeg_28964_n_173 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_173);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_27),
.Y(n_50)
);

BUFx8_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_44),
.Y(n_58)
);

BUFx16f_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_0),
.Y(n_61)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_15),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_5),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_49),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_10),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_35),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx10_ASAP7_75t_L g69 ( 
.A(n_12),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_9),
.Y(n_70)
);

BUFx16f_ASAP7_75t_L g71 ( 
.A(n_3),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_42),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_3),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_0),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

NOR3xp33_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_21),
.C(n_48),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_51),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_59),
.Y(n_77)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_61),
.B(n_1),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_83),
.Y(n_94)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_79),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_1),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_80),
.B(n_51),
.Y(n_100)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_73),
.B(n_2),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_84),
.Y(n_90)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_85),
.A2(n_70),
.B1(n_71),
.B2(n_66),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_86),
.A2(n_87),
.B1(n_68),
.B2(n_55),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_79),
.A2(n_71),
.B1(n_60),
.B2(n_66),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_92),
.Y(n_103)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_91),
.Y(n_110)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_57),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_95),
.B(n_62),
.Y(n_113)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_98),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_53),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_59),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_118),
.C(n_62),
.Y(n_131)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_90),
.Y(n_104)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_50),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_106),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_96),
.A2(n_68),
.B1(n_55),
.B2(n_75),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_107),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_108),
.A2(n_114),
.B(n_106),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_100),
.B(n_69),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_120),
.Y(n_130)
);

AND2x4_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_69),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_111),
.A2(n_4),
.B(n_6),
.Y(n_139)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_90),
.Y(n_112)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_116),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_69),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_115),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_88),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_98),
.Y(n_117)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_89),
.B(n_54),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_119),
.B(n_110),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_56),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_92),
.B(n_58),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_2),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g122 ( 
.A1(n_91),
.A2(n_72),
.B1(n_67),
.B2(n_65),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_122),
.A2(n_63),
.B1(n_99),
.B2(n_62),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_134),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_129),
.A2(n_137),
.B1(n_138),
.B2(n_13),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_133),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_114),
.Y(n_134)
);

INVxp67_ASAP7_75t_SL g135 ( 
.A(n_102),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_135),
.Y(n_153)
);

OAI32xp33_ASAP7_75t_L g136 ( 
.A1(n_103),
.A2(n_22),
.A3(n_46),
.B1(n_40),
.B2(n_39),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_136),
.B(n_16),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_103),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_139),
.A2(n_11),
.B(n_12),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_111),
.A2(n_20),
.B1(n_37),
.B2(n_36),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_140),
.A2(n_142),
.B1(n_8),
.B2(n_9),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_111),
.A2(n_19),
.B1(n_34),
.B2(n_33),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_7),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_143),
.B(n_144),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_109),
.B(n_8),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_145),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_123),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_147),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_135),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_148),
.A2(n_151),
.B(n_152),
.Y(n_163)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_141),
.Y(n_150)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_125),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_11),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_131),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_161),
.A2(n_153),
.B1(n_132),
.B2(n_140),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_127),
.C(n_126),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_162),
.A2(n_154),
.B1(n_142),
.B2(n_153),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_165),
.C(n_139),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_163),
.A2(n_159),
.B1(n_132),
.B2(n_145),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_166),
.B(n_162),
.Y(n_167)
);

AOI322xp5_ASAP7_75t_L g169 ( 
.A1(n_167),
.A2(n_168),
.A3(n_160),
.B1(n_165),
.B2(n_136),
.C1(n_161),
.C2(n_157),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_169),
.B(n_151),
.Y(n_170)
);

AOI322xp5_ASAP7_75t_L g171 ( 
.A1(n_170),
.A2(n_158),
.A3(n_124),
.B1(n_23),
.B2(n_24),
.C1(n_26),
.C2(n_17),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_18),
.C(n_28),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_29),
.Y(n_173)
);


endmodule