module real_jpeg_33937_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_657;
wire n_643;
wire n_656;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_669;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_679;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_666;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_685;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_680;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_678;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_578;
wire n_328;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_682;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_684;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_673;
wire n_631;
wire n_175;
wire n_338;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_411;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_615;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_670;
wire n_589;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_638;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_572;
wire n_155;
wire n_586;
wire n_405;
wire n_412;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_667;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_683;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_677;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_675;
wire n_138;
wire n_662;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_681;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_660;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_0),
.Y(n_84)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_0),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_0),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_0),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_0),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_1),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_2),
.A2(n_179),
.B1(n_180),
.B2(n_183),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g179 ( 
.A(n_2),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g426 ( 
.A1(n_2),
.A2(n_179),
.B1(n_197),
.B2(n_427),
.Y(n_426)
);

AOI22xp33_ASAP7_75t_SL g488 ( 
.A1(n_2),
.A2(n_179),
.B1(n_489),
.B2(n_494),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_3),
.A2(n_145),
.B1(n_149),
.B2(n_150),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_3),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_3),
.A2(n_149),
.B1(n_239),
.B2(n_240),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_3),
.A2(n_149),
.B1(n_358),
.B2(n_360),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_3),
.A2(n_149),
.B1(n_454),
.B2(n_456),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g676 ( 
.A(n_4),
.Y(n_676)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_5),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_5),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_5),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_6),
.Y(n_107)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_6),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_7),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_7),
.Y(n_330)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_7),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_8),
.A2(n_86),
.B1(n_90),
.B2(n_92),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_8),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_8),
.A2(n_92),
.B1(n_197),
.B2(n_200),
.Y(n_196)
);

OAI22x1_ASAP7_75t_L g600 ( 
.A1(n_8),
.A2(n_92),
.B1(n_601),
.B2(n_603),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_L g654 ( 
.A1(n_8),
.A2(n_92),
.B1(n_655),
.B2(n_658),
.Y(n_654)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_9),
.A2(n_76),
.B1(n_79),
.B2(n_80),
.Y(n_75)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_9),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_9),
.A2(n_79),
.B1(n_268),
.B2(n_270),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g622 ( 
.A1(n_9),
.A2(n_79),
.B1(n_377),
.B2(n_623),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_L g663 ( 
.A1(n_9),
.A2(n_79),
.B1(n_229),
.B2(n_658),
.Y(n_663)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_10),
.A2(n_54),
.B1(n_58),
.B2(n_59),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_10),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_10),
.A2(n_58),
.B1(n_113),
.B2(n_117),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g325 ( 
.A1(n_10),
.A2(n_58),
.B1(n_326),
.B2(n_331),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g588 ( 
.A1(n_10),
.A2(n_58),
.B1(n_589),
.B2(n_593),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_11),
.B(n_150),
.Y(n_317)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_11),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_11),
.B(n_154),
.Y(n_414)
);

OAI32xp33_ASAP7_75t_L g434 ( 
.A1(n_11),
.A2(n_427),
.A3(n_435),
.B1(n_440),
.B2(n_446),
.Y(n_434)
);

AOI22xp33_ASAP7_75t_SL g469 ( 
.A1(n_11),
.A2(n_344),
.B1(n_371),
.B2(n_470),
.Y(n_469)
);

OAI21xp33_ASAP7_75t_L g554 ( 
.A1(n_11),
.A2(n_93),
.B(n_498),
.Y(n_554)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_12),
.Y(n_71)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_12),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_13),
.A2(n_228),
.B1(n_229),
.B2(n_230),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_13),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_13),
.A2(n_228),
.B1(n_377),
.B2(n_379),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_13),
.A2(n_228),
.B1(n_475),
.B2(n_478),
.Y(n_474)
);

AOI22xp33_ASAP7_75t_SL g509 ( 
.A1(n_13),
.A2(n_228),
.B1(n_510),
.B2(n_513),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_14),
.Y(n_675)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_14),
.B(n_673),
.Y(n_685)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_15),
.A2(n_31),
.B1(n_35),
.B2(n_36),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_15),
.A2(n_35),
.B1(n_210),
.B2(n_213),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_15),
.A2(n_35),
.B1(n_256),
.B2(n_260),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_15),
.A2(n_35),
.B1(n_314),
.B2(n_615),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_16),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_16),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_17),
.A2(n_136),
.B1(n_139),
.B2(n_140),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_17),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_17),
.A2(n_139),
.B1(n_219),
.B2(n_224),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_17),
.A2(n_139),
.B1(n_284),
.B2(n_287),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_17),
.A2(n_139),
.B1(n_407),
.B2(n_411),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_18),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_18),
.Y(n_124)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_18),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_18),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_671),
.B(n_683),
.Y(n_19)
);

AOI31xp33_ASAP7_75t_L g683 ( 
.A1(n_20),
.A2(n_672),
.A3(n_684),
.B(n_685),
.Y(n_683)
);

AO21x2_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_580),
.B(n_665),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_415),
.B(n_572),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_349),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g572 ( 
.A1(n_23),
.A2(n_573),
.B(n_575),
.Y(n_572)
);

OA21x2_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_246),
.B(n_292),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_24),
.B(n_246),
.Y(n_579)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_25),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_187),
.C(n_204),
.Y(n_25)
);

INVxp33_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_27),
.B(n_187),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_98),
.Y(n_27)
);

INVxp67_ASAP7_75t_SL g248 ( 
.A(n_28),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_74),
.Y(n_28)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_29),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_42),
.B1(n_53),
.B2(n_63),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_30),
.A2(n_42),
.B1(n_63),
.B2(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_33),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_41),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_41),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_42),
.A2(n_53),
.B1(n_63),
.B2(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_42),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_42),
.A2(n_63),
.B1(n_426),
.B2(n_474),
.Y(n_473)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_64),
.Y(n_63)
);

OAI22x1_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_46),
.B1(n_50),
.B2(n_51),
.Y(n_43)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

BUFx2_ASAP7_75t_SL g512 ( 
.A(n_44),
.Y(n_512)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_45),
.Y(n_215)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_45),
.Y(n_493)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx4f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_55),
.Y(n_224)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_57),
.Y(n_273)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_63),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_63),
.Y(n_425)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_67),
.B1(n_70),
.B2(n_72),
.Y(n_64)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_65),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_66),
.Y(n_199)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_66),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_66),
.Y(n_363)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_66),
.Y(n_548)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_70),
.Y(n_540)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp33_ASAP7_75t_SL g541 ( 
.A(n_73),
.B(n_371),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_74),
.A2(n_299),
.B1(n_300),
.B2(n_301),
.Y(n_298)
);

INVxp67_ASAP7_75t_SL g301 ( 
.A(n_74),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_83),
.B1(n_85),
.B2(n_93),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_75),
.A2(n_189),
.B(n_190),
.Y(n_188)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_76),
.Y(n_455)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_77),
.Y(n_538)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_78),
.Y(n_212)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx4f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_85),
.A2(n_93),
.B1(n_208),
.B2(n_216),
.Y(n_207)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_90),
.Y(n_456)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_91),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_91),
.Y(n_497)
);

OA22x2_ASAP7_75t_L g402 ( 
.A1(n_93),
.A2(n_325),
.B1(n_403),
.B2(n_406),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_93),
.A2(n_488),
.B(n_498),
.Y(n_487)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_94),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_94),
.A2(n_209),
.B1(n_324),
.B2(n_332),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_94),
.B(n_453),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_94),
.A2(n_332),
.B1(n_508),
.B2(n_515),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.Y(n_94)
);

INVx5_ASAP7_75t_L g514 ( 
.A(n_95),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_142),
.B1(n_185),
.B2(n_186),
.Y(n_98)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_99),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_112),
.B1(n_121),
.B2(n_135),
.Y(n_99)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_100),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_100),
.B(n_238),
.Y(n_347)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_122),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_105),
.B1(n_108),
.B2(n_110),
.Y(n_101)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_102),
.Y(n_527)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g430 ( 
.A(n_104),
.Y(n_430)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_107),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_107),
.Y(n_127)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g445 ( 
.A(n_111),
.Y(n_445)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_112),
.A2(n_121),
.B1(n_254),
.B2(n_255),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g113 ( 
.A(n_114),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_116),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g164 ( 
.A(n_116),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_116),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_116),
.Y(n_265)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_121),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_121),
.B(n_376),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_121),
.B(n_238),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_SL g599 ( 
.A1(n_121),
.A2(n_254),
.B1(n_255),
.B2(n_600),
.Y(n_599)
);

AO22x2_ASAP7_75t_L g621 ( 
.A1(n_121),
.A2(n_254),
.B1(n_600),
.B2(n_622),
.Y(n_621)
);

OAI21xp33_ASAP7_75t_SL g650 ( 
.A1(n_121),
.A2(n_254),
.B(n_622),
.Y(n_650)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_125),
.B1(n_128),
.B2(n_132),
.Y(n_122)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_123),
.Y(n_239)
);

INVx5_ASAP7_75t_L g378 ( 
.A(n_123),
.Y(n_378)
);

INVx4_ASAP7_75t_L g380 ( 
.A(n_123),
.Y(n_380)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_124),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_124),
.Y(n_472)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_133),
.Y(n_141)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_133),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g138 ( 
.A(n_134),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_134),
.Y(n_608)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_135),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_142),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_165),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_143),
.B(n_165),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_143),
.B(n_366),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_154),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_144),
.B(n_166),
.Y(n_281)
);

INVx3_ASAP7_75t_SL g145 ( 
.A(n_146),
.Y(n_145)
);

INVx4_ASAP7_75t_SL g146 ( 
.A(n_147),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_148),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_148),
.Y(n_286)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_152),
.Y(n_234)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_152),
.Y(n_618)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g290 ( 
.A(n_153),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_153),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g592 ( 
.A(n_153),
.Y(n_592)
);

AO22x1_ASAP7_75t_L g226 ( 
.A1(n_154),
.A2(n_166),
.B1(n_178),
.B2(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_154),
.B(n_283),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_154),
.B(n_227),
.Y(n_336)
);

BUFx2_ASAP7_75t_L g587 ( 
.A(n_154),
.Y(n_587)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_155),
.B(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_159),
.B1(n_162),
.B2(n_163),
.Y(n_155)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_157),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_158),
.Y(n_162)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_158),
.Y(n_174)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_158),
.Y(n_322)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_160),
.Y(n_242)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_161),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_161),
.Y(n_442)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_162),
.Y(n_312)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_178),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_166),
.B(n_367),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g586 ( 
.A(n_166),
.Y(n_586)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_173),
.B1(n_175),
.B2(n_177),
.Y(n_167)
);

INVx2_ASAP7_75t_SL g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_171),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx4_ASAP7_75t_L g370 ( 
.A(n_176),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_176),
.Y(n_594)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_179),
.A2(n_340),
.B(n_343),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_179),
.B(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx4_ASAP7_75t_SL g181 ( 
.A(n_182),
.Y(n_181)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_183),
.Y(n_229)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_186),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_195),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_188),
.B(n_195),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_188),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g552 ( 
.A1(n_190),
.A2(n_452),
.B(n_509),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_190),
.B(n_371),
.Y(n_556)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_191),
.Y(n_216)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_196),
.Y(n_276)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g359 ( 
.A(n_199),
.Y(n_359)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_205),
.B(n_294),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_225),
.C(n_235),
.Y(n_205)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_206),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_217),
.Y(n_206)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_207),
.Y(n_383)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_217),
.Y(n_384)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_218),
.Y(n_364)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx4f_ASAP7_75t_SL g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_223),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_226),
.B(n_236),
.Y(n_303)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_231),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

OAI22x1_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_243),
.B1(n_244),
.B2(n_245),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_241),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_243),
.A2(n_339),
.B(n_347),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g468 ( 
.A1(n_243),
.A2(n_347),
.B(n_469),
.Y(n_468)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_245),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_245),
.A2(n_399),
.B(n_400),
.Y(n_398)
);

NOR2xp67_ASAP7_75t_R g486 ( 
.A(n_245),
.B(n_371),
.Y(n_486)
);

NOR2xp67_ASAP7_75t_L g577 ( 
.A(n_246),
.B(n_578),
.Y(n_577)
);

XOR2x2_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_251),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g634 ( 
.A(n_247),
.B(n_635),
.C(n_636),
.Y(n_634)
);

MAJx2_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.C(n_250),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_277),
.Y(n_251)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_252),
.Y(n_636)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_266),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_253),
.B(n_266),
.Y(n_630)
);

AOI21x1_ASAP7_75t_L g373 ( 
.A1(n_254),
.A2(n_374),
.B(n_375),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g256 ( 
.A(n_257),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_259),
.Y(n_439)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_264),
.Y(n_310)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_274),
.B1(n_275),
.B2(n_276),
.Y(n_266)
);

OA21x2_ASAP7_75t_L g596 ( 
.A1(n_267),
.A2(n_274),
.B(n_275),
.Y(n_596)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVxp67_ASAP7_75t_SL g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_274),
.A2(n_275),
.B1(n_357),
.B2(n_364),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_274),
.B(n_357),
.Y(n_431)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_274),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_275),
.B(n_357),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_275),
.B(n_544),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_277),
.Y(n_635)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

OAI21xp33_ASAP7_75t_L g632 ( 
.A1(n_278),
.A2(n_280),
.B(n_291),
.Y(n_632)
);

XNOR2x1_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_291),
.Y(n_279)
);

NAND2x1_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_281),
.B(n_336),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_SL g585 ( 
.A1(n_283),
.A2(n_586),
.B1(n_587),
.B2(n_588),
.Y(n_585)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_295),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g576 ( 
.A(n_293),
.B(n_295),
.Y(n_576)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_305),
.B(n_348),
.Y(n_295)
);

NOR2xp67_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_302),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_297),
.B(n_302),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_297),
.A2(n_298),
.B1(n_302),
.B2(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_302),
.Y(n_387)
);

XNOR2x1_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_305),
.B(n_386),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_334),
.C(n_337),
.Y(n_305)
);

INVxp67_ASAP7_75t_SL g306 ( 
.A(n_307),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_307),
.B(n_354),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_323),
.Y(n_307)
);

XOR2x2_ASAP7_75t_L g395 ( 
.A(n_308),
.B(n_323),
.Y(n_395)
);

AOI32xp33_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_311),
.A3(n_313),
.B1(n_317),
.B2(n_318),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx11_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

BUFx12f_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_317),
.Y(n_372)
);

NAND2xp33_ASAP7_75t_SL g318 ( 
.A(n_319),
.B(n_321),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_329),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx6_ASAP7_75t_L g410 ( 
.A(n_330),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_330),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_334),
.A2(n_335),
.B1(n_337),
.B2(n_338),
.Y(n_354)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_339),
.Y(n_374)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_342),
.Y(n_341)
);

INVx5_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx8_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_350),
.A2(n_385),
.B(n_388),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_350),
.B(n_385),
.C(n_574),
.Y(n_573)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_355),
.C(n_381),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_353),
.B(n_391),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_355),
.B(n_382),
.Y(n_391)
);

MAJx2_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_365),
.C(n_373),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_356),
.B(n_373),
.Y(n_394)
);

INVx2_ASAP7_75t_SL g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_363),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_365),
.B(n_394),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_368),
.A2(n_371),
.B(n_372),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g368 ( 
.A(n_369),
.Y(n_368)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_370),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_371),
.B(n_447),
.Y(n_446)
);

OAI21xp33_ASAP7_75t_SL g544 ( 
.A1(n_371),
.A2(n_541),
.B(n_545),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_SL g551 ( 
.A(n_371),
.B(n_484),
.Y(n_551)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_376),
.Y(n_399)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx3_ASAP7_75t_SL g379 ( 
.A(n_380),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_384),
.Y(n_382)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_390),
.B(n_392),
.Y(n_389)
);

OR2x2_ASAP7_75t_L g574 ( 
.A(n_390),
.B(n_392),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_395),
.C(n_396),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_393),
.B(n_458),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_395),
.A2(n_396),
.B1(n_397),
.B2(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_SL g459 ( 
.A(n_395),
.Y(n_459)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_401),
.C(n_414),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_398),
.B(n_422),
.Y(n_421)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_402),
.B(n_414),
.Y(n_422)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

BUFx4f_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g448 ( 
.A1(n_406),
.A2(n_449),
.B(n_452),
.Y(n_448)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

OAI21x1_ASAP7_75t_SL g416 ( 
.A1(n_417),
.A2(n_460),
.B(n_570),
.Y(n_416)
);

AND2x4_ASAP7_75t_SL g417 ( 
.A(n_418),
.B(n_457),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_419),
.B(n_571),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_423),
.C(n_432),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_421),
.B(n_464),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g464 ( 
.A1(n_423),
.A2(n_424),
.B1(n_433),
.B2(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

OAI21xp33_ASAP7_75t_SL g424 ( 
.A1(n_425),
.A2(n_426),
.B(n_431),
.Y(n_424)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx4_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_431),
.B(n_543),
.Y(n_542)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_433),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_448),
.Y(n_433)
);

XOR2x2_ASAP7_75t_L g467 ( 
.A(n_434),
.B(n_448),
.Y(n_467)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_443),
.Y(n_440)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_441),
.Y(n_602)
);

BUFx3_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

HB1xp67_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

BUFx3_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_451),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_453),
.B(n_499),
.Y(n_498)
);

INVx1_ASAP7_75t_SL g454 ( 
.A(n_455),
.Y(n_454)
);

INVxp67_ASAP7_75t_SL g571 ( 
.A(n_457),
.Y(n_571)
);

AOI21x1_ASAP7_75t_L g460 ( 
.A1(n_461),
.A2(n_504),
.B(n_569),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_479),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_463),
.B(n_466),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_463),
.B(n_466),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_468),
.C(n_473),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_467),
.B(n_481),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_468),
.B(n_473),
.Y(n_481)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_474),
.A2(n_484),
.B(n_485),
.Y(n_483)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx3_ASAP7_75t_SL g476 ( 
.A(n_477),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_480),
.B(n_482),
.Y(n_479)
);

OR2x2_ASAP7_75t_L g567 ( 
.A(n_480),
.B(n_482),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_486),
.C(n_487),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_483),
.B(n_486),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_L g564 ( 
.A(n_487),
.B(n_565),
.Y(n_564)
);

INVxp67_ASAP7_75t_L g515 ( 
.A(n_488),
.Y(n_515)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx4_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

INVx4_ASAP7_75t_L g492 ( 
.A(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

OAI211xp5_ASAP7_75t_SL g504 ( 
.A1(n_505),
.A2(n_563),
.B(n_567),
.C(n_568),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_506),
.A2(n_549),
.B(n_562),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_516),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_507),
.B(n_516),
.Y(n_562)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_517),
.B(n_542),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_517),
.B(n_542),
.Y(n_566)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_518),
.A2(n_524),
.B(n_533),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_525),
.B(n_528),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

BUFx2_ASAP7_75t_L g526 ( 
.A(n_527),
.Y(n_526)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_534),
.A2(n_539),
.B(n_541),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_546),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

INVx4_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

OAI21xp5_ASAP7_75t_SL g549 ( 
.A1(n_550),
.A2(n_553),
.B(n_561),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_551),
.B(n_552),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_551),
.B(n_552),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_554),
.B(n_555),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_SL g555 ( 
.A(n_556),
.B(n_557),
.Y(n_555)
);

INVx1_ASAP7_75t_SL g557 ( 
.A(n_558),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_559),
.Y(n_558)
);

HB1xp67_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

NOR2x1_ASAP7_75t_L g563 ( 
.A(n_564),
.B(n_566),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_564),
.B(n_566),
.Y(n_568)
);

OAI21xp5_ASAP7_75t_L g575 ( 
.A1(n_576),
.A2(n_577),
.B(n_579),
.Y(n_575)
);

NOR3xp33_ASAP7_75t_L g580 ( 
.A(n_581),
.B(n_639),
.C(n_661),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_582),
.B(n_633),
.Y(n_581)
);

A2O1A1Ixp33_ASAP7_75t_L g667 ( 
.A1(n_582),
.A2(n_640),
.B(n_668),
.C(n_669),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_583),
.B(n_626),
.Y(n_582)
);

NOR2x1_ASAP7_75t_L g669 ( 
.A(n_583),
.B(n_626),
.Y(n_669)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_584),
.B(n_609),
.Y(n_583)
);

INVxp67_ASAP7_75t_SL g644 ( 
.A(n_584),
.Y(n_644)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_585),
.B(n_595),
.C(n_597),
.Y(n_584)
);

XOR2xp5_ASAP7_75t_L g609 ( 
.A(n_585),
.B(n_610),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_L g627 ( 
.A(n_585),
.B(n_628),
.Y(n_627)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_585),
.Y(n_643)
);

INVx1_ASAP7_75t_SL g613 ( 
.A(n_586),
.Y(n_613)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_587),
.Y(n_619)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_587),
.A2(n_652),
.B1(n_653),
.B2(n_654),
.Y(n_651)
);

AOI22x1_ASAP7_75t_L g662 ( 
.A1(n_587),
.A2(n_653),
.B1(n_654),
.B2(n_663),
.Y(n_662)
);

OAI21xp5_ASAP7_75t_L g680 ( 
.A1(n_587),
.A2(n_653),
.B(n_663),
.Y(n_680)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_588),
.Y(n_612)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_590),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_591),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_592),
.Y(n_591)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_594),
.Y(n_593)
);

INVx3_ASAP7_75t_SL g657 ( 
.A(n_594),
.Y(n_657)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_595),
.Y(n_647)
);

HB1xp67_ASAP7_75t_L g595 ( 
.A(n_596),
.Y(n_595)
);

XOR2xp5_ASAP7_75t_L g620 ( 
.A(n_596),
.B(n_621),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g628 ( 
.A1(n_596),
.A2(n_598),
.B1(n_599),
.B2(n_629),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_596),
.Y(n_629)
);

HB1xp67_ASAP7_75t_L g597 ( 
.A(n_598),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_599),
.Y(n_598)
);

INVx1_ASAP7_75t_SL g601 ( 
.A(n_602),
.Y(n_601)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_604),
.Y(n_603)
);

HB1xp67_ASAP7_75t_L g604 ( 
.A(n_605),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_606),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_607),
.Y(n_606)
);

INVx4_ASAP7_75t_L g607 ( 
.A(n_608),
.Y(n_607)
);

HB1xp67_ASAP7_75t_L g642 ( 
.A(n_610),
.Y(n_642)
);

XNOR2xp5_ASAP7_75t_L g610 ( 
.A(n_611),
.B(n_620),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g646 ( 
.A(n_611),
.B(n_621),
.C(n_647),
.Y(n_646)
);

OAI22xp5_ASAP7_75t_SL g611 ( 
.A1(n_612),
.A2(n_613),
.B1(n_614),
.B2(n_619),
.Y(n_611)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_613),
.Y(n_653)
);

INVxp67_ASAP7_75t_L g652 ( 
.A(n_614),
.Y(n_652)
);

INVx1_ASAP7_75t_SL g615 ( 
.A(n_616),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_617),
.Y(n_616)
);

HB1xp67_ASAP7_75t_L g617 ( 
.A(n_618),
.Y(n_617)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_624),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_625),
.Y(n_624)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_627),
.B(n_630),
.C(n_631),
.Y(n_626)
);

XNOR2x1_ASAP7_75t_L g638 ( 
.A(n_627),
.B(n_630),
.Y(n_638)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_632),
.Y(n_631)
);

XNOR2xp5_ASAP7_75t_L g637 ( 
.A(n_632),
.B(n_638),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_634),
.B(n_637),
.Y(n_633)
);

NOR2xp67_ASAP7_75t_L g668 ( 
.A(n_634),
.B(n_637),
.Y(n_668)
);

INVxp67_ASAP7_75t_SL g639 ( 
.A(n_640),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_641),
.B(n_645),
.Y(n_640)
);

OR2x2_ASAP7_75t_L g666 ( 
.A(n_641),
.B(n_645),
.Y(n_666)
);

MAJIxp5_ASAP7_75t_L g641 ( 
.A(n_642),
.B(n_643),
.C(n_644),
.Y(n_641)
);

XNOR2xp5_ASAP7_75t_L g645 ( 
.A(n_646),
.B(n_648),
.Y(n_645)
);

MAJIxp5_ASAP7_75t_L g664 ( 
.A(n_646),
.B(n_649),
.C(n_651),
.Y(n_664)
);

XNOR2xp5_ASAP7_75t_L g648 ( 
.A(n_649),
.B(n_651),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_650),
.Y(n_649)
);

INVxp67_ASAP7_75t_L g655 ( 
.A(n_656),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_657),
.Y(n_656)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_659),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_660),
.Y(n_659)
);

A2O1A1Ixp33_ASAP7_75t_L g665 ( 
.A1(n_661),
.A2(n_666),
.B(n_667),
.C(n_670),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_662),
.B(n_664),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_662),
.B(n_664),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_662),
.B(n_679),
.Y(n_678)
);

CKINVDCx16_ASAP7_75t_R g682 ( 
.A(n_662),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_672),
.B(n_677),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_673),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_674),
.B(n_676),
.Y(n_673)
);

CKINVDCx20_ASAP7_75t_R g674 ( 
.A(n_675),
.Y(n_674)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_677),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_678),
.B(n_681),
.Y(n_677)
);

CKINVDCx20_ASAP7_75t_R g679 ( 
.A(n_680),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_680),
.B(n_682),
.Y(n_681)
);


endmodule