module real_jpeg_7600_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_166;
wire n_176;
wire n_288;
wire n_215;
wire n_221;
wire n_249;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_276;
wire n_163;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_65;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_80;
wire n_32;
wire n_20;
wire n_228;
wire n_74;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_259;
wire n_225;
wire n_103;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_279;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_216;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_269;
wire n_253;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_1),
.Y(n_77)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_1),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_1),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_2),
.A2(n_20),
.B1(n_25),
.B2(n_26),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_2),
.A2(n_25),
.B1(n_95),
.B2(n_98),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_2),
.A2(n_25),
.B1(n_234),
.B2(n_236),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_3),
.B(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_3),
.A2(n_81),
.B1(n_85),
.B2(n_86),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_3),
.Y(n_85)
);

O2A1O1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_3),
.A2(n_102),
.B(n_104),
.C(n_110),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_3),
.A2(n_85),
.B1(n_121),
.B2(n_125),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_3),
.B(n_76),
.C(n_147),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_3),
.B(n_28),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_3),
.B(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_3),
.B(n_128),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_3),
.A2(n_59),
.B1(n_85),
.B2(n_277),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_4),
.A2(n_53),
.B1(n_57),
.B2(n_58),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_4),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_4),
.A2(n_57),
.B1(n_137),
.B2(n_139),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_4),
.A2(n_57),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_4),
.A2(n_57),
.B1(n_226),
.B2(n_228),
.Y(n_225)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_6),
.Y(n_79)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_6),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_6),
.Y(n_250)
);

BUFx5_ASAP7_75t_L g64 ( 
.A(n_7),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_7),
.Y(n_69)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_7),
.Y(n_160)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_7),
.Y(n_185)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_9),
.Y(n_161)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_9),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_9),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_9),
.Y(n_181)
);

BUFx5_ASAP7_75t_L g189 ( 
.A(n_9),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_9),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_10),
.A2(n_76),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_10),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_11),
.Y(n_130)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_11),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g147 ( 
.A(n_11),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_11),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_206),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_204),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_150),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_15),
.B(n_150),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_100),
.C(n_115),
.Y(n_15)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_16),
.B(n_285),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_60),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_17),
.B(n_61),
.C(n_71),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_41),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_28),
.Y(n_18)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_19),
.Y(n_198)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g278 ( 
.A(n_22),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_27),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_28),
.B(n_52),
.Y(n_199)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_33),
.B1(n_35),
.B2(n_38),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_32),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_34),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_34),
.Y(n_124)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_34),
.Y(n_126)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_34),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_34),
.Y(n_238)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_35),
.Y(n_235)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_37),
.Y(n_141)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_42),
.B(n_52),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_42),
.B(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_43),
.B(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

AO22x1_ASAP7_75t_SL g63 ( 
.A1(n_47),
.A2(n_64),
.B1(n_65),
.B2(n_67),
.Y(n_63)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp33_ASAP7_75t_SL g166 ( 
.A(n_51),
.B(n_64),
.Y(n_166)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_54),
.Y(n_157)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_70),
.B2(n_71),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NOR2x1_ASAP7_75t_L g179 ( 
.A(n_63),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_63),
.B(n_191),
.Y(n_190)
);

INVx6_ASAP7_75t_SL g65 ( 
.A(n_66),
.Y(n_65)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_69),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_90),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_72),
.B(n_248),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_80),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_73),
.A2(n_80),
.B(n_113),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_73),
.B(n_94),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_73),
.B(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_78),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_77),
.Y(n_132)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_77),
.Y(n_229)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_80),
.Y(n_222)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

OAI21xp33_ASAP7_75t_L g104 ( 
.A1(n_85),
.A2(n_105),
.B(n_107),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_85),
.B(n_164),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_85),
.A2(n_163),
.B(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_86),
.Y(n_170)
);

INVx4_ASAP7_75t_SL g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_90),
.B(n_224),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_94),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_93),
.Y(n_172)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_93),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_96),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_97),
.Y(n_131)
);

BUFx8_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g257 ( 
.A(n_99),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_100),
.A2(n_115),
.B1(n_116),
.B2(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_100),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_112),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_101),
.A2(n_112),
.B1(n_280),
.B2(n_281),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_101),
.Y(n_281)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_109),
.Y(n_214)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_112),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_114),
.B(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_135),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_119),
.B(n_127),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_119),
.A2(n_127),
.B(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_120),
.B(n_142),
.Y(n_218)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_126),
.Y(n_149)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NOR2x1_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_128),
.B(n_136),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_128),
.B(n_233),
.Y(n_232)
);

AO22x1_ASAP7_75t_SL g128 ( 
.A1(n_129),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_131),
.Y(n_227)
);

BUFx5_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_135),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_142),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_138),
.Y(n_145)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_142),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_142),
.B(n_233),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_146),
.B1(n_148),
.B2(n_149),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx4_ASAP7_75t_SL g146 ( 
.A(n_147),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_174),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_154),
.B2(n_155),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_167),
.Y(n_155)
);

AOI32xp33_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_158),
.A3(n_161),
.B1(n_162),
.B2(n_166),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVxp33_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_164),
.Y(n_193)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_171),
.B(n_173),
.Y(n_167)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_173),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_194),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_190),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_186),
.B2(n_188),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_200),
.B1(n_201),
.B2(n_203),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_195),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_199),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_199),
.B(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_283),
.B(n_288),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_267),
.B(n_282),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_242),
.B(n_266),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_219),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_210),
.B(n_219),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_216),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_211),
.A2(n_212),
.B1(n_216),
.B2(n_245),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_215),
.Y(n_212)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_216),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_217),
.B(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_230),
.Y(n_219)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_220),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_223),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_249),
.Y(n_248)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_230)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_231),
.Y(n_240)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_239),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_239),
.B(n_240),
.C(n_269),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_252),
.B(n_265),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_246),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_244),
.B(n_246),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_251),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_261),
.B(n_264),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_260),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_258),
.Y(n_254)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_256),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_263),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_270),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_270),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_279),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_274),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_274),
.C(n_279),
.Y(n_287)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_284),
.B(n_287),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_287),
.Y(n_288)
);


endmodule