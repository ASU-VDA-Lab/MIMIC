module fake_jpeg_13183_n_532 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_532);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_532;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

INVx6_ASAP7_75t_SL g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx16f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_18),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_15),
.B(n_16),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_1),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

BUFx16f_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_12),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_8),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_59),
.Y(n_136)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_60),
.B(n_72),
.Y(n_125)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_61),
.Y(n_166)
);

HAxp5_ASAP7_75t_SL g62 ( 
.A(n_20),
.B(n_42),
.CON(n_62),
.SN(n_62)
);

AOI21xp33_ASAP7_75t_L g150 ( 
.A1(n_62),
.A2(n_86),
.B(n_30),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_63),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_40),
.A2(n_17),
.B1(n_16),
.B2(n_13),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_64),
.A2(n_41),
.B1(n_26),
.B2(n_55),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_65),
.Y(n_170)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx5_ASAP7_75t_L g151 ( 
.A(n_66),
.Y(n_151)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_67),
.Y(n_155)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_68),
.Y(n_141)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_69),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_70),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_40),
.B(n_18),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_71),
.B(n_91),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_36),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_73),
.Y(n_184)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_74),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_19),
.B(n_18),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_75),
.B(n_100),
.Y(n_195)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_76),
.Y(n_197)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_77),
.B(n_80),
.Y(n_131)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_78),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_79),
.Y(n_201)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

BUFx10_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_81),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_82),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_83),
.Y(n_154)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_57),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_84),
.B(n_109),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_31),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_85),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_35),
.B(n_13),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_87),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_88),
.Y(n_158)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_89),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_90),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_19),
.B(n_17),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_92),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_93),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_33),
.Y(n_94)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_94),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_27),
.B(n_12),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_95),
.B(n_104),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_96),
.Y(n_171)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_33),
.Y(n_98)
);

INVx8_ASAP7_75t_L g183 ( 
.A(n_98),
.Y(n_183)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_32),
.Y(n_99)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_27),
.B(n_0),
.Y(n_100)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_42),
.Y(n_101)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_101),
.Y(n_187)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

BUFx12_ASAP7_75t_L g148 ( 
.A(n_102),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_53),
.Y(n_103)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_103),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_28),
.B(n_1),
.Y(n_104)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_105),
.Y(n_147)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_106),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_28),
.B(n_12),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_107),
.B(n_115),
.Y(n_202)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_29),
.Y(n_108)
);

INVx6_ASAP7_75t_SL g175 ( 
.A(n_108),
.Y(n_175)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_34),
.Y(n_109)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_42),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_110),
.Y(n_192)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_51),
.Y(n_111)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_111),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_44),
.B(n_2),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_116),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_53),
.Y(n_113)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_113),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_32),
.Y(n_114)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_114),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_44),
.B(n_10),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_34),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_53),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_117),
.B(n_118),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_32),
.Y(n_118)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_32),
.Y(n_119)
);

INVx11_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_24),
.B(n_3),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_121),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_24),
.B(n_5),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_32),
.Y(n_122)
);

INVx2_ASAP7_75t_R g181 ( 
.A(n_122),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_26),
.B(n_5),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_123),
.B(n_124),
.Y(n_161)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_29),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_62),
.A2(n_42),
.B1(n_22),
.B2(n_53),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_129),
.A2(n_130),
.B1(n_156),
.B2(n_177),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_76),
.A2(n_22),
.B1(n_29),
.B2(n_45),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_100),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_133),
.B(n_169),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_61),
.A2(n_45),
.B1(n_22),
.B2(n_58),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_137),
.A2(n_138),
.B1(n_142),
.B2(n_165),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_117),
.A2(n_45),
.B1(n_56),
.B2(n_50),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_86),
.A2(n_45),
.B1(n_49),
.B2(n_48),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_140),
.A2(n_180),
.B1(n_36),
.B2(n_9),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_113),
.A2(n_38),
.B1(n_56),
.B2(n_50),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_63),
.A2(n_58),
.B1(n_38),
.B2(n_30),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_149),
.A2(n_204),
.B1(n_10),
.B2(n_202),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_150),
.B(n_162),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_101),
.A2(n_55),
.B1(n_39),
.B2(n_49),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_75),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_159),
.B(n_168),
.Y(n_233)
);

AND2x2_ASAP7_75t_SL g162 ( 
.A(n_99),
.B(n_6),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_65),
.A2(n_79),
.B1(n_82),
.B2(n_103),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_104),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_81),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_66),
.B(n_41),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_172),
.B(n_174),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_81),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_176),
.B(n_194),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_110),
.A2(n_48),
.B1(n_39),
.B2(n_37),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_70),
.A2(n_37),
.B1(n_54),
.B2(n_21),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_178),
.A2(n_203),
.B1(n_185),
.B2(n_158),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_70),
.A2(n_102),
.B1(n_93),
.B2(n_98),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_83),
.A2(n_54),
.B1(n_21),
.B2(n_36),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_185),
.A2(n_36),
.B1(n_8),
.B2(n_9),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_93),
.A2(n_37),
.B(n_54),
.Y(n_186)
);

O2A1O1Ixp33_ASAP7_75t_L g252 ( 
.A1(n_186),
.A2(n_126),
.B(n_180),
.C(n_192),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_74),
.B(n_54),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_102),
.B(n_21),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_196),
.B(n_198),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_94),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_108),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_199),
.B(n_151),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_108),
.A2(n_21),
.B1(n_7),
.B2(n_8),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_71),
.A2(n_36),
.B1(n_7),
.B2(n_8),
.Y(n_204)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_175),
.Y(n_206)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_206),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_207),
.A2(n_215),
.B1(n_234),
.B2(n_252),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_133),
.B(n_6),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_208),
.B(n_211),
.Y(n_276)
);

INVx3_ASAP7_75t_SL g210 ( 
.A(n_175),
.Y(n_210)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_210),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_162),
.B(n_6),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_213),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_162),
.B(n_10),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_216),
.B(n_228),
.Y(n_281)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_132),
.Y(n_219)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_219),
.Y(n_283)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_134),
.Y(n_220)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_220),
.Y(n_285)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_190),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g319 ( 
.A(n_221),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_132),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_222),
.Y(n_293)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_128),
.Y(n_223)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_223),
.Y(n_287)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_134),
.Y(n_224)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_224),
.Y(n_325)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_136),
.Y(n_225)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_225),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_136),
.B(n_10),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_226),
.B(n_248),
.C(n_199),
.Y(n_278)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_128),
.Y(n_227)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_227),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_191),
.B(n_161),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_125),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_229),
.B(n_231),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_135),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_230),
.B(n_247),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_131),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_151),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_232),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_195),
.A2(n_152),
.B1(n_140),
.B2(n_164),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_186),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_235),
.B(n_240),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_171),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_236),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_139),
.B(n_184),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_237),
.B(n_245),
.Y(n_288)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_171),
.Y(n_238)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_238),
.Y(n_300)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_179),
.Y(n_241)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_241),
.Y(n_305)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_179),
.Y(n_242)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_242),
.Y(n_316)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_145),
.Y(n_243)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_243),
.Y(n_318)
);

OA22x2_ASAP7_75t_L g244 ( 
.A1(n_169),
.A2(n_176),
.B1(n_127),
.B2(n_200),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_244),
.A2(n_254),
.B1(n_261),
.B2(n_267),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_155),
.B(n_184),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_158),
.Y(n_246)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_246),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_135),
.Y(n_247)
);

AND2x2_ASAP7_75t_SL g248 ( 
.A(n_181),
.B(n_155),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_145),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_249),
.B(n_250),
.Y(n_302)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_193),
.Y(n_250)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_190),
.Y(n_251)
);

INVx6_ASAP7_75t_L g315 ( 
.A(n_251),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_148),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_253),
.B(n_259),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_167),
.Y(n_256)
);

INVx3_ASAP7_75t_SL g309 ( 
.A(n_256),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_144),
.A2(n_142),
.B1(n_138),
.B2(n_137),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_257),
.A2(n_260),
.B1(n_269),
.B2(n_274),
.Y(n_286)
);

AO22x1_ASAP7_75t_L g258 ( 
.A1(n_127),
.A2(n_189),
.B1(n_200),
.B2(n_163),
.Y(n_258)
);

A2O1A1Ixp33_ASAP7_75t_L g307 ( 
.A1(n_258),
.A2(n_192),
.B(n_197),
.C(n_148),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_148),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_146),
.A2(n_182),
.B1(n_154),
.B2(n_189),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_160),
.A2(n_165),
.B1(n_141),
.B2(n_143),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_160),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_262),
.B(n_265),
.Y(n_303)
);

BUFx2_ASAP7_75t_SL g263 ( 
.A(n_205),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_263),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_181),
.B(n_193),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_264),
.B(n_272),
.Y(n_290)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_205),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_141),
.B(n_143),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_266),
.B(n_268),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_173),
.A2(n_188),
.B1(n_147),
.B2(n_153),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_147),
.B(n_188),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_173),
.A2(n_153),
.B1(n_157),
.B2(n_187),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_166),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_270),
.B(n_273),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_166),
.A2(n_146),
.B1(n_182),
.B2(n_154),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g313 ( 
.A1(n_271),
.A2(n_207),
.B1(n_250),
.B2(n_243),
.Y(n_313)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_163),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_126),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_157),
.A2(n_187),
.B1(n_163),
.B2(n_183),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_217),
.B(n_126),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_277),
.B(n_311),
.C(n_248),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_SL g364 ( 
.A(n_278),
.B(n_299),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_214),
.A2(n_167),
.B1(n_170),
.B2(n_201),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_279),
.A2(n_308),
.B1(n_310),
.B2(n_286),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_239),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_284),
.B(n_321),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_208),
.B(n_183),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_295),
.B(n_304),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_211),
.B(n_170),
.Y(n_304)
);

O2A1O1Ixp33_ASAP7_75t_L g338 ( 
.A1(n_307),
.A2(n_244),
.B(n_258),
.C(n_272),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_214),
.A2(n_197),
.B1(n_201),
.B2(n_235),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_209),
.A2(n_212),
.B1(n_255),
.B2(n_273),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_217),
.B(n_228),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_233),
.B(n_218),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_312),
.B(n_326),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_313),
.A2(n_242),
.B1(n_241),
.B2(n_227),
.Y(n_330)
);

BUFx24_ASAP7_75t_SL g314 ( 
.A(n_229),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_314),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_264),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_245),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_323),
.B(n_246),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_237),
.B(n_219),
.Y(n_326)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_318),
.Y(n_328)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_328),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_296),
.A2(n_217),
.B(n_252),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g368 ( 
.A1(n_329),
.A2(n_353),
.B(n_338),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_330),
.A2(n_346),
.B1(n_351),
.B2(n_275),
.Y(n_372)
);

INVx1_ASAP7_75t_SL g331 ( 
.A(n_320),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_331),
.B(n_333),
.Y(n_376)
);

A2O1A1Ixp33_ASAP7_75t_L g332 ( 
.A1(n_278),
.A2(n_216),
.B(n_226),
.C(n_248),
.Y(n_332)
);

A2O1A1Ixp33_ASAP7_75t_L g397 ( 
.A1(n_332),
.A2(n_334),
.B(n_358),
.C(n_340),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_301),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_334),
.B(n_362),
.Y(n_390)
);

OAI21xp33_ASAP7_75t_L g335 ( 
.A1(n_321),
.A2(n_226),
.B(n_244),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_335),
.A2(n_336),
.B(n_352),
.Y(n_398)
);

AOI22x1_ASAP7_75t_SL g336 ( 
.A1(n_308),
.A2(n_244),
.B1(n_206),
.B2(n_271),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_323),
.B(n_223),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_337),
.B(n_342),
.Y(n_374)
);

O2A1O1Ixp33_ASAP7_75t_L g379 ( 
.A1(n_338),
.A2(n_317),
.B(n_300),
.C(n_297),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_288),
.B(n_249),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_288),
.B(n_290),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_343),
.B(n_349),
.Y(n_395)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_318),
.Y(n_344)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_344),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_281),
.B(n_265),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_345),
.B(n_350),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_294),
.A2(n_270),
.B1(n_251),
.B2(n_225),
.Y(n_346)
);

OA22x2_ASAP7_75t_SL g347 ( 
.A1(n_307),
.A2(n_258),
.B1(n_210),
.B2(n_221),
.Y(n_347)
);

A2O1A1Ixp33_ASAP7_75t_SL g391 ( 
.A1(n_347),
.A2(n_357),
.B(n_285),
.C(n_325),
.Y(n_391)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_283),
.Y(n_348)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_348),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_290),
.B(n_295),
.Y(n_349)
);

INVxp33_ASAP7_75t_L g350 ( 
.A(n_298),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_294),
.A2(n_256),
.B1(n_232),
.B2(n_238),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_352),
.B(n_354),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g353 ( 
.A1(n_310),
.A2(n_259),
.B(n_262),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_284),
.B(n_236),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_281),
.B(n_220),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_355),
.B(n_358),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_324),
.B(n_224),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_356),
.B(n_364),
.Y(n_386)
);

AO22x1_ASAP7_75t_SL g357 ( 
.A1(n_279),
.A2(n_289),
.B1(n_283),
.B2(n_305),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_276),
.B(n_304),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_359),
.A2(n_365),
.B1(n_297),
.B2(n_300),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_311),
.B(n_276),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_360),
.B(n_363),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_306),
.A2(n_291),
.B(n_302),
.Y(n_361)
);

OR2x2_ASAP7_75t_L g378 ( 
.A(n_361),
.B(n_275),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_277),
.B(n_316),
.C(n_305),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_303),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_291),
.A2(n_316),
.B1(n_299),
.B2(n_287),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_287),
.B(n_282),
.C(n_293),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_366),
.B(n_292),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_359),
.A2(n_320),
.B1(n_293),
.B2(n_280),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_367),
.A2(n_370),
.B1(n_373),
.B2(n_381),
.Y(n_401)
);

AO21x1_ASAP7_75t_L g404 ( 
.A1(n_368),
.A2(n_391),
.B(n_347),
.Y(n_404)
);

INVx13_ASAP7_75t_L g369 ( 
.A(n_347),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_369),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_343),
.A2(n_280),
.B1(n_309),
.B2(n_319),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_341),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_371),
.B(n_388),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_372),
.A2(n_380),
.B1(n_348),
.B2(n_354),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_349),
.A2(n_309),
.B1(n_319),
.B2(n_315),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_378),
.A2(n_393),
.B(n_379),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_379),
.B(n_398),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_351),
.A2(n_319),
.B1(n_315),
.B2(n_309),
.Y(n_380)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_328),
.Y(n_383)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_383),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_342),
.A2(n_322),
.B1(n_292),
.B2(n_317),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_385),
.A2(n_389),
.B1(n_346),
.B2(n_330),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g389 ( 
.A1(n_336),
.A2(n_322),
.B1(n_285),
.B2(n_325),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_353),
.A2(n_329),
.B(n_338),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_341),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_394),
.B(n_376),
.Y(n_416)
);

A2O1A1O1Ixp25_ASAP7_75t_L g407 ( 
.A1(n_397),
.A2(n_355),
.B(n_362),
.C(n_360),
.D(n_332),
.Y(n_407)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_344),
.Y(n_399)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_399),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_368),
.A2(n_357),
.B1(n_340),
.B2(n_337),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_400),
.A2(n_419),
.B1(n_421),
.B2(n_379),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_371),
.B(n_394),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_403),
.B(n_415),
.Y(n_428)
);

INVx1_ASAP7_75t_SL g432 ( 
.A(n_404),
.Y(n_432)
);

XNOR2x1_ASAP7_75t_L g406 ( 
.A(n_390),
.B(n_364),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_406),
.B(n_409),
.C(n_411),
.Y(n_437)
);

OA21x2_ASAP7_75t_SL g441 ( 
.A1(n_407),
.A2(n_397),
.B(n_374),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_390),
.B(n_366),
.C(n_333),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_386),
.B(n_361),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_412),
.B(n_381),
.Y(n_429)
);

MAJx2_ASAP7_75t_L g413 ( 
.A(n_386),
.B(n_332),
.C(n_356),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_413),
.B(n_417),
.Y(n_447)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_383),
.Y(n_414)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_414),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_387),
.B(n_339),
.Y(n_415)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_416),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_388),
.B(n_395),
.C(n_387),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_389),
.A2(n_357),
.B1(n_336),
.B2(n_345),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_418),
.A2(n_391),
.B1(n_372),
.B2(n_396),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_393),
.A2(n_357),
.B1(n_365),
.B2(n_347),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_398),
.A2(n_369),
.B(n_391),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_420),
.A2(n_427),
.B(n_391),
.Y(n_434)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_376),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_422),
.B(n_375),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_395),
.B(n_331),
.C(n_339),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_423),
.B(n_385),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_374),
.B(n_327),
.Y(n_424)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_424),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_425),
.A2(n_378),
.B(n_375),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_369),
.A2(n_391),
.B(n_378),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_429),
.A2(n_419),
.B1(n_400),
.B2(n_426),
.Y(n_457)
);

CKINVDCx16_ASAP7_75t_R g430 ( 
.A(n_416),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_430),
.B(n_431),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_410),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_410),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_433),
.Y(n_459)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_434),
.Y(n_453)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_425),
.Y(n_435)
);

NAND2xp33_ASAP7_75t_SL g470 ( 
.A(n_435),
.B(n_436),
.Y(n_470)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_438),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_420),
.A2(n_391),
.B(n_382),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_439),
.B(n_448),
.Y(n_465)
);

XNOR2x1_ASAP7_75t_L g463 ( 
.A(n_441),
.B(n_442),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_403),
.B(n_382),
.Y(n_443)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_443),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_444),
.A2(n_445),
.B1(n_450),
.B2(n_452),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_418),
.A2(n_396),
.B1(n_397),
.B2(n_380),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_424),
.B(n_367),
.Y(n_448)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_405),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_451),
.B(n_413),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_404),
.A2(n_377),
.B1(n_384),
.B2(n_392),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_437),
.B(n_409),
.C(n_406),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_455),
.B(n_456),
.C(n_472),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_437),
.B(n_417),
.C(n_411),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_457),
.A2(n_458),
.B1(n_464),
.B2(n_442),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_444),
.A2(n_426),
.B1(n_410),
.B2(n_415),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_445),
.A2(n_427),
.B1(n_401),
.B2(n_423),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_447),
.B(n_408),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_466),
.B(n_467),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_447),
.B(n_407),
.Y(n_467)
);

NOR3xp33_ASAP7_75t_SL g468 ( 
.A(n_449),
.B(n_405),
.C(n_377),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_468),
.B(n_430),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_447),
.B(n_401),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_469),
.B(n_471),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_437),
.B(n_370),
.Y(n_472)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_473),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_466),
.B(n_451),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_475),
.B(n_477),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_472),
.B(n_435),
.C(n_441),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_478),
.B(n_482),
.Y(n_499)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_468),
.Y(n_479)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_479),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_462),
.A2(n_452),
.B1(n_429),
.B2(n_432),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_480),
.A2(n_485),
.B1(n_487),
.B2(n_464),
.Y(n_495)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_460),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_481),
.B(n_483),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_456),
.B(n_433),
.C(n_431),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_459),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_469),
.B(n_436),
.C(n_432),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_484),
.B(n_467),
.C(n_463),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_459),
.A2(n_432),
.B1(n_449),
.B2(n_446),
.Y(n_485)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_461),
.Y(n_487)
);

CKINVDCx16_ASAP7_75t_R g489 ( 
.A(n_485),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_489),
.B(n_495),
.Y(n_502)
);

AO22x1_ASAP7_75t_L g491 ( 
.A1(n_483),
.A2(n_453),
.B1(n_446),
.B2(n_458),
.Y(n_491)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_491),
.Y(n_503)
);

A2O1A1Ixp33_ASAP7_75t_SL g492 ( 
.A1(n_477),
.A2(n_434),
.B(n_439),
.C(n_470),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_492),
.B(n_496),
.C(n_498),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_476),
.B(n_455),
.C(n_463),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_497),
.B(n_486),
.Y(n_506)
);

A2O1A1Ixp33_ASAP7_75t_SL g498 ( 
.A1(n_480),
.A2(n_465),
.B(n_457),
.C(n_454),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_490),
.A2(n_450),
.B1(n_440),
.B2(n_448),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_501),
.B(n_506),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_499),
.A2(n_482),
.B(n_497),
.Y(n_504)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_504),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_496),
.B(n_476),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_505),
.B(n_507),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_494),
.B(n_474),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_493),
.B(n_428),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g514 ( 
.A1(n_508),
.A2(n_440),
.B(n_414),
.Y(n_514)
);

OAI321xp33_ASAP7_75t_L g509 ( 
.A1(n_492),
.A2(n_428),
.A3(n_443),
.B1(n_438),
.B2(n_484),
.C(n_478),
.Y(n_509)
);

AOI322xp5_ASAP7_75t_L g516 ( 
.A1(n_509),
.A2(n_498),
.A3(n_471),
.B1(n_492),
.B2(n_486),
.C1(n_474),
.C2(n_373),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_500),
.B(n_488),
.Y(n_510)
);

OR2x2_ASAP7_75t_L g523 ( 
.A(n_510),
.B(n_512),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_503),
.A2(n_491),
.B1(n_498),
.B2(n_492),
.Y(n_512)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_514),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_516),
.B(n_517),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_502),
.B(n_498),
.C(n_509),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_510),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_518),
.B(n_519),
.Y(n_526)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_515),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_513),
.B(n_508),
.C(n_402),
.Y(n_521)
);

OR2x2_ASAP7_75t_L g525 ( 
.A(n_521),
.B(n_514),
.Y(n_525)
);

NOR3xp33_ASAP7_75t_L g524 ( 
.A(n_522),
.B(n_517),
.C(n_511),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_524),
.A2(n_527),
.B(n_512),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_525),
.B(n_511),
.C(n_520),
.Y(n_528)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_523),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_SL g530 ( 
.A1(n_528),
.A2(n_529),
.B(n_526),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_530),
.B(n_402),
.C(n_392),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_531),
.A2(n_384),
.B(n_399),
.Y(n_532)
);


endmodule