module fake_aes_11108_n_39 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_39);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_39;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
NOR2x1_ASAP7_75t_L g11 ( .A(n_6), .B(n_1), .Y(n_11) );
NAND2xp33_ASAP7_75t_L g12 ( .A(n_1), .B(n_0), .Y(n_12) );
BUFx6f_ASAP7_75t_L g13 ( .A(n_2), .Y(n_13) );
AND2x2_ASAP7_75t_L g14 ( .A(n_8), .B(n_2), .Y(n_14) );
AND2x2_ASAP7_75t_L g15 ( .A(n_6), .B(n_7), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_0), .Y(n_16) );
NAND2xp33_ASAP7_75t_L g17 ( .A(n_13), .B(n_3), .Y(n_17) );
BUFx4f_ASAP7_75t_SL g18 ( .A(n_14), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_16), .B(n_3), .Y(n_19) );
AOI22xp33_ASAP7_75t_L g20 ( .A1(n_16), .A2(n_4), .B1(n_5), .B2(n_7), .Y(n_20) );
NAND2x1p5_ASAP7_75t_L g21 ( .A(n_19), .B(n_14), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_18), .B(n_14), .Y(n_22) );
OAI21x1_ASAP7_75t_SL g23 ( .A1(n_20), .A2(n_19), .B(n_11), .Y(n_23) );
AND2x2_ASAP7_75t_L g24 ( .A(n_21), .B(n_15), .Y(n_24) );
AND2x2_ASAP7_75t_L g25 ( .A(n_21), .B(n_15), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_24), .Y(n_26) );
NOR3xp33_ASAP7_75t_SL g27 ( .A(n_24), .B(n_22), .C(n_23), .Y(n_27) );
NAND3xp33_ASAP7_75t_SL g28 ( .A(n_27), .B(n_25), .C(n_12), .Y(n_28) );
OAI22xp5_ASAP7_75t_L g29 ( .A1(n_26), .A2(n_11), .B1(n_13), .B2(n_17), .Y(n_29) );
NAND3xp33_ASAP7_75t_SL g30 ( .A(n_29), .B(n_26), .C(n_5), .Y(n_30) );
INVx2_ASAP7_75t_SL g31 ( .A(n_28), .Y(n_31) );
NOR2x1_ASAP7_75t_SL g32 ( .A(n_28), .B(n_13), .Y(n_32) );
OAI22xp5_ASAP7_75t_L g33 ( .A1(n_31), .A2(n_13), .B1(n_8), .B2(n_9), .Y(n_33) );
INVx2_ASAP7_75t_L g34 ( .A(n_31), .Y(n_34) );
NAND3xp33_ASAP7_75t_L g35 ( .A(n_30), .B(n_13), .C(n_9), .Y(n_35) );
INVxp67_ASAP7_75t_L g36 ( .A(n_34), .Y(n_36) );
AOI22xp5_ASAP7_75t_L g37 ( .A1(n_33), .A2(n_13), .B1(n_32), .B2(n_4), .Y(n_37) );
INVx1_ASAP7_75t_L g38 ( .A(n_36), .Y(n_38) );
AOI22xp5_ASAP7_75t_L g39 ( .A1(n_38), .A2(n_35), .B1(n_37), .B2(n_10), .Y(n_39) );
endmodule