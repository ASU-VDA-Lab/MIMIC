module fake_jpeg_9066_n_204 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_204);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_204;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_3),
.B(n_5),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_1),
.B(n_4),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_28),
.B(n_0),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_32),
.Y(n_43)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_36),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_1),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_27),
.Y(n_47)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_27),
.Y(n_45)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_33),
.A2(n_19),
.B1(n_18),
.B2(n_21),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_39),
.A2(n_41),
.B1(n_46),
.B2(n_38),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_30),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_19),
.B1(n_18),
.B2(n_21),
.Y(n_41)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

AO22x1_ASAP7_75t_SL g46 ( 
.A1(n_34),
.A2(n_22),
.B1(n_25),
.B2(n_15),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_47),
.B(n_35),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_37),
.A2(n_19),
.B1(n_17),
.B2(n_23),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_31),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_17),
.Y(n_49)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_46),
.A2(n_36),
.B1(n_19),
.B2(n_17),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_52),
.A2(n_57),
.B1(n_51),
.B2(n_36),
.Y(n_87)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_53),
.B(n_55),
.Y(n_78)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_64),
.Y(n_86)
);

AND2x4_ASAP7_75t_SL g58 ( 
.A(n_46),
.B(n_38),
.Y(n_58)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_58),
.A2(n_60),
.B(n_61),
.C(n_69),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_59),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_SL g60 ( 
.A1(n_48),
.A2(n_34),
.B(n_38),
.C(n_30),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_32),
.Y(n_61)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_63),
.B(n_75),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_32),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_67),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_40),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_70),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_27),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_35),
.Y(n_71)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_23),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_26),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_73),
.B(n_76),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_44),
.B(n_31),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_40),
.B(n_24),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_81),
.B(n_82),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_42),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_54),
.B(n_24),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_83),
.B(n_89),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_61),
.B(n_40),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_93),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_87),
.A2(n_94),
.B1(n_95),
.B2(n_16),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_74),
.B(n_23),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_61),
.B(n_22),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_53),
.A2(n_36),
.B1(n_51),
.B2(n_39),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_58),
.A2(n_41),
.B1(n_51),
.B2(n_34),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_69),
.B(n_26),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_97),
.B(n_89),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_98),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_25),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_99),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_58),
.C(n_57),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_90),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_55),
.Y(n_102)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_104),
.Y(n_126)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_91),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_86),
.B(n_56),
.Y(n_105)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_78),
.A2(n_60),
.B1(n_72),
.B2(n_69),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_106),
.A2(n_113),
.B1(n_117),
.B2(n_84),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_26),
.Y(n_108)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_78),
.A2(n_60),
.B1(n_72),
.B2(n_34),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_109),
.A2(n_120),
.B1(n_92),
.B2(n_97),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_96),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_122),
.Y(n_135)
);

NOR4xp25_ASAP7_75t_L g112 ( 
.A(n_81),
.B(n_60),
.C(n_13),
.D(n_12),
.Y(n_112)
);

A2O1A1O1Ixp25_ASAP7_75t_L g142 ( 
.A1(n_112),
.A2(n_121),
.B(n_20),
.C(n_15),
.D(n_83),
.Y(n_142)
);

AO21x2_ASAP7_75t_L g113 ( 
.A1(n_95),
.A2(n_65),
.B(n_25),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_96),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_115),
.B(n_116),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_79),
.A2(n_16),
.B1(n_22),
.B2(n_25),
.Y(n_117)
);

INVxp33_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_80),
.Y(n_136)
);

OAI21x1_ASAP7_75t_SL g121 ( 
.A1(n_79),
.A2(n_22),
.B(n_20),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_93),
.Y(n_123)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_125),
.A2(n_140),
.B(n_142),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_118),
.B(n_90),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_133),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_128),
.B(n_114),
.C(n_122),
.Y(n_144)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_107),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_129),
.B(n_130),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_77),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_132),
.A2(n_113),
.B1(n_117),
.B2(n_109),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_118),
.B(n_121),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_136),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_107),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_137),
.B(n_139),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_113),
.A2(n_92),
.B1(n_88),
.B2(n_85),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_138),
.A2(n_104),
.B1(n_103),
.B2(n_111),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_110),
.B(n_88),
.Y(n_139)
);

AOI21x1_ASAP7_75t_L g140 ( 
.A1(n_113),
.A2(n_77),
.B(n_20),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_100),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_143),
.B(n_144),
.C(n_153),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_145),
.B(n_146),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_126),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_133),
.C(n_123),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_151),
.B(n_156),
.C(n_150),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_113),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_135),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_155),
.B(n_134),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_132),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_157),
.A2(n_124),
.B(n_141),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_140),
.A2(n_119),
.B1(n_15),
.B2(n_98),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_158),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_169)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_159),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_148),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_160),
.A2(n_165),
.B(n_168),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_138),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_162),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_129),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_163),
.B(n_153),
.Y(n_174)
);

OA21x2_ASAP7_75t_SL g164 ( 
.A1(n_150),
.A2(n_142),
.B(n_131),
.Y(n_164)
);

AOI31xp67_ASAP7_75t_L g180 ( 
.A1(n_164),
.A2(n_154),
.A3(n_144),
.B(n_13),
.Y(n_180)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_147),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_149),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_167),
.A2(n_169),
.B1(n_149),
.B2(n_152),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_151),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_161),
.B(n_170),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_177),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_173),
.B(n_174),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_166),
.A2(n_165),
.B1(n_162),
.B2(n_156),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_176),
.A2(n_159),
.B(n_4),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_161),
.B(n_143),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_179),
.B(n_168),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_180),
.A2(n_6),
.B(n_7),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_184),
.C(n_187),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_182),
.A2(n_6),
.B(n_7),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_176),
.B(n_12),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_2),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_186),
.B(n_8),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_175),
.A2(n_5),
.B(n_6),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_188),
.B(n_8),
.Y(n_191)
);

OAI221xp5_ASAP7_75t_L g189 ( 
.A1(n_184),
.A2(n_171),
.B1(n_177),
.B2(n_172),
.C(n_179),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_189),
.B(n_193),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_190),
.B(n_9),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_191),
.B(n_192),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_188),
.B(n_185),
.Y(n_192)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_196),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_194),
.B(n_183),
.C(n_10),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_197),
.Y(n_199)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_195),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_201),
.A2(n_9),
.B1(n_175),
.B2(n_200),
.Y(n_203)
);

AO22x1_ASAP7_75t_L g202 ( 
.A1(n_199),
.A2(n_198),
.B1(n_10),
.B2(n_11),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_202),
.B(n_203),
.Y(n_204)
);


endmodule