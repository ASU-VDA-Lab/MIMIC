module real_jpeg_17828_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_578;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_594;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_586;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_588;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_SL g20 ( 
.A(n_0),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_0),
.B(n_22),
.Y(n_21)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_1),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_1),
.Y(n_104)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_1),
.Y(n_460)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_2),
.Y(n_135)
);

BUFx5_ASAP7_75t_L g138 ( 
.A(n_2),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_2),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_2),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_3),
.A2(n_272),
.B1(n_273),
.B2(n_274),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_3),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_3),
.A2(n_273),
.B1(n_301),
.B2(n_304),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g470 ( 
.A1(n_3),
.A2(n_273),
.B1(n_471),
.B2(n_474),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_3),
.A2(n_273),
.B1(n_530),
.B2(n_532),
.Y(n_529)
);

OAI32xp33_ASAP7_75t_L g309 ( 
.A1(n_4),
.A2(n_310),
.A3(n_313),
.B1(n_316),
.B2(n_320),
.Y(n_309)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_4),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g375 ( 
.A1(n_4),
.A2(n_319),
.B1(n_376),
.B2(n_379),
.Y(n_375)
);

OAI32xp33_ASAP7_75t_L g397 ( 
.A1(n_4),
.A2(n_310),
.A3(n_313),
.B1(n_316),
.B2(n_320),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_4),
.B(n_27),
.Y(n_406)
);

OAI32xp33_ASAP7_75t_L g440 ( 
.A1(n_4),
.A2(n_441),
.A3(n_445),
.B1(n_449),
.B2(n_452),
.Y(n_440)
);

AOI22xp33_ASAP7_75t_SL g478 ( 
.A1(n_4),
.A2(n_310),
.B1(n_319),
.B2(n_479),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_4),
.B(n_94),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_4),
.B(n_567),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_4),
.B(n_236),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_5),
.A2(n_78),
.B1(n_79),
.B2(n_81),
.Y(n_77)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_5),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_5),
.A2(n_81),
.B1(n_165),
.B2(n_168),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_5),
.A2(n_81),
.B1(n_226),
.B2(n_230),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_5),
.A2(n_81),
.B1(n_218),
.B2(n_337),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_6),
.A2(n_70),
.B1(n_72),
.B2(n_73),
.Y(n_69)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_6),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_6),
.A2(n_73),
.B1(n_184),
.B2(n_187),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_6),
.A2(n_73),
.B1(n_265),
.B2(n_269),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g329 ( 
.A1(n_6),
.A2(n_73),
.B1(n_330),
.B2(n_331),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_7),
.A2(n_44),
.B1(n_47),
.B2(n_48),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_7),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_7),
.A2(n_47),
.B1(n_86),
.B2(n_89),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_7),
.A2(n_47),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_7),
.A2(n_47),
.B1(n_255),
.B2(n_259),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_8),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_8),
.A2(n_37),
.B1(n_121),
.B2(n_124),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_8),
.A2(n_37),
.B1(n_153),
.B2(n_155),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_8),
.A2(n_37),
.B1(n_218),
.B2(n_219),
.Y(n_217)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_9),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_9),
.Y(n_216)
);

BUFx5_ASAP7_75t_L g252 ( 
.A(n_9),
.Y(n_252)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_10),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_10),
.Y(n_102)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_10),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_10),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_10),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_10),
.Y(n_229)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_10),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g507 ( 
.A(n_10),
.Y(n_507)
);

AOI22xp33_ASAP7_75t_L g342 ( 
.A1(n_11),
.A2(n_272),
.B1(n_343),
.B2(n_344),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_11),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_SL g400 ( 
.A1(n_11),
.A2(n_343),
.B1(n_401),
.B2(n_404),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_11),
.A2(n_343),
.B1(n_519),
.B2(n_524),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g557 ( 
.A1(n_11),
.A2(n_343),
.B1(n_558),
.B2(n_562),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_13),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_14),
.A2(n_19),
.B(n_21),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_15),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_15),
.Y(n_137)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_15),
.Y(n_212)
);

BUFx4f_ASAP7_75t_L g258 ( 
.A(n_15),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_16),
.Y(n_348)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx8_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g323 ( 
.A(n_17),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_594),
.Y(n_22)
);

OAI221xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_60),
.B1(n_63),
.B2(n_292),
.C(n_588),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_24),
.B(n_60),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_25),
.B(n_291),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_25),
.B(n_291),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_42),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_26),
.A2(n_51),
.B(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_36),
.Y(n_26)
);

OR2x6_ASAP7_75t_L g51 ( 
.A(n_27),
.B(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_27),
.B(n_43),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_27),
.A2(n_50),
.B1(n_341),
.B2(n_345),
.Y(n_340)
);

AO22x2_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_30),
.B1(n_33),
.B2(n_34),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_31),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_31),
.Y(n_307)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_31),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_32),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_32),
.Y(n_126)
);

INVx2_ASAP7_75t_SL g171 ( 
.A(n_33),
.Y(n_171)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_33),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_33),
.Y(n_455)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_38),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_39),
.Y(n_274)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g344 ( 
.A(n_41),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_42),
.A2(n_61),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_50),
.Y(n_42)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_44),
.Y(n_272)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx8_ASAP7_75t_L g315 ( 
.A(n_45),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g50 ( 
.A(n_51),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_51),
.A2(n_61),
.B(n_62),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_51),
.A2(n_61),
.B1(n_69),
.B2(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_51),
.A2(n_62),
.B(n_239),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_51),
.A2(n_77),
.B(n_239),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_51),
.A2(n_61),
.B1(n_271),
.B2(n_346),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_51),
.A2(n_61),
.B1(n_342),
.B2(n_375),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_54),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_55),
.Y(n_380)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND3xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_282),
.C(n_290),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_240),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_L g589 ( 
.A1(n_65),
.A2(n_590),
.B(n_591),
.Y(n_589)
);

NOR2xp67_ASAP7_75t_SL g65 ( 
.A(n_66),
.B(n_174),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_66),
.B(n_174),
.Y(n_591)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_162),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_74),
.B1(n_75),
.B2(n_161),
.Y(n_67)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_68),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_68),
.B(n_127),
.C(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_68),
.A2(n_161),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_68),
.B(n_75),
.C(n_162),
.Y(n_283)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_82),
.Y(n_75)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_76),
.Y(n_289)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_127),
.B2(n_160),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_83),
.B(n_160),
.C(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

AO21x1_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_92),
.B(n_118),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_85),
.B(n_94),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_85),
.Y(n_277)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_88),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_90),
.Y(n_481)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_91),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_92),
.A2(n_164),
.B(n_172),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_92),
.A2(n_94),
.B1(n_164),
.B2(n_182),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_92),
.A2(n_94),
.B(n_287),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_92),
.A2(n_118),
.B(n_299),
.Y(n_298)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_93),
.A2(n_119),
.B1(n_183),
.B2(n_277),
.Y(n_276)
);

OAI21x1_ASAP7_75t_L g366 ( 
.A1(n_93),
.A2(n_120),
.B(n_173),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_93),
.A2(n_119),
.B1(n_300),
.B2(n_382),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_93),
.A2(n_119),
.B1(n_382),
.B2(n_400),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_93),
.A2(n_119),
.B1(n_400),
.B2(n_478),
.Y(n_477)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_105),
.Y(n_93)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_94),
.Y(n_119)
);

AO22x2_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_99),
.B1(n_102),
.B2(n_103),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_100),
.Y(n_197)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_102),
.Y(n_194)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_104),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_109),
.B1(n_113),
.B2(n_116),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_111),
.Y(n_167)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_120),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_120),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_123),
.Y(n_386)
);

INVxp67_ASAP7_75t_SL g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_126),
.Y(n_188)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_127),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_127),
.B(n_163),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_139),
.B(n_151),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_128),
.B(n_264),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_128),
.A2(n_139),
.B1(n_515),
.B2(n_518),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_128),
.A2(n_139),
.B1(n_465),
.B2(n_518),
.Y(n_538)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_129),
.B(n_152),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_129),
.A2(n_225),
.B1(n_234),
.B2(n_263),
.Y(n_262)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_130),
.B(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_130),
.Y(n_236)
);

OA22x2_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_134),
.B1(n_136),
.B2(n_138),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_133),
.Y(n_500)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_134),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_137),
.Y(n_218)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_137),
.Y(n_261)
);

INVx4_ASAP7_75t_L g565 ( 
.A(n_137),
.Y(n_565)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_138),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_139),
.B(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_139),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_139),
.A2(n_190),
.B(n_486),
.Y(n_485)
);

OAI22xp33_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_144),
.B1(n_145),
.B2(n_149),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_142),
.Y(n_154)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_149),
.Y(n_475)
);

BUFx12f_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_150),
.Y(n_451)
);

INVx4_ASAP7_75t_L g517 ( 
.A(n_150),
.Y(n_517)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_152),
.A2(n_234),
.B(n_235),
.Y(n_373)
);

OAI32xp33_ASAP7_75t_L g495 ( 
.A1(n_153),
.A2(n_496),
.A3(n_501),
.B1(n_505),
.B2(n_508),
.Y(n_495)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_158),
.Y(n_473)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_179),
.C(n_198),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_176),
.A2(n_179),
.B1(n_180),
.B2(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_176),
.Y(n_281)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_177),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

OAI21xp33_ASAP7_75t_L g245 ( 
.A1(n_180),
.A2(n_181),
.B(n_189),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_189),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_186),
.Y(n_303)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

INVxp33_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_192),
.B(n_363),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_193),
.B(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_198),
.A2(n_199),
.B1(n_279),
.B2(n_280),
.Y(n_278)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

AOI21xp33_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_222),
.B(n_237),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_200),
.A2(n_201),
.B1(n_237),
.B2(n_238),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_200),
.A2(n_201),
.B1(n_224),
.B2(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

NOR2x1_ASAP7_75t_R g223 ( 
.A(n_201),
.B(n_224),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_208),
.B(n_217),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_206),
.Y(n_361)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_207),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_208),
.B(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_208),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g528 ( 
.A1(n_208),
.A2(n_529),
.B(n_536),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_208),
.A2(n_319),
.B1(n_556),
.B2(n_557),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_208),
.A2(n_544),
.B1(n_557),
.B2(n_570),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_213),
.Y(n_208)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_210),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_211),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_212),
.Y(n_333)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_213),
.Y(n_556)
);

INVx6_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx4_ASAP7_75t_L g567 ( 
.A(n_215),
.Y(n_567)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_217),
.B(n_250),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_217),
.Y(n_462)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_221),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XNOR2x1_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_243),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_224),
.Y(n_416)
);

OA21x2_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_234),
.B(n_235),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx4_ASAP7_75t_L g467 ( 
.A(n_228),
.Y(n_467)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_229),
.Y(n_469)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_230),
.Y(n_269)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_233),
.Y(n_268)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_233),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_234),
.A2(n_464),
.B1(n_470),
.B2(n_476),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_236),
.Y(n_476)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_278),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_241),
.B(n_278),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_244),
.C(n_246),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_242),
.A2(n_244),
.B1(n_245),
.B2(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_242),
.Y(n_427)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_246),
.B(n_426),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_270),
.C(n_275),
.Y(n_246)
);

XNOR2x1_ASAP7_75t_L g417 ( 
.A(n_247),
.B(n_418),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_262),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g367 ( 
.A(n_248),
.B(n_262),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_253),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_249),
.Y(n_536)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_253),
.A2(n_329),
.B(n_408),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_254),
.B(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_255),
.Y(n_330)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_258),
.Y(n_547)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_258),
.Y(n_561)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_268),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_268),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_270),
.B(n_276),
.Y(n_418)
);

INVx5_ASAP7_75t_L g350 ( 
.A(n_274),
.Y(n_350)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g588 ( 
.A1(n_282),
.A2(n_290),
.B(n_589),
.C(n_592),
.D(n_593),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_283),
.B(n_284),
.Y(n_592)
);

BUFx24_ASAP7_75t_SL g595 ( 
.A(n_284),
.Y(n_595)
);

FAx1_ASAP7_75t_SL g284 ( 
.A(n_285),
.B(n_286),
.CI(n_288),
.CON(n_284),
.SN(n_284)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_285),
.B(n_286),
.C(n_288),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_429),
.Y(n_293)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g294 ( 
.A1(n_295),
.A2(n_411),
.B(n_420),
.C(n_421),
.D(n_428),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_369),
.C(n_391),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_296),
.B(n_369),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_352),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_297),
.B(n_353),
.C(n_368),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_308),
.C(n_340),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_298),
.B(n_340),
.Y(n_371)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx3_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_308),
.B(n_371),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_327),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx8_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_319),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g449 ( 
.A(n_319),
.B(n_450),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_319),
.B(n_506),
.Y(n_505)
);

OAI21xp33_ASAP7_75t_SL g515 ( 
.A1(n_319),
.A2(n_505),
.B(n_516),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_324),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx4_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_327),
.B(n_397),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_328),
.A2(n_329),
.B1(n_334),
.B2(n_336),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_328),
.A2(n_336),
.B(n_357),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_328),
.A2(n_357),
.B(n_462),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_328),
.A2(n_334),
.B1(n_543),
.B2(n_550),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_332),
.Y(n_562)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_333),
.Y(n_512)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_333),
.Y(n_535)
);

INVx6_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx4_ASAP7_75t_L g347 ( 
.A(n_344),
.Y(n_347)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_347),
.A2(n_348),
.B1(n_349),
.B2(n_351),
.Y(n_346)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_348),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_SL g382 ( 
.A1(n_348),
.A2(n_351),
.B1(n_383),
.B2(n_387),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_348),
.A2(n_351),
.B1(n_466),
.B2(n_468),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_348),
.A2(n_351),
.B1(n_545),
.B2(n_548),
.Y(n_544)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g352 ( 
.A1(n_353),
.A2(n_354),
.B1(n_367),
.B2(n_368),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_364),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_355),
.B(n_365),
.C(n_366),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_362),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_356),
.B(n_362),
.Y(n_390)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx4_ASAP7_75t_SL g408 ( 
.A(n_361),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_366),
.Y(n_364)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_367),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_372),
.C(n_390),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_370),
.B(n_410),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_372),
.B(n_390),
.Y(n_410)
);

MAJx2_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_374),
.C(n_381),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_373),
.B(n_381),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_374),
.B(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_385),
.Y(n_403)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_386),
.Y(n_404)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_409),
.Y(n_391)
);

OR2x2_ASAP7_75t_L g433 ( 
.A(n_392),
.B(n_409),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_395),
.C(n_398),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_393),
.B(n_584),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_SL g584 ( 
.A1(n_395),
.A2(n_396),
.B1(n_398),
.B2(n_585),
.Y(n_584)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_398),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_405),
.C(n_407),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_SL g488 ( 
.A(n_399),
.B(n_489),
.Y(n_488)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_406),
.B(n_407),
.Y(n_489)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_411),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_413),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_412),
.B(n_413),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_419),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_417),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_415),
.B(n_417),
.C(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_419),
.Y(n_424)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

NOR3xp33_ASAP7_75t_L g430 ( 
.A(n_422),
.B(n_431),
.C(n_434),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_425),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_423),
.B(n_425),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_435),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_432),
.B(n_433),
.Y(n_431)
);

OAI21x1_ASAP7_75t_L g435 ( 
.A1(n_436),
.A2(n_582),
.B(n_587),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_437),
.A2(n_491),
.B(n_581),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_482),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_SL g581 ( 
.A(n_438),
.B(n_482),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_439),
.B(n_463),
.C(n_477),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g577 ( 
.A(n_439),
.B(n_578),
.Y(n_577)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_461),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_440),
.B(n_461),
.Y(n_484)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_456),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_463),
.B(n_477),
.Y(n_578)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx4_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_470),
.Y(n_486)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx8_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_483),
.A2(n_487),
.B1(n_488),
.B2(n_490),
.Y(n_482)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_483),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_485),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g586 ( 
.A(n_484),
.B(n_485),
.C(n_487),
.Y(n_586)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_492),
.A2(n_576),
.B(n_580),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_493),
.A2(n_540),
.B(n_575),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_527),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_494),
.B(n_527),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_513),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_495),
.A2(n_513),
.B1(n_514),
.B2(n_552),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_495),
.Y(n_552)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

BUFx2_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

BUFx2_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx8_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_509),
.B(n_510),
.Y(n_508)
);

BUFx2_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

BUFx2_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_528),
.B(n_537),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_528),
.B(n_538),
.C(n_539),
.Y(n_579)
);

INVxp67_ASAP7_75t_L g550 ( 
.A(n_529),
.Y(n_550)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_538),
.B(n_539),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_SL g540 ( 
.A1(n_541),
.A2(n_553),
.B(n_574),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_542),
.B(n_551),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_542),
.B(n_551),
.Y(n_574)
);

INVxp67_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

INVx1_ASAP7_75t_SL g545 ( 
.A(n_546),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

BUFx2_ASAP7_75t_L g549 ( 
.A(n_547),
.Y(n_549)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_554),
.A2(n_568),
.B(n_573),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_555),
.B(n_563),
.Y(n_554)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_559),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_564),
.B(n_566),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_565),
.Y(n_564)
);

INVx5_ASAP7_75t_L g571 ( 
.A(n_567),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_569),
.B(n_572),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_569),
.B(n_572),
.Y(n_573)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_571),
.Y(n_570)
);

NOR2xp67_ASAP7_75t_SL g576 ( 
.A(n_577),
.B(n_579),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_577),
.B(n_579),
.Y(n_580)
);

NOR2xp67_ASAP7_75t_SL g582 ( 
.A(n_583),
.B(n_586),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_583),
.B(n_586),
.Y(n_587)
);


endmodule