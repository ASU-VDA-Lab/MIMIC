module fake_netlist_6_2909_n_595 (n_52, n_16, n_1, n_91, n_119, n_46, n_18, n_21, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_127, n_125, n_77, n_106, n_92, n_42, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_17, n_23, n_20, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_122, n_45, n_34, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_41, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_595);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_18;
input n_21;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_127;
input n_125;
input n_77;
input n_106;
input n_92;
input n_42;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_17;
input n_23;
input n_20;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_122;
input n_45;
input n_34;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_41;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_595;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_507;
wire n_580;
wire n_209;
wire n_367;
wire n_465;
wire n_590;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_148;
wire n_226;
wire n_208;
wire n_161;
wire n_462;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_578;
wire n_144;
wire n_365;
wire n_168;
wire n_384;
wire n_297;
wire n_524;
wire n_342;
wire n_358;
wire n_160;
wire n_449;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_142;
wire n_143;
wire n_382;
wire n_180;
wire n_557;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_400;
wire n_140;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_327;
wire n_369;
wire n_280;
wire n_287;
wire n_353;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_461;
wire n_141;
wire n_383;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_222;
wire n_179;
wire n_248;
wire n_300;
wire n_517;
wire n_229;
wire n_542;
wire n_305;
wire n_532;
wire n_173;
wire n_535;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_183;
wire n_510;
wire n_375;
wire n_338;
wire n_522;
wire n_466;
wire n_506;
wire n_360;
wire n_235;
wire n_536;
wire n_147;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_344;
wire n_581;
wire n_428;
wire n_432;
wire n_167;
wire n_174;
wire n_516;
wire n_153;
wire n_525;
wire n_156;
wire n_491;
wire n_145;
wire n_133;
wire n_371;
wire n_567;
wire n_189;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_197;
wire n_137;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_155;
wire n_529;
wire n_445;
wire n_425;
wire n_454;
wire n_218;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_172;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_196;
wire n_402;
wire n_352;
wire n_478;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_374;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_185;
wire n_348;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_163;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_154;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_279;
wire n_252;
wire n_228;
wire n_565;
wire n_594;
wire n_356;
wire n_577;
wire n_166;
wire n_184;
wire n_552;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_323;
wire n_393;
wire n_411;
wire n_503;
wire n_152;
wire n_513;
wire n_321;
wire n_331;
wire n_227;
wire n_570;
wire n_406;
wire n_483;
wire n_204;
wire n_482;
wire n_474;
wire n_527;
wire n_261;
wire n_420;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_164;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_150;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_505;
wire n_240;
wire n_139;
wire n_319;
wire n_134;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_311;
wire n_403;
wire n_253;
wire n_583;
wire n_136;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_159;
wire n_157;
wire n_162;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_560;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_146;
wire n_318;
wire n_303;
wire n_511;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_582;
wire n_199;
wire n_138;
wire n_266;
wire n_296;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_439;
wire n_158;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_453;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_149;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_251;
wire n_301;
wire n_274;
wire n_151;
wire n_412;
wire n_267;
wire n_438;
wire n_339;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_422;
wire n_135;
wire n_165;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_528;
wire n_391;
wire n_457;
wire n_364;
wire n_385;
wire n_295;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_379;
wire n_170;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_194;
wire n_171;
wire n_192;
wire n_169;
wire n_283;

INVx1_ASAP7_75t_L g133 ( 
.A(n_53),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_18),
.Y(n_134)
);

CKINVDCx5p33_ASAP7_75t_R g135 ( 
.A(n_46),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_42),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_15),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_25),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_30),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_88),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_49),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_72),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_78),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_22),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_55),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_15),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_57),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_97),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_104),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_69),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_92),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_87),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_8),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_40),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_41),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_76),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_26),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_115),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_52),
.Y(n_161)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_77),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_24),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_64),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_93),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_27),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_81),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_131),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_14),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_91),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_94),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_28),
.Y(n_172)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_10),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_84),
.Y(n_174)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_32),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_43),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_23),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_111),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_100),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_85),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_107),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_127),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_2),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_126),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_51),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_122),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_70),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_99),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_38),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_83),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_110),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_39),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_128),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_50),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_137),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_169),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_148),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_183),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_162),
.B(n_0),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_138),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_138),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_167),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_194),
.B(n_1),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_135),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_133),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_140),
.Y(n_206)
);

NOR2xp67_ASAP7_75t_L g207 ( 
.A(n_134),
.B(n_1),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_141),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_142),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_175),
.B(n_2),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_144),
.Y(n_211)
);

INVxp67_ASAP7_75t_SL g212 ( 
.A(n_146),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_151),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_143),
.Y(n_214)
);

INVxp67_ASAP7_75t_SL g215 ( 
.A(n_152),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_167),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_136),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_139),
.B(n_147),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_136),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_154),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_168),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_170),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_145),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_155),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_149),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_150),
.Y(n_226)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_139),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_153),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_173),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_156),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_147),
.B(n_3),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_174),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_180),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_179),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_178),
.B(n_3),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_157),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_227),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_217),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_227),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_224),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_197),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_4),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_223),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_205),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_227),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_208),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_212),
.B(n_134),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_219),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_195),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_196),
.Y(n_250)
);

BUFx8_ASAP7_75t_L g251 ( 
.A(n_211),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_213),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_220),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_235),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_228),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_221),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_219),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_215),
.B(n_171),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_222),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_197),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_232),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_230),
.A2(n_178),
.B1(n_177),
.B2(n_181),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_234),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_233),
.Y(n_264)
);

OA21x2_ASAP7_75t_L g265 ( 
.A1(n_218),
.A2(n_189),
.B(n_192),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_204),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_229),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_231),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_198),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_210),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_199),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_206),
.B(n_158),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_200),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_203),
.Y(n_274)
);

AND2x4_ASAP7_75t_L g275 ( 
.A(n_207),
.B(n_180),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_209),
.Y(n_276)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_200),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_214),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_201),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_236),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_225),
.Y(n_281)
);

AND2x4_ASAP7_75t_L g282 ( 
.A(n_225),
.B(n_180),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_226),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_226),
.Y(n_284)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_240),
.B(n_198),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_201),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_202),
.Y(n_287)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_237),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_244),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_202),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g291 ( 
.A1(n_268),
.A2(n_180),
.B1(n_182),
.B2(n_187),
.Y(n_291)
);

AO21x2_ASAP7_75t_L g292 ( 
.A1(n_272),
.A2(n_216),
.B(n_193),
.Y(n_292)
);

AND2x4_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_159),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_246),
.Y(n_294)
);

AND2x6_ASAP7_75t_L g295 ( 
.A(n_282),
.B(n_182),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_256),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_278),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_259),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_216),
.Y(n_299)
);

AND2x6_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_182),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_280),
.B(n_191),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g302 ( 
.A(n_254),
.Y(n_302)
);

INVx2_ASAP7_75t_SL g303 ( 
.A(n_277),
.Y(n_303)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_237),
.Y(n_304)
);

AND2x6_ASAP7_75t_L g305 ( 
.A(n_276),
.B(n_182),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_L g306 ( 
.A1(n_268),
.A2(n_187),
.B1(n_188),
.B2(n_190),
.Y(n_306)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_239),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_264),
.B(n_274),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_L g309 ( 
.A1(n_270),
.A2(n_187),
.B1(n_186),
.B2(n_185),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_258),
.B(n_160),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_261),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_255),
.B(n_161),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_263),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_249),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_249),
.Y(n_315)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_239),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_270),
.A2(n_166),
.B1(n_184),
.B2(n_176),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_276),
.B(n_163),
.Y(n_318)
);

INVx2_ASAP7_75t_SL g319 ( 
.A(n_277),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_274),
.B(n_164),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_254),
.B(n_187),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_250),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_252),
.Y(n_323)
);

INVx5_ASAP7_75t_L g324 ( 
.A(n_254),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_254),
.B(n_165),
.Y(n_325)
);

OR2x6_ASAP7_75t_L g326 ( 
.A(n_281),
.B(n_4),
.Y(n_326)
);

OA22x2_ASAP7_75t_L g327 ( 
.A1(n_271),
.A2(n_172),
.B1(n_6),
.B2(n_7),
.Y(n_327)
);

AND2x4_ASAP7_75t_L g328 ( 
.A(n_247),
.B(n_19),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_253),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_254),
.B(n_132),
.Y(n_330)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_253),
.Y(n_331)
);

AND2x6_ASAP7_75t_L g332 ( 
.A(n_274),
.B(n_20),
.Y(n_332)
);

OR2x2_ASAP7_75t_L g333 ( 
.A(n_267),
.B(n_5),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g334 ( 
.A(n_273),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_245),
.Y(n_335)
);

INVx2_ASAP7_75t_SL g336 ( 
.A(n_277),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_245),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_281),
.B(n_6),
.Y(n_338)
);

BUFx3_ASAP7_75t_L g339 ( 
.A(n_266),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_266),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_265),
.B(n_247),
.Y(n_341)
);

INVx4_ASAP7_75t_L g342 ( 
.A(n_275),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_283),
.B(n_284),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_284),
.B(n_8),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_288),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_325),
.A2(n_265),
.B(n_275),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_328),
.B(n_265),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_328),
.B(n_265),
.Y(n_348)
);

INVxp67_ASAP7_75t_SL g349 ( 
.A(n_302),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_288),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_302),
.B(n_275),
.Y(n_351)
);

BUFx12f_ASAP7_75t_L g352 ( 
.A(n_297),
.Y(n_352)
);

AND2x6_ASAP7_75t_SL g353 ( 
.A(n_286),
.B(n_242),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_302),
.B(n_278),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_290),
.B(n_241),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_304),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_332),
.Y(n_357)
);

NOR2xp67_ASAP7_75t_SL g358 ( 
.A(n_324),
.B(n_260),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_314),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_299),
.B(n_269),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_299),
.B(n_310),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_L g362 ( 
.A1(n_327),
.A2(n_262),
.B1(n_242),
.B2(n_251),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_285),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_L g364 ( 
.A1(n_327),
.A2(n_251),
.B1(n_273),
.B2(n_257),
.Y(n_364)
);

INVx2_ASAP7_75t_SL g365 ( 
.A(n_293),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_315),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_318),
.B(n_251),
.Y(n_367)
);

NAND2xp33_ASAP7_75t_SL g368 ( 
.A(n_309),
.B(n_306),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_324),
.B(n_21),
.Y(n_369)
);

OR2x6_ASAP7_75t_L g370 ( 
.A(n_326),
.B(n_243),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_324),
.B(n_29),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_324),
.B(n_31),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_303),
.B(n_255),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_342),
.B(n_33),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_287),
.B(n_238),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_342),
.B(n_34),
.Y(n_376)
);

INVx2_ASAP7_75t_SL g377 ( 
.A(n_293),
.Y(n_377)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_326),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_322),
.Y(n_379)
);

OR2x2_ASAP7_75t_L g380 ( 
.A(n_334),
.B(n_9),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_325),
.B(n_35),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_343),
.B(n_9),
.Y(n_382)
);

AOI22xp33_ASAP7_75t_L g383 ( 
.A1(n_341),
.A2(n_257),
.B1(n_248),
.B2(n_238),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_301),
.B(n_36),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_319),
.B(n_336),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_341),
.A2(n_248),
.B(n_71),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_309),
.B(n_11),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_289),
.B(n_73),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_339),
.B(n_11),
.Y(n_389)
);

OR2x2_ASAP7_75t_L g390 ( 
.A(n_334),
.B(n_308),
.Y(n_390)
);

OR2x2_ASAP7_75t_L g391 ( 
.A(n_333),
.B(n_12),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_306),
.B(n_12),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_296),
.B(n_74),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_298),
.B(n_75),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_311),
.B(n_68),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_313),
.B(n_79),
.Y(n_396)
);

INVx2_ASAP7_75t_SL g397 ( 
.A(n_340),
.Y(n_397)
);

OR2x6_ASAP7_75t_L g398 ( 
.A(n_326),
.B(n_13),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_344),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_321),
.B(n_67),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_321),
.B(n_80),
.Y(n_401)
);

NOR2xp67_ASAP7_75t_L g402 ( 
.A(n_312),
.B(n_130),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_294),
.Y(n_403)
);

NAND2x1_ASAP7_75t_L g404 ( 
.A(n_332),
.B(n_66),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g405 ( 
.A(n_344),
.Y(n_405)
);

CKINVDCx8_ASAP7_75t_R g406 ( 
.A(n_353),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_360),
.B(n_292),
.Y(n_407)
);

INVx6_ASAP7_75t_L g408 ( 
.A(n_352),
.Y(n_408)
);

INVx4_ASAP7_75t_L g409 ( 
.A(n_357),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_399),
.B(n_292),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_363),
.B(n_317),
.Y(n_411)
);

NAND2xp33_ASAP7_75t_SL g412 ( 
.A(n_367),
.B(n_338),
.Y(n_412)
);

BUFx2_ASAP7_75t_L g413 ( 
.A(n_370),
.Y(n_413)
);

NAND3xp33_ASAP7_75t_SL g414 ( 
.A(n_383),
.B(n_317),
.C(n_291),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_405),
.B(n_330),
.Y(n_415)
);

NOR3xp33_ASAP7_75t_SL g416 ( 
.A(n_355),
.B(n_320),
.C(n_330),
.Y(n_416)
);

INVx2_ASAP7_75t_SL g417 ( 
.A(n_390),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_359),
.Y(n_418)
);

O2A1O1Ixp33_ASAP7_75t_L g419 ( 
.A1(n_387),
.A2(n_392),
.B(n_386),
.C(n_399),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_363),
.B(n_323),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_361),
.B(n_329),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_405),
.B(n_335),
.Y(n_422)
);

NAND3xp33_ASAP7_75t_L g423 ( 
.A(n_368),
.B(n_331),
.C(n_291),
.Y(n_423)
);

INVx2_ASAP7_75t_SL g424 ( 
.A(n_380),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_366),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_379),
.Y(n_426)
);

NAND2x1p5_ASAP7_75t_L g427 ( 
.A(n_357),
.B(n_316),
.Y(n_427)
);

INVxp33_ASAP7_75t_SL g428 ( 
.A(n_375),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_397),
.B(n_337),
.Y(n_429)
);

BUFx2_ASAP7_75t_L g430 ( 
.A(n_370),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_403),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_347),
.B(n_316),
.Y(n_432)
);

INVx3_ASAP7_75t_SL g433 ( 
.A(n_370),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_348),
.B(n_307),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_354),
.Y(n_435)
);

BUFx10_ASAP7_75t_L g436 ( 
.A(n_382),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_373),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_357),
.Y(n_438)
);

BUFx4f_ASAP7_75t_L g439 ( 
.A(n_398),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_R g440 ( 
.A(n_365),
.B(n_300),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_R g441 ( 
.A(n_377),
.B(n_300),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_378),
.B(n_385),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_357),
.Y(n_443)
);

NOR2x1_ASAP7_75t_SL g444 ( 
.A(n_443),
.B(n_381),
.Y(n_444)
);

AO31x2_ASAP7_75t_L g445 ( 
.A1(n_407),
.A2(n_346),
.A3(n_382),
.B(n_400),
.Y(n_445)
);

OAI21x1_ASAP7_75t_L g446 ( 
.A1(n_432),
.A2(n_374),
.B(n_376),
.Y(n_446)
);

OAI21x1_ASAP7_75t_L g447 ( 
.A1(n_432),
.A2(n_401),
.B(n_351),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g448 ( 
.A1(n_434),
.A2(n_349),
.B(n_384),
.Y(n_448)
);

NOR2x1_ASAP7_75t_SL g449 ( 
.A(n_443),
.B(n_388),
.Y(n_449)
);

OAI21x1_ASAP7_75t_L g450 ( 
.A1(n_434),
.A2(n_369),
.B(n_371),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_415),
.A2(n_372),
.B(n_393),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g452 ( 
.A1(n_415),
.A2(n_394),
.B(n_395),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_425),
.Y(n_453)
);

HAxp5_ASAP7_75t_L g454 ( 
.A(n_406),
.B(n_383),
.CON(n_454),
.SN(n_454)
);

BUFx2_ASAP7_75t_L g455 ( 
.A(n_413),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_419),
.A2(n_396),
.B(n_404),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_421),
.A2(n_356),
.B(n_345),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_422),
.B(n_364),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_423),
.A2(n_410),
.B(n_411),
.Y(n_459)
);

OAI21x1_ASAP7_75t_L g460 ( 
.A1(n_427),
.A2(n_350),
.B(n_304),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_418),
.Y(n_461)
);

AOI221xp5_ASAP7_75t_L g462 ( 
.A1(n_414),
.A2(n_362),
.B1(n_364),
.B2(n_389),
.C(n_391),
.Y(n_462)
);

OAI21x1_ASAP7_75t_L g463 ( 
.A1(n_427),
.A2(n_378),
.B(n_332),
.Y(n_463)
);

OAI21x1_ASAP7_75t_L g464 ( 
.A1(n_431),
.A2(n_332),
.B(n_358),
.Y(n_464)
);

NAND2x1p5_ASAP7_75t_L g465 ( 
.A(n_409),
.B(n_402),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_424),
.Y(n_466)
);

AOI21x1_ASAP7_75t_SL g467 ( 
.A1(n_410),
.A2(n_332),
.B(n_305),
.Y(n_467)
);

BUFx2_ASAP7_75t_L g468 ( 
.A(n_430),
.Y(n_468)
);

O2A1O1Ixp5_ASAP7_75t_L g469 ( 
.A1(n_412),
.A2(n_305),
.B(n_300),
.C(n_295),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_426),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_409),
.Y(n_471)
);

NOR4xp25_ASAP7_75t_L g472 ( 
.A(n_422),
.B(n_362),
.C(n_398),
.D(n_16),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_461),
.B(n_438),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_458),
.B(n_428),
.Y(n_474)
);

OAI21x1_ASAP7_75t_L g475 ( 
.A1(n_467),
.A2(n_429),
.B(n_420),
.Y(n_475)
);

AOI221xp5_ASAP7_75t_L g476 ( 
.A1(n_472),
.A2(n_435),
.B1(n_417),
.B2(n_442),
.C(n_437),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_459),
.B(n_443),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g478 ( 
.A(n_455),
.Y(n_478)
);

OAI21x1_ASAP7_75t_L g479 ( 
.A1(n_467),
.A2(n_416),
.B(n_436),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_453),
.B(n_436),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_470),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_462),
.A2(n_439),
.B1(n_398),
.B2(n_433),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_468),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_466),
.Y(n_484)
);

OAI21x1_ASAP7_75t_L g485 ( 
.A1(n_447),
.A2(n_441),
.B(n_440),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_463),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_460),
.Y(n_487)
);

OA21x2_ASAP7_75t_L g488 ( 
.A1(n_446),
.A2(n_305),
.B(n_295),
.Y(n_488)
);

OA21x2_ASAP7_75t_L g489 ( 
.A1(n_448),
.A2(n_305),
.B(n_295),
.Y(n_489)
);

OA21x2_ASAP7_75t_L g490 ( 
.A1(n_448),
.A2(n_305),
.B(n_295),
.Y(n_490)
);

OAI21x1_ASAP7_75t_L g491 ( 
.A1(n_450),
.A2(n_300),
.B(n_89),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_471),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_471),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_454),
.B(n_408),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_457),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_474),
.B(n_465),
.Y(n_496)
);

AOI22xp33_ASAP7_75t_L g497 ( 
.A1(n_476),
.A2(n_456),
.B1(n_452),
.B2(n_457),
.Y(n_497)
);

INVx8_ASAP7_75t_L g498 ( 
.A(n_473),
.Y(n_498)
);

AO31x2_ASAP7_75t_L g499 ( 
.A1(n_495),
.A2(n_456),
.A3(n_451),
.B(n_444),
.Y(n_499)
);

OAI221xp5_ASAP7_75t_L g500 ( 
.A1(n_476),
.A2(n_451),
.B1(n_408),
.B2(n_469),
.C(n_445),
.Y(n_500)
);

AOI22xp33_ASAP7_75t_L g501 ( 
.A1(n_482),
.A2(n_464),
.B1(n_445),
.B2(n_18),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_481),
.Y(n_502)
);

OAI22xp33_ASAP7_75t_L g503 ( 
.A1(n_484),
.A2(n_449),
.B1(n_445),
.B2(n_16),
.Y(n_503)
);

BUFx2_ASAP7_75t_L g504 ( 
.A(n_478),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g505 ( 
.A(n_478),
.Y(n_505)
);

OA21x2_ASAP7_75t_L g506 ( 
.A1(n_491),
.A2(n_17),
.B(n_37),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_480),
.B(n_17),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g508 ( 
.A1(n_483),
.A2(n_44),
.B1(n_45),
.B2(n_47),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_483),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_494),
.B(n_48),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_481),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_495),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_492),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_L g514 ( 
.A1(n_477),
.A2(n_129),
.B1(n_56),
.B2(n_58),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_L g515 ( 
.A1(n_473),
.A2(n_54),
.B1(n_59),
.B2(n_60),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_473),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_493),
.B(n_125),
.Y(n_517)
);

NOR2xp67_ASAP7_75t_L g518 ( 
.A(n_492),
.B(n_61),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_492),
.Y(n_519)
);

AND2x4_ASAP7_75t_L g520 ( 
.A(n_504),
.B(n_479),
.Y(n_520)
);

AOI33xp33_ASAP7_75t_L g521 ( 
.A1(n_497),
.A2(n_486),
.A3(n_487),
.B1(n_479),
.B2(n_475),
.B3(n_86),
.Y(n_521)
);

NAND2x1_ASAP7_75t_L g522 ( 
.A(n_512),
.B(n_487),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g523 ( 
.A1(n_496),
.A2(n_487),
.B1(n_490),
.B2(n_489),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_L g524 ( 
.A1(n_514),
.A2(n_507),
.B1(n_510),
.B2(n_515),
.Y(n_524)
);

NAND4xp25_ASAP7_75t_L g525 ( 
.A(n_507),
.B(n_491),
.C(n_63),
.D(n_65),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_502),
.Y(n_526)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_497),
.A2(n_485),
.B(n_489),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_509),
.B(n_62),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_505),
.B(n_82),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_516),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g531 ( 
.A1(n_514),
.A2(n_490),
.B1(n_489),
.B2(n_488),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_501),
.A2(n_90),
.B1(n_95),
.B2(n_96),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_500),
.A2(n_98),
.B1(n_101),
.B2(n_105),
.Y(n_533)
);

OAI222xp33_ASAP7_75t_L g534 ( 
.A1(n_508),
.A2(n_106),
.B1(n_108),
.B2(n_109),
.C1(n_112),
.C2(n_113),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_501),
.A2(n_114),
.B1(n_116),
.B2(n_117),
.Y(n_535)
);

OAI322xp33_ASAP7_75t_L g536 ( 
.A1(n_503),
.A2(n_118),
.A3(n_119),
.B1(n_120),
.B2(n_121),
.C1(n_123),
.C2(n_124),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_L g537 ( 
.A1(n_517),
.A2(n_516),
.B1(n_511),
.B2(n_498),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_526),
.Y(n_538)
);

OR2x2_ASAP7_75t_L g539 ( 
.A(n_523),
.B(n_499),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_520),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_520),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_522),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_524),
.B(n_513),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_530),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_521),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_530),
.B(n_537),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_529),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_531),
.Y(n_548)
);

HB1xp67_ASAP7_75t_L g549 ( 
.A(n_525),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_527),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_544),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_538),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_540),
.Y(n_553)
);

AOI211xp5_ASAP7_75t_SL g554 ( 
.A1(n_549),
.A2(n_536),
.B(n_534),
.C(n_535),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_544),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_547),
.B(n_528),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_541),
.Y(n_557)
);

CKINVDCx14_ASAP7_75t_R g558 ( 
.A(n_547),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_557),
.B(n_548),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_552),
.B(n_548),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_552),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_555),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_558),
.B(n_547),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_553),
.B(n_551),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_553),
.B(n_550),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_561),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_560),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_565),
.B(n_555),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_562),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_564),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_567),
.B(n_556),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_566),
.Y(n_572)
);

OR2x2_ASAP7_75t_L g573 ( 
.A(n_568),
.B(n_559),
.Y(n_573)
);

NOR2xp67_ASAP7_75t_R g574 ( 
.A(n_570),
.B(n_545),
.Y(n_574)
);

NAND2x1_ASAP7_75t_L g575 ( 
.A(n_569),
.B(n_564),
.Y(n_575)
);

OR2x2_ASAP7_75t_L g576 ( 
.A(n_573),
.B(n_568),
.Y(n_576)
);

INVxp33_ASAP7_75t_L g577 ( 
.A(n_574),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_572),
.Y(n_578)
);

O2A1O1Ixp33_ASAP7_75t_L g579 ( 
.A1(n_577),
.A2(n_554),
.B(n_575),
.C(n_525),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_578),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_580),
.B(n_571),
.Y(n_581)
);

AND3x1_ASAP7_75t_L g582 ( 
.A(n_581),
.B(n_579),
.C(n_563),
.Y(n_582)
);

NOR3xp33_ASAP7_75t_SL g583 ( 
.A(n_582),
.B(n_532),
.C(n_546),
.Y(n_583)
);

AOI21xp5_ASAP7_75t_L g584 ( 
.A1(n_583),
.A2(n_576),
.B(n_565),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_584),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_585),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_586),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_L g588 ( 
.A1(n_587),
.A2(n_533),
.B1(n_551),
.B2(n_543),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_588),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_589),
.Y(n_590)
);

AOI22xp5_ASAP7_75t_L g591 ( 
.A1(n_590),
.A2(n_518),
.B1(n_551),
.B2(n_542),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_591),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_SL g593 ( 
.A1(n_592),
.A2(n_506),
.B1(n_516),
.B2(n_519),
.Y(n_593)
);

AOI221xp5_ASAP7_75t_L g594 ( 
.A1(n_593),
.A2(n_499),
.B1(n_519),
.B2(n_539),
.C(n_586),
.Y(n_594)
);

AOI211xp5_ASAP7_75t_L g595 ( 
.A1(n_594),
.A2(n_519),
.B(n_539),
.C(n_499),
.Y(n_595)
);


endmodule