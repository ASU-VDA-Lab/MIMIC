module fake_jpeg_30912_n_486 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_486);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_486;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_378;
wire n_132;
wire n_133;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_10),
.B(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_13),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_50),
.Y(n_103)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_56),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_31),
.B(n_15),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_57),
.B(n_87),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_31),
.A2(n_15),
.B1(n_1),
.B2(n_2),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_58),
.A2(n_49),
.B1(n_32),
.B2(n_28),
.Y(n_140)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_62),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_19),
.B(n_0),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_63),
.B(n_67),
.Y(n_116)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_64),
.Y(n_108)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_65),
.Y(n_137)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_66),
.Y(n_122)
);

HAxp5_ASAP7_75t_SL g67 ( 
.A(n_45),
.B(n_0),
.CON(n_67),
.SN(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_27),
.B(n_2),
.C(n_3),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_68),
.B(n_32),
.C(n_36),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_69),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_70),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_35),
.Y(n_71)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_71),
.Y(n_146)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_73),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_19),
.B(n_2),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_74),
.B(n_17),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_75),
.Y(n_147)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_76),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_16),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_77),
.Y(n_107)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g129 ( 
.A(n_79),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_80),
.Y(n_111)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_30),
.Y(n_81)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_82),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_83),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_84),
.Y(n_141)
);

INVx6_ASAP7_75t_SL g85 ( 
.A(n_42),
.Y(n_85)
);

CKINVDCx9p33_ASAP7_75t_R g125 ( 
.A(n_85),
.Y(n_125)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_86),
.Y(n_149)
);

INVx6_ASAP7_75t_SL g87 ( 
.A(n_47),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g135 ( 
.A(n_88),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_89),
.Y(n_142)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_21),
.Y(n_90)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_90),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_17),
.Y(n_91)
);

NAND2xp33_ASAP7_75t_SL g152 ( 
.A(n_91),
.B(n_92),
.Y(n_152)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_21),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_93),
.B(n_95),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_24),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_97),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_22),
.Y(n_96)
);

BUFx12_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_65),
.A2(n_21),
.B1(n_24),
.B2(n_48),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_99),
.A2(n_73),
.B1(n_88),
.B2(n_84),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_64),
.A2(n_24),
.B1(n_21),
.B2(n_49),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_104),
.A2(n_133),
.B1(n_140),
.B2(n_20),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_50),
.A2(n_25),
.B1(n_39),
.B2(n_38),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_110),
.A2(n_143),
.B1(n_18),
.B2(n_41),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_89),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_121),
.B(n_126),
.Y(n_171)
);

AOI21xp33_ASAP7_75t_L g123 ( 
.A1(n_67),
.A2(n_23),
.B(n_48),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_123),
.B(n_145),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_91),
.B(n_25),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_131),
.B(n_138),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_69),
.A2(n_24),
.B1(n_32),
.B2(n_49),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_77),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_134),
.B(n_150),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_96),
.B(n_17),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_55),
.A2(n_28),
.B1(n_39),
.B2(n_38),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_59),
.B(n_37),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_79),
.B(n_36),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_151),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_131),
.B(n_20),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_153),
.B(n_154),
.Y(n_210)
);

O2A1O1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_152),
.A2(n_52),
.B(n_37),
.C(n_29),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_116),
.A2(n_81),
.B1(n_29),
.B2(n_60),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_155),
.B(n_164),
.Y(n_219)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_100),
.Y(n_156)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_156),
.Y(n_215)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_116),
.A2(n_56),
.B1(n_95),
.B2(n_93),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_157),
.A2(n_161),
.B1(n_163),
.B2(n_172),
.Y(n_211)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_112),
.Y(n_158)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_158),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_124),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_159),
.B(n_160),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_138),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_122),
.Y(n_162)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_162),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_99),
.A2(n_75),
.B1(n_83),
.B2(n_70),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_L g164 ( 
.A1(n_109),
.A2(n_62),
.B(n_78),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_23),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_165),
.B(n_196),
.Y(n_214)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_144),
.Y(n_166)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_166),
.Y(n_207)
);

AND2x2_ASAP7_75t_SL g168 ( 
.A(n_149),
.B(n_54),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_168),
.B(n_107),
.C(n_111),
.Y(n_234)
);

NAND2xp33_ASAP7_75t_SL g169 ( 
.A(n_125),
.B(n_97),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_169),
.B(n_177),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_137),
.A2(n_61),
.B1(n_71),
.B2(n_53),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_170),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_133),
.A2(n_80),
.B1(n_23),
.B2(n_41),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_108),
.Y(n_173)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_173),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_174),
.A2(n_147),
.B1(n_146),
.B2(n_132),
.Y(n_237)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_139),
.Y(n_176)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_176),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g177 ( 
.A(n_106),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_115),
.Y(n_178)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_178),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_103),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_179),
.Y(n_216)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_113),
.Y(n_181)
);

INVx3_ASAP7_75t_SL g231 ( 
.A(n_181),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_119),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_182),
.B(n_184),
.Y(n_240)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_106),
.Y(n_183)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_183),
.Y(n_248)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_127),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_103),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_185),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_137),
.A2(n_20),
.B1(n_48),
.B2(n_41),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_118),
.A2(n_18),
.B1(n_46),
.B2(n_43),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_104),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_197),
.Y(n_205)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_127),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_190),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_128),
.A2(n_18),
.B1(n_72),
.B2(n_46),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_191),
.A2(n_192),
.B1(n_111),
.B2(n_107),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_118),
.A2(n_46),
.B1(n_43),
.B2(n_26),
.Y(n_192)
);

INVx4_ASAP7_75t_SL g193 ( 
.A(n_112),
.Y(n_193)
);

INVx6_ASAP7_75t_SL g222 ( 
.A(n_193),
.Y(n_222)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_117),
.Y(n_194)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_194),
.Y(n_239)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_117),
.Y(n_195)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_195),
.Y(n_236)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_98),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_119),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_117),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_198),
.B(n_203),
.Y(n_209)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_136),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_199),
.Y(n_225)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_135),
.Y(n_201)
);

INVx6_ASAP7_75t_L g213 ( 
.A(n_201),
.Y(n_213)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_141),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_202),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_114),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_218),
.B(n_234),
.Y(n_260)
);

BUFx8_ASAP7_75t_L g220 ( 
.A(n_198),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_220),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_165),
.B(n_105),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_247),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_175),
.B(n_129),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_227),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_159),
.B(n_129),
.Y(n_227)
);

MAJx2_ASAP7_75t_L g228 ( 
.A(n_167),
.B(n_102),
.C(n_129),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_228),
.B(n_33),
.C(n_22),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_171),
.B(n_98),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_230),
.B(n_232),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_167),
.B(n_102),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_187),
.A2(n_128),
.B1(n_105),
.B2(n_120),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_233),
.A2(n_241),
.B1(n_242),
.B2(n_243),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_237),
.A2(n_142),
.B1(n_197),
.B2(n_196),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_180),
.B(n_101),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_101),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_200),
.A2(n_120),
.B1(n_130),
.B2(n_147),
.Y(n_241)
);

OAI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_154),
.A2(n_180),
.B1(n_155),
.B2(n_162),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_160),
.A2(n_130),
.B1(n_146),
.B2(n_135),
.Y(n_243)
);

A2O1A1Ixp33_ASAP7_75t_L g244 ( 
.A1(n_153),
.A2(n_176),
.B(n_172),
.C(n_168),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_244),
.A2(n_168),
.B(n_177),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_166),
.B(n_135),
.Y(n_247)
);

AND2x2_ASAP7_75t_SL g321 ( 
.A(n_250),
.B(n_215),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_214),
.B(n_163),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_254),
.B(n_281),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_223),
.B(n_156),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_255),
.B(n_263),
.Y(n_290)
);

OAI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_244),
.A2(n_219),
.B1(n_210),
.B2(n_211),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_257),
.A2(n_266),
.B1(n_272),
.B2(n_275),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_209),
.Y(n_258)
);

INVx13_ASAP7_75t_L g291 ( 
.A(n_258),
.Y(n_291)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_225),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_259),
.Y(n_314)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_206),
.Y(n_261)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_261),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_262),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_214),
.B(n_182),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_210),
.B(n_178),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_264),
.B(n_274),
.Y(n_294)
);

NOR3xp33_ASAP7_75t_SL g265 ( 
.A(n_235),
.B(n_203),
.C(n_193),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_265),
.B(n_220),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_205),
.A2(n_184),
.B(n_190),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_267),
.A2(n_231),
.B(n_217),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_219),
.A2(n_173),
.B(n_183),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_268),
.A2(n_269),
.B(n_273),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_219),
.A2(n_194),
.B(n_195),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_206),
.Y(n_270)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_270),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_212),
.A2(n_161),
.B1(n_202),
.B2(n_199),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_271),
.A2(n_282),
.B1(n_284),
.B2(n_278),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_211),
.A2(n_185),
.B1(n_179),
.B2(n_132),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_221),
.A2(n_76),
.B(n_201),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_240),
.B(n_181),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_237),
.A2(n_142),
.B1(n_158),
.B2(n_43),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_225),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_276),
.B(n_285),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_228),
.B(n_101),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_277),
.B(n_221),
.C(n_208),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_241),
.B(n_3),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_278),
.B(n_279),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_224),
.B(n_26),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_233),
.A2(n_33),
.B1(n_22),
.B2(n_6),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_280),
.B(n_283),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_212),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_221),
.A2(n_33),
.B1(n_22),
.B2(n_8),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_218),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_234),
.B(n_5),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_247),
.B(n_9),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_286),
.B(n_287),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_207),
.B(n_9),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_229),
.Y(n_288)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_288),
.Y(n_305)
);

XNOR2x1_ASAP7_75t_L g351 ( 
.A(n_292),
.B(n_213),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_243),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_295),
.B(n_301),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_260),
.B(n_217),
.C(n_245),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_296),
.B(n_322),
.C(n_324),
.Y(n_352)
);

CKINVDCx14_ASAP7_75t_R g349 ( 
.A(n_297),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_258),
.B(n_236),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_299),
.B(n_300),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_251),
.B(n_252),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_281),
.B(n_222),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_274),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_303),
.B(n_311),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_306),
.A2(n_272),
.B1(n_266),
.B2(n_264),
.Y(n_330)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_261),
.Y(n_309)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_309),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g339 ( 
.A1(n_310),
.A2(n_319),
.B(n_321),
.Y(n_339)
);

INVx13_ASAP7_75t_L g311 ( 
.A(n_256),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_260),
.B(n_222),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_313),
.B(n_216),
.C(n_246),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_251),
.B(n_236),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_315),
.B(n_239),
.Y(n_353)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_270),
.Y(n_317)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_317),
.Y(n_334)
);

MAJx2_ASAP7_75t_L g318 ( 
.A(n_260),
.B(n_220),
.C(n_231),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_318),
.B(n_250),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_268),
.B(n_204),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_262),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_320),
.B(n_302),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_263),
.B(n_215),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_249),
.B(n_204),
.C(n_248),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_288),
.Y(n_325)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_325),
.Y(n_340)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_309),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_326),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_304),
.A2(n_267),
.B(n_269),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_328),
.A2(n_304),
.B(n_319),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_317),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_329),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_330),
.B(n_332),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_311),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_331),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_323),
.A2(n_253),
.B1(n_271),
.B2(n_249),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_323),
.A2(n_253),
.B1(n_282),
.B2(n_254),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_333),
.B(n_338),
.Y(n_375)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_335),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_336),
.B(n_350),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_312),
.A2(n_254),
.B1(n_255),
.B2(n_284),
.Y(n_338)
);

A2O1A1O1Ixp25_ASAP7_75t_L g341 ( 
.A1(n_294),
.A2(n_252),
.B(n_273),
.C(n_265),
.D(n_286),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_341),
.B(n_351),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_306),
.A2(n_275),
.B1(n_280),
.B2(n_285),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_342),
.B(n_347),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_312),
.A2(n_287),
.B1(n_279),
.B2(n_256),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_343),
.A2(n_302),
.B1(n_320),
.B2(n_319),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_290),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_345),
.Y(n_385)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_293),
.Y(n_346)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_346),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_290),
.A2(n_276),
.B1(n_283),
.B2(n_216),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_294),
.B(n_259),
.Y(n_348)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_348),
.Y(n_362)
);

MAJx2_ASAP7_75t_L g350 ( 
.A(n_289),
.B(n_213),
.C(n_239),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_353),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_316),
.B(n_248),
.Y(n_354)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_354),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_308),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_356),
.B(n_307),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_357),
.B(n_318),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_352),
.B(n_289),
.C(n_301),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_360),
.B(n_363),
.C(n_374),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_352),
.B(n_313),
.C(n_296),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g394 ( 
.A1(n_364),
.A2(n_339),
.B(n_348),
.Y(n_394)
);

CKINVDCx14_ASAP7_75t_R g386 ( 
.A(n_365),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_356),
.B(n_316),
.Y(n_366)
);

CKINVDCx14_ASAP7_75t_R g401 ( 
.A(n_366),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_368),
.A2(n_328),
.B1(n_330),
.B2(n_342),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_371),
.B(n_372),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_355),
.B(n_292),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_344),
.Y(n_373)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_373),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_355),
.B(n_322),
.C(n_321),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_335),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_377),
.B(n_384),
.Y(n_402)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_327),
.Y(n_381)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_381),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_345),
.B(n_307),
.Y(n_382)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_382),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_349),
.B(n_298),
.Y(n_384)
);

NAND4xp25_ASAP7_75t_L g388 ( 
.A(n_383),
.B(n_331),
.C(n_341),
.D(n_291),
.Y(n_388)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_388),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_385),
.A2(n_332),
.B1(n_333),
.B2(n_338),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_389),
.A2(n_409),
.B1(n_358),
.B2(n_367),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_SL g413 ( 
.A(n_390),
.B(n_394),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_363),
.B(n_350),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_391),
.B(n_392),
.Y(n_417)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_374),
.B(n_351),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_372),
.B(n_336),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_395),
.B(n_403),
.Y(n_418)
);

NOR2x1_ASAP7_75t_SL g396 ( 
.A(n_384),
.B(n_337),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_396),
.A2(n_366),
.B1(n_365),
.B2(n_378),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_373),
.B(n_324),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_398),
.B(n_405),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_SL g399 ( 
.A(n_370),
.B(n_369),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_SL g422 ( 
.A(n_399),
.B(n_310),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_371),
.B(n_339),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_360),
.B(n_321),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_404),
.B(n_380),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_383),
.Y(n_405)
);

FAx1_ASAP7_75t_SL g407 ( 
.A(n_370),
.B(n_369),
.CI(n_375),
.CON(n_407),
.SN(n_407)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_407),
.Y(n_428)
);

NOR3xp33_ASAP7_75t_L g408 ( 
.A(n_385),
.B(n_291),
.C(n_354),
.Y(n_408)
);

INVxp67_ASAP7_75t_SL g425 ( 
.A(n_408),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_359),
.A2(n_347),
.B1(n_295),
.B2(n_340),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_397),
.B(n_357),
.C(n_368),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_410),
.B(n_414),
.C(n_416),
.Y(n_430)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_411),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_386),
.A2(n_359),
.B1(n_362),
.B2(n_358),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_412),
.A2(n_424),
.B1(n_389),
.B2(n_400),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_397),
.B(n_375),
.C(n_364),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_387),
.B(n_380),
.C(n_362),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_419),
.B(n_427),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_393),
.A2(n_376),
.B(n_382),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_420),
.A2(n_415),
.B(n_424),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_421),
.B(n_427),
.Y(n_431)
);

XNOR2x1_ASAP7_75t_L g429 ( 
.A(n_422),
.B(n_403),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_401),
.A2(n_367),
.B1(n_381),
.B2(n_378),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_423),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_406),
.A2(n_361),
.B1(n_379),
.B2(n_340),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_391),
.B(n_361),
.Y(n_427)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_429),
.B(n_441),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_L g432 ( 
.A1(n_426),
.A2(n_402),
.B(n_394),
.Y(n_432)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_432),
.Y(n_452)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_433),
.Y(n_455)
);

MAJx2_ASAP7_75t_L g434 ( 
.A(n_414),
.B(n_428),
.C(n_410),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_434),
.B(n_439),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_416),
.B(n_387),
.C(n_395),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_435),
.B(n_436),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_417),
.B(n_392),
.C(n_404),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_417),
.B(n_409),
.C(n_399),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_438),
.B(n_440),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_419),
.B(n_407),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_413),
.B(n_407),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_443),
.A2(n_334),
.B1(n_422),
.B2(n_346),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_442),
.B(n_412),
.Y(n_446)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_446),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_437),
.A2(n_425),
.B1(n_379),
.B2(n_327),
.Y(n_448)
);

AOI322xp5_ASAP7_75t_L g462 ( 
.A1(n_448),
.A2(n_456),
.A3(n_418),
.B1(n_314),
.B2(n_246),
.C1(n_33),
.C2(n_14),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_430),
.B(n_413),
.Y(n_450)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_450),
.Y(n_458)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_451),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_437),
.A2(n_334),
.B1(n_325),
.B2(n_305),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_453),
.B(n_12),
.Y(n_465)
);

OR2x2_ASAP7_75t_L g454 ( 
.A(n_431),
.B(n_314),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g459 ( 
.A1(n_454),
.A2(n_429),
.B(n_431),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_430),
.A2(n_434),
.B1(n_438),
.B2(n_435),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_459),
.B(n_462),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_444),
.B(n_436),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_460),
.B(n_466),
.Y(n_475)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_452),
.Y(n_461)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_461),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_444),
.B(n_418),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_463),
.B(n_464),
.Y(n_471)
);

CKINVDCx16_ASAP7_75t_R g464 ( 
.A(n_455),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_465),
.B(n_467),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_450),
.B(n_12),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_L g470 ( 
.A1(n_458),
.A2(n_445),
.B(n_447),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_470),
.A2(n_449),
.B(n_12),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_461),
.B(n_446),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_472),
.A2(n_459),
.B(n_454),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_460),
.A2(n_457),
.B(n_466),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_473),
.A2(n_469),
.B(n_471),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_474),
.B(n_465),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_476),
.B(n_478),
.Y(n_482)
);

NOR2xp67_ASAP7_75t_SL g477 ( 
.A(n_468),
.B(n_449),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_477),
.A2(n_479),
.B(n_480),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_478),
.A2(n_475),
.B(n_472),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_483),
.B(n_12),
.C(n_14),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_484),
.B(n_482),
.Y(n_485)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_485),
.B(n_481),
.Y(n_486)
);


endmodule