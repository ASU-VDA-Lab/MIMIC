module real_jpeg_1335_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_1),
.A2(n_23),
.B1(n_27),
.B2(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_1),
.Y(n_66)
);

BUFx4f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_3),
.B(n_34),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_3),
.A2(n_51),
.B1(n_52),
.B2(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_3),
.Y(n_57)
);

O2A1O1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_3),
.A2(n_4),
.B(n_51),
.C(n_70),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_3),
.B(n_23),
.C(n_26),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_3),
.A2(n_18),
.B1(n_19),
.B2(n_57),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_3),
.B(n_40),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_3),
.B(n_82),
.Y(n_97)
);

AO22x2_ASAP7_75t_L g34 ( 
.A1(n_4),
.A2(n_18),
.B1(n_19),
.B2(n_35),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

O2A1O1Ixp33_ASAP7_75t_L g50 ( 
.A1(n_4),
.A2(n_34),
.B(n_51),
.C(n_55),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_4),
.B(n_51),
.Y(n_55)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_7),
.A2(n_18),
.B1(n_19),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_7),
.A2(n_23),
.B1(n_27),
.B2(n_32),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_7),
.A2(n_32),
.B1(n_51),
.B2(n_52),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_8),
.A2(n_23),
.B1(n_27),
.B2(n_42),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_8),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_8),
.A2(n_18),
.B1(n_19),
.B2(n_42),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_9),
.A2(n_18),
.B1(n_19),
.B2(n_21),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_9),
.A2(n_21),
.B1(n_23),
.B2(n_27),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_73),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_71),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_46),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_14),
.B(n_46),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_33),
.C(n_36),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_15),
.A2(n_16),
.B1(n_33),
.B2(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_22),
.B(n_28),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_17),
.A2(n_22),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_L g30 ( 
.A1(n_18),
.A2(n_19),
.B1(n_25),
.B2(n_26),
.Y(n_30)
);

OAI21xp33_ASAP7_75t_L g70 ( 
.A1(n_18),
.A2(n_35),
.B(n_57),
.Y(n_70)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_19),
.B(n_78),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_22),
.Y(n_82)
);

OA22x2_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_22)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_23),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_23),
.B(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_31),
.B(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_36),
.A2(n_37),
.B1(n_84),
.B2(n_86),
.Y(n_83)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_41),
.B(n_43),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_38),
.B(n_45),
.Y(n_68)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_38),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_38),
.A2(n_39),
.B1(n_41),
.B2(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_45),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_39),
.A2(n_65),
.B(n_67),
.Y(n_64)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_40),
.A2(n_68),
.B(n_96),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_44),
.A2(n_57),
.B(n_93),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_63),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_60),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_56),
.B(n_58),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_61),
.A2(n_80),
.B(n_81),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_69),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_87),
.B(n_105),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_83),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_83),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_76),
.A2(n_77),
.B1(n_79),
.B2(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_79),
.Y(n_103)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_84),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_99),
.B(n_104),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_94),
.B(n_98),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_92),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_95),
.B(n_97),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_97),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_102),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_100),
.B(n_102),
.Y(n_104)
);


endmodule