module fake_aes_12629_n_680 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_680);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_680;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
NOR2xp67_ASAP7_75t_L g81 ( .A(n_48), .B(n_80), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_5), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_10), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_27), .Y(n_84) );
INVx2_ASAP7_75t_L g85 ( .A(n_54), .Y(n_85) );
INVxp33_ASAP7_75t_L g86 ( .A(n_75), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_64), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_55), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_22), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_44), .Y(n_90) );
INVx2_ASAP7_75t_L g91 ( .A(n_71), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_52), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_50), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_58), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_0), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_41), .Y(n_96) );
NOR2xp67_ASAP7_75t_L g97 ( .A(n_66), .B(n_74), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_42), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_40), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_51), .Y(n_100) );
INVxp67_ASAP7_75t_SL g101 ( .A(n_12), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_11), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_25), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_72), .Y(n_104) );
HB1xp67_ASAP7_75t_L g105 ( .A(n_30), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_31), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_69), .Y(n_107) );
INVx1_ASAP7_75t_SL g108 ( .A(n_24), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_53), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_36), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_14), .Y(n_111) );
BUFx10_ASAP7_75t_L g112 ( .A(n_45), .Y(n_112) );
INVxp33_ASAP7_75t_SL g113 ( .A(n_49), .Y(n_113) );
INVxp67_ASAP7_75t_L g114 ( .A(n_16), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_73), .Y(n_115) );
INVxp67_ASAP7_75t_SL g116 ( .A(n_76), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_65), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_61), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_0), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_84), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_84), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_87), .Y(n_122) );
OA21x2_ASAP7_75t_L g123 ( .A1(n_87), .A2(n_109), .B(n_100), .Y(n_123) );
AOI22xp5_ASAP7_75t_L g124 ( .A1(n_82), .A2(n_119), .B1(n_83), .B2(n_95), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_89), .Y(n_125) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_85), .Y(n_126) );
OAI22xp5_ASAP7_75t_SL g127 ( .A1(n_101), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_89), .Y(n_128) );
OA21x2_ASAP7_75t_L g129 ( .A1(n_90), .A2(n_38), .B(n_79), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_90), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_92), .Y(n_131) );
BUFx3_ASAP7_75t_L g132 ( .A(n_85), .Y(n_132) );
AND2x4_ASAP7_75t_L g133 ( .A(n_82), .B(n_1), .Y(n_133) );
OAI21x1_ASAP7_75t_L g134 ( .A1(n_85), .A2(n_39), .B(n_78), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_105), .B(n_2), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_91), .Y(n_136) );
OAI22xp5_ASAP7_75t_L g137 ( .A1(n_83), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_137) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_91), .Y(n_138) );
OAI21x1_ASAP7_75t_L g139 ( .A1(n_91), .A2(n_43), .B(n_77), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_120), .B(n_92), .Y(n_140) );
INVx3_ASAP7_75t_L g141 ( .A(n_132), .Y(n_141) );
BUFx2_ASAP7_75t_L g142 ( .A(n_135), .Y(n_142) );
AND2x2_ASAP7_75t_L g143 ( .A(n_120), .B(n_112), .Y(n_143) );
INVx5_ASAP7_75t_L g144 ( .A(n_126), .Y(n_144) );
INVx3_ASAP7_75t_L g145 ( .A(n_132), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_136), .Y(n_146) );
AOI22xp33_ASAP7_75t_L g147 ( .A1(n_121), .A2(n_95), .B1(n_102), .B2(n_111), .Y(n_147) );
OR2x2_ASAP7_75t_L g148 ( .A(n_135), .B(n_114), .Y(n_148) );
AOI22xp33_ASAP7_75t_L g149 ( .A1(n_121), .A2(n_102), .B1(n_111), .B2(n_119), .Y(n_149) );
AOI22xp33_ASAP7_75t_L g150 ( .A1(n_122), .A2(n_113), .B1(n_109), .B2(n_96), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_133), .B(n_96), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_122), .B(n_100), .Y(n_152) );
INVxp67_ASAP7_75t_SL g153 ( .A(n_125), .Y(n_153) );
AOI22xp33_ASAP7_75t_L g154 ( .A1(n_125), .A2(n_104), .B1(n_103), .B2(n_107), .Y(n_154) );
AOI22xp33_ASAP7_75t_L g155 ( .A1(n_128), .A2(n_104), .B1(n_103), .B2(n_107), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_128), .B(n_110), .Y(n_156) );
NOR2x1p5_ASAP7_75t_L g157 ( .A(n_133), .B(n_116), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_136), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_134), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_130), .B(n_86), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_136), .Y(n_161) );
AOI22xp33_ASAP7_75t_L g162 ( .A1(n_130), .A2(n_110), .B1(n_117), .B2(n_93), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_131), .B(n_93), .Y(n_163) );
INVx4_ASAP7_75t_L g164 ( .A(n_133), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_126), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_126), .Y(n_166) );
INVx4_ASAP7_75t_L g167 ( .A(n_133), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_126), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_136), .Y(n_169) );
A2O1A1Ixp33_ASAP7_75t_L g170 ( .A1(n_153), .A2(n_131), .B(n_132), .C(n_124), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_142), .B(n_124), .Y(n_171) );
OR2x2_ASAP7_75t_L g172 ( .A(n_142), .B(n_137), .Y(n_172) );
AOI22xp5_ASAP7_75t_L g173 ( .A1(n_157), .A2(n_127), .B1(n_137), .B2(n_123), .Y(n_173) );
INVxp67_ASAP7_75t_SL g174 ( .A(n_153), .Y(n_174) );
HB1xp67_ASAP7_75t_L g175 ( .A(n_142), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_141), .Y(n_176) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_157), .A2(n_127), .B1(n_123), .B2(n_112), .Y(n_177) );
AOI22xp5_ASAP7_75t_L g178 ( .A1(n_143), .A2(n_123), .B1(n_112), .B2(n_117), .Y(n_178) );
NOR3xp33_ASAP7_75t_L g179 ( .A(n_143), .B(n_108), .C(n_115), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_141), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_143), .B(n_123), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_141), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_148), .B(n_123), .Y(n_183) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_159), .Y(n_184) );
NOR3x1_ASAP7_75t_L g185 ( .A(n_148), .B(n_139), .C(n_134), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_160), .B(n_88), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_141), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_141), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_148), .B(n_112), .Y(n_189) );
AO22x1_ASAP7_75t_L g190 ( .A1(n_151), .A2(n_117), .B1(n_99), .B2(n_93), .Y(n_190) );
AND2x2_ASAP7_75t_L g191 ( .A(n_160), .B(n_134), .Y(n_191) );
INVx2_ASAP7_75t_SL g192 ( .A(n_164), .Y(n_192) );
AND2x2_ASAP7_75t_L g193 ( .A(n_164), .B(n_139), .Y(n_193) );
INVxp67_ASAP7_75t_SL g194 ( .A(n_145), .Y(n_194) );
INVx3_ASAP7_75t_L g195 ( .A(n_164), .Y(n_195) );
INVxp67_ASAP7_75t_SL g196 ( .A(n_145), .Y(n_196) );
AOI22xp33_ASAP7_75t_L g197 ( .A1(n_151), .A2(n_126), .B1(n_138), .B2(n_136), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_151), .B(n_139), .Y(n_198) );
NOR3xp33_ASAP7_75t_L g199 ( .A(n_140), .B(n_94), .C(n_98), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_164), .B(n_106), .Y(n_200) );
OR2x6_ASAP7_75t_L g201 ( .A(n_164), .B(n_129), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_167), .B(n_118), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_151), .B(n_129), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_151), .B(n_99), .Y(n_204) );
AOI22xp33_ASAP7_75t_L g205 ( .A1(n_167), .A2(n_126), .B1(n_136), .B2(n_138), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_167), .B(n_99), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_167), .B(n_145), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_167), .B(n_97), .Y(n_208) );
NOR3xp33_ASAP7_75t_L g209 ( .A(n_171), .B(n_140), .C(n_152), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_198), .A2(n_159), .B(n_152), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g211 ( .A1(n_198), .A2(n_159), .B(n_156), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_181), .B(n_159), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_175), .B(n_150), .Y(n_213) );
NOR3xp33_ASAP7_75t_L g214 ( .A(n_172), .B(n_156), .C(n_163), .Y(n_214) );
O2A1O1Ixp5_ASAP7_75t_L g215 ( .A1(n_190), .A2(n_145), .B(n_163), .C(n_166), .Y(n_215) );
O2A1O1Ixp5_ASAP7_75t_L g216 ( .A1(n_190), .A2(n_145), .B(n_168), .C(n_166), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_203), .A2(n_159), .B(n_129), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_174), .B(n_150), .Y(n_218) );
OAI21xp5_ASAP7_75t_L g219 ( .A1(n_203), .A2(n_162), .B(n_154), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_181), .A2(n_159), .B(n_129), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_183), .B(n_159), .Y(n_221) );
OR2x6_ASAP7_75t_SL g222 ( .A(n_172), .B(n_147), .Y(n_222) );
OA22x2_ASAP7_75t_L g223 ( .A1(n_173), .A2(n_154), .B1(n_155), .B2(n_147), .Y(n_223) );
AOI22xp5_ASAP7_75t_L g224 ( .A1(n_189), .A2(n_149), .B1(n_155), .B2(n_162), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_184), .Y(n_225) );
AO21x1_ASAP7_75t_L g226 ( .A1(n_191), .A2(n_169), .B(n_146), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_183), .B(n_149), .Y(n_227) );
AND2x2_ASAP7_75t_L g228 ( .A(n_177), .B(n_173), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_176), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g230 ( .A(n_177), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_178), .B(n_159), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_193), .A2(n_129), .B(n_146), .Y(n_232) );
AOI21x1_ASAP7_75t_L g233 ( .A1(n_193), .A2(n_169), .B(n_158), .Y(n_233) );
AND2x4_ASAP7_75t_L g234 ( .A(n_179), .B(n_81), .Y(n_234) );
O2A1O1Ixp33_ASAP7_75t_L g235 ( .A1(n_170), .A2(n_161), .B(n_158), .C(n_165), .Y(n_235) );
NAND2x1p5_ASAP7_75t_L g236 ( .A(n_195), .B(n_138), .Y(n_236) );
AOI22xp33_ASAP7_75t_L g237 ( .A1(n_191), .A2(n_138), .B1(n_126), .B2(n_161), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_186), .B(n_4), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_178), .B(n_6), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_207), .A2(n_168), .B(n_166), .Y(n_240) );
BUFx2_ASAP7_75t_L g241 ( .A(n_239), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_212), .A2(n_184), .B(n_206), .Y(n_242) );
OAI22xp5_ASAP7_75t_L g243 ( .A1(n_230), .A2(n_204), .B1(n_200), .B2(n_202), .Y(n_243) );
AOI22xp5_ASAP7_75t_L g244 ( .A1(n_230), .A2(n_199), .B1(n_192), .B2(n_195), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_212), .A2(n_184), .B(n_201), .Y(n_245) );
OR2x2_ASAP7_75t_L g246 ( .A(n_213), .B(n_194), .Y(n_246) );
OAI21x1_ASAP7_75t_L g247 ( .A1(n_220), .A2(n_208), .B(n_197), .Y(n_247) );
BUFx8_ASAP7_75t_L g248 ( .A(n_228), .Y(n_248) );
AOI21x1_ASAP7_75t_L g249 ( .A1(n_217), .A2(n_201), .B(n_165), .Y(n_249) );
OAI21x1_ASAP7_75t_L g250 ( .A1(n_232), .A2(n_205), .B(n_185), .Y(n_250) );
OR2x2_ASAP7_75t_L g251 ( .A(n_218), .B(n_196), .Y(n_251) );
BUFx3_ASAP7_75t_L g252 ( .A(n_236), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_229), .Y(n_253) );
AO31x2_ASAP7_75t_L g254 ( .A1(n_226), .A2(n_211), .A3(n_210), .B(n_238), .Y(n_254) );
OAI21x1_ASAP7_75t_L g255 ( .A1(n_231), .A2(n_185), .B(n_168), .Y(n_255) );
OAI22xp33_ASAP7_75t_L g256 ( .A1(n_222), .A2(n_195), .B1(n_201), .B2(n_188), .Y(n_256) );
OAI21xp5_ASAP7_75t_L g257 ( .A1(n_221), .A2(n_188), .B(n_176), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_223), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_223), .Y(n_259) );
A2O1A1Ixp33_ASAP7_75t_L g260 ( .A1(n_238), .A2(n_219), .B(n_209), .C(n_214), .Y(n_260) );
AO21x2_ASAP7_75t_L g261 ( .A1(n_231), .A2(n_165), .B(n_187), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_221), .A2(n_184), .B(n_240), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_260), .A2(n_201), .B(n_225), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_260), .A2(n_201), .B(n_225), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_253), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_253), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_251), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_246), .Y(n_268) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_252), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_245), .A2(n_235), .B(n_184), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g271 ( .A1(n_262), .A2(n_227), .B(n_216), .Y(n_271) );
AOI21xp5_ASAP7_75t_L g272 ( .A1(n_242), .A2(n_237), .B(n_215), .Y(n_272) );
OAI21x1_ASAP7_75t_L g273 ( .A1(n_249), .A2(n_233), .B(n_236), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_241), .B(n_222), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_246), .Y(n_275) );
AO31x2_ASAP7_75t_L g276 ( .A1(n_258), .A2(n_187), .A3(n_182), .B(n_180), .Y(n_276) );
INVxp67_ASAP7_75t_L g277 ( .A(n_248), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_251), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_259), .Y(n_279) );
AO21x2_ASAP7_75t_L g280 ( .A1(n_255), .A2(n_234), .B(n_224), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_254), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_241), .B(n_234), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_248), .B(n_234), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_248), .B(n_182), .Y(n_284) );
BUFx3_ASAP7_75t_L g285 ( .A(n_269), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_266), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_281), .Y(n_287) );
OR2x6_ASAP7_75t_L g288 ( .A(n_263), .B(n_255), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_266), .B(n_254), .Y(n_289) );
INVx1_ASAP7_75t_SL g290 ( .A(n_265), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_279), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_279), .Y(n_292) );
INVxp33_ASAP7_75t_SL g293 ( .A(n_284), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_281), .Y(n_294) );
OR2x2_ASAP7_75t_L g295 ( .A(n_274), .B(n_254), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_267), .B(n_254), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_276), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_276), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_276), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_276), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_276), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_267), .B(n_254), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_280), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_278), .B(n_252), .Y(n_304) );
BUFx6f_ASAP7_75t_L g305 ( .A(n_273), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_278), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_280), .Y(n_307) );
INVx8_ASAP7_75t_L g308 ( .A(n_277), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_280), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_268), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_275), .B(n_261), .Y(n_311) );
INVx3_ASAP7_75t_L g312 ( .A(n_273), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_264), .Y(n_313) );
BUFx2_ASAP7_75t_SL g314 ( .A(n_270), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_271), .Y(n_315) );
AO21x2_ASAP7_75t_L g316 ( .A1(n_272), .A2(n_256), .B(n_250), .Y(n_316) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_290), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_289), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_287), .Y(n_319) );
OR2x2_ASAP7_75t_L g320 ( .A(n_295), .B(n_282), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_289), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_287), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_289), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_291), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_287), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_296), .B(n_261), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_296), .B(n_261), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_294), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_302), .B(n_283), .Y(n_329) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_290), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_302), .B(n_243), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_291), .Y(n_332) );
INVxp67_ASAP7_75t_L g333 ( .A(n_286), .Y(n_333) );
BUFx2_ASAP7_75t_L g334 ( .A(n_285), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_311), .B(n_250), .Y(n_335) );
OR2x2_ASAP7_75t_L g336 ( .A(n_295), .B(n_257), .Y(n_336) );
OR2x2_ASAP7_75t_L g337 ( .A(n_311), .B(n_138), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_311), .B(n_138), .Y(n_338) );
HB1xp67_ASAP7_75t_L g339 ( .A(n_285), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_292), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_306), .B(n_286), .Y(n_341) );
INVx3_ASAP7_75t_L g342 ( .A(n_305), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_294), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_292), .Y(n_344) );
INVx2_ASAP7_75t_SL g345 ( .A(n_285), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_298), .Y(n_346) );
AOI22xp33_ASAP7_75t_L g347 ( .A1(n_293), .A2(n_244), .B1(n_247), .B2(n_180), .Y(n_347) );
INVx4_ASAP7_75t_L g348 ( .A(n_308), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_297), .Y(n_349) );
INVxp67_ASAP7_75t_SL g350 ( .A(n_298), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_297), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_298), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_299), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_301), .Y(n_354) );
BUFx2_ASAP7_75t_L g355 ( .A(n_312), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_306), .B(n_247), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_310), .B(n_7), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_301), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_310), .B(n_7), .Y(n_359) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_299), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_299), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_300), .B(n_8), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_300), .Y(n_363) );
AND2x4_ASAP7_75t_L g364 ( .A(n_300), .B(n_47), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_315), .Y(n_365) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_312), .Y(n_366) );
NOR2xp33_ASAP7_75t_R g367 ( .A(n_308), .B(n_8), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_315), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_303), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_349), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_349), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_351), .Y(n_372) );
AND2x4_ASAP7_75t_L g373 ( .A(n_318), .B(n_312), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_351), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_321), .B(n_307), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_321), .B(n_307), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_354), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_323), .B(n_303), .Y(n_378) );
BUFx3_ASAP7_75t_L g379 ( .A(n_334), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_323), .B(n_309), .Y(n_380) );
INVxp67_ASAP7_75t_L g381 ( .A(n_339), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_346), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_335), .B(n_309), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_324), .Y(n_384) );
INVxp67_ASAP7_75t_SL g385 ( .A(n_317), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_329), .B(n_304), .Y(n_386) );
AND2x4_ASAP7_75t_L g387 ( .A(n_354), .B(n_312), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_335), .B(n_303), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_358), .Y(n_389) );
OR2x2_ASAP7_75t_L g390 ( .A(n_320), .B(n_309), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_329), .B(n_320), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_326), .B(n_316), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_324), .B(n_304), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_326), .B(n_316), .Y(n_394) );
OR2x2_ASAP7_75t_L g395 ( .A(n_317), .B(n_313), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_356), .B(n_316), .Y(n_396) );
INVxp67_ASAP7_75t_SL g397 ( .A(n_330), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_356), .B(n_316), .Y(n_398) );
INVx3_ASAP7_75t_R g399 ( .A(n_364), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_338), .B(n_313), .Y(n_400) );
AND2x4_ASAP7_75t_SL g401 ( .A(n_348), .B(n_308), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_358), .Y(n_402) );
INVx1_ASAP7_75t_SL g403 ( .A(n_334), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_346), .Y(n_404) );
AND2x4_ASAP7_75t_L g405 ( .A(n_345), .B(n_288), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_338), .B(n_288), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_332), .B(n_288), .Y(n_407) );
OR2x2_ASAP7_75t_L g408 ( .A(n_330), .B(n_288), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_346), .Y(n_409) );
BUFx2_ASAP7_75t_L g410 ( .A(n_345), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_332), .B(n_288), .Y(n_411) );
NOR2xp67_ASAP7_75t_L g412 ( .A(n_348), .B(n_9), .Y(n_412) );
INVxp67_ASAP7_75t_SL g413 ( .A(n_360), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_340), .Y(n_414) );
INVxp67_ASAP7_75t_SL g415 ( .A(n_360), .Y(n_415) );
AND2x4_ASAP7_75t_L g416 ( .A(n_345), .B(n_288), .Y(n_416) );
INVx2_ASAP7_75t_SL g417 ( .A(n_348), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_352), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_340), .B(n_305), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_344), .B(n_305), .Y(n_420) );
NOR2x1_ASAP7_75t_L g421 ( .A(n_348), .B(n_305), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_344), .Y(n_422) );
OR2x2_ASAP7_75t_L g423 ( .A(n_331), .B(n_305), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_368), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_368), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_341), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_331), .B(n_308), .Y(n_427) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_337), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_341), .B(n_308), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_352), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_361), .B(n_305), .Y(n_431) );
INVxp67_ASAP7_75t_L g432 ( .A(n_357), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_361), .Y(n_433) );
INVx3_ASAP7_75t_L g434 ( .A(n_355), .Y(n_434) );
OR2x2_ASAP7_75t_L g435 ( .A(n_327), .B(n_305), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_363), .B(n_314), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_363), .B(n_314), .Y(n_437) );
INVx2_ASAP7_75t_SL g438 ( .A(n_319), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_333), .B(n_308), .Y(n_439) );
AND2x4_ASAP7_75t_SL g440 ( .A(n_364), .B(n_362), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_327), .B(n_9), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_352), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_353), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_319), .B(n_10), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_319), .B(n_11), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_353), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_365), .Y(n_447) );
OR2x2_ASAP7_75t_L g448 ( .A(n_391), .B(n_333), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_381), .B(n_362), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_386), .B(n_336), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_432), .B(n_336), .Y(n_451) );
AND2x4_ASAP7_75t_L g452 ( .A(n_373), .B(n_355), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_384), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_382), .Y(n_454) );
AND2x4_ASAP7_75t_L g455 ( .A(n_373), .B(n_366), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_414), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_422), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_428), .B(n_350), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_390), .B(n_322), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_441), .B(n_357), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_382), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_370), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_371), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_403), .B(n_322), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_371), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_404), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_426), .B(n_365), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_390), .B(n_322), .Y(n_468) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_413), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_372), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_393), .B(n_365), .Y(n_471) );
NOR2x1_ASAP7_75t_L g472 ( .A(n_412), .B(n_359), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_404), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_392), .B(n_353), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_423), .B(n_343), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_417), .B(n_367), .Y(n_476) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_427), .B(n_359), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_383), .B(n_343), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_383), .B(n_343), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_388), .B(n_325), .Y(n_480) );
INVx1_ASAP7_75t_SL g481 ( .A(n_401), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_388), .B(n_325), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_423), .B(n_325), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_372), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_374), .Y(n_485) );
INVxp67_ASAP7_75t_L g486 ( .A(n_410), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_406), .B(n_328), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_409), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_406), .B(n_328), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_374), .Y(n_490) );
INVxp67_ASAP7_75t_SL g491 ( .A(n_415), .Y(n_491) );
NAND2x1_ASAP7_75t_L g492 ( .A(n_417), .B(n_364), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_392), .B(n_369), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_394), .B(n_369), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_385), .B(n_328), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_377), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_418), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_394), .B(n_369), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_396), .B(n_366), .Y(n_499) );
OAI332xp33_ASAP7_75t_L g500 ( .A1(n_395), .A2(n_12), .A3(n_13), .B1(n_14), .B2(n_15), .B3(n_16), .C1(n_17), .C2(n_18), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_377), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_396), .B(n_342), .Y(n_502) );
INVxp67_ASAP7_75t_L g503 ( .A(n_410), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_379), .B(n_364), .Y(n_504) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_438), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_389), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_389), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_397), .B(n_342), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_402), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_379), .B(n_342), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_375), .B(n_347), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_375), .B(n_342), .Y(n_512) );
INVx2_ASAP7_75t_SL g513 ( .A(n_421), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_378), .B(n_13), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_418), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_378), .B(n_15), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_440), .B(n_17), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_402), .Y(n_518) );
AND2x4_ASAP7_75t_SL g519 ( .A(n_405), .B(n_19), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_438), .B(n_19), .Y(n_520) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_430), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_424), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_430), .Y(n_523) );
OR2x2_ASAP7_75t_L g524 ( .A(n_435), .B(n_20), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_376), .B(n_20), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_424), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_425), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_442), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_425), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_433), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_433), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_453), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_487), .B(n_407), .Y(n_533) );
NAND3xp33_ASAP7_75t_SL g534 ( .A(n_476), .B(n_439), .C(n_445), .Y(n_534) );
AND2x4_ASAP7_75t_SL g535 ( .A(n_452), .B(n_405), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_450), .B(n_398), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_456), .Y(n_537) );
OAI22xp33_ASAP7_75t_L g538 ( .A1(n_481), .A2(n_429), .B1(n_408), .B2(n_434), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_489), .B(n_407), .Y(n_539) );
NAND2xp33_ASAP7_75t_SL g540 ( .A(n_492), .B(n_399), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_457), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_448), .B(n_435), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_499), .B(n_411), .Y(n_543) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_476), .A2(n_411), .B1(n_401), .B2(n_373), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_462), .Y(n_545) );
NAND3xp33_ASAP7_75t_SL g546 ( .A(n_517), .B(n_445), .C(n_444), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_463), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_465), .Y(n_548) );
NAND2x1p5_ASAP7_75t_L g549 ( .A(n_472), .B(n_444), .Y(n_549) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_469), .Y(n_550) );
AND2x4_ASAP7_75t_L g551 ( .A(n_455), .B(n_452), .Y(n_551) );
OAI32xp33_ASAP7_75t_L g552 ( .A1(n_469), .A2(n_408), .A3(n_434), .B1(n_395), .B2(n_399), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_499), .B(n_416), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_454), .Y(n_554) );
OAI31xp67_ASAP7_75t_L g555 ( .A1(n_500), .A2(n_446), .A3(n_443), .B(n_442), .Y(n_555) );
AND2x4_ASAP7_75t_L g556 ( .A(n_455), .B(n_405), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_451), .B(n_380), .Y(n_557) );
INVxp67_ASAP7_75t_L g558 ( .A(n_505), .Y(n_558) );
INVxp67_ASAP7_75t_SL g559 ( .A(n_491), .Y(n_559) );
NAND2x1p5_ASAP7_75t_L g560 ( .A(n_520), .B(n_416), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_461), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_461), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_470), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_493), .B(n_416), .Y(n_564) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_521), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_484), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_485), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_490), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_494), .B(n_440), .Y(n_569) );
AND2x4_ASAP7_75t_L g570 ( .A(n_455), .B(n_387), .Y(n_570) );
OR2x2_ASAP7_75t_L g571 ( .A(n_494), .B(n_400), .Y(n_571) );
OAI22xp33_ASAP7_75t_L g572 ( .A1(n_514), .A2(n_434), .B1(n_447), .B2(n_443), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_498), .B(n_419), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_496), .Y(n_574) );
NOR2xp33_ASAP7_75t_SL g575 ( .A(n_519), .B(n_437), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_501), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_498), .B(n_420), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_506), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_502), .B(n_420), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_502), .B(n_387), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_507), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_466), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_509), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_474), .B(n_387), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_474), .B(n_447), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_466), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_518), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_478), .B(n_437), .Y(n_588) );
NAND2x1p5_ASAP7_75t_L g589 ( .A(n_504), .B(n_436), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g590 ( .A(n_477), .B(n_436), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_479), .B(n_431), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_480), .B(n_431), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_473), .Y(n_593) );
INVx1_ASAP7_75t_SL g594 ( .A(n_519), .Y(n_594) );
OAI21xp33_ASAP7_75t_L g595 ( .A1(n_486), .A2(n_446), .B(n_21), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_477), .B(n_21), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_482), .B(n_23), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_522), .Y(n_598) );
OAI322xp33_ASAP7_75t_L g599 ( .A1(n_590), .A2(n_516), .A3(n_524), .B1(n_460), .B2(n_525), .C1(n_503), .C2(n_486), .Y(n_599) );
OAI21xp33_ASAP7_75t_SL g600 ( .A1(n_559), .A2(n_491), .B(n_513), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_550), .Y(n_601) );
INVxp67_ASAP7_75t_SL g602 ( .A(n_550), .Y(n_602) );
INVxp67_ASAP7_75t_L g603 ( .A(n_575), .Y(n_603) );
O2A1O1Ixp33_ASAP7_75t_SL g604 ( .A1(n_594), .A2(n_503), .B(n_505), .C(n_513), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_532), .Y(n_605) );
INVxp67_ASAP7_75t_L g606 ( .A(n_565), .Y(n_606) );
AOI31xp33_ASAP7_75t_L g607 ( .A1(n_549), .A2(n_460), .A3(n_449), .B(n_458), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_536), .B(n_471), .Y(n_608) );
OA21x2_ASAP7_75t_L g609 ( .A1(n_559), .A2(n_512), .B(n_467), .Y(n_609) );
OAI21xp5_ASAP7_75t_SL g610 ( .A1(n_534), .A2(n_452), .B(n_511), .Y(n_610) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_565), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_590), .B(n_464), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_557), .B(n_529), .Y(n_613) );
OAI21xp5_ASAP7_75t_L g614 ( .A1(n_595), .A2(n_521), .B(n_508), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_537), .Y(n_615) );
AOI21xp5_ASAP7_75t_SL g616 ( .A1(n_534), .A2(n_495), .B(n_510), .Y(n_616) );
OAI21xp5_ASAP7_75t_L g617 ( .A1(n_546), .A2(n_549), .B(n_558), .Y(n_617) );
OAI22xp33_ASAP7_75t_L g618 ( .A1(n_544), .A2(n_459), .B1(n_468), .B2(n_531), .Y(n_618) );
OAI22xp5_ASAP7_75t_L g619 ( .A1(n_589), .A2(n_475), .B1(n_483), .B2(n_530), .Y(n_619) );
NAND2xp5_ASAP7_75t_SL g620 ( .A(n_540), .B(n_528), .Y(n_620) );
OA22x2_ASAP7_75t_L g621 ( .A1(n_535), .A2(n_526), .B1(n_527), .B2(n_528), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_541), .Y(n_622) );
BUFx3_ASAP7_75t_L g623 ( .A(n_551), .Y(n_623) );
OR2x2_ASAP7_75t_L g624 ( .A(n_571), .B(n_523), .Y(n_624) );
INVx1_ASAP7_75t_SL g625 ( .A(n_542), .Y(n_625) );
AOI211xp5_ASAP7_75t_L g626 ( .A1(n_538), .A2(n_515), .B(n_497), .C(n_488), .Y(n_626) );
OR4x1_ASAP7_75t_L g627 ( .A(n_555), .B(n_26), .C(n_28), .D(n_29), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_556), .A2(n_144), .B1(n_33), .B2(n_34), .Y(n_628) );
A2O1A1Ixp33_ASAP7_75t_SL g629 ( .A1(n_596), .A2(n_32), .B(n_35), .C(n_37), .Y(n_629) );
OAI21xp5_ASAP7_75t_SL g630 ( .A1(n_538), .A2(n_46), .B(n_56), .Y(n_630) );
OAI21xp5_ASAP7_75t_SL g631 ( .A1(n_572), .A2(n_57), .B(n_59), .Y(n_631) );
NAND2xp5_ASAP7_75t_SL g632 ( .A(n_600), .B(n_551), .Y(n_632) );
OAI221xp5_ASAP7_75t_L g633 ( .A1(n_610), .A2(n_560), .B1(n_589), .B2(n_584), .C(n_547), .Y(n_633) );
AOI222xp33_ASAP7_75t_L g634 ( .A1(n_617), .A2(n_552), .B1(n_563), .B2(n_578), .C1(n_568), .C2(n_567), .Y(n_634) );
AOI221xp5_ASAP7_75t_SL g635 ( .A1(n_607), .A2(n_585), .B1(n_553), .B2(n_580), .C(n_564), .Y(n_635) );
O2A1O1Ixp33_ASAP7_75t_L g636 ( .A1(n_630), .A2(n_560), .B(n_576), .C(n_587), .Y(n_636) );
AOI211xp5_ASAP7_75t_SL g637 ( .A1(n_630), .A2(n_597), .B(n_551), .C(n_556), .Y(n_637) );
INVx2_ASAP7_75t_SL g638 ( .A(n_623), .Y(n_638) );
AOI21xp5_ASAP7_75t_L g639 ( .A1(n_604), .A2(n_556), .B(n_570), .Y(n_639) );
AND3x1_ASAP7_75t_L g640 ( .A(n_610), .B(n_569), .C(n_588), .Y(n_640) );
OA21x2_ASAP7_75t_L g641 ( .A1(n_603), .A2(n_593), .B(n_586), .Y(n_641) );
INVxp67_ASAP7_75t_L g642 ( .A(n_602), .Y(n_642) );
AOI322xp5_ASAP7_75t_L g643 ( .A1(n_625), .A2(n_543), .A3(n_573), .B1(n_577), .B2(n_533), .C1(n_539), .C2(n_579), .Y(n_643) );
OAI21xp5_ASAP7_75t_SL g644 ( .A1(n_631), .A2(n_570), .B(n_598), .Y(n_644) );
AOI21xp5_ASAP7_75t_L g645 ( .A1(n_616), .A2(n_570), .B(n_545), .Y(n_645) );
AOI22xp5_ASAP7_75t_L g646 ( .A1(n_621), .A2(n_574), .B1(n_548), .B2(n_583), .Y(n_646) );
O2A1O1Ixp33_ASAP7_75t_L g647 ( .A1(n_631), .A2(n_581), .B(n_566), .C(n_593), .Y(n_647) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_619), .A2(n_591), .B1(n_592), .B2(n_582), .Y(n_648) );
INVx2_ASAP7_75t_L g649 ( .A(n_609), .Y(n_649) );
AOI222xp33_ASAP7_75t_L g650 ( .A1(n_614), .A2(n_562), .B1(n_561), .B2(n_554), .C1(n_144), .C2(n_67), .Y(n_650) );
AND4x1_ASAP7_75t_L g651 ( .A(n_626), .B(n_60), .C(n_62), .D(n_63), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_618), .A2(n_144), .B1(n_68), .B2(n_70), .Y(n_652) );
AOI221xp5_ASAP7_75t_L g653 ( .A1(n_599), .A2(n_627), .B1(n_605), .B2(n_622), .C(n_615), .Y(n_653) );
OAI221xp5_ASAP7_75t_L g654 ( .A1(n_606), .A2(n_609), .B1(n_611), .B2(n_613), .C(n_612), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_601), .B(n_608), .Y(n_655) );
AOI221xp5_ASAP7_75t_SL g656 ( .A1(n_624), .A2(n_607), .B1(n_603), .B2(n_617), .C(n_599), .Y(n_656) );
AOI211xp5_ASAP7_75t_L g657 ( .A1(n_629), .A2(n_600), .B(n_610), .C(n_616), .Y(n_657) );
O2A1O1Ixp5_ASAP7_75t_L g658 ( .A1(n_628), .A2(n_617), .B(n_620), .C(n_599), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_655), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_653), .B(n_656), .Y(n_660) );
AND4x1_ASAP7_75t_L g661 ( .A(n_637), .B(n_657), .C(n_658), .D(n_634), .Y(n_661) );
NAND2xp5_ASAP7_75t_SL g662 ( .A(n_640), .B(n_645), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_632), .B(n_642), .Y(n_663) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_654), .B(n_638), .Y(n_664) );
OAI211xp5_ASAP7_75t_L g665 ( .A1(n_660), .A2(n_644), .B(n_634), .C(n_650), .Y(n_665) );
NAND2x1p5_ASAP7_75t_L g666 ( .A(n_661), .B(n_651), .Y(n_666) );
NAND2x1p5_ASAP7_75t_L g667 ( .A(n_662), .B(n_639), .Y(n_667) );
NOR3xp33_ASAP7_75t_L g668 ( .A(n_663), .B(n_636), .C(n_633), .Y(n_668) );
AND2x4_ASAP7_75t_L g669 ( .A(n_668), .B(n_659), .Y(n_669) );
BUFx2_ASAP7_75t_L g670 ( .A(n_666), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_665), .B(n_664), .Y(n_671) );
INVx2_ASAP7_75t_L g672 ( .A(n_670), .Y(n_672) );
INVx2_ASAP7_75t_L g673 ( .A(n_669), .Y(n_673) );
AOI22xp5_ASAP7_75t_L g674 ( .A1(n_672), .A2(n_671), .B1(n_669), .B2(n_667), .Y(n_674) );
OAI22xp5_ASAP7_75t_L g675 ( .A1(n_673), .A2(n_649), .B1(n_646), .B2(n_648), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_674), .Y(n_676) );
AOI21xp5_ASAP7_75t_L g677 ( .A1(n_676), .A2(n_675), .B(n_647), .Y(n_677) );
OAI21xp5_ASAP7_75t_L g678 ( .A1(n_677), .A2(n_635), .B(n_643), .Y(n_678) );
OR2x2_ASAP7_75t_SL g679 ( .A(n_678), .B(n_641), .Y(n_679) );
AOI21xp33_ASAP7_75t_SL g680 ( .A1(n_679), .A2(n_650), .B(n_652), .Y(n_680) );
endmodule