module real_aes_9221_n_286 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_286);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_286;
wire n_480;
wire n_476;
wire n_758;
wire n_887;
wire n_436;
wire n_599;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_905;
wire n_357;
wire n_673;
wire n_386;
wire n_792;
wire n_518;
wire n_635;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_900;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_857;
wire n_461;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_815;
wire n_519;
wire n_638;
wire n_564;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_462;
wire n_289;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_356;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_906;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_505;
wire n_527;
wire n_769;
wire n_434;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_296;
wire n_702;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_723;
wire n_662;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_907;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_290;
wire n_365;
wire n_526;
wire n_637;
wire n_899;
wire n_692;
wire n_544;
wire n_789;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_741;
wire n_314;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_456;
wire n_717;
wire n_359;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_839;
wire n_639;
wire n_587;
wire n_546;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_652;
wire n_703;
wire n_500;
wire n_601;
wire n_307;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_SL g829 ( .A1(n_0), .A2(n_262), .B1(n_808), .B2(n_830), .Y(n_829) );
AOI22xp33_ASAP7_75t_SL g876 ( .A1(n_1), .A2(n_247), .B1(n_759), .B2(n_877), .Y(n_876) );
AOI22xp33_ASAP7_75t_SL g878 ( .A1(n_2), .A2(n_127), .B1(n_423), .B2(n_568), .Y(n_878) );
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_3), .A2(n_102), .B1(n_388), .B2(n_418), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_4), .B(n_449), .Y(n_774) );
AOI22xp5_ASAP7_75t_SL g809 ( .A1(n_5), .A2(n_71), .B1(n_384), .B2(n_414), .Y(n_809) );
CKINVDCx20_ASAP7_75t_R g701 ( .A(n_6), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_7), .A2(n_27), .B1(n_589), .B2(n_627), .Y(n_721) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_8), .A2(n_216), .B1(n_410), .B2(n_414), .Y(n_409) );
AOI22xp33_ASAP7_75t_SL g548 ( .A1(n_9), .A2(n_115), .B1(n_337), .B2(n_549), .Y(n_548) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_10), .A2(n_182), .B1(n_392), .B2(n_394), .Y(n_391) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_11), .A2(n_181), .B1(n_418), .B2(n_679), .Y(n_678) );
AOI211xp5_ASAP7_75t_L g561 ( .A1(n_12), .A2(n_562), .B(n_563), .C(n_569), .Y(n_561) );
XOR2x2_ASAP7_75t_L g513 ( .A(n_13), .B(n_514), .Y(n_513) );
AOI22xp33_ASAP7_75t_SL g880 ( .A1(n_14), .A2(n_229), .B1(n_412), .B2(n_506), .Y(n_880) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_15), .Y(n_739) );
OA22x2_ASAP7_75t_L g401 ( .A1(n_16), .A2(n_402), .B1(n_403), .B2(n_450), .Y(n_401) );
CKINVDCx20_ASAP7_75t_R g402 ( .A(n_16), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_17), .A2(n_29), .B1(n_379), .B2(n_499), .Y(n_498) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_18), .A2(n_196), .B1(n_502), .B2(n_517), .Y(n_516) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_19), .Y(n_486) );
AOI22xp33_ASAP7_75t_SL g406 ( .A1(n_20), .A2(n_241), .B1(n_394), .B2(n_407), .Y(n_406) );
AOI22xp33_ASAP7_75t_SL g551 ( .A1(n_21), .A2(n_270), .B1(n_438), .B2(n_441), .Y(n_551) );
AOI22xp33_ASAP7_75t_SL g575 ( .A1(n_22), .A2(n_152), .B1(n_456), .B2(n_503), .Y(n_575) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_23), .Y(n_769) );
OA22x2_ASAP7_75t_L g477 ( .A1(n_24), .A2(n_478), .B1(n_479), .B2(n_511), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_24), .Y(n_478) );
AOI22xp33_ASAP7_75t_SL g778 ( .A1(n_25), .A2(n_202), .B1(n_472), .B2(n_503), .Y(n_778) );
CKINVDCx20_ASAP7_75t_R g636 ( .A(n_26), .Y(n_636) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_28), .A2(n_239), .B1(n_505), .B2(n_506), .Y(n_504) );
AOI22xp33_ASAP7_75t_SL g819 ( .A1(n_30), .A2(n_157), .B1(n_741), .B2(n_794), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g902 ( .A1(n_31), .A2(n_159), .B1(n_741), .B2(n_794), .Y(n_902) );
CKINVDCx20_ASAP7_75t_R g547 ( .A(n_32), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g753 ( .A1(n_33), .A2(n_45), .B1(n_379), .B2(n_683), .Y(n_753) );
AOI22xp5_ASAP7_75t_L g461 ( .A1(n_34), .A2(n_276), .B1(n_462), .B2(n_463), .Y(n_461) );
AOI22xp5_ASAP7_75t_SL g807 ( .A1(n_35), .A2(n_280), .B1(n_558), .B2(n_808), .Y(n_807) );
AO22x2_ASAP7_75t_L g311 ( .A1(n_36), .A2(n_97), .B1(n_312), .B2(n_313), .Y(n_311) );
INVx1_ASAP7_75t_L g853 ( .A(n_36), .Y(n_853) );
CKINVDCx20_ASAP7_75t_R g631 ( .A(n_37), .Y(n_631) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_38), .A2(n_245), .B1(n_419), .B2(n_502), .C(n_653), .Y(n_652) );
AOI22xp5_ASAP7_75t_L g770 ( .A1(n_39), .A2(n_46), .B1(n_441), .B2(n_616), .Y(n_770) );
AOI22xp33_ASAP7_75t_SL g835 ( .A1(n_40), .A2(n_76), .B1(n_394), .B2(n_836), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_41), .A2(n_111), .B1(n_418), .B2(n_419), .Y(n_417) );
AOI222xp33_ASAP7_75t_L g666 ( .A1(n_42), .A2(n_123), .B1(n_175), .B2(n_549), .C1(n_667), .C2(n_668), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g443 ( .A1(n_43), .A2(n_47), .B1(n_444), .B2(n_447), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g650 ( .A(n_44), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g672 ( .A1(n_48), .A2(n_673), .B1(n_702), .B2(n_703), .Y(n_672) );
INVx1_ASAP7_75t_L g702 ( .A(n_48), .Y(n_702) );
AOI22xp5_ASAP7_75t_SL g803 ( .A1(n_49), .A2(n_155), .B1(n_562), .B2(n_638), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g612 ( .A1(n_50), .A2(n_67), .B1(n_613), .B2(n_614), .Y(n_612) );
AOI22xp33_ASAP7_75t_L g584 ( .A1(n_51), .A2(n_278), .B1(n_432), .B2(n_439), .Y(n_584) );
AOI222xp33_ASAP7_75t_L g722 ( .A1(n_52), .A2(n_142), .B1(n_209), .B2(n_429), .C1(n_613), .C2(n_614), .Y(n_722) );
AOI22xp33_ASAP7_75t_SL g422 ( .A1(n_53), .A2(n_139), .B1(n_423), .B2(n_425), .Y(n_422) );
AO22x2_ASAP7_75t_L g315 ( .A1(n_54), .A2(n_100), .B1(n_312), .B2(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g854 ( .A(n_54), .Y(n_854) );
AOI22xp33_ASAP7_75t_SL g781 ( .A1(n_55), .A2(n_138), .B1(n_392), .B2(n_500), .Y(n_781) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_56), .A2(n_204), .B1(n_384), .B2(n_388), .Y(n_383) );
AOI22xp33_ASAP7_75t_SL g373 ( .A1(n_57), .A2(n_117), .B1(n_374), .B2(n_379), .Y(n_373) );
CKINVDCx20_ASAP7_75t_R g687 ( .A(n_58), .Y(n_687) );
CKINVDCx20_ASAP7_75t_R g901 ( .A(n_59), .Y(n_901) );
CKINVDCx20_ASAP7_75t_R g611 ( .A(n_60), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_61), .B(n_697), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_62), .A2(n_285), .B1(n_389), .B2(n_527), .Y(n_576) );
CKINVDCx20_ASAP7_75t_R g862 ( .A(n_63), .Y(n_862) );
AOI22xp33_ASAP7_75t_SL g823 ( .A1(n_64), .A2(n_91), .B1(n_824), .B2(n_826), .Y(n_823) );
CKINVDCx20_ASAP7_75t_R g661 ( .A(n_65), .Y(n_661) );
CKINVDCx20_ASAP7_75t_R g618 ( .A(n_66), .Y(n_618) );
XNOR2xp5_ASAP7_75t_L g542 ( .A(n_68), .B(n_543), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_69), .A2(n_251), .B1(n_638), .B2(n_677), .Y(n_720) );
OAI22xp5_ASAP7_75t_L g813 ( .A1(n_70), .A2(n_814), .B1(n_815), .B2(n_838), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_70), .Y(n_814) );
AOI22xp33_ASAP7_75t_SL g718 ( .A1(n_72), .A2(n_151), .B1(n_439), .B2(n_463), .Y(n_718) );
CKINVDCx20_ASAP7_75t_R g473 ( .A(n_73), .Y(n_473) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_74), .A2(n_254), .B1(n_508), .B2(n_524), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g482 ( .A(n_75), .Y(n_482) );
AOI22xp33_ASAP7_75t_L g471 ( .A1(n_77), .A2(n_203), .B1(n_366), .B2(n_472), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g894 ( .A(n_78), .Y(n_894) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_79), .B(n_466), .Y(n_465) );
AOI221xp5_ASAP7_75t_L g643 ( .A1(n_80), .A2(n_156), .B1(n_364), .B2(n_644), .C(n_646), .Y(n_643) );
INVx1_ASAP7_75t_L g537 ( .A(n_81), .Y(n_537) );
AOI221xp5_ASAP7_75t_L g658 ( .A1(n_82), .A2(n_160), .B1(n_531), .B2(n_659), .C(n_660), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_83), .A2(n_179), .B1(n_509), .B2(n_527), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_84), .A2(n_230), .B1(n_508), .B2(n_509), .Y(n_507) );
AOI22xp33_ASAP7_75t_SL g800 ( .A1(n_85), .A2(n_263), .B1(n_533), .B2(n_801), .Y(n_800) );
CKINVDCx20_ASAP7_75t_R g619 ( .A(n_86), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_87), .A2(n_171), .B1(n_421), .B2(n_456), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_88), .A2(n_269), .B1(n_338), .B2(n_539), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g433 ( .A(n_89), .Y(n_433) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_90), .A2(n_642), .B1(n_669), .B2(n_670), .Y(n_641) );
INVx1_ASAP7_75t_L g669 ( .A(n_90), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_92), .A2(n_221), .B1(n_442), .B2(n_533), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g525 ( .A1(n_93), .A2(n_141), .B1(n_526), .B2(n_527), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_94), .A2(n_173), .B1(n_683), .B2(n_684), .Y(n_682) );
CKINVDCx20_ASAP7_75t_R g492 ( .A(n_95), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g699 ( .A(n_96), .Y(n_699) );
CKINVDCx20_ASAP7_75t_R g590 ( .A(n_98), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_99), .A2(n_145), .B1(n_384), .B2(n_751), .Y(n_750) );
AOI22xp33_ASAP7_75t_SL g363 ( .A1(n_101), .A2(n_195), .B1(n_364), .B2(n_369), .Y(n_363) );
NAND2xp5_ASAP7_75t_SL g799 ( .A(n_103), .B(n_717), .Y(n_799) );
AOI22xp33_ASAP7_75t_SL g559 ( .A1(n_104), .A2(n_268), .B1(n_407), .B2(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g294 ( .A(n_105), .Y(n_294) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_106), .A2(n_208), .B1(n_374), .B2(n_657), .Y(n_891) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_107), .Y(n_747) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_108), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g655 ( .A(n_109), .Y(n_655) );
CKINVDCx20_ASAP7_75t_R g334 ( .A(n_110), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_112), .A2(n_201), .B1(n_421), .B2(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g292 ( .A(n_113), .Y(n_292) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_114), .A2(n_226), .B1(n_488), .B2(n_489), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_116), .A2(n_131), .B1(n_625), .B2(n_711), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_118), .B(n_568), .Y(n_567) );
CKINVDCx20_ASAP7_75t_R g664 ( .A(n_119), .Y(n_664) );
CKINVDCx20_ASAP7_75t_R g896 ( .A(n_120), .Y(n_896) );
CKINVDCx20_ASAP7_75t_R g342 ( .A(n_121), .Y(n_342) );
CKINVDCx20_ASAP7_75t_R g609 ( .A(n_122), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g890 ( .A1(n_124), .A2(n_205), .B1(n_506), .B2(n_836), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g906 ( .A1(n_125), .A2(n_249), .B1(n_773), .B2(n_907), .Y(n_906) );
CKINVDCx20_ASAP7_75t_R g873 ( .A(n_126), .Y(n_873) );
AOI22xp33_ASAP7_75t_SL g831 ( .A1(n_128), .A2(n_129), .B1(n_568), .B2(n_832), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_130), .A2(n_147), .B1(n_439), .B2(n_539), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_132), .A2(n_224), .B1(n_623), .B2(n_625), .Y(n_622) );
AOI22xp33_ASAP7_75t_SL g437 ( .A1(n_133), .A2(n_161), .B1(n_438), .B2(n_441), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_134), .A2(n_244), .B1(n_557), .B2(n_757), .Y(n_756) );
AOI22xp33_ASAP7_75t_SL g793 ( .A1(n_135), .A2(n_187), .B1(n_616), .B2(n_794), .Y(n_793) );
AOI22xp33_ASAP7_75t_SL g552 ( .A1(n_136), .A2(n_232), .B1(n_466), .B2(n_553), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_137), .A2(n_178), .B1(n_503), .B2(n_713), .Y(n_712) );
AOI22xp33_ASAP7_75t_SL g454 ( .A1(n_140), .A2(n_225), .B1(n_375), .B2(n_393), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_143), .B(n_741), .Y(n_740) );
XOR2x2_ASAP7_75t_L g301 ( .A(n_144), .B(n_302), .Y(n_301) );
CKINVDCx20_ASAP7_75t_R g689 ( .A(n_146), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g881 ( .A1(n_148), .A2(n_227), .B1(n_388), .B2(n_882), .Y(n_881) );
CKINVDCx20_ASAP7_75t_R g872 ( .A(n_149), .Y(n_872) );
XNOR2x2_ASAP7_75t_L g886 ( .A(n_150), .B(n_887), .Y(n_886) );
CKINVDCx20_ASAP7_75t_R g914 ( .A(n_150), .Y(n_914) );
INVx2_ASAP7_75t_L g295 ( .A(n_153), .Y(n_295) );
CKINVDCx20_ASAP7_75t_R g792 ( .A(n_154), .Y(n_792) );
CKINVDCx20_ASAP7_75t_R g897 ( .A(n_158), .Y(n_897) );
INVx1_ASAP7_75t_L g783 ( .A(n_162), .Y(n_783) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_163), .B(n_449), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_164), .B(n_530), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_165), .A2(n_279), .B1(n_374), .B2(n_627), .Y(n_626) );
AND2x6_ASAP7_75t_L g291 ( .A(n_166), .B(n_292), .Y(n_291) );
HB1xp67_ASAP7_75t_L g847 ( .A(n_166), .Y(n_847) );
AO22x2_ASAP7_75t_L g321 ( .A1(n_167), .A2(n_236), .B1(n_312), .B2(n_316), .Y(n_321) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_168), .A2(n_220), .B1(n_502), .B2(n_503), .Y(n_501) );
XOR2xp5_ASAP7_75t_L g856 ( .A(n_169), .B(n_857), .Y(n_856) );
CKINVDCx20_ASAP7_75t_R g322 ( .A(n_170), .Y(n_322) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_172), .Y(n_744) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_174), .A2(n_266), .B1(n_462), .B2(n_463), .Y(n_580) );
AOI22xp33_ASAP7_75t_SL g904 ( .A1(n_176), .A2(n_246), .B1(n_826), .B2(n_905), .Y(n_904) );
AOI22xp5_ASAP7_75t_SL g804 ( .A1(n_177), .A2(n_234), .B1(n_520), .B2(n_805), .Y(n_804) );
CKINVDCx20_ASAP7_75t_R g654 ( .A(n_180), .Y(n_654) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_183), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g865 ( .A(n_184), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_185), .A2(n_223), .B1(n_345), .B2(n_439), .Y(n_468) );
NAND2xp5_ASAP7_75t_SL g822 ( .A(n_186), .B(n_717), .Y(n_822) );
CKINVDCx20_ASAP7_75t_R g893 ( .A(n_188), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_189), .B(n_773), .Y(n_772) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_190), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_191), .A2(n_284), .B1(n_530), .B2(n_531), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g647 ( .A(n_192), .Y(n_647) );
AO22x2_ASAP7_75t_L g319 ( .A1(n_193), .A2(n_253), .B1(n_312), .B2(n_313), .Y(n_319) );
CKINVDCx20_ASAP7_75t_R g695 ( .A(n_194), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_197), .A2(n_282), .B1(n_366), .B2(n_589), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g779 ( .A1(n_198), .A2(n_231), .B1(n_366), .B2(n_412), .Y(n_779) );
AOI22xp5_ASAP7_75t_L g518 ( .A1(n_199), .A2(n_267), .B1(n_519), .B2(n_520), .Y(n_518) );
NAND2xp5_ASAP7_75t_SL g821 ( .A(n_200), .B(n_553), .Y(n_821) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_206), .Y(n_715) );
INVx1_ASAP7_75t_L g810 ( .A(n_207), .Y(n_810) );
CKINVDCx20_ASAP7_75t_R g867 ( .A(n_210), .Y(n_867) );
CKINVDCx20_ASAP7_75t_R g353 ( .A(n_211), .Y(n_353) );
CKINVDCx20_ASAP7_75t_R g564 ( .A(n_212), .Y(n_564) );
AOI22xp33_ASAP7_75t_SL g555 ( .A1(n_213), .A2(n_248), .B1(n_556), .B2(n_557), .Y(n_555) );
AOI22xp33_ASAP7_75t_SL g586 ( .A1(n_214), .A2(n_281), .B1(n_392), .B2(n_587), .Y(n_586) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_215), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_217), .A2(n_250), .B1(n_384), .B2(n_677), .Y(n_676) );
AOI22xp33_ASAP7_75t_SL g837 ( .A1(n_218), .A2(n_219), .B1(n_414), .B2(n_524), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_222), .B(n_449), .Y(n_583) );
CKINVDCx20_ASAP7_75t_R g639 ( .A(n_228), .Y(n_639) );
CKINVDCx20_ASAP7_75t_R g607 ( .A(n_233), .Y(n_607) );
AOI22x1_ASAP7_75t_L g734 ( .A1(n_235), .A2(n_735), .B1(n_760), .B2(n_761), .Y(n_734) );
INVx1_ASAP7_75t_L g760 ( .A(n_235), .Y(n_760) );
NOR2xp33_ASAP7_75t_L g851 ( .A(n_236), .B(n_852), .Y(n_851) );
CKINVDCx20_ASAP7_75t_R g305 ( .A(n_237), .Y(n_305) );
CKINVDCx20_ASAP7_75t_R g430 ( .A(n_238), .Y(n_430) );
CKINVDCx20_ASAP7_75t_R g579 ( .A(n_240), .Y(n_579) );
CKINVDCx20_ASAP7_75t_R g570 ( .A(n_242), .Y(n_570) );
AOI22xp33_ASAP7_75t_SL g470 ( .A1(n_243), .A2(n_283), .B1(n_386), .B2(n_395), .Y(n_470) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_252), .Y(n_459) );
INVx1_ASAP7_75t_L g850 ( .A(n_253), .Y(n_850) );
CKINVDCx20_ASAP7_75t_R g349 ( .A(n_255), .Y(n_349) );
CKINVDCx20_ASAP7_75t_R g435 ( .A(n_256), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_257), .B(n_344), .Y(n_343) );
OA22x2_ASAP7_75t_L g599 ( .A1(n_258), .A2(n_600), .B1(n_601), .B2(n_602), .Y(n_599) );
CKINVDCx16_ASAP7_75t_R g600 ( .A(n_258), .Y(n_600) );
CKINVDCx20_ASAP7_75t_R g818 ( .A(n_259), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_260), .B(n_717), .Y(n_716) );
CKINVDCx20_ASAP7_75t_R g629 ( .A(n_261), .Y(n_629) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_264), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g861 ( .A(n_265), .Y(n_861) );
INVx1_ASAP7_75t_L g312 ( .A(n_271), .Y(n_312) );
INVx1_ASAP7_75t_L g314 ( .A(n_271), .Y(n_314) );
CKINVDCx20_ASAP7_75t_R g693 ( .A(n_272), .Y(n_693) );
CKINVDCx20_ASAP7_75t_R g723 ( .A(n_273), .Y(n_723) );
CKINVDCx20_ASAP7_75t_R g869 ( .A(n_274), .Y(n_869) );
AOI211xp5_ASAP7_75t_L g286 ( .A1(n_275), .A2(n_287), .B(n_296), .C(n_855), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_277), .B(n_798), .Y(n_797) );
CKINVDCx20_ASAP7_75t_R g287 ( .A(n_288), .Y(n_287) );
CKINVDCx20_ASAP7_75t_R g288 ( .A(n_289), .Y(n_288) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x4_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
HB1xp67_ASAP7_75t_L g846 ( .A(n_292), .Y(n_846) );
OAI21xp5_ASAP7_75t_L g912 ( .A1(n_293), .A2(n_845), .B(n_913), .Y(n_912) );
AND2x2_ASAP7_75t_L g293 ( .A(n_294), .B(n_295), .Y(n_293) );
AOI221xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_596), .B1(n_840), .B2(n_841), .C(n_842), .Y(n_296) );
INVx1_ASAP7_75t_L g840 ( .A(n_297), .Y(n_840) );
AOI22xp5_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_299), .B1(n_475), .B2(n_595), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_301), .B1(n_397), .B2(n_398), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_361), .Y(n_302) );
NOR3xp33_ASAP7_75t_L g303 ( .A(n_304), .B(n_328), .C(n_348), .Y(n_303) );
OAI22xp5_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_306), .B1(n_322), .B2(n_323), .Y(n_304) );
INVx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
BUFx6f_ASAP7_75t_L g493 ( .A(n_308), .Y(n_493) );
BUFx3_ASAP7_75t_L g688 ( .A(n_308), .Y(n_688) );
OR2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_317), .Y(n_308) );
INVx2_ASAP7_75t_L g387 ( .A(n_309), .Y(n_387) );
OR2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_315), .Y(n_309) );
AND2x2_ASAP7_75t_L g327 ( .A(n_310), .B(n_315), .Y(n_327) );
AND2x2_ASAP7_75t_L g368 ( .A(n_310), .B(n_347), .Y(n_368) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AND2x2_ASAP7_75t_L g331 ( .A(n_311), .B(n_315), .Y(n_331) );
AND2x2_ASAP7_75t_L g341 ( .A(n_311), .B(n_321), .Y(n_341) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g316 ( .A(n_314), .Y(n_316) );
INVx2_ASAP7_75t_L g347 ( .A(n_315), .Y(n_347) );
INVx1_ASAP7_75t_L g381 ( .A(n_315), .Y(n_381) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NAND2x1p5_ASAP7_75t_L g326 ( .A(n_318), .B(n_327), .Y(n_326) );
AND2x4_ASAP7_75t_L g390 ( .A(n_318), .B(n_368), .Y(n_390) );
AND2x4_ASAP7_75t_L g446 ( .A(n_318), .B(n_387), .Y(n_446) );
AND2x6_ASAP7_75t_L g449 ( .A(n_318), .B(n_327), .Y(n_449) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx1_ASAP7_75t_L g333 ( .A(n_319), .Y(n_333) );
INVx1_ASAP7_75t_L g340 ( .A(n_319), .Y(n_340) );
INVx1_ASAP7_75t_L g360 ( .A(n_319), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_319), .B(n_321), .Y(n_372) );
AND2x2_ASAP7_75t_L g332 ( .A(n_320), .B(n_333), .Y(n_332) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g378 ( .A(n_321), .B(n_360), .Y(n_378) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
BUFx3_ASAP7_75t_L g608 ( .A(n_325), .Y(n_608) );
OAI22xp5_ASAP7_75t_SL g860 ( .A1(n_325), .A2(n_493), .B1(n_861), .B2(n_862), .Y(n_860) );
BUFx3_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g496 ( .A(n_326), .Y(n_496) );
AND2x2_ASAP7_75t_L g377 ( .A(n_327), .B(n_378), .Y(n_377) );
AND2x4_ASAP7_75t_L g393 ( .A(n_327), .B(n_332), .Y(n_393) );
NAND2xp5_ASAP7_75t_SL g566 ( .A(n_327), .B(n_378), .Y(n_566) );
OAI221xp5_ASAP7_75t_L g328 ( .A1(n_329), .A2(n_334), .B1(n_335), .B2(n_342), .C(n_343), .Y(n_328) );
OAI21xp33_ASAP7_75t_L g485 ( .A1(n_329), .A2(n_486), .B(n_487), .Y(n_485) );
OAI221xp5_ASAP7_75t_L g737 ( .A1(n_329), .A2(n_694), .B1(n_738), .B2(n_739), .C(n_740), .Y(n_737) );
OAI21xp5_ASAP7_75t_L g768 ( .A1(n_329), .A2(n_769), .B(n_770), .Y(n_768) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
BUFx6f_ASAP7_75t_L g429 ( .A(n_330), .Y(n_429) );
INVx4_ASAP7_75t_L g460 ( .A(n_330), .Y(n_460) );
BUFx3_ASAP7_75t_L g536 ( .A(n_330), .Y(n_536) );
INVx2_ASAP7_75t_SL g866 ( .A(n_330), .Y(n_866) );
INVx2_ASAP7_75t_L g900 ( .A(n_330), .Y(n_900) );
AND2x6_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
INVx1_ASAP7_75t_L g357 ( .A(n_331), .Y(n_357) );
AND2x4_ASAP7_75t_L g442 ( .A(n_331), .B(n_359), .Y(n_442) );
AND2x2_ASAP7_75t_L g367 ( .A(n_332), .B(n_368), .Y(n_367) );
AND2x6_ASAP7_75t_L g386 ( .A(n_332), .B(n_387), .Y(n_386) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
BUFx3_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g490 ( .A(n_337), .Y(n_490) );
BUFx2_ASAP7_75t_L g697 ( .A(n_337), .Y(n_697) );
BUFx6f_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g434 ( .A(n_338), .Y(n_434) );
BUFx6f_ASAP7_75t_L g462 ( .A(n_338), .Y(n_462) );
BUFx12f_ASAP7_75t_L g616 ( .A(n_338), .Y(n_616) );
AND2x4_ASAP7_75t_L g338 ( .A(n_339), .B(n_341), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g346 ( .A(n_340), .B(n_347), .Y(n_346) );
AND2x4_ASAP7_75t_L g345 ( .A(n_341), .B(n_346), .Y(n_345) );
NAND2x1p5_ASAP7_75t_L g351 ( .A(n_341), .B(n_352), .Y(n_351) );
AND2x4_ASAP7_75t_L g439 ( .A(n_341), .B(n_440), .Y(n_439) );
BUFx2_ASAP7_75t_L g613 ( .A(n_344), .Y(n_613) );
INVx4_ASAP7_75t_L g795 ( .A(n_344), .Y(n_795) );
BUFx6f_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
BUFx4f_ASAP7_75t_SL g432 ( .A(n_345), .Y(n_432) );
BUFx6f_ASAP7_75t_L g488 ( .A(n_345), .Y(n_488) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_345), .Y(n_539) );
INVx1_ASAP7_75t_L g352 ( .A(n_347), .Y(n_352) );
OAI22xp5_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_350), .B1(n_353), .B2(n_354), .Y(n_348) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g481 ( .A1(n_351), .A2(n_482), .B1(n_483), .B2(n_484), .Y(n_481) );
OAI22xp33_ASAP7_75t_SL g617 ( .A1(n_351), .A2(n_354), .B1(n_618), .B2(n_619), .Y(n_617) );
INVx4_ASAP7_75t_L g663 ( .A(n_351), .Y(n_663) );
BUFx3_ASAP7_75t_L g871 ( .A(n_351), .Y(n_871) );
AND2x2_ASAP7_75t_L g456 ( .A(n_352), .B(n_371), .Y(n_456) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_354), .A2(n_699), .B1(n_700), .B2(n_701), .Y(n_698) );
OAI22xp5_ASAP7_75t_SL g870 ( .A1(n_354), .A2(n_871), .B1(n_872), .B2(n_873), .Y(n_870) );
INVx2_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx2_ASAP7_75t_L g484 ( .A(n_355), .Y(n_484) );
CKINVDCx16_ASAP7_75t_R g355 ( .A(n_356), .Y(n_355) );
BUFx2_ASAP7_75t_L g665 ( .A(n_356), .Y(n_665) );
OR2x6_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_362), .B(n_382), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_363), .B(n_373), .Y(n_362) );
INVx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx3_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
BUFx3_ASAP7_75t_L g418 ( .A(n_366), .Y(n_418) );
BUFx6f_ASAP7_75t_L g836 ( .A(n_366), .Y(n_836) );
BUFx3_ASAP7_75t_L g877 ( .A(n_366), .Y(n_877) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
BUFx2_ASAP7_75t_SL g508 ( .A(n_367), .Y(n_508) );
BUFx2_ASAP7_75t_SL g562 ( .A(n_367), .Y(n_562) );
INVx2_ASAP7_75t_L g624 ( .A(n_367), .Y(n_624) );
AND2x4_ASAP7_75t_L g370 ( .A(n_368), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g396 ( .A(n_368), .B(n_378), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_368), .B(n_378), .Y(n_634) );
BUFx2_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g408 ( .A(n_370), .Y(n_408) );
BUFx3_ASAP7_75t_L g472 ( .A(n_370), .Y(n_472) );
BUFx2_ASAP7_75t_SL g506 ( .A(n_370), .Y(n_506) );
BUFx3_ASAP7_75t_L g527 ( .A(n_370), .Y(n_527) );
BUFx3_ASAP7_75t_L g711 ( .A(n_370), .Y(n_711) );
BUFx2_ASAP7_75t_L g808 ( .A(n_370), .Y(n_808) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OR2x6_ASAP7_75t_L g380 ( .A(n_372), .B(n_381), .Y(n_380) );
BUFx6f_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g424 ( .A(n_375), .Y(n_424) );
BUFx2_ASAP7_75t_L g805 ( .A(n_375), .Y(n_805) );
INVx4_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx5_ASAP7_75t_L g500 ( .A(n_376), .Y(n_500) );
INVx2_ASAP7_75t_L g519 ( .A(n_376), .Y(n_519) );
INVx3_ASAP7_75t_L g589 ( .A(n_376), .Y(n_589) );
BUFx3_ASAP7_75t_L g833 ( .A(n_376), .Y(n_833) );
INVx8_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_SL g425 ( .A(n_380), .Y(n_425) );
INVx6_ASAP7_75t_SL g521 ( .A(n_380), .Y(n_521) );
INVx1_ASAP7_75t_SL g568 ( .A(n_380), .Y(n_568) );
INVx1_ASAP7_75t_L g440 ( .A(n_381), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_383), .B(n_391), .Y(n_382) );
INVx2_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
INVx4_ASAP7_75t_L g505 ( .A(n_385), .Y(n_505) );
INVx4_ASAP7_75t_L g524 ( .A(n_385), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g569 ( .A(n_385), .B(n_570), .Y(n_569) );
INVx11_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx11_ASAP7_75t_L g413 ( .A(n_386), .Y(n_413) );
BUFx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
BUFx3_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_390), .Y(n_421) );
INVx2_ASAP7_75t_L g510 ( .A(n_390), .Y(n_510) );
BUFx3_ASAP7_75t_L g526 ( .A(n_390), .Y(n_526) );
BUFx3_ASAP7_75t_L g638 ( .A(n_390), .Y(n_638) );
BUFx3_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx6_ASAP7_75t_L g415 ( .A(n_393), .Y(n_415) );
BUFx3_ASAP7_75t_L g556 ( .A(n_393), .Y(n_556) );
BUFx3_ASAP7_75t_L g759 ( .A(n_393), .Y(n_759) );
BUFx4f_ASAP7_75t_SL g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g883 ( .A(n_395), .Y(n_883) );
BUFx3_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
BUFx3_ASAP7_75t_L g503 ( .A(n_396), .Y(n_503) );
BUFx3_ASAP7_75t_L g517 ( .A(n_396), .Y(n_517) );
BUFx3_ASAP7_75t_L g558 ( .A(n_396), .Y(n_558) );
INVx1_ASAP7_75t_SL g397 ( .A(n_398), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AOI22xp5_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_401), .B1(n_451), .B2(n_474), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g450 ( .A(n_403), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_404), .B(n_426), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_405), .B(n_416), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_406), .B(n_409), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_408), .A2(n_636), .B1(n_637), .B2(n_639), .Y(n_635) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
OAI22xp5_ASAP7_75t_L g892 ( .A1(n_411), .A2(n_420), .B1(n_893), .B2(n_894), .Y(n_892) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx5_ASAP7_75t_SL g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_SL g587 ( .A(n_413), .Y(n_587) );
INVx2_ASAP7_75t_L g625 ( .A(n_413), .Y(n_625) );
INVx4_ASAP7_75t_L g649 ( .A(n_413), .Y(n_649) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g502 ( .A(n_415), .Y(n_502) );
INVx3_ASAP7_75t_L g677 ( .A(n_415), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g895 ( .A1(n_415), .A2(n_632), .B1(n_896), .B2(n_897), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_417), .B(n_422), .Y(n_416) );
INVx4_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx3_ASAP7_75t_L g830 ( .A(n_420), .Y(n_830) );
INVx4_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx3_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g426 ( .A(n_427), .B(n_436), .Y(n_426) );
OAI222xp33_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_430), .B1(n_431), .B2(n_433), .C1(n_434), .C2(n_435), .Y(n_427) );
INVx2_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g546 ( .A(n_429), .Y(n_546) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_437), .B(n_443), .Y(n_436) );
BUFx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
BUFx3_ASAP7_75t_L g533 ( .A(n_439), .Y(n_533) );
INVx1_ASAP7_75t_L g825 ( .A(n_439), .Y(n_825) );
BUFx3_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
BUFx6f_ASAP7_75t_L g463 ( .A(n_442), .Y(n_463) );
BUFx2_ASAP7_75t_SL g801 ( .A(n_442), .Y(n_801) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx5_ASAP7_75t_L g466 ( .A(n_445), .Y(n_466) );
INVx2_ASAP7_75t_L g530 ( .A(n_445), .Y(n_530) );
INVx2_ASAP7_75t_L g773 ( .A(n_445), .Y(n_773) );
INVx4_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_SL g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_SL g798 ( .A(n_448), .Y(n_798) );
INVx1_ASAP7_75t_SL g448 ( .A(n_449), .Y(n_448) );
BUFx4f_ASAP7_75t_L g531 ( .A(n_449), .Y(n_531) );
BUFx2_ASAP7_75t_L g553 ( .A(n_449), .Y(n_553) );
BUFx2_ASAP7_75t_L g907 ( .A(n_449), .Y(n_907) );
INVx3_ASAP7_75t_L g474 ( .A(n_451), .Y(n_474) );
XOR2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_473), .Y(n_451) );
NAND3x1_ASAP7_75t_SL g452 ( .A(n_453), .B(n_457), .C(n_469), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
NOR2x1_ASAP7_75t_L g457 ( .A(n_458), .B(n_464), .Y(n_457) );
OAI21xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_460), .B(n_461), .Y(n_458) );
OAI21xp5_ASAP7_75t_L g578 ( .A1(n_460), .A2(n_579), .B(n_580), .Y(n_578) );
INVx4_ASAP7_75t_L g667 ( .A(n_460), .Y(n_667) );
BUFx2_ASAP7_75t_L g692 ( .A(n_460), .Y(n_692) );
OAI21xp5_ASAP7_75t_SL g791 ( .A1(n_460), .A2(n_792), .B(n_793), .Y(n_791) );
BUFx4f_ASAP7_75t_L g741 ( .A(n_462), .Y(n_741) );
INVx1_ASAP7_75t_SL g827 ( .A(n_463), .Y(n_827) );
NAND3xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_467), .C(n_468), .Y(n_464) );
BUFx6f_ASAP7_75t_L g717 ( .A(n_466), .Y(n_717) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_471), .Y(n_469) );
INVx2_ASAP7_75t_L g752 ( .A(n_472), .Y(n_752) );
INVx1_ASAP7_75t_L g595 ( .A(n_475), .Y(n_595) );
AOI22xp5_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_477), .B1(n_512), .B2(n_594), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g511 ( .A(n_479), .Y(n_511) );
NAND2x1_ASAP7_75t_L g479 ( .A(n_480), .B(n_497), .Y(n_479) );
NOR3xp33_ASAP7_75t_SL g480 ( .A(n_481), .B(n_485), .C(n_491), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g745 ( .A1(n_484), .A2(n_700), .B1(n_746), .B2(n_747), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g694 ( .A(n_488), .Y(n_694) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
OAI22xp5_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_493), .B1(n_494), .B2(n_495), .Y(n_491) );
INVx1_ASAP7_75t_L g606 ( .A(n_493), .Y(n_606) );
OA211x2_ASAP7_75t_L g714 ( .A1(n_495), .A2(n_715), .B(n_716), .C(n_718), .Y(n_714) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g690 ( .A(n_496), .Y(n_690) );
AND4x1_ASAP7_75t_L g497 ( .A(n_498), .B(n_501), .C(n_504), .D(n_507), .Y(n_497) );
BUFx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
BUFx6f_ASAP7_75t_L g683 ( .A(n_500), .Y(n_683) );
INVx2_ASAP7_75t_L g630 ( .A(n_502), .Y(n_630) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g594 ( .A(n_512), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_540), .B1(n_541), .B2(n_593), .Y(n_512) );
INVx1_ASAP7_75t_SL g593 ( .A(n_513), .Y(n_593) );
NOR4xp75_ASAP7_75t_L g514 ( .A(n_515), .B(n_522), .C(n_528), .D(n_534), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_516), .B(n_518), .Y(n_515) );
BUFx3_ASAP7_75t_L g679 ( .A(n_517), .Y(n_679) );
BUFx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
BUFx2_ASAP7_75t_L g627 ( .A(n_521), .Y(n_627) );
BUFx2_ASAP7_75t_L g657 ( .A(n_521), .Y(n_657) );
BUFx4f_ASAP7_75t_SL g684 ( .A(n_521), .Y(n_684) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_523), .B(n_525), .Y(n_522) );
BUFx2_ASAP7_75t_L g560 ( .A(n_526), .Y(n_560) );
INVx1_ASAP7_75t_L g651 ( .A(n_527), .Y(n_651) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_529), .B(n_532), .Y(n_528) );
BUFx2_ASAP7_75t_L g659 ( .A(n_530), .Y(n_659) );
OAI21xp5_ASAP7_75t_SL g534 ( .A1(n_535), .A2(n_537), .B(n_538), .Y(n_534) );
OAI21xp33_ASAP7_75t_SL g610 ( .A1(n_535), .A2(n_611), .B(n_612), .Y(n_610) );
INVx3_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_539), .Y(n_549) );
INVx1_ASAP7_75t_SL g540 ( .A(n_541), .Y(n_540) );
OAI22x1_ASAP7_75t_L g541 ( .A1(n_542), .A2(n_571), .B1(n_591), .B2(n_592), .Y(n_541) );
INVx1_ASAP7_75t_L g591 ( .A(n_542), .Y(n_591) );
NAND3x1_ASAP7_75t_L g543 ( .A(n_544), .B(n_554), .C(n_561), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_545), .B(n_550), .Y(n_544) );
OAI21xp5_ASAP7_75t_SL g545 ( .A1(n_546), .A2(n_547), .B(n_548), .Y(n_545) );
OAI21xp5_ASAP7_75t_SL g817 ( .A1(n_546), .A2(n_818), .B(n_819), .Y(n_817) );
INVx2_ASAP7_75t_SL g864 ( .A(n_549), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
AND2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_559), .Y(n_554) );
BUFx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g645 ( .A(n_558), .Y(n_645) );
OAI21xp33_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_565), .B(n_567), .Y(n_563) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_565), .A2(n_654), .B1(n_655), .B2(n_656), .Y(n_653) );
BUFx2_ASAP7_75t_R g565 ( .A(n_566), .Y(n_565) );
INVx1_ASAP7_75t_L g592 ( .A(n_571), .Y(n_592) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
XOR2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_590), .Y(n_572) );
NAND3x1_ASAP7_75t_L g573 ( .A(n_574), .B(n_577), .C(n_585), .Y(n_573) );
AND2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
NOR2x1_ASAP7_75t_L g577 ( .A(n_578), .B(n_581), .Y(n_577) );
NAND3xp33_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .C(n_584), .Y(n_581) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_588), .Y(n_585) );
INVx1_ASAP7_75t_L g841 ( .A(n_596), .Y(n_841) );
XOR2xp5_ASAP7_75t_L g596 ( .A(n_597), .B(n_729), .Y(n_596) );
AOI22xp5_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_640), .B1(n_727), .B2(n_728), .Y(n_597) );
INVx2_ASAP7_75t_L g727 ( .A(n_598), .Y(n_727) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_620), .Y(n_602) );
NOR3xp33_ASAP7_75t_L g603 ( .A(n_604), .B(n_610), .C(n_617), .Y(n_603) );
OAI22xp5_ASAP7_75t_SL g604 ( .A1(n_605), .A2(n_607), .B1(n_608), .B2(n_609), .Y(n_604) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx3_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
BUFx4f_ASAP7_75t_SL g668 ( .A(n_616), .Y(n_668) );
NOR3xp33_ASAP7_75t_L g620 ( .A(n_621), .B(n_628), .C(n_635), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_622), .B(n_626), .Y(n_621) );
INVx3_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx3_ASAP7_75t_L g713 ( .A(n_624), .Y(n_713) );
OAI22xp5_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_630), .B1(n_631), .B2(n_632), .Y(n_628) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g728 ( .A(n_640), .Y(n_728) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_671), .B1(n_725), .B2(n_726), .Y(n_640) );
INVx1_ASAP7_75t_L g725 ( .A(n_641), .Y(n_725) );
INVx1_ASAP7_75t_L g670 ( .A(n_642), .Y(n_670) );
AND4x2_ASAP7_75t_L g642 ( .A(n_643), .B(n_652), .C(n_658), .D(n_666), .Y(n_642) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_647), .A2(n_648), .B1(n_650), .B2(n_651), .Y(n_646) );
INVx1_ASAP7_75t_SL g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
OAI22xp5_ASAP7_75t_L g660 ( .A1(n_661), .A2(n_662), .B1(n_664), .B2(n_665), .Y(n_660) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx3_ASAP7_75t_SL g700 ( .A(n_663), .Y(n_700) );
INVx1_ASAP7_75t_L g726 ( .A(n_671), .Y(n_726) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_704), .B1(n_705), .B2(n_724), .Y(n_671) );
INVx1_ASAP7_75t_L g724 ( .A(n_672), .Y(n_724) );
INVx1_ASAP7_75t_SL g703 ( .A(n_673), .Y(n_703) );
AND2x2_ASAP7_75t_SL g673 ( .A(n_674), .B(n_685), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g674 ( .A(n_675), .B(n_680), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_676), .B(n_678), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_681), .B(n_682), .Y(n_680) );
NOR3xp33_ASAP7_75t_L g685 ( .A(n_686), .B(n_691), .C(n_698), .Y(n_685) );
OAI22xp5_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_688), .B1(n_689), .B2(n_690), .Y(n_686) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_688), .A2(n_690), .B1(n_743), .B2(n_744), .Y(n_742) );
OAI221xp5_ASAP7_75t_L g691 ( .A1(n_692), .A2(n_693), .B1(n_694), .B2(n_695), .C(n_696), .Y(n_691) );
INVx1_ASAP7_75t_L g704 ( .A(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
XOR2x2_ASAP7_75t_L g707 ( .A(n_708), .B(n_723), .Y(n_707) );
NAND4xp75_ASAP7_75t_L g708 ( .A(n_709), .B(n_714), .C(n_719), .D(n_722), .Y(n_708) );
AND2x2_ASAP7_75t_L g709 ( .A(n_710), .B(n_712), .Y(n_709) );
AND2x2_ASAP7_75t_L g719 ( .A(n_720), .B(n_721), .Y(n_719) );
XNOR2xp5_ASAP7_75t_L g729 ( .A(n_730), .B(n_785), .Y(n_729) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
AOI22xp5_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_762), .B1(n_763), .B2(n_784), .Y(n_733) );
INVx1_ASAP7_75t_L g784 ( .A(n_734), .Y(n_784) );
INVx2_ASAP7_75t_SL g761 ( .A(n_735), .Y(n_761) );
AND2x4_ASAP7_75t_L g735 ( .A(n_736), .B(n_748), .Y(n_735) );
NOR3xp33_ASAP7_75t_SL g736 ( .A(n_737), .B(n_742), .C(n_745), .Y(n_736) );
INVx1_ASAP7_75t_L g868 ( .A(n_741), .Y(n_868) );
NOR2x1_ASAP7_75t_L g748 ( .A(n_749), .B(n_754), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_750), .B(n_753), .Y(n_749) );
INVx2_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_755), .B(n_756), .Y(n_754) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx3_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx2_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
XOR2x2_ASAP7_75t_L g765 ( .A(n_766), .B(n_783), .Y(n_765) );
NAND2x1p5_ASAP7_75t_L g766 ( .A(n_767), .B(n_776), .Y(n_766) );
NOR2xp33_ASAP7_75t_L g767 ( .A(n_768), .B(n_771), .Y(n_767) );
NAND3xp33_ASAP7_75t_L g771 ( .A(n_772), .B(n_774), .C(n_775), .Y(n_771) );
NOR2x1_ASAP7_75t_L g776 ( .A(n_777), .B(n_780), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_778), .B(n_779), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_781), .B(n_782), .Y(n_780) );
AOI22xp5_ASAP7_75t_L g785 ( .A1(n_786), .A2(n_787), .B1(n_811), .B2(n_839), .Y(n_785) );
INVx2_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
HB1xp67_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
XOR2x2_ASAP7_75t_L g788 ( .A(n_789), .B(n_810), .Y(n_788) );
NAND3x1_ASAP7_75t_L g789 ( .A(n_790), .B(n_802), .C(n_806), .Y(n_789) );
NOR2x1_ASAP7_75t_L g790 ( .A(n_791), .B(n_796), .Y(n_790) );
INVx3_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
NAND3xp33_ASAP7_75t_L g796 ( .A(n_797), .B(n_799), .C(n_800), .Y(n_796) );
AND2x2_ASAP7_75t_L g802 ( .A(n_803), .B(n_804), .Y(n_802) );
AND2x2_ASAP7_75t_L g806 ( .A(n_807), .B(n_809), .Y(n_806) );
INVx2_ASAP7_75t_L g839 ( .A(n_811), .Y(n_839) );
BUFx2_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g838 ( .A(n_815), .Y(n_838) );
NAND3x1_ASAP7_75t_L g815 ( .A(n_816), .B(n_828), .C(n_834), .Y(n_815) );
NOR2x1_ASAP7_75t_L g816 ( .A(n_817), .B(n_820), .Y(n_816) );
NAND3xp33_ASAP7_75t_L g820 ( .A(n_821), .B(n_822), .C(n_823), .Y(n_820) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g905 ( .A(n_825), .Y(n_905) );
INVx2_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
AND2x2_ASAP7_75t_L g828 ( .A(n_829), .B(n_831), .Y(n_828) );
INVx3_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
AND2x2_ASAP7_75t_L g834 ( .A(n_835), .B(n_837), .Y(n_834) );
INVx2_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
NOR2x1_ASAP7_75t_L g843 ( .A(n_844), .B(n_848), .Y(n_843) );
OR2x2_ASAP7_75t_SL g910 ( .A(n_844), .B(n_849), .Y(n_910) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_845), .B(n_847), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_845), .B(n_885), .Y(n_884) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g913 ( .A(n_846), .B(n_885), .Y(n_913) );
CKINVDCx16_ASAP7_75t_R g885 ( .A(n_847), .Y(n_885) );
CKINVDCx20_ASAP7_75t_R g848 ( .A(n_849), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g849 ( .A(n_850), .B(n_851), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_853), .B(n_854), .Y(n_852) );
OAI222xp33_ASAP7_75t_L g855 ( .A1(n_856), .A2(n_884), .B1(n_886), .B2(n_908), .C1(n_911), .C2(n_914), .Y(n_855) );
HB1xp67_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
AND2x2_ASAP7_75t_L g858 ( .A(n_859), .B(n_874), .Y(n_858) );
NOR3xp33_ASAP7_75t_L g859 ( .A(n_860), .B(n_863), .C(n_870), .Y(n_859) );
OAI222xp33_ASAP7_75t_L g863 ( .A1(n_864), .A2(n_865), .B1(n_866), .B2(n_867), .C1(n_868), .C2(n_869), .Y(n_863) );
NOR2xp33_ASAP7_75t_L g874 ( .A(n_875), .B(n_879), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_876), .B(n_878), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g879 ( .A(n_880), .B(n_881), .Y(n_879) );
INVx1_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
NAND2xp5_ASAP7_75t_SL g887 ( .A(n_888), .B(n_898), .Y(n_887) );
NOR3xp33_ASAP7_75t_L g888 ( .A(n_889), .B(n_892), .C(n_895), .Y(n_888) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_890), .B(n_891), .Y(n_889) );
NOR2xp33_ASAP7_75t_L g898 ( .A(n_899), .B(n_903), .Y(n_898) );
OAI21xp5_ASAP7_75t_SL g899 ( .A1(n_900), .A2(n_901), .B(n_902), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g903 ( .A(n_904), .B(n_906), .Y(n_903) );
CKINVDCx20_ASAP7_75t_R g908 ( .A(n_909), .Y(n_908) );
CKINVDCx20_ASAP7_75t_R g909 ( .A(n_910), .Y(n_909) );
CKINVDCx16_ASAP7_75t_R g911 ( .A(n_912), .Y(n_911) );
endmodule