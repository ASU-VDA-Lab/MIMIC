module fake_jpeg_23515_n_259 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_259);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_259;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

INVx2_ASAP7_75t_SL g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_18),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_34),
.B(n_35),
.Y(n_43)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_20),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_40),
.Y(n_46)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_42),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_40),
.A2(n_30),
.B1(n_28),
.B2(n_32),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_47),
.A2(n_52),
.B(n_33),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_32),
.C(n_31),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_39),
.C(n_35),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_34),
.B(n_21),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_49),
.B(n_51),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_34),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_50),
.A2(n_19),
.B1(n_30),
.B2(n_32),
.Y(n_56)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_40),
.A2(n_19),
.B1(n_30),
.B2(n_17),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_24),
.Y(n_54)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_24),
.Y(n_55)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_56),
.A2(n_72),
.B1(n_80),
.B2(n_81),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_42),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_57),
.B(n_61),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVxp67_ASAP7_75t_SL g97 ( 
.A(n_59),
.Y(n_97)
);

NOR4xp25_ASAP7_75t_SL g60 ( 
.A(n_49),
.B(n_34),
.C(n_36),
.D(n_15),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_60),
.A2(n_25),
.B(n_23),
.C(n_27),
.Y(n_98)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_54),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_65),
.B(n_68),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_21),
.Y(n_66)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_55),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_34),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_69),
.B(n_76),
.Y(n_86)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_71),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_41),
.A2(n_19),
.B1(n_16),
.B2(n_17),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_21),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_73),
.B(n_79),
.Y(n_95)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx13_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_46),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_75),
.B(n_45),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_37),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_77),
.B(n_85),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_20),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_41),
.A2(n_19),
.B1(n_16),
.B2(n_24),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_48),
.B(n_35),
.C(n_36),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_76),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_89),
.A2(n_90),
.B1(n_92),
.B2(n_22),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_65),
.B(n_29),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_68),
.B(n_29),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_71),
.A2(n_80),
.B1(n_78),
.B2(n_84),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_94),
.A2(n_100),
.B1(n_106),
.B2(n_58),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_98),
.A2(n_69),
.B(n_83),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_38),
.C(n_25),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_77),
.A2(n_50),
.B1(n_48),
.B2(n_33),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_67),
.B(n_45),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_102),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_67),
.B(n_45),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_58),
.B(n_51),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_38),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_75),
.A2(n_37),
.B1(n_16),
.B2(n_17),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_111),
.A2(n_64),
.B(n_102),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_86),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_113),
.A2(n_119),
.B1(n_121),
.B2(n_133),
.Y(n_147)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_117),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_115),
.A2(n_123),
.B(n_124),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_110),
.B(n_61),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_116),
.Y(n_155)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_88),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_125),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_87),
.A2(n_69),
.B1(n_19),
.B2(n_82),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_103),
.A2(n_70),
.B1(n_74),
.B2(n_37),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_120),
.A2(n_126),
.B1(n_109),
.B2(n_108),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_107),
.A2(n_85),
.B1(n_27),
.B2(n_23),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_110),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_122),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_94),
.A2(n_62),
.B(n_59),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_88),
.A2(n_29),
.B(n_22),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_97),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_98),
.A2(n_38),
.B1(n_22),
.B2(n_26),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_101),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_129),
.Y(n_150)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_106),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_131),
.Y(n_160)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_95),
.Y(n_132)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_132),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_87),
.A2(n_57),
.B1(n_38),
.B2(n_26),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_95),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_134),
.B(n_136),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_135),
.B(n_96),
.C(n_25),
.Y(n_162)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_90),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_25),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_R g139 ( 
.A(n_112),
.B(n_86),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_139),
.A2(n_151),
.B(n_127),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_113),
.A2(n_107),
.B1(n_99),
.B2(n_100),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_140),
.B(n_146),
.Y(n_183)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_120),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_141),
.B(n_149),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_144),
.B(n_162),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_119),
.A2(n_107),
.B1(n_86),
.B2(n_91),
.Y(n_146)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_136),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_130),
.A2(n_93),
.B1(n_92),
.B2(n_57),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_123),
.A2(n_93),
.B1(n_108),
.B2(n_109),
.Y(n_153)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_153),
.Y(n_166)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_154),
.B(n_157),
.Y(n_187)
);

OA21x2_ASAP7_75t_L g156 ( 
.A1(n_133),
.A2(n_26),
.B(n_109),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_156),
.A2(n_158),
.B(n_20),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_115),
.A2(n_20),
.B(n_25),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_164),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_118),
.A2(n_96),
.B1(n_104),
.B2(n_27),
.Y(n_161)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_161),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_163),
.C(n_141),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_96),
.C(n_63),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_165),
.A2(n_170),
.B(n_176),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_126),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_167),
.A2(n_148),
.B(n_156),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_131),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_168),
.B(n_181),
.Y(n_203)
);

NAND5xp2_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_160),
.C(n_142),
.D(n_158),
.E(n_150),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_145),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_171),
.B(n_172),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_143),
.B(n_137),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_154),
.B(n_114),
.Y(n_173)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_173),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_155),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_174),
.Y(n_191)
);

NAND5xp2_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_159),
.C(n_146),
.D(n_152),
.E(n_151),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_134),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_177),
.B(n_179),
.Y(n_198)
);

NOR4xp25_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_125),
.C(n_124),
.D(n_129),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_20),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_164),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_180),
.B(n_186),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_25),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_157),
.C(n_138),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_23),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_166),
.A2(n_153),
.B1(n_148),
.B2(n_138),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_188),
.A2(n_202),
.B1(n_175),
.B2(n_184),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_190),
.B(n_204),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g192 ( 
.A(n_187),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_192),
.B(n_167),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_194),
.C(n_195),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_185),
.B(n_156),
.C(n_104),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_104),
.C(n_25),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_199),
.Y(n_205)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_180),
.A2(n_27),
.B1(n_23),
.B2(n_20),
.Y(n_202)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_206),
.Y(n_222)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_198),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_208),
.B(n_209),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_177),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_193),
.A2(n_183),
.B(n_173),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_203),
.C(n_190),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_200),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_211),
.A2(n_214),
.B1(n_215),
.B2(n_219),
.Y(n_220)
);

NOR2xp67_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_176),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_212),
.B(n_218),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_194),
.A2(n_197),
.B1(n_195),
.B2(n_170),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_201),
.A2(n_165),
.B(n_169),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_168),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_217),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_204),
.B(n_181),
.Y(n_217)
);

AOI322xp5_ASAP7_75t_SL g218 ( 
.A1(n_189),
.A2(n_167),
.A3(n_186),
.B1(n_169),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_224),
.B(n_226),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_215),
.B(n_188),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_227),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_202),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_207),
.C(n_217),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_213),
.B(n_191),
.C(n_2),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_229),
.A2(n_211),
.B(n_207),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_0),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_230),
.B(n_3),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_9),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_232),
.B(n_233),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_3),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_229),
.B(n_223),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_234),
.B(n_9),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_220),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_8),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_222),
.A2(n_226),
.B1(n_227),
.B2(n_221),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_237),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_221),
.A2(n_5),
.B(n_6),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_238),
.A2(n_14),
.B(n_11),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_236),
.C(n_12),
.Y(n_250)
);

OAI21x1_ASAP7_75t_L g241 ( 
.A1(n_238),
.A2(n_7),
.B(n_8),
.Y(n_241)
);

AND2x4_ASAP7_75t_SL g247 ( 
.A(n_241),
.B(n_246),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_243),
.B(n_244),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_245),
.B(n_10),
.Y(n_248)
);

AO21x1_ASAP7_75t_L g253 ( 
.A1(n_248),
.A2(n_249),
.B(n_11),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_243),
.A2(n_239),
.B(n_235),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_250),
.A2(n_242),
.B(n_12),
.Y(n_252)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_252),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_253),
.A2(n_254),
.B1(n_251),
.B2(n_13),
.Y(n_255)
);

A2O1A1Ixp33_ASAP7_75t_SL g254 ( 
.A1(n_247),
.A2(n_11),
.B(n_13),
.C(n_14),
.Y(n_254)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_255),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_257),
.B(n_256),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_258),
.B(n_14),
.Y(n_259)
);


endmodule