module real_jpeg_20482_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_268;
wire n_42;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_258;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_216;
wire n_202;
wire n_167;
wire n_128;
wire n_179;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_256;
wire n_101;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_0),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_0),
.A2(n_30),
.B1(n_36),
.B2(n_37),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_1),
.A2(n_64),
.B1(n_70),
.B2(n_75),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_1),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_1),
.A2(n_52),
.B1(n_54),
.B2(n_75),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_1),
.A2(n_36),
.B1(n_37),
.B2(n_75),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_75),
.Y(n_218)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_2),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_3),
.A2(n_64),
.B1(n_70),
.B2(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_3),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_3),
.A2(n_52),
.B1(n_54),
.B2(n_92),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_3),
.A2(n_36),
.B1(n_37),
.B2(n_92),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_92),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_4),
.Y(n_140)
);

AOI21xp33_ASAP7_75t_L g141 ( 
.A1(n_4),
.A2(n_52),
.B(n_142),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_4),
.A2(n_64),
.B1(n_70),
.B2(n_140),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_4),
.B(n_73),
.Y(n_190)
);

A2O1A1O1Ixp25_ASAP7_75t_L g201 ( 
.A1(n_4),
.A2(n_36),
.B(n_40),
.C(n_202),
.D(n_203),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_4),
.B(n_36),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_4),
.B(n_58),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_4),
.A2(n_25),
.B(n_217),
.Y(n_234)
);

A2O1A1O1Ixp25_ASAP7_75t_L g247 ( 
.A1(n_4),
.A2(n_54),
.B(n_55),
.C(n_151),
.D(n_248),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_4),
.B(n_54),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_5),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_5),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_5),
.A2(n_36),
.B1(n_37),
.B2(n_53),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_5),
.A2(n_53),
.B1(n_64),
.B2(n_70),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_53),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_6),
.B(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_6),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_6),
.A2(n_26),
.B1(n_145),
.B2(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_6),
.B(n_218),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_7),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_35)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_7),
.A2(n_38),
.B1(n_52),
.B2(n_54),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_38),
.Y(n_145)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_9),
.A2(n_36),
.B1(n_37),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_46),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_9),
.A2(n_46),
.B1(n_52),
.B2(n_54),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_10),
.A2(n_64),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_10),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_10),
.A2(n_52),
.B1(n_54),
.B2(n_71),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_71),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_10),
.A2(n_36),
.B1(n_37),
.B2(n_71),
.Y(n_246)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_12),
.A2(n_33),
.B1(n_36),
.B2(n_37),
.Y(n_108)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

INVx13_ASAP7_75t_L g66 ( 
.A(n_14),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_14),
.A2(n_52),
.B1(n_54),
.B2(n_66),
.Y(n_68)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_127),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_125),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_100),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_20),
.B(n_100),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_76),
.C(n_83),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_21),
.A2(n_22),
.B1(n_76),
.B2(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_48),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_23),
.B(n_50),
.C(n_61),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_34),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_24),
.B(n_34),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_25),
.A2(n_32),
.B(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_25),
.A2(n_29),
.B1(n_31),
.B2(n_86),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_25),
.A2(n_31),
.B1(n_86),
.B2(n_144),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_25),
.A2(n_216),
.B(n_217),
.Y(n_215)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_26),
.A2(n_222),
.B1(n_224),
.B2(n_225),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_26),
.B(n_218),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_27),
.A2(n_28),
.B1(n_41),
.B2(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_27),
.B(n_41),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_27),
.B(n_236),
.Y(n_235)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_28),
.A2(n_42),
.B1(n_206),
.B2(n_207),
.Y(n_205)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_31),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_39),
.B1(n_45),
.B2(n_47),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_35),
.A2(n_39),
.B1(n_47),
.B2(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_36),
.A2(n_37),
.B1(n_56),
.B2(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_36),
.B(n_56),
.Y(n_254)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

O2A1O1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_37),
.A2(n_41),
.B(n_42),
.C(n_43),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_41),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_37),
.A2(n_57),
.B1(n_253),
.B2(n_254),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_39),
.A2(n_45),
.B1(n_47),
.B2(n_81),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_39),
.A2(n_47),
.B1(n_214),
.B2(n_246),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_39),
.A2(n_246),
.B(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_40),
.A2(n_43),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_40),
.B(n_167),
.Y(n_166)
);

CKINVDCx9p33_ASAP7_75t_R g44 ( 
.A(n_41),
.Y(n_44)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_47),
.A2(n_88),
.B(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_47),
.B(n_168),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_47),
.A2(n_166),
.B(n_214),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_47),
.B(n_140),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_61),
.B2(n_62),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_55),
.B1(n_58),
.B2(n_60),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_51),
.Y(n_95)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_SL g55 ( 
.A1(n_52),
.A2(n_56),
.B(n_57),
.C(n_58),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_56),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_55),
.B(n_98),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_55),
.A2(n_58),
.B1(n_60),
.B2(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_55),
.Y(n_149)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_69),
.B(n_72),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_63),
.A2(n_68),
.B1(n_69),
.B2(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_63),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_66),
.B(n_67),
.C(n_68),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_66),
.Y(n_67)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_64),
.A2(n_66),
.B(n_140),
.C(n_141),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_66),
.Y(n_142)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_68),
.A2(n_119),
.B(n_120),
.Y(n_118)
);

OAI21xp33_ASAP7_75t_L g136 ( 
.A1(n_68),
.A2(n_91),
.B(n_120),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_72),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_74),
.B(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_76),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_78),
.B1(n_80),
.B2(n_82),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_77),
.A2(n_78),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_78),
.B(n_80),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_79),
.A2(n_223),
.B(n_232),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_79),
.B(n_140),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_79),
.A2(n_232),
.B(n_256),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_80),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_81),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_83),
.B(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_89),
.C(n_93),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_84),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_87),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_85),
.B(n_87),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_89),
.A2(n_90),
.B1(n_93),
.B2(n_94),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_96),
.B(n_97),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_96),
.B(n_99),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_96),
.A2(n_148),
.B1(n_149),
.B2(n_174),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_96),
.A2(n_97),
.B(n_174),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_123),
.B2(n_124),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_112),
.B2(n_113),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_109),
.B(n_111),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_105),
.B(n_109),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_116),
.B2(n_122),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_116),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_121),
.A2(n_170),
.B(n_171),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g124 ( 
.A(n_123),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_155),
.B(n_280),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_152),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_129),
.B(n_152),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.C(n_133),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_130),
.B(n_132),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_133),
.A2(n_134),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_137),
.C(n_146),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_135),
.A2(n_136),
.B1(n_146),
.B2(n_147),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_143),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_138),
.A2(n_139),
.B1(n_143),
.B2(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_143),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B(n_150),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_194),
.Y(n_155)
);

INVxp33_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

AOI21xp33_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_178),
.B(n_193),
.Y(n_157)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_158),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_175),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_159),
.B(n_175),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.C(n_163),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_163),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_169),
.C(n_172),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_164),
.A2(n_165),
.B1(n_172),
.B2(n_173),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_183),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_179),
.B(n_181),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_184),
.C(n_186),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_182),
.B(n_275),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_184),
.A2(n_186),
.B1(n_187),
.B2(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_184),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_187),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_190),
.C(n_191),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_188),
.A2(n_189),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_190),
.B(n_191),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_192),
.Y(n_256)
);

NOR3xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_278),
.C(n_279),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_272),
.B(n_277),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_259),
.B(n_271),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_240),
.B(n_258),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_219),
.B(n_239),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_208),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_200),
.B(n_208),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_204),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_201),
.A2(n_204),
.B1(n_205),
.B2(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_201),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_202),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_203),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_215),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_211),
.B1(n_212),
.B2(n_213),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_210),
.B(n_213),
.C(n_215),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_216),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_228),
.B(n_238),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_226),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_221),
.B(n_226),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_233),
.B(n_237),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_230),
.B(n_231),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_241),
.B(n_242),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_251),
.B2(n_257),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_245),
.A2(n_247),
.B1(n_249),
.B2(n_250),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_245),
.Y(n_250)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_247),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_247),
.B(n_250),
.C(n_257),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_248),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_251),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_255),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_255),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_261),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_260),
.B(n_261),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_265),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_267),
.C(n_269),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_263),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_269),
.B2(n_270),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_266),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_267),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_273),
.B(n_274),
.Y(n_277)
);


endmodule