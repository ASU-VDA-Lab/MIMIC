module fake_jpeg_8858_n_206 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_206);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_1),
.B(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_SL g20 ( 
.A(n_2),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_20),
.Y(n_33)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_39),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_19),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_40),
.B(n_41),
.Y(n_45)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_43),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_17),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx4f_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_16),
.Y(n_54)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_35),
.A2(n_21),
.B1(n_25),
.B2(n_29),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_55),
.A2(n_59),
.B1(n_23),
.B2(n_29),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_32),
.Y(n_56)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_56),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_58),
.B(n_22),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_35),
.A2(n_21),
.B1(n_17),
.B2(n_19),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_22),
.Y(n_61)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_62),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_33),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_34),
.B(n_23),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_64),
.A2(n_26),
.B(n_27),
.C(n_28),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_55),
.A2(n_43),
.B1(n_21),
.B2(n_38),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_65),
.A2(n_83),
.B1(n_60),
.B2(n_51),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_67),
.A2(n_28),
.B(n_31),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_69),
.Y(n_89)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_50),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_73),
.B(n_75),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_58),
.B(n_44),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_81),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_45),
.B(n_31),
.Y(n_80)
);

AOI32xp33_ASAP7_75t_L g87 ( 
.A1(n_80),
.A2(n_64),
.A3(n_46),
.B1(n_44),
.B2(n_60),
.Y(n_87)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_61),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_85),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_53),
.A2(n_43),
.B1(n_30),
.B2(n_42),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_53),
.A2(n_26),
.B1(n_24),
.B2(n_18),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_84),
.A2(n_50),
.B1(n_33),
.B2(n_42),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_54),
.B(n_0),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_27),
.Y(n_120)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_88),
.B(n_97),
.Y(n_109)
);

AND2x2_ASAP7_75t_SL g90 ( 
.A(n_70),
.B(n_52),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_90),
.A2(n_107),
.B(n_79),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_93),
.A2(n_102),
.B1(n_106),
.B2(n_69),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_82),
.B(n_47),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_96),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_47),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_95),
.B(n_76),
.Y(n_113)
);

AO22x1_ASAP7_75t_L g96 ( 
.A1(n_74),
.A2(n_34),
.B1(n_49),
.B2(n_33),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_105),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_74),
.B(n_64),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_103),
.Y(n_122)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_101),
.B(n_104),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_24),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_70),
.A2(n_50),
.B1(n_28),
.B2(n_31),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_108),
.B(n_113),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_110),
.A2(n_116),
.B(n_117),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_88),
.A2(n_79),
.B1(n_76),
.B2(n_71),
.Y(n_111)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_111),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_95),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_114),
.B(n_115),
.Y(n_143)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_92),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_92),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_86),
.A2(n_66),
.B(n_27),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_118),
.A2(n_90),
.B(n_107),
.Y(n_135)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_119),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_106),
.C(n_110),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_97),
.A2(n_66),
.B1(n_33),
.B2(n_57),
.Y(n_125)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_125),
.Y(n_132)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_90),
.Y(n_126)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_126),
.Y(n_139)
);

OAI21xp33_ASAP7_75t_L g127 ( 
.A1(n_109),
.A2(n_86),
.B(n_99),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_127),
.A2(n_135),
.B(n_27),
.Y(n_159)
);

NOR4xp25_ASAP7_75t_L g129 ( 
.A(n_116),
.B(n_103),
.C(n_87),
.D(n_101),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_130),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_123),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_133),
.B(n_136),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_90),
.C(n_100),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_144),
.C(n_118),
.Y(n_145)
);

NAND3xp33_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_94),
.C(n_100),
.Y(n_136)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_111),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_141),
.Y(n_150)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

NAND3xp33_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_94),
.C(n_96),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_112),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_105),
.C(n_104),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_147),
.C(n_151),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_128),
.A2(n_117),
.B1(n_114),
.B2(n_121),
.Y(n_146)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_146),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_120),
.C(n_126),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_128),
.A2(n_93),
.B1(n_124),
.B2(n_115),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_148),
.A2(n_158),
.B1(n_132),
.B2(n_139),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_96),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g153 ( 
.A(n_138),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_153),
.B(n_156),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_112),
.C(n_78),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_39),
.C(n_63),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_159),
.Y(n_165)
);

INVxp33_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_157),
.A2(n_131),
.B(n_135),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_140),
.A2(n_119),
.B1(n_24),
.B2(n_18),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_163),
.A2(n_166),
.B(n_150),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_164),
.A2(n_169),
.B1(n_63),
.B2(n_62),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_152),
.A2(n_139),
.B(n_132),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_156),
.B(n_141),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_167),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_134),
.C(n_78),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_170),
.C(n_172),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_157),
.A2(n_18),
.B1(n_57),
.B2(n_39),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_149),
.B(n_39),
.C(n_36),
.Y(n_170)
);

AOI322xp5_ASAP7_75t_L g171 ( 
.A1(n_149),
.A2(n_36),
.A3(n_39),
.B1(n_12),
.B2(n_15),
.C1(n_14),
.C2(n_13),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_154),
.Y(n_177)
);

MAJx2_ASAP7_75t_L g186 ( 
.A(n_174),
.B(n_3),
.C(n_4),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_166),
.A2(n_151),
.B(n_145),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_175),
.A2(n_180),
.B(n_3),
.Y(n_190)
);

INVxp67_ASAP7_75t_SL g176 ( 
.A(n_162),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_176),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_179),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_160),
.A2(n_1),
.B(n_2),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_165),
.A2(n_13),
.B1(n_12),
.B2(n_5),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_181),
.B(n_182),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_168),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_178),
.B(n_161),
.C(n_172),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_183),
.B(n_189),
.C(n_62),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_180),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_184),
.A2(n_190),
.B(n_173),
.Y(n_191)
);

MAJx2_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_7),
.C(n_8),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_63),
.C(n_62),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_191),
.B(n_196),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_187),
.A2(n_176),
.B1(n_5),
.B2(n_6),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_193),
.C(n_195),
.Y(n_200)
);

OAI21xp33_ASAP7_75t_L g194 ( 
.A1(n_189),
.A2(n_4),
.B(n_5),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_194),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_6),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_188),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_199),
.B(n_183),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_203),
.C(n_9),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_198),
.Y(n_202)
);

AOI21x1_ASAP7_75t_L g204 ( 
.A1(n_202),
.A2(n_197),
.B(n_7),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_186),
.C(n_8),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_204),
.B(n_205),
.Y(n_206)
);


endmodule