module fake_jpeg_1171_n_615 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_615);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_615;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_18),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx11_ASAP7_75t_SL g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_6),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_11),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx24_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

BUFx6f_ASAP7_75t_SL g54 ( 
.A(n_10),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

BUFx16f_ASAP7_75t_L g56 ( 
.A(n_7),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_5),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_56),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_59),
.B(n_78),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_26),
.B(n_17),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_60),
.B(n_67),
.Y(n_133)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g156 ( 
.A(n_61),
.Y(n_156)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_62),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_64),
.Y(n_131)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_66),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_26),
.B(n_17),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_68),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_69),
.Y(n_128)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_70),
.Y(n_138)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_71),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_72),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_22),
.B(n_0),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_73),
.B(n_76),
.Y(n_151)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_74),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_75),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_22),
.B(n_0),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_29),
.B(n_0),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_77),
.B(n_86),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_24),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_79),
.Y(n_147)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_80),
.Y(n_158)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_81),
.Y(n_141)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_82),
.Y(n_135)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_83),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_21),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_84),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_85),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_29),
.B(n_0),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_87),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_24),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_88),
.B(n_89),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_33),
.B(n_1),
.Y(n_89)
);

INVx13_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_90),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_91),
.Y(n_142)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_23),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_92),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_24),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_93),
.B(n_103),
.Y(n_175)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_37),
.Y(n_94)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_94),
.Y(n_191)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_25),
.Y(n_95)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_95),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_40),
.Y(n_96)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_96),
.Y(n_185)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_97),
.Y(n_202)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_42),
.Y(n_98)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_98),
.Y(n_143)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_99),
.Y(n_182)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_40),
.Y(n_100)
);

INVx3_ASAP7_75t_SL g169 ( 
.A(n_100),
.Y(n_169)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_101),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_41),
.Y(n_102)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_102),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_32),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_33),
.Y(n_104)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_104),
.Y(n_178)
);

INVx8_ASAP7_75t_L g105 ( 
.A(n_25),
.Y(n_105)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_105),
.Y(n_183)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_106),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_46),
.Y(n_107)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_107),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_32),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_108),
.B(n_112),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_41),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_109),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_34),
.B(n_15),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_110),
.B(n_117),
.Y(n_148)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_111),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_41),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_53),
.Y(n_113)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_113),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_53),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_114),
.B(n_46),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_115),
.Y(n_213)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_31),
.Y(n_116)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_116),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_35),
.B(n_1),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_31),
.Y(n_118)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_118),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_39),
.B(n_2),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_2),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_45),
.Y(n_120)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_120),
.Y(n_161)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_35),
.Y(n_121)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_121),
.Y(n_215)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_58),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_122),
.Y(n_197)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_48),
.Y(n_123)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_123),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_45),
.Y(n_124)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_124),
.Y(n_160)
);

BUFx12_ASAP7_75t_L g125 ( 
.A(n_46),
.Y(n_125)
);

BUFx16f_ASAP7_75t_L g194 ( 
.A(n_125),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_51),
.Y(n_126)
);

INVx8_ASAP7_75t_L g173 ( 
.A(n_126),
.Y(n_173)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_48),
.Y(n_127)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_127),
.Y(n_165)
);

INVx11_ASAP7_75t_L g140 ( 
.A(n_72),
.Y(n_140)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_140),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_100),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_146),
.B(n_170),
.Y(n_219)
);

INVx11_ASAP7_75t_L g150 ( 
.A(n_72),
.Y(n_150)
);

BUFx10_ASAP7_75t_L g239 ( 
.A(n_150),
.Y(n_239)
);

BUFx12_ASAP7_75t_L g155 ( 
.A(n_61),
.Y(n_155)
);

CKINVDCx12_ASAP7_75t_R g231 ( 
.A(n_155),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_159),
.B(n_164),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_97),
.B(n_52),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_120),
.A2(n_58),
.B1(n_51),
.B2(n_39),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_166),
.A2(n_198),
.B1(n_9),
.B2(n_11),
.Y(n_286)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_68),
.Y(n_168)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_168),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_99),
.Y(n_170)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_63),
.Y(n_172)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_172),
.Y(n_250)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_64),
.Y(n_174)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_174),
.Y(n_261)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_66),
.Y(n_176)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_176),
.Y(n_272)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_75),
.Y(n_177)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_177),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_121),
.B(n_52),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_180),
.B(n_199),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_84),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_181),
.B(n_193),
.Y(n_223)
);

OAI21xp33_ASAP7_75t_L g184 ( 
.A1(n_90),
.A2(n_44),
.B(n_43),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_184),
.A2(n_214),
.B(n_111),
.Y(n_227)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_85),
.Y(n_187)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_187),
.Y(n_276)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_91),
.Y(n_192)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_192),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_96),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_126),
.A2(n_54),
.B1(n_44),
.B2(n_43),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_69),
.B(n_2),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_102),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_200),
.B(n_201),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_113),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_205),
.B(n_12),
.Y(n_287)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_122),
.Y(n_209)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_209),
.Y(n_222)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_109),
.Y(n_210)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_210),
.Y(n_233)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_115),
.Y(n_211)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_211),
.Y(n_257)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_124),
.Y(n_212)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_212),
.Y(n_281)
);

NAND2x1_ASAP7_75t_L g214 ( 
.A(n_82),
.B(n_54),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_130),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_216),
.Y(n_310)
);

INVx6_ASAP7_75t_L g217 ( 
.A(n_130),
.Y(n_217)
);

INVx8_ASAP7_75t_L g322 ( 
.A(n_217),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_131),
.Y(n_218)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_218),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_157),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_221),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_131),
.Y(n_224)
);

INVx4_ASAP7_75t_L g326 ( 
.A(n_224),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_157),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g344 ( 
.A(n_225),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_186),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_226),
.B(n_232),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_227),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_147),
.A2(n_106),
.B1(n_83),
.B2(n_80),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_228),
.A2(n_268),
.B1(n_282),
.B2(n_285),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_129),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_230),
.B(n_156),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_194),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_148),
.B(n_3),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_234),
.B(n_251),
.Y(n_302)
);

CKINVDCx9p33_ASAP7_75t_R g235 ( 
.A(n_129),
.Y(n_235)
);

INVx11_ASAP7_75t_L g320 ( 
.A(n_235),
.Y(n_320)
);

INVx6_ASAP7_75t_L g237 ( 
.A(n_189),
.Y(n_237)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_237),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_179),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_238),
.B(n_254),
.Y(n_298)
);

NAND2xp33_ASAP7_75t_SL g240 ( 
.A(n_152),
.B(n_125),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g346 ( 
.A1(n_240),
.A2(n_252),
.B(n_230),
.Y(n_346)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_136),
.Y(n_241)
);

BUFx3_ASAP7_75t_L g337 ( 
.A(n_241),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_171),
.A2(n_105),
.B1(n_95),
.B2(n_92),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_242),
.A2(n_247),
.B1(n_259),
.B2(n_266),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_189),
.Y(n_244)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_244),
.Y(n_292)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_135),
.Y(n_245)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_245),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_188),
.B(n_61),
.C(n_79),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_246),
.B(n_248),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_151),
.A2(n_125),
.B1(n_50),
.B2(n_47),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_196),
.B(n_134),
.C(n_138),
.Y(n_248)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_135),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_249),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_151),
.B(n_3),
.Y(n_251)
);

OR2x4_ASAP7_75t_L g252 ( 
.A(n_184),
.B(n_50),
.Y(n_252)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_195),
.Y(n_253)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_253),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_179),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_167),
.B(n_3),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_255),
.B(n_264),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_175),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_256),
.B(n_258),
.Y(n_319)
);

NOR3xp33_ASAP7_75t_L g258 ( 
.A(n_133),
.B(n_167),
.C(n_171),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_165),
.A2(n_175),
.B1(n_132),
.B2(n_137),
.Y(n_259)
);

INVx8_ASAP7_75t_L g260 ( 
.A(n_156),
.Y(n_260)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_260),
.Y(n_294)
);

INVx4_ASAP7_75t_SL g262 ( 
.A(n_194),
.Y(n_262)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_262),
.Y(n_296)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_128),
.Y(n_263)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_263),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_133),
.B(n_4),
.Y(n_264)
);

INVx2_ASAP7_75t_SL g265 ( 
.A(n_215),
.Y(n_265)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_265),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_L g266 ( 
.A1(n_198),
.A2(n_50),
.B1(n_47),
.B2(n_27),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_214),
.B(n_5),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_267),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_147),
.A2(n_50),
.B1(n_47),
.B2(n_27),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_178),
.B(n_139),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_269),
.B(n_280),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_191),
.A2(n_47),
.B1(n_27),
.B2(n_8),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_270),
.A2(n_169),
.B1(n_154),
.B2(n_197),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_195),
.Y(n_271)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_271),
.Y(n_315)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_153),
.Y(n_274)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_274),
.Y(n_317)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_183),
.Y(n_275)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_275),
.Y(n_323)
);

INVx2_ASAP7_75t_SL g277 ( 
.A(n_182),
.Y(n_277)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_277),
.Y(n_332)
);

INVx8_ASAP7_75t_L g279 ( 
.A(n_156),
.Y(n_279)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_279),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_141),
.B(n_144),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_203),
.A2(n_27),
.B1(n_7),
.B2(n_8),
.Y(n_282)
);

OR2x2_ASAP7_75t_SL g283 ( 
.A(n_158),
.B(n_6),
.Y(n_283)
);

NOR2x1_ASAP7_75t_L g327 ( 
.A(n_283),
.B(n_128),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_203),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_284),
.B(n_287),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_163),
.A2(n_6),
.B1(n_9),
.B2(n_11),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_286),
.A2(n_162),
.B1(n_145),
.B2(n_160),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_204),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_288),
.Y(n_303)
);

INVx6_ASAP7_75t_L g289 ( 
.A(n_204),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_289),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_291),
.B(n_327),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_236),
.B(n_143),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_299),
.B(n_276),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_242),
.A2(n_169),
.B1(n_190),
.B2(n_206),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_301),
.A2(n_330),
.B1(n_333),
.B2(n_338),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_252),
.A2(n_207),
.B1(n_161),
.B2(n_173),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_304),
.A2(n_314),
.B1(n_334),
.B2(n_307),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_L g305 ( 
.A1(n_223),
.A2(n_278),
.B1(n_202),
.B2(n_266),
.Y(n_305)
);

OA22x2_ASAP7_75t_L g386 ( 
.A1(n_305),
.A2(n_312),
.B1(n_343),
.B2(n_334),
.Y(n_386)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_307),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_L g312 ( 
.A1(n_229),
.A2(n_219),
.B1(n_149),
.B2(n_235),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_267),
.A2(n_207),
.B1(n_173),
.B2(n_161),
.Y(n_314)
);

OAI22xp33_ASAP7_75t_L g365 ( 
.A1(n_318),
.A2(n_282),
.B1(n_285),
.B2(n_277),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_259),
.A2(n_206),
.B1(n_142),
.B2(n_190),
.Y(n_330)
);

OAI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_228),
.A2(n_182),
.B1(n_208),
.B2(n_185),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_255),
.A2(n_213),
.B1(n_208),
.B2(n_185),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_241),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_335),
.B(n_336),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_263),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_268),
.A2(n_142),
.B1(n_13),
.B2(n_15),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_SL g339 ( 
.A1(n_274),
.A2(n_155),
.B1(n_13),
.B2(n_15),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_SL g357 ( 
.A1(n_339),
.A2(n_262),
.B1(n_243),
.B2(n_265),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_248),
.B(n_12),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_342),
.B(n_347),
.Y(n_359)
);

AOI22x1_ASAP7_75t_L g343 ( 
.A1(n_240),
.A2(n_12),
.B1(n_283),
.B2(n_275),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_346),
.A2(n_220),
.B(n_273),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_222),
.B(n_281),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_348),
.A2(n_365),
.B1(n_371),
.B2(n_379),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_297),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_351),
.B(n_353),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_304),
.B(n_246),
.Y(n_352)
);

CKINVDCx14_ASAP7_75t_R g417 ( 
.A(n_352),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_344),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_293),
.Y(n_354)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_354),
.Y(n_410)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_313),
.Y(n_355)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_355),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_325),
.B(n_257),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_356),
.B(n_358),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_357),
.Y(n_415)
);

AO22x2_ASAP7_75t_L g358 ( 
.A1(n_308),
.A2(n_290),
.B1(n_250),
.B2(n_261),
.Y(n_358)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_313),
.Y(n_360)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_360),
.Y(n_423)
);

INVx13_ASAP7_75t_L g361 ( 
.A(n_320),
.Y(n_361)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_361),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_362),
.B(n_368),
.Y(n_411)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_317),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_363),
.B(n_364),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_319),
.B(n_233),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_321),
.B(n_245),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_367),
.B(n_369),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_325),
.B(n_272),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_298),
.B(n_249),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_293),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_370),
.B(n_378),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_329),
.A2(n_217),
.B1(n_253),
.B2(n_237),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_373),
.A2(n_388),
.B(n_389),
.Y(n_421)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_317),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_374),
.B(n_376),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_329),
.B(n_343),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_SL g408 ( 
.A(n_375),
.B(n_385),
.Y(n_408)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_323),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_296),
.B(n_279),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_377),
.B(n_380),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_328),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_299),
.A2(n_289),
.B1(n_218),
.B2(n_224),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_323),
.Y(n_380)
);

OAI22xp33_ASAP7_75t_L g381 ( 
.A1(n_300),
.A2(n_216),
.B1(n_288),
.B2(n_271),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_381),
.A2(n_301),
.B1(n_338),
.B2(n_303),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_308),
.A2(n_244),
.B1(n_243),
.B2(n_260),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_382),
.A2(n_366),
.B1(n_372),
.B2(n_360),
.Y(n_422)
);

BUFx2_ASAP7_75t_L g383 ( 
.A(n_295),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_383),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_316),
.B(n_239),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_384),
.B(n_386),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_343),
.B(n_231),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_296),
.B(n_239),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_387),
.A2(n_390),
.B(n_373),
.Y(n_413)
);

AND2x6_ASAP7_75t_L g388 ( 
.A(n_346),
.B(n_239),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_332),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_332),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_316),
.B(n_327),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_391),
.B(n_327),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_394),
.B(n_368),
.Y(n_435)
);

INVx1_ASAP7_75t_SL g444 ( 
.A(n_395),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_385),
.A2(n_307),
.B(n_336),
.Y(n_396)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_396),
.A2(n_398),
.B(n_400),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_352),
.A2(n_330),
.B1(n_340),
.B2(n_309),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_397),
.A2(n_404),
.B1(n_386),
.B2(n_358),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_385),
.A2(n_335),
.B(n_294),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_349),
.A2(n_345),
.B(n_294),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_352),
.A2(n_340),
.B1(n_309),
.B2(n_314),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_349),
.A2(n_320),
.B(n_345),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_406),
.A2(n_412),
.B(n_424),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_391),
.A2(n_291),
.B1(n_303),
.B2(n_341),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_407),
.B(n_426),
.Y(n_441)
);

OA21x2_ASAP7_75t_L g409 ( 
.A1(n_349),
.A2(n_331),
.B(n_311),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_409),
.B(n_428),
.Y(n_451)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_375),
.A2(n_328),
.B(n_306),
.Y(n_412)
);

CKINVDCx16_ASAP7_75t_R g457 ( 
.A(n_413),
.Y(n_457)
);

AOI22xp33_ASAP7_75t_L g443 ( 
.A1(n_422),
.A2(n_417),
.B1(n_425),
.B2(n_402),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_375),
.A2(n_306),
.B(n_311),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_366),
.A2(n_324),
.B1(n_341),
.B2(n_315),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g439 ( 
.A1(n_425),
.A2(n_350),
.B1(n_378),
.B2(n_355),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_384),
.A2(n_315),
.B1(n_292),
.B2(n_326),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_382),
.A2(n_292),
.B1(n_295),
.B2(n_326),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_427),
.A2(n_379),
.B1(n_383),
.B2(n_374),
.Y(n_459)
);

OAI32xp33_ASAP7_75t_L g428 ( 
.A1(n_362),
.A2(n_324),
.A3(n_302),
.B1(n_331),
.B2(n_322),
.Y(n_428)
);

AOI22xp33_ASAP7_75t_SL g429 ( 
.A1(n_415),
.A2(n_371),
.B1(n_348),
.B2(n_372),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_429),
.Y(n_471)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_405),
.Y(n_430)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_430),
.Y(n_465)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_405),
.Y(n_431)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_431),
.Y(n_468)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_418),
.Y(n_432)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_432),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_403),
.B(n_351),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_433),
.B(n_437),
.Y(n_469)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_418),
.Y(n_434)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_434),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_435),
.B(n_396),
.Y(n_483)
);

OR2x2_ASAP7_75t_L g436 ( 
.A(n_409),
.B(n_386),
.Y(n_436)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_436),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_403),
.B(n_353),
.Y(n_437)
);

AOI22xp33_ASAP7_75t_L g481 ( 
.A1(n_439),
.A2(n_450),
.B1(n_459),
.B2(n_461),
.Y(n_481)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_414),
.Y(n_440)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_440),
.Y(n_491)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_414),
.Y(n_442)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_442),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_443),
.A2(n_404),
.B1(n_392),
.B2(n_395),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_401),
.B(n_380),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_SL g474 ( 
.A(n_445),
.B(n_453),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_SL g446 ( 
.A(n_401),
.B(n_356),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_446),
.B(n_448),
.Y(n_462)
);

OR2x4_ASAP7_75t_L g447 ( 
.A(n_419),
.B(n_388),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g472 ( 
.A(n_447),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g448 ( 
.A(n_393),
.B(n_359),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_416),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_SL g452 ( 
.A1(n_422),
.A2(n_390),
.B1(n_389),
.B2(n_383),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_452),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_393),
.B(n_363),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_454),
.A2(n_455),
.B1(n_409),
.B2(n_407),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_419),
.A2(n_392),
.B1(n_417),
.B2(n_397),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_416),
.B(n_376),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_456),
.B(n_458),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_SL g458 ( 
.A(n_411),
.B(n_302),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_423),
.B(n_354),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_460),
.B(n_410),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_398),
.Y(n_461)
);

BUFx24_ASAP7_75t_SL g463 ( 
.A(n_448),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_463),
.B(n_466),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_435),
.B(n_394),
.C(n_408),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_464),
.B(n_470),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_446),
.B(n_337),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_457),
.B(n_408),
.C(n_421),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_456),
.B(n_411),
.Y(n_476)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_476),
.Y(n_498)
);

NOR4xp25_ASAP7_75t_L g477 ( 
.A(n_430),
.B(n_413),
.C(n_408),
.D(n_423),
.Y(n_477)
);

OR2x2_ASAP7_75t_L g520 ( 
.A(n_477),
.B(n_479),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_445),
.B(n_402),
.Y(n_478)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_478),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_483),
.B(n_455),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_450),
.B(n_337),
.Y(n_484)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_484),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_485),
.A2(n_489),
.B1(n_457),
.B2(n_451),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_458),
.B(n_426),
.Y(n_486)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_486),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_487),
.A2(n_444),
.B1(n_436),
.B2(n_434),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_433),
.B(n_421),
.Y(n_488)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_488),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_443),
.A2(n_400),
.B1(n_424),
.B2(n_412),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_431),
.B(n_409),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_490),
.B(n_432),
.Y(n_502)
);

AOI22xp33_ASAP7_75t_SL g494 ( 
.A1(n_471),
.A2(n_444),
.B1(n_454),
.B2(n_439),
.Y(n_494)
);

OAI22xp33_ASAP7_75t_SL g530 ( 
.A1(n_494),
.A2(n_471),
.B1(n_480),
.B2(n_475),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_496),
.B(n_502),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_469),
.Y(n_497)
);

AOI22xp33_ASAP7_75t_L g531 ( 
.A1(n_497),
.A2(n_506),
.B1(n_515),
.B2(n_516),
.Y(n_531)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_499),
.A2(n_501),
.B1(n_513),
.B2(n_518),
.Y(n_527)
);

INVx1_ASAP7_75t_SL g500 ( 
.A(n_491),
.Y(n_500)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_500),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_487),
.A2(n_436),
.B1(n_444),
.B2(n_451),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_470),
.B(n_447),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_503),
.B(n_510),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_465),
.B(n_437),
.Y(n_505)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_505),
.Y(n_543)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_491),
.Y(n_506)
);

OAI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_507),
.A2(n_517),
.B1(n_482),
.B2(n_473),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_464),
.B(n_447),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_SL g511 ( 
.A(n_483),
.B(n_451),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_511),
.B(n_386),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_SL g513 ( 
.A1(n_481),
.A2(n_451),
.B1(n_441),
.B2(n_461),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_465),
.B(n_453),
.Y(n_514)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_514),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_462),
.A2(n_441),
.B1(n_459),
.B2(n_406),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_468),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_485),
.A2(n_449),
.B1(n_438),
.B2(n_427),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_482),
.A2(n_449),
.B1(n_438),
.B2(n_442),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g519 ( 
.A1(n_472),
.A2(n_406),
.B(n_428),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_SL g535 ( 
.A1(n_519),
.A2(n_492),
.B(n_440),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_493),
.B(n_472),
.C(n_473),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_521),
.B(n_524),
.Y(n_549)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_523),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_508),
.B(n_469),
.Y(n_524)
);

AOI21xp33_ASAP7_75t_L g525 ( 
.A1(n_512),
.A2(n_467),
.B(n_474),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_525),
.B(n_520),
.Y(n_546)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_519),
.A2(n_490),
.B(n_489),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_L g560 ( 
.A1(n_526),
.A2(n_535),
.B(n_537),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_495),
.B(n_476),
.Y(n_529)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_529),
.Y(n_557)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_530),
.B(n_539),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_493),
.B(n_468),
.C(n_480),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_532),
.B(n_533),
.C(n_536),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_510),
.B(n_475),
.C(n_478),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_514),
.B(n_460),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g544 ( 
.A(n_534),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_503),
.B(n_410),
.C(n_492),
.Y(n_536)
);

OAI21xp5_ASAP7_75t_L g537 ( 
.A1(n_518),
.A2(n_420),
.B(n_399),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_511),
.B(n_420),
.C(n_370),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_541),
.B(n_502),
.C(n_500),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_496),
.B(n_381),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_542),
.B(n_517),
.Y(n_547)
);

OR2x2_ASAP7_75t_L g574 ( 
.A(n_546),
.B(n_555),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_L g566 ( 
.A(n_547),
.B(n_553),
.Y(n_566)
);

INVx13_ASAP7_75t_L g548 ( 
.A(n_531),
.Y(n_548)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_548),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_527),
.A2(n_520),
.B1(n_509),
.B2(n_498),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_L g569 ( 
.A1(n_552),
.A2(n_556),
.B1(n_558),
.B2(n_526),
.Y(n_569)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_538),
.Y(n_554)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_554),
.Y(n_563)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_543),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_540),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_L g558 ( 
.A1(n_527),
.A2(n_507),
.B1(n_504),
.B2(n_505),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_532),
.B(n_513),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g573 ( 
.A(n_559),
.B(n_539),
.Y(n_573)
);

BUFx12_ASAP7_75t_L g561 ( 
.A(n_535),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_561),
.B(n_358),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_551),
.B(n_536),
.C(n_528),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_564),
.B(n_565),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_551),
.B(n_528),
.C(n_533),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_545),
.A2(n_523),
.B1(n_501),
.B2(n_542),
.Y(n_567)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_567),
.Y(n_583)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_559),
.B(n_521),
.C(n_522),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_568),
.B(n_570),
.Y(n_587)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_569),
.Y(n_585)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_553),
.B(n_522),
.C(n_541),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_557),
.B(n_544),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_571),
.B(n_572),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_544),
.B(n_537),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_573),
.B(n_566),
.Y(n_588)
);

OAI21xp5_ASAP7_75t_SL g575 ( 
.A1(n_549),
.A2(n_506),
.B(n_399),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_575),
.B(n_554),
.Y(n_578)
);

OAI21xp33_ASAP7_75t_L g580 ( 
.A1(n_576),
.A2(n_555),
.B(n_556),
.Y(n_580)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_562),
.Y(n_577)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_577),
.Y(n_589)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_578),
.Y(n_593)
);

INVxp67_ASAP7_75t_L g579 ( 
.A(n_565),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_579),
.B(n_580),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_566),
.B(n_545),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_581),
.B(n_570),
.Y(n_595)
);

OAI221xp5_ASAP7_75t_SL g582 ( 
.A1(n_574),
.A2(n_561),
.B1(n_560),
.B2(n_548),
.C(n_550),
.Y(n_582)
);

O2A1O1Ixp33_ASAP7_75t_L g594 ( 
.A1(n_582),
.A2(n_560),
.B(n_561),
.C(n_563),
.Y(n_594)
);

INVxp33_ASAP7_75t_L g591 ( 
.A(n_588),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_587),
.B(n_564),
.C(n_574),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_590),
.B(n_595),
.Y(n_599)
);

AOI21xp5_ASAP7_75t_L g598 ( 
.A1(n_594),
.A2(n_596),
.B(n_585),
.Y(n_598)
);

OR2x2_ASAP7_75t_L g596 ( 
.A(n_584),
.B(n_567),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_586),
.B(n_568),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_597),
.B(n_547),
.Y(n_602)
);

NOR3xp33_ASAP7_75t_L g606 ( 
.A(n_598),
.B(n_601),
.C(n_602),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_591),
.B(n_588),
.C(n_583),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_600),
.B(n_603),
.Y(n_607)
);

AO21x1_ASAP7_75t_L g601 ( 
.A1(n_591),
.A2(n_580),
.B(n_573),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_593),
.B(n_550),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_592),
.B(n_596),
.C(n_589),
.Y(n_604)
);

XOR2xp5_ASAP7_75t_L g605 ( 
.A(n_604),
.B(n_358),
.Y(n_605)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_605),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g608 ( 
.A(n_599),
.B(n_310),
.C(n_365),
.Y(n_608)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_608),
.Y(n_610)
);

OAI311xp33_ASAP7_75t_L g611 ( 
.A1(n_609),
.A2(n_607),
.A3(n_606),
.B1(n_603),
.C1(n_358),
.Y(n_611)
);

XOR2xp5_ASAP7_75t_L g612 ( 
.A(n_611),
.B(n_610),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_612),
.B(n_310),
.Y(n_613)
);

AOI221xp5_ASAP7_75t_L g614 ( 
.A1(n_613),
.A2(n_310),
.B1(n_322),
.B2(n_361),
.C(n_584),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_614),
.B(n_322),
.Y(n_615)
);


endmodule