module fake_jpeg_7168_n_340 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx4_ASAP7_75t_SL g33 ( 
.A(n_9),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_39),
.Y(n_49)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

OR2x2_ASAP7_75t_SL g40 ( 
.A(n_17),
.B(n_18),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_44),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx8_ASAP7_75t_SL g46 ( 
.A(n_22),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_31),
.Y(n_62)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_50),
.B(n_51),
.Y(n_94)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_48),
.A2(n_24),
.B1(n_32),
.B2(n_18),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_53),
.A2(n_67),
.B1(n_27),
.B2(n_33),
.Y(n_98)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_58),
.B(n_60),
.Y(n_99)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_24),
.Y(n_61)
);

NAND3xp33_ASAP7_75t_L g90 ( 
.A(n_61),
.B(n_15),
.C(n_16),
.Y(n_90)
);

INVxp33_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_65),
.Y(n_76)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_44),
.A2(n_17),
.B1(n_31),
.B2(n_34),
.Y(n_67)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_71),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_41),
.B(n_19),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_34),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g73 ( 
.A(n_66),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_73),
.B(n_78),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_79),
.A2(n_88),
.B1(n_92),
.B2(n_96),
.Y(n_113)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_80),
.A2(n_30),
.B1(n_22),
.B2(n_20),
.Y(n_128)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_83),
.Y(n_114)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_84),
.B(n_86),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_87),
.Y(n_103)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_89),
.Y(n_101)
);

OAI21xp33_ASAP7_75t_SL g109 ( 
.A1(n_90),
.A2(n_98),
.B(n_53),
.Y(n_109)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx3_ASAP7_75t_SL g116 ( 
.A(n_91),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_50),
.A2(n_33),
.B1(n_21),
.B2(n_19),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_55),
.A2(n_33),
.B1(n_27),
.B2(n_21),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_93),
.A2(n_33),
.B1(n_49),
.B2(n_57),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_61),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_112),
.Y(n_130)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

INVx11_ASAP7_75t_L g143 ( 
.A(n_104),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_98),
.A2(n_51),
.B1(n_58),
.B2(n_68),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_105),
.A2(n_107),
.B1(n_121),
.B2(n_124),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_94),
.A2(n_68),
.B1(n_54),
.B2(n_57),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_76),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_108),
.B(n_118),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_109),
.A2(n_115),
.B1(n_128),
.B2(n_96),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_67),
.Y(n_112)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_99),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_73),
.Y(n_142)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_85),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_120),
.B(n_84),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_79),
.A2(n_72),
.B1(n_65),
.B2(n_64),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_99),
.B(n_43),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_28),
.C(n_29),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_77),
.A2(n_20),
.B(n_35),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_123),
.A2(n_25),
.B(n_80),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_88),
.A2(n_69),
.B1(n_20),
.B2(n_35),
.Y(n_124)
);

AOI22x1_ASAP7_75t_L g126 ( 
.A1(n_97),
.A2(n_45),
.B1(n_42),
.B2(n_35),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_126),
.A2(n_91),
.B1(n_81),
.B2(n_86),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_95),
.B(n_35),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_120),
.Y(n_154)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_116),
.Y(n_129)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_129),
.Y(n_162)
);

O2A1O1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_126),
.A2(n_97),
.B(n_28),
.C(n_29),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_131),
.A2(n_134),
.B1(n_139),
.B2(n_103),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_102),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_132),
.B(n_135),
.C(n_105),
.Y(n_161)
);

AND2x6_ASAP7_75t_L g133 ( 
.A(n_126),
.B(n_15),
.Y(n_133)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_133),
.Y(n_156)
);

O2A1O1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_115),
.A2(n_28),
.B(n_29),
.C(n_25),
.Y(n_134)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_137),
.B(n_140),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_138),
.A2(n_146),
.B(n_25),
.Y(n_175)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_142),
.B(n_117),
.Y(n_176)
);

AND2x6_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_14),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_144),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_145),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_119),
.B(n_0),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_L g178 ( 
.A1(n_147),
.A2(n_111),
.B1(n_101),
.B2(n_106),
.Y(n_178)
);

CKINVDCx10_ASAP7_75t_R g148 ( 
.A(n_116),
.Y(n_148)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_106),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_150),
.Y(n_181)
);

INVx13_ASAP7_75t_L g150 ( 
.A(n_100),
.Y(n_150)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_100),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_84),
.Y(n_184)
);

INVx6_ASAP7_75t_L g152 ( 
.A(n_100),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_152),
.Y(n_171)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_153),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_154),
.B(n_127),
.Y(n_157)
);

INVx4_ASAP7_75t_SL g155 ( 
.A(n_104),
.Y(n_155)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_155),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_157),
.B(n_158),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_112),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_107),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_159),
.B(n_129),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_160),
.A2(n_137),
.B1(n_138),
.B2(n_155),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_132),
.C(n_133),
.Y(n_187)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_143),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_166),
.B(n_150),
.Y(n_195)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_154),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_174),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_141),
.A2(n_113),
.B1(n_123),
.B2(n_78),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_169),
.A2(n_170),
.B1(n_129),
.B2(n_155),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_141),
.A2(n_83),
.B1(n_110),
.B2(n_108),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_140),
.A2(n_124),
.B1(n_125),
.B2(n_103),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_172),
.A2(n_180),
.B1(n_143),
.B2(n_152),
.Y(n_207)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_175),
.A2(n_177),
.B1(n_178),
.B2(n_182),
.Y(n_196)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_176),
.B(n_183),
.Y(n_205)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_136),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_130),
.A2(n_117),
.B1(n_111),
.B2(n_73),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_136),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_142),
.B(n_95),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_184),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_186),
.A2(n_207),
.B1(n_150),
.B2(n_101),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_187),
.B(n_188),
.C(n_197),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_146),
.Y(n_188)
);

NAND3xp33_ASAP7_75t_L g189 ( 
.A(n_176),
.B(n_144),
.C(n_177),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_189),
.B(n_194),
.Y(n_220)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_173),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_190),
.B(n_198),
.Y(n_239)
);

A2O1A1Ixp33_ASAP7_75t_L g191 ( 
.A1(n_158),
.A2(n_146),
.B(n_131),
.C(n_134),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_191),
.B(n_175),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_192),
.A2(n_169),
.B1(n_171),
.B2(n_164),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_181),
.Y(n_194)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_195),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_75),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_179),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_199),
.A2(n_165),
.B(n_164),
.Y(n_229)
);

AND2x6_ASAP7_75t_L g201 ( 
.A(n_156),
.B(n_75),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_201),
.Y(n_225)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_157),
.Y(n_202)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_202),
.Y(n_226)
);

AND2x6_ASAP7_75t_L g203 ( 
.A(n_156),
.B(n_74),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_203),
.A2(n_209),
.B(n_167),
.Y(n_215)
);

XNOR2x1_ASAP7_75t_SL g204 ( 
.A(n_168),
.B(n_74),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_204),
.B(n_89),
.Y(n_234)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_170),
.Y(n_206)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_206),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_151),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_208),
.B(n_210),
.Y(n_213)
);

AND2x6_ASAP7_75t_L g209 ( 
.A(n_156),
.B(n_74),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_183),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_172),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_211),
.B(n_212),
.Y(n_216)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_166),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_174),
.Y(n_214)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_214),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_215),
.A2(n_221),
.B(n_227),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_193),
.Y(n_217)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_217),
.Y(n_250)
);

OR2x2_ASAP7_75t_L g218 ( 
.A(n_205),
.B(n_167),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_218),
.B(n_231),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_219),
.A2(n_190),
.B1(n_185),
.B2(n_212),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_207),
.A2(n_160),
.B1(n_163),
.B2(n_171),
.Y(n_223)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_223),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_188),
.B(n_187),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_230),
.C(n_236),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_199),
.A2(n_159),
.B(n_163),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_229),
.B(n_234),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_193),
.B(n_159),
.C(n_165),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g231 ( 
.A(n_196),
.B(n_149),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_200),
.B(n_162),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_232),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_208),
.B(n_162),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_233),
.B(n_237),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_197),
.B(n_84),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_201),
.A2(n_14),
.B(n_13),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_238),
.A2(n_225),
.B1(n_191),
.B2(n_215),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_192),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_242),
.B(n_253),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_225),
.A2(n_199),
.B1(n_209),
.B2(n_203),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_243),
.A2(n_216),
.B1(n_213),
.B2(n_226),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_239),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_244),
.B(n_233),
.Y(n_271)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_245),
.Y(n_264)
);

XNOR2x2_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_214),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_248),
.A2(n_214),
.B1(n_226),
.B2(n_227),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_252),
.A2(n_223),
.B1(n_235),
.B2(n_221),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_30),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_222),
.B(n_30),
.Y(n_254)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_254),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_219),
.A2(n_14),
.B1(n_1),
.B2(n_2),
.Y(n_255)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_255),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_228),
.B(n_0),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_257),
.B(n_259),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_235),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_258),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_228),
.B(n_0),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_1),
.C(n_2),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_260),
.B(n_262),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_229),
.B(n_2),
.C(n_3),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_256),
.Y(n_263)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_263),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_267),
.Y(n_289)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_248),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_275),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_271),
.B(n_274),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_272),
.A2(n_261),
.B1(n_262),
.B2(n_232),
.Y(n_287)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_256),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_244),
.B(n_252),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_251),
.A2(n_238),
.B1(n_216),
.B2(n_217),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_277),
.A2(n_278),
.B1(n_280),
.B2(n_250),
.Y(n_281)
);

FAx1_ASAP7_75t_SL g279 ( 
.A(n_241),
.B(n_213),
.CI(n_218),
.CON(n_279),
.SN(n_279)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_3),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_249),
.A2(n_231),
.B1(n_222),
.B2(n_220),
.Y(n_280)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_281),
.Y(n_300)
);

INVx13_ASAP7_75t_L g283 ( 
.A(n_271),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_263),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_246),
.C(n_242),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_288),
.C(n_293),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_270),
.A2(n_247),
.B1(n_240),
.B2(n_241),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_285),
.A2(n_294),
.B1(n_4),
.B2(n_5),
.Y(n_306)
);

NOR2xp67_ASAP7_75t_SL g286 ( 
.A(n_279),
.B(n_243),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_286),
.B(n_6),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_287),
.B(n_279),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_246),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_264),
.A2(n_261),
.B1(n_253),
.B2(n_260),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_265),
.Y(n_301)
);

AOI322xp5_ASAP7_75t_SL g292 ( 
.A1(n_280),
.A2(n_259),
.A3(n_257),
.B1(n_5),
.B2(n_6),
.C1(n_7),
.C2(n_8),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_292),
.A2(n_268),
.B(n_273),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_272),
.B(n_278),
.Y(n_293)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_296),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_267),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_297),
.B(n_299),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_302),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_301),
.B(n_309),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_274),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_266),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_305),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_4),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_307),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_289),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_282),
.B(n_6),
.C(n_7),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_8),
.C(n_9),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_297),
.A2(n_289),
.B(n_295),
.Y(n_311)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_311),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_300),
.A2(n_283),
.B1(n_287),
.B2(n_291),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_314),
.B(n_308),
.Y(n_327)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_317),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_304),
.A2(n_10),
.B(n_11),
.Y(n_319)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_319),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_315),
.B(n_304),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_320),
.B(n_317),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_301),
.Y(n_321)
);

CKINVDCx14_ASAP7_75t_R g328 ( 
.A(n_321),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_318),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_322),
.B(n_327),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_310),
.A2(n_309),
.B(n_299),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_316),
.Y(n_330)
);

A2O1A1O1Ixp25_ASAP7_75t_L g333 ( 
.A1(n_330),
.A2(n_331),
.B(n_327),
.C(n_323),
.D(n_326),
.Y(n_333)
);

AOI31xp67_ASAP7_75t_L g331 ( 
.A1(n_324),
.A2(n_316),
.A3(n_314),
.B(n_312),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_332),
.B(n_10),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_333),
.B(n_334),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_329),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_328),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_337),
.A2(n_10),
.B(n_11),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_11),
.Y(n_339)
);

OAI311xp33_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_11),
.A3(n_12),
.B1(n_331),
.C1(n_338),
.Y(n_340)
);


endmodule