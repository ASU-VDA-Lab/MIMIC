module fake_aes_12446_n_721 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_721);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_721;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_476;
wire n_384;
wire n_227;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_167;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_649;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_159;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_SL g107 ( .A(n_70), .Y(n_107) );
BUFx6f_ASAP7_75t_L g108 ( .A(n_75), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_56), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_28), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_10), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_65), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_86), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_103), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_44), .Y(n_115) );
CKINVDCx16_ASAP7_75t_R g116 ( .A(n_25), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_79), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_50), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_8), .Y(n_119) );
INVxp33_ASAP7_75t_L g120 ( .A(n_11), .Y(n_120) );
INVxp67_ASAP7_75t_SL g121 ( .A(n_20), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_77), .Y(n_122) );
BUFx2_ASAP7_75t_L g123 ( .A(n_73), .Y(n_123) );
BUFx2_ASAP7_75t_SL g124 ( .A(n_78), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_84), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_34), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_59), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_35), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_66), .Y(n_129) );
BUFx2_ASAP7_75t_L g130 ( .A(n_0), .Y(n_130) );
INVx1_ASAP7_75t_SL g131 ( .A(n_15), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_62), .Y(n_132) );
INVxp33_ASAP7_75t_L g133 ( .A(n_57), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_52), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_37), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_81), .Y(n_136) );
NOR2xp67_ASAP7_75t_L g137 ( .A(n_64), .B(n_5), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_38), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_36), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_89), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_42), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_53), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_46), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_106), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_41), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_23), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_1), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_17), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_4), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_24), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_94), .Y(n_151) );
BUFx12f_ASAP7_75t_L g152 ( .A(n_123), .Y(n_152) );
BUFx8_ASAP7_75t_L g153 ( .A(n_123), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_130), .B(n_120), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_136), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_108), .Y(n_156) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_108), .B(n_146), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_136), .Y(n_158) );
INVx6_ASAP7_75t_L g159 ( .A(n_108), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_108), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_122), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_151), .Y(n_162) );
AND2x2_ASAP7_75t_L g163 ( .A(n_130), .B(n_0), .Y(n_163) );
BUFx8_ASAP7_75t_L g164 ( .A(n_108), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_146), .Y(n_165) );
INVxp67_ASAP7_75t_L g166 ( .A(n_111), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_146), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_151), .Y(n_168) );
AND2x4_ASAP7_75t_L g169 ( .A(n_122), .B(n_1), .Y(n_169) );
HB1xp67_ASAP7_75t_L g170 ( .A(n_148), .Y(n_170) );
INVx3_ASAP7_75t_L g171 ( .A(n_169), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_153), .B(n_116), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_169), .Y(n_173) );
INVx3_ASAP7_75t_L g174 ( .A(n_169), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_155), .B(n_145), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_169), .Y(n_176) );
NAND3xp33_ASAP7_75t_L g177 ( .A(n_155), .B(n_150), .C(n_132), .Y(n_177) );
INVx2_ASAP7_75t_SL g178 ( .A(n_164), .Y(n_178) );
INVx2_ASAP7_75t_SL g179 ( .A(n_153), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_152), .B(n_133), .Y(n_180) );
INVx3_ASAP7_75t_L g181 ( .A(n_161), .Y(n_181) );
INVx1_ASAP7_75t_SL g182 ( .A(n_170), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_158), .B(n_145), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_161), .Y(n_184) );
OR2x6_ASAP7_75t_L g185 ( .A(n_163), .B(n_124), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_160), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_160), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_160), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_160), .Y(n_189) );
AND2x2_ASAP7_75t_L g190 ( .A(n_154), .B(n_148), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_153), .B(n_113), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_158), .Y(n_192) );
NAND3xp33_ASAP7_75t_L g193 ( .A(n_162), .B(n_128), .C(n_109), .Y(n_193) );
INVx2_ASAP7_75t_L g194 ( .A(n_160), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_165), .Y(n_195) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_152), .B(n_110), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_192), .Y(n_197) );
INVx3_ASAP7_75t_L g198 ( .A(n_171), .Y(n_198) );
OR2x2_ASAP7_75t_SL g199 ( .A(n_179), .B(n_153), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_192), .Y(n_200) );
AND3x1_ASAP7_75t_L g201 ( .A(n_179), .B(n_163), .C(n_168), .Y(n_201) );
AOI22xp33_ASAP7_75t_L g202 ( .A1(n_185), .A2(n_168), .B1(n_162), .B2(n_164), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_171), .Y(n_203) );
INVxp67_ASAP7_75t_SL g204 ( .A(n_178), .Y(n_204) );
NAND2xp33_ASAP7_75t_L g205 ( .A(n_178), .B(n_113), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_178), .B(n_114), .Y(n_206) );
O2A1O1Ixp5_ASAP7_75t_L g207 ( .A1(n_171), .A2(n_157), .B(n_125), .C(n_126), .Y(n_207) );
BUFx12f_ASAP7_75t_L g208 ( .A(n_185), .Y(n_208) );
AND2x4_ASAP7_75t_L g209 ( .A(n_185), .B(n_166), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_171), .Y(n_210) );
AND2x6_ASAP7_75t_SL g211 ( .A(n_180), .B(n_119), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_182), .B(n_114), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_190), .B(n_115), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_181), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_174), .Y(n_215) );
BUFx8_ASAP7_75t_L g216 ( .A(n_190), .Y(n_216) );
INVxp33_ASAP7_75t_L g217 ( .A(n_196), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_182), .B(n_115), .Y(n_218) );
BUFx12f_ASAP7_75t_L g219 ( .A(n_185), .Y(n_219) );
NAND3xp33_ASAP7_75t_L g220 ( .A(n_177), .B(n_164), .C(n_117), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_173), .B(n_129), .Y(n_221) );
AOI22xp5_ASAP7_75t_L g222 ( .A1(n_185), .A2(n_112), .B1(n_121), .B2(n_149), .Y(n_222) );
INVxp67_ASAP7_75t_L g223 ( .A(n_172), .Y(n_223) );
INVx3_ASAP7_75t_L g224 ( .A(n_174), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_173), .B(n_129), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_181), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_176), .B(n_134), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_181), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_176), .B(n_134), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_174), .B(n_138), .Y(n_230) );
OR2x6_ASAP7_75t_L g231 ( .A(n_208), .B(n_191), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_197), .A2(n_174), .B(n_175), .Y(n_232) );
INVx2_ASAP7_75t_L g233 ( .A(n_197), .Y(n_233) );
OAI22xp33_ASAP7_75t_L g234 ( .A1(n_222), .A2(n_183), .B1(n_175), .B2(n_131), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_197), .A2(n_183), .B(n_177), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_217), .B(n_193), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_198), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_209), .B(n_184), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_209), .B(n_213), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_200), .A2(n_193), .B(n_184), .Y(n_240) );
AND2x2_ASAP7_75t_L g241 ( .A(n_209), .B(n_181), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_198), .Y(n_242) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_208), .Y(n_243) );
AOI22xp33_ASAP7_75t_L g244 ( .A1(n_209), .A2(n_164), .B1(n_147), .B2(n_124), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_200), .A2(n_118), .B(n_140), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_221), .B(n_138), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_200), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_203), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_198), .Y(n_249) );
NOR2xp33_ASAP7_75t_L g250 ( .A(n_223), .B(n_141), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_225), .B(n_141), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_198), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_203), .A2(n_143), .B(n_139), .Y(n_253) );
AND2x4_ASAP7_75t_L g254 ( .A(n_201), .B(n_137), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_210), .A2(n_135), .B(n_127), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g256 ( .A1(n_210), .A2(n_195), .B(n_194), .Y(n_256) );
A2O1A1Ixp33_ASAP7_75t_L g257 ( .A1(n_215), .A2(n_224), .B(n_202), .C(n_227), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_229), .B(n_142), .Y(n_258) );
HB1xp67_ASAP7_75t_L g259 ( .A(n_216), .Y(n_259) );
NAND2x1p5_ASAP7_75t_L g260 ( .A(n_224), .B(n_146), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_224), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_234), .B(n_216), .Y(n_262) );
O2A1O1Ixp33_ASAP7_75t_L g263 ( .A1(n_257), .A2(n_218), .B(n_212), .C(n_230), .Y(n_263) );
O2A1O1Ixp33_ASAP7_75t_SL g264 ( .A1(n_257), .A2(n_220), .B(n_215), .C(n_206), .Y(n_264) );
INVx3_ASAP7_75t_L g265 ( .A(n_233), .Y(n_265) );
OAI21x1_ASAP7_75t_L g266 ( .A1(n_260), .A2(n_207), .B(n_201), .Y(n_266) );
NAND2xp33_ASAP7_75t_L g267 ( .A(n_243), .B(n_222), .Y(n_267) );
OAI21xp5_ASAP7_75t_L g268 ( .A1(n_235), .A2(n_224), .B(n_220), .Y(n_268) );
AO32x2_ASAP7_75t_L g269 ( .A1(n_254), .A2(n_199), .A3(n_211), .B1(n_219), .B2(n_208), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_232), .A2(n_204), .B(n_205), .Y(n_270) );
OAI21x1_ASAP7_75t_L g271 ( .A1(n_260), .A2(n_228), .B(n_226), .Y(n_271) );
BUFx6f_ASAP7_75t_L g272 ( .A(n_243), .Y(n_272) );
NAND2xp5_ASAP7_75t_SL g273 ( .A(n_243), .B(n_216), .Y(n_273) );
INVx1_ASAP7_75t_SL g274 ( .A(n_259), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_241), .Y(n_275) );
OAI21x1_ASAP7_75t_L g276 ( .A1(n_260), .A2(n_228), .B(n_226), .Y(n_276) );
OAI22xp5_ASAP7_75t_L g277 ( .A1(n_238), .A2(n_219), .B1(n_199), .B2(n_226), .Y(n_277) );
NOR2x1_ASAP7_75t_SL g278 ( .A(n_243), .B(n_219), .Y(n_278) );
OAI21x1_ASAP7_75t_L g279 ( .A1(n_240), .A2(n_228), .B(n_214), .Y(n_279) );
OA21x2_ASAP7_75t_L g280 ( .A1(n_245), .A2(n_214), .B(n_167), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_239), .B(n_216), .Y(n_281) );
AO31x2_ASAP7_75t_L g282 ( .A1(n_233), .A2(n_156), .A3(n_167), .B(n_214), .Y(n_282) );
AOI21xp5_ASAP7_75t_L g283 ( .A1(n_247), .A2(n_188), .B(n_195), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_247), .B(n_142), .Y(n_284) );
AND2x2_ASAP7_75t_L g285 ( .A(n_241), .B(n_144), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_265), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_265), .Y(n_287) );
OAI21x1_ASAP7_75t_L g288 ( .A1(n_279), .A2(n_256), .B(n_248), .Y(n_288) );
OAI21xp5_ASAP7_75t_L g289 ( .A1(n_263), .A2(n_236), .B(n_255), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_265), .Y(n_290) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_274), .Y(n_291) );
OAI21x1_ASAP7_75t_L g292 ( .A1(n_279), .A2(n_248), .B(n_253), .Y(n_292) );
OAI21x1_ASAP7_75t_L g293 ( .A1(n_271), .A2(n_276), .B(n_268), .Y(n_293) );
AO31x2_ASAP7_75t_L g294 ( .A1(n_277), .A2(n_167), .A3(n_156), .B(n_261), .Y(n_294) );
OA21x2_ASAP7_75t_L g295 ( .A1(n_271), .A2(n_254), .B(n_156), .Y(n_295) );
INVx1_ASAP7_75t_SL g296 ( .A(n_272), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_262), .B(n_243), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_281), .B(n_211), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_275), .Y(n_299) );
A2O1A1Ixp33_ASAP7_75t_L g300 ( .A1(n_267), .A2(n_254), .B(n_244), .C(n_251), .Y(n_300) );
A2O1A1Ixp33_ASAP7_75t_L g301 ( .A1(n_267), .A2(n_246), .B(n_258), .C(n_237), .Y(n_301) );
OAI21xp5_ASAP7_75t_L g302 ( .A1(n_270), .A2(n_250), .B(n_242), .Y(n_302) );
OAI21x1_ASAP7_75t_L g303 ( .A1(n_276), .A2(n_261), .B(n_252), .Y(n_303) );
NAND2x1p5_ASAP7_75t_L g304 ( .A(n_272), .B(n_249), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_282), .Y(n_305) );
OAI21x1_ASAP7_75t_L g306 ( .A1(n_266), .A2(n_252), .B(n_249), .Y(n_306) );
AND2x4_ASAP7_75t_L g307 ( .A(n_278), .B(n_231), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_305), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_305), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_286), .Y(n_310) );
BUFx2_ASAP7_75t_L g311 ( .A(n_307), .Y(n_311) );
AO21x2_ASAP7_75t_L g312 ( .A1(n_301), .A2(n_264), .B(n_266), .Y(n_312) );
BUFx2_ASAP7_75t_L g313 ( .A(n_307), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_288), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g315 ( .A(n_298), .B(n_273), .Y(n_315) );
AND2x4_ASAP7_75t_L g316 ( .A(n_286), .B(n_272), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_288), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_306), .Y(n_318) );
CKINVDCx5p33_ASAP7_75t_R g319 ( .A(n_291), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_299), .B(n_284), .Y(n_320) );
NAND2x1p5_ASAP7_75t_L g321 ( .A(n_307), .B(n_272), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_287), .Y(n_322) );
INVx2_ASAP7_75t_SL g323 ( .A(n_307), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_287), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_306), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_293), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_290), .Y(n_327) );
HB1xp67_ASAP7_75t_L g328 ( .A(n_297), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_290), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_299), .B(n_284), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_293), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_295), .Y(n_332) );
AO21x2_ASAP7_75t_L g333 ( .A1(n_302), .A2(n_289), .B(n_300), .Y(n_333) );
BUFx3_ASAP7_75t_L g334 ( .A(n_304), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_308), .B(n_295), .Y(n_335) );
OR2x2_ASAP7_75t_L g336 ( .A(n_308), .B(n_295), .Y(n_336) );
INVx3_ASAP7_75t_L g337 ( .A(n_334), .Y(n_337) );
INVx1_ASAP7_75t_SL g338 ( .A(n_311), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_314), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_309), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_309), .B(n_295), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_314), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_332), .B(n_294), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_332), .B(n_294), .Y(n_344) );
OAI21x1_ASAP7_75t_L g345 ( .A1(n_318), .A2(n_292), .B(n_303), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_310), .Y(n_346) );
OAI222xp33_ASAP7_75t_L g347 ( .A1(n_311), .A2(n_231), .B1(n_296), .B2(n_304), .C1(n_269), .C2(n_285), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_314), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_317), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_333), .B(n_294), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_330), .A2(n_231), .B1(n_272), .B2(n_304), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_310), .B(n_294), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_322), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_317), .Y(n_354) );
OR2x6_ASAP7_75t_L g355 ( .A(n_313), .B(n_292), .Y(n_355) );
BUFx3_ASAP7_75t_L g356 ( .A(n_321), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_322), .Y(n_357) );
INVx5_ASAP7_75t_L g358 ( .A(n_334), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_324), .Y(n_359) );
BUFx2_ASAP7_75t_L g360 ( .A(n_313), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_324), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_315), .A2(n_285), .B1(n_231), .B2(n_280), .Y(n_362) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_328), .Y(n_363) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_317), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_327), .B(n_294), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_327), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_329), .B(n_282), .Y(n_367) );
INVx2_ASAP7_75t_SL g368 ( .A(n_334), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_329), .B(n_282), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_318), .Y(n_370) );
BUFx2_ASAP7_75t_L g371 ( .A(n_321), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_333), .B(n_282), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_320), .B(n_282), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_333), .B(n_303), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_320), .B(n_278), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_318), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_325), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_330), .B(n_280), .Y(n_378) );
AND2x4_ASAP7_75t_L g379 ( .A(n_355), .B(n_326), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_340), .B(n_333), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_340), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_335), .B(n_326), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_346), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_346), .B(n_323), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_335), .B(n_326), .Y(n_385) );
INVxp67_ASAP7_75t_SL g386 ( .A(n_364), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_335), .B(n_331), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_370), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_370), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_353), .B(n_323), .Y(n_390) );
INVxp67_ASAP7_75t_SL g391 ( .A(n_364), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_370), .Y(n_392) );
BUFx2_ASAP7_75t_SL g393 ( .A(n_358), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_372), .B(n_331), .Y(n_394) );
NOR2x1_ASAP7_75t_L g395 ( .A(n_347), .B(n_316), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_353), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_372), .B(n_331), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_372), .B(n_325), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_341), .B(n_325), .Y(n_399) );
AND2x4_ASAP7_75t_SL g400 ( .A(n_337), .B(n_316), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_357), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_357), .B(n_359), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_351), .A2(n_319), .B1(n_316), .B2(n_312), .Y(n_403) );
AND3x2_ASAP7_75t_L g404 ( .A(n_371), .B(n_316), .C(n_269), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_359), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_375), .B(n_2), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_361), .B(n_312), .Y(n_407) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_363), .Y(n_408) );
NOR2xp33_ASAP7_75t_SL g409 ( .A(n_347), .B(n_321), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_341), .B(n_312), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_376), .Y(n_411) );
OR2x2_ASAP7_75t_L g412 ( .A(n_363), .B(n_312), .Y(n_412) );
CKINVDCx14_ASAP7_75t_R g413 ( .A(n_360), .Y(n_413) );
INVx3_ASAP7_75t_L g414 ( .A(n_355), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_376), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_351), .A2(n_146), .B1(n_280), .B2(n_269), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_376), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_361), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_352), .B(n_165), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_366), .B(n_280), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_375), .B(n_2), .Y(n_421) );
BUFx2_ASAP7_75t_L g422 ( .A(n_355), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_352), .B(n_165), .Y(n_423) );
AND2x4_ASAP7_75t_L g424 ( .A(n_355), .B(n_165), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_365), .B(n_165), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_377), .Y(n_426) );
INVxp67_ASAP7_75t_SL g427 ( .A(n_377), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_377), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_366), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_365), .B(n_3), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_373), .B(n_3), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_339), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_373), .B(n_4), .Y(n_433) );
NAND2xp5_ASAP7_75t_SL g434 ( .A(n_358), .B(n_144), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_350), .B(n_5), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_336), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_339), .Y(n_437) );
AND2x4_ASAP7_75t_L g438 ( .A(n_355), .B(n_21), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_350), .B(n_6), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_350), .B(n_6), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_343), .B(n_7), .Y(n_441) );
OR2x2_ASAP7_75t_L g442 ( .A(n_360), .B(n_7), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_339), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_367), .B(n_8), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_408), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_408), .Y(n_446) );
INVx2_ASAP7_75t_SL g447 ( .A(n_400), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_381), .Y(n_448) );
OR2x2_ASAP7_75t_L g449 ( .A(n_441), .B(n_338), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_436), .B(n_380), .Y(n_450) );
OR2x2_ASAP7_75t_L g451 ( .A(n_441), .B(n_338), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_413), .B(n_368), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_381), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_430), .B(n_368), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_430), .B(n_368), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_419), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_436), .B(n_336), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_383), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_383), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_435), .B(n_337), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_406), .B(n_9), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_396), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_380), .B(n_367), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_396), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_435), .B(n_337), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_439), .B(n_337), .Y(n_466) );
INVx4_ASAP7_75t_L g467 ( .A(n_438), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_439), .B(n_369), .Y(n_468) );
NOR2xp67_ASAP7_75t_L g469 ( .A(n_414), .B(n_358), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_401), .B(n_369), .Y(n_470) );
INVxp67_ASAP7_75t_SL g471 ( .A(n_386), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_401), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_405), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_419), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_405), .Y(n_475) );
NAND4xp25_ASAP7_75t_L g476 ( .A(n_421), .B(n_362), .C(n_374), .D(n_378), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_423), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_418), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_440), .B(n_371), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_423), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_418), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_429), .B(n_343), .Y(n_482) );
INVx1_ASAP7_75t_SL g483 ( .A(n_393), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_429), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_398), .B(n_378), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_398), .B(n_440), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_425), .B(n_355), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_402), .Y(n_488) );
NOR2x1_ASAP7_75t_L g489 ( .A(n_393), .B(n_356), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_402), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_399), .B(n_343), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_425), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_388), .Y(n_493) );
NAND2x1_ASAP7_75t_L g494 ( .A(n_438), .B(n_344), .Y(n_494) );
BUFx3_ASAP7_75t_L g495 ( .A(n_400), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g496 ( .A1(n_409), .A2(n_344), .B1(n_356), .B2(n_374), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_394), .B(n_344), .Y(n_497) );
AND2x4_ASAP7_75t_L g498 ( .A(n_414), .B(n_358), .Y(n_498) );
AND2x4_ASAP7_75t_L g499 ( .A(n_414), .B(n_358), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_384), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_410), .B(n_374), .Y(n_501) );
INVx2_ASAP7_75t_SL g502 ( .A(n_400), .Y(n_502) );
AND3x2_ASAP7_75t_L g503 ( .A(n_409), .B(n_354), .C(n_349), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_438), .B(n_358), .Y(n_504) );
NOR2x1_ASAP7_75t_L g505 ( .A(n_442), .B(n_356), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_399), .B(n_342), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_384), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_410), .B(n_342), .Y(n_508) );
HB1xp67_ASAP7_75t_L g509 ( .A(n_386), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_390), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_394), .B(n_342), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_390), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_397), .B(n_358), .Y(n_513) );
AND2x4_ASAP7_75t_SL g514 ( .A(n_438), .B(n_348), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_431), .B(n_9), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_412), .B(n_348), .Y(n_516) );
OR2x6_ASAP7_75t_L g517 ( .A(n_395), .B(n_345), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_397), .B(n_348), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_442), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_431), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_412), .B(n_349), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_382), .B(n_349), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_388), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_382), .B(n_354), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_385), .B(n_354), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_433), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_433), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_445), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_509), .Y(n_529) );
A2O1A1Ixp33_ASAP7_75t_L g530 ( .A1(n_494), .A2(n_395), .B(n_414), .C(n_422), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_450), .B(n_407), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_446), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_491), .B(n_391), .Y(n_533) );
AND2x4_ASAP7_75t_L g534 ( .A(n_467), .B(n_422), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_504), .A2(n_391), .B(n_420), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_497), .B(n_385), .Y(n_536) );
NOR2xp33_ASAP7_75t_L g537 ( .A(n_520), .B(n_444), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_486), .B(n_387), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_450), .B(n_407), .Y(n_539) );
INVxp67_ASAP7_75t_SL g540 ( .A(n_509), .Y(n_540) );
INVx2_ASAP7_75t_SL g541 ( .A(n_452), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_488), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_460), .B(n_387), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_506), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_490), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_511), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_493), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_448), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_500), .B(n_388), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_465), .B(n_424), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g551 ( .A1(n_476), .A2(n_461), .B1(n_515), .B2(n_505), .Y(n_551) );
AND2x4_ASAP7_75t_L g552 ( .A(n_467), .B(n_424), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_523), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_453), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_507), .B(n_389), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_510), .B(n_389), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_466), .B(n_424), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_512), .B(n_501), .Y(n_558) );
INVxp67_ASAP7_75t_L g559 ( .A(n_471), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_479), .B(n_424), .Y(n_560) );
NAND5xp2_ASAP7_75t_L g561 ( .A(n_515), .B(n_403), .C(n_416), .D(n_444), .E(n_404), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_458), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_501), .B(n_389), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_454), .B(n_379), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_459), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_462), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_485), .B(n_427), .Y(n_567) );
INVx2_ASAP7_75t_SL g568 ( .A(n_495), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_455), .B(n_379), .Y(n_569) );
HB1xp67_ASAP7_75t_L g570 ( .A(n_471), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_524), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_463), .B(n_392), .Y(n_572) );
INVxp67_ASAP7_75t_L g573 ( .A(n_526), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_463), .B(n_392), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_508), .B(n_427), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_518), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_508), .B(n_420), .Y(n_577) );
INVx2_ASAP7_75t_SL g578 ( .A(n_489), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_464), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_468), .B(n_379), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_472), .Y(n_581) );
NAND2xp5_ASAP7_75t_SL g582 ( .A(n_483), .B(n_379), .Y(n_582) );
OR2x2_ASAP7_75t_L g583 ( .A(n_449), .B(n_392), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_487), .B(n_404), .Y(n_584) );
NAND2xp5_ASAP7_75t_SL g585 ( .A(n_483), .B(n_411), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_473), .Y(n_586) );
OR2x2_ASAP7_75t_L g587 ( .A(n_451), .B(n_411), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_527), .B(n_411), .Y(n_588) );
NAND2x1p5_ASAP7_75t_L g589 ( .A(n_469), .B(n_434), .Y(n_589) );
NAND2x2_ASAP7_75t_L g590 ( .A(n_447), .B(n_269), .Y(n_590) );
INVxp67_ASAP7_75t_SL g591 ( .A(n_516), .Y(n_591) );
HB1xp67_ASAP7_75t_L g592 ( .A(n_522), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_475), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_478), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_481), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_484), .Y(n_596) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_522), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_513), .B(n_415), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_502), .B(n_415), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_482), .Y(n_600) );
AOI211xp5_ASAP7_75t_L g601 ( .A1(n_476), .A2(n_443), .B(n_437), .C(n_432), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_482), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_457), .B(n_415), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_470), .Y(n_604) );
NAND2x1_ASAP7_75t_L g605 ( .A(n_578), .B(n_517), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_600), .B(n_519), .Y(n_606) );
AOI21xp5_ASAP7_75t_L g607 ( .A1(n_535), .A2(n_517), .B(n_514), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_588), .Y(n_608) );
NOR3xp33_ASAP7_75t_L g609 ( .A(n_561), .B(n_470), .C(n_521), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_588), .Y(n_610) );
CKINVDCx16_ASAP7_75t_R g611 ( .A(n_568), .Y(n_611) );
OAI322xp33_ASAP7_75t_L g612 ( .A1(n_551), .A2(n_496), .A3(n_525), .B1(n_521), .B2(n_516), .C1(n_474), .C2(n_456), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_580), .B(n_498), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_536), .B(n_498), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_592), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_543), .B(n_499), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_564), .B(n_499), .Y(n_617) );
INVxp67_ASAP7_75t_SL g618 ( .A(n_570), .Y(n_618) );
OAI22xp5_ASAP7_75t_L g619 ( .A1(n_590), .A2(n_517), .B1(n_477), .B2(n_492), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_602), .B(n_525), .Y(n_620) );
AOI32xp33_ASAP7_75t_L g621 ( .A1(n_601), .A2(n_480), .A3(n_503), .B1(n_443), .B2(n_437), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_569), .B(n_503), .Y(n_622) );
OR2x2_ASAP7_75t_L g623 ( .A(n_567), .B(n_417), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_573), .B(n_10), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_604), .B(n_417), .Y(n_625) );
AOI222xp33_ASAP7_75t_L g626 ( .A1(n_537), .A2(n_443), .B1(n_437), .B2(n_432), .C1(n_428), .C2(n_426), .Y(n_626) );
INVx2_ASAP7_75t_SL g627 ( .A(n_541), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_592), .Y(n_628) );
AOI21xp33_ASAP7_75t_SL g629 ( .A1(n_530), .A2(n_11), .B(n_12), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_591), .B(n_417), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_552), .A2(n_432), .B1(n_428), .B2(n_426), .Y(n_631) );
INVx3_ASAP7_75t_L g632 ( .A(n_552), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_597), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_591), .B(n_426), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_597), .B(n_428), .Y(n_635) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_589), .A2(n_269), .B1(n_159), .B2(n_107), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_542), .Y(n_637) );
OAI221xp5_ASAP7_75t_L g638 ( .A1(n_573), .A2(n_159), .B1(n_13), .B2(n_14), .C(n_15), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_558), .B(n_345), .Y(n_639) );
AOI32xp33_ASAP7_75t_L g640 ( .A1(n_540), .A2(n_345), .A3(n_13), .B1(n_14), .B2(n_16), .Y(n_640) );
AOI21xp5_ASAP7_75t_L g641 ( .A1(n_535), .A2(n_283), .B(n_16), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_561), .A2(n_159), .B1(n_194), .B2(n_189), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_545), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_575), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_558), .B(n_159), .Y(n_645) );
AOI32xp33_ASAP7_75t_L g646 ( .A1(n_540), .A2(n_12), .A3(n_17), .B1(n_18), .B2(n_19), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_538), .B(n_584), .Y(n_647) );
INVx1_ASAP7_75t_SL g648 ( .A(n_529), .Y(n_648) );
NAND2x1_ASAP7_75t_L g649 ( .A(n_534), .B(n_18), .Y(n_649) );
NAND2x1p5_ASAP7_75t_L g650 ( .A(n_534), .B(n_19), .Y(n_650) );
OAI322xp33_ASAP7_75t_L g651 ( .A1(n_559), .A2(n_20), .A3(n_195), .B1(n_194), .B2(n_189), .C1(n_188), .C2(n_187), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_595), .Y(n_652) );
NAND2xp5_ASAP7_75t_SL g653 ( .A(n_559), .B(n_189), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_528), .Y(n_654) );
AOI221x1_ASAP7_75t_L g655 ( .A1(n_629), .A2(n_532), .B1(n_539), .B2(n_531), .C(n_596), .Y(n_655) );
OAI32xp33_ASAP7_75t_L g656 ( .A1(n_611), .A2(n_589), .A3(n_533), .B1(n_582), .B2(n_577), .Y(n_656) );
OAI221xp5_ASAP7_75t_L g657 ( .A1(n_621), .A2(n_531), .B1(n_539), .B2(n_572), .C(n_574), .Y(n_657) );
OAI21xp33_ASAP7_75t_L g658 ( .A1(n_609), .A2(n_574), .B(n_572), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_645), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_608), .Y(n_660) );
OAI221xp5_ASAP7_75t_L g661 ( .A1(n_642), .A2(n_563), .B1(n_548), .B2(n_562), .C(n_594), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_626), .B(n_563), .Y(n_662) );
AND2x2_ASAP7_75t_L g663 ( .A(n_632), .B(n_544), .Y(n_663) );
OAI22xp33_ASAP7_75t_L g664 ( .A1(n_632), .A2(n_571), .B1(n_576), .B2(n_585), .Y(n_664) );
O2A1O1Ixp33_ASAP7_75t_L g665 ( .A1(n_649), .A2(n_549), .B(n_555), .C(n_556), .Y(n_665) );
AOI222xp33_ASAP7_75t_L g666 ( .A1(n_624), .A2(n_565), .B1(n_581), .B2(n_566), .C1(n_593), .C2(n_554), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_610), .Y(n_667) );
OAI322xp33_ASAP7_75t_L g668 ( .A1(n_607), .A2(n_583), .A3(n_587), .B1(n_603), .B2(n_579), .C1(n_586), .C2(n_556), .Y(n_668) );
NAND4xp25_ASAP7_75t_SL g669 ( .A(n_640), .B(n_646), .C(n_626), .D(n_622), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_627), .A2(n_560), .B1(n_550), .B2(n_557), .Y(n_670) );
AOI21xp5_ASAP7_75t_L g671 ( .A1(n_636), .A2(n_549), .B(n_555), .Y(n_671) );
OAI21xp5_ASAP7_75t_SL g672 ( .A1(n_650), .A2(n_599), .B(n_598), .Y(n_672) );
AOI221xp5_ASAP7_75t_SL g673 ( .A1(n_612), .A2(n_546), .B1(n_547), .B2(n_553), .C(n_188), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_637), .Y(n_674) );
AOI221xp5_ASAP7_75t_L g675 ( .A1(n_612), .A2(n_186), .B1(n_187), .B2(n_27), .C(n_29), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g676 ( .A1(n_650), .A2(n_187), .B1(n_186), .B2(n_30), .Y(n_676) );
OAI22xp33_ASAP7_75t_L g677 ( .A1(n_605), .A2(n_186), .B1(n_26), .B2(n_31), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_643), .Y(n_678) );
OAI22xp5_ASAP7_75t_L g679 ( .A1(n_647), .A2(n_22), .B1(n_32), .B2(n_33), .Y(n_679) );
OAI322xp33_ASAP7_75t_L g680 ( .A1(n_618), .A2(n_39), .A3(n_40), .B1(n_43), .B2(n_45), .C1(n_47), .C2(n_48), .Y(n_680) );
OAI21xp33_ASAP7_75t_SL g681 ( .A1(n_614), .A2(n_49), .B(n_51), .Y(n_681) );
AOI31xp33_ASAP7_75t_L g682 ( .A1(n_619), .A2(n_54), .A3(n_55), .B(n_58), .Y(n_682) );
NAND3xp33_ASAP7_75t_SL g683 ( .A(n_675), .B(n_641), .C(n_638), .Y(n_683) );
OAI21xp5_ASAP7_75t_L g684 ( .A1(n_673), .A2(n_653), .B(n_631), .Y(n_684) );
AOI21xp5_ASAP7_75t_L g685 ( .A1(n_665), .A2(n_630), .B(n_634), .Y(n_685) );
AOI222xp33_ASAP7_75t_L g686 ( .A1(n_658), .A2(n_628), .B1(n_615), .B2(n_633), .C1(n_606), .C2(n_648), .Y(n_686) );
O2A1O1Ixp5_ASAP7_75t_L g687 ( .A1(n_656), .A2(n_654), .B(n_639), .C(n_651), .Y(n_687) );
AOI322xp5_ASAP7_75t_L g688 ( .A1(n_662), .A2(n_644), .A3(n_616), .B1(n_648), .B2(n_613), .C1(n_620), .C2(n_617), .Y(n_688) );
INVx2_ASAP7_75t_SL g689 ( .A(n_663), .Y(n_689) );
OAI211xp5_ASAP7_75t_L g690 ( .A1(n_681), .A2(n_652), .B(n_625), .C(n_623), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_669), .A2(n_635), .B1(n_651), .B2(n_63), .Y(n_691) );
INVxp67_ASAP7_75t_SL g692 ( .A(n_664), .Y(n_692) );
AOI221xp5_ASAP7_75t_L g693 ( .A1(n_668), .A2(n_60), .B1(n_61), .B2(n_67), .C(n_68), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_659), .B(n_69), .Y(n_694) );
XOR2x2_ASAP7_75t_L g695 ( .A(n_657), .B(n_71), .Y(n_695) );
AOI21xp5_ASAP7_75t_L g696 ( .A1(n_672), .A2(n_72), .B(n_74), .Y(n_696) );
NAND5xp2_ASAP7_75t_L g697 ( .A(n_691), .B(n_675), .C(n_666), .D(n_671), .E(n_661), .Y(n_697) );
NOR3xp33_ASAP7_75t_L g698 ( .A(n_687), .B(n_680), .C(n_677), .Y(n_698) );
OAI221xp5_ASAP7_75t_SL g699 ( .A1(n_688), .A2(n_692), .B1(n_690), .B2(n_686), .C(n_693), .Y(n_699) );
AOI322xp5_ASAP7_75t_L g700 ( .A1(n_683), .A2(n_670), .A3(n_660), .B1(n_667), .B2(n_678), .C1(n_674), .C2(n_655), .Y(n_700) );
NOR2x1p5_ASAP7_75t_L g701 ( .A(n_694), .B(n_682), .Y(n_701) );
OAI211xp5_ASAP7_75t_L g702 ( .A1(n_684), .A2(n_671), .B(n_679), .C(n_676), .Y(n_702) );
AND2x2_ASAP7_75t_L g703 ( .A(n_689), .B(n_76), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_703), .Y(n_704) );
NOR3xp33_ASAP7_75t_SL g705 ( .A(n_699), .B(n_696), .C(n_685), .Y(n_705) );
NAND4xp25_ASAP7_75t_L g706 ( .A(n_698), .B(n_695), .C(n_82), .D(n_83), .Y(n_706) );
AND2x2_ASAP7_75t_SL g707 ( .A(n_697), .B(n_80), .Y(n_707) );
OAI221xp5_ASAP7_75t_L g708 ( .A1(n_705), .A2(n_702), .B1(n_700), .B2(n_701), .C(n_90), .Y(n_708) );
NAND4xp75_ASAP7_75t_L g709 ( .A(n_707), .B(n_85), .C(n_87), .D(n_88), .Y(n_709) );
NOR2x1_ASAP7_75t_L g710 ( .A(n_706), .B(n_91), .Y(n_710) );
NAND4xp75_ASAP7_75t_L g711 ( .A(n_710), .B(n_704), .C(n_93), .D(n_95), .Y(n_711) );
INVx3_ASAP7_75t_L g712 ( .A(n_709), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_712), .Y(n_713) );
INVx2_ASAP7_75t_SL g714 ( .A(n_711), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_713), .B(n_708), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g716 ( .A1(n_714), .A2(n_92), .B1(n_96), .B2(n_97), .Y(n_716) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_715), .Y(n_717) );
AND2x2_ASAP7_75t_L g718 ( .A(n_717), .B(n_716), .Y(n_718) );
NAND2xp5_ASAP7_75t_SL g719 ( .A(n_718), .B(n_105), .Y(n_719) );
AOI22x1_ASAP7_75t_L g720 ( .A1(n_719), .A2(n_98), .B1(n_99), .B2(n_100), .Y(n_720) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_720), .A2(n_101), .B1(n_102), .B2(n_104), .Y(n_721) );
endmodule