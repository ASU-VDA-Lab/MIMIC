module fake_aes_5086_n_442 (n_117, n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_115, n_97, n_80, n_107, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_16, n_13, n_113, n_95, n_120, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_111, n_79, n_38, n_64, n_46, n_31, n_58, n_118, n_32, n_0, n_84, n_112, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_110, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_109, n_93, n_51, n_96, n_39, n_442);
input n_117;
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_115;
input n_97;
input n_80;
input n_107;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_16;
input n_13;
input n_113;
input n_95;
input n_120;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_111;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_118;
input n_32;
input n_0;
input n_84;
input n_112;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_110;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_51;
input n_96;
input n_39;
output n_442;
wire n_361;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_125;
wire n_431;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_229;
wire n_336;
wire n_348;
wire n_252;
wire n_152;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_131;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_231;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_141;
wire n_167;
wire n_171;
wire n_196;
wire n_192;
wire n_312;
wire n_137;
wire n_277;
wire n_367;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_417;
wire n_241;
wire n_238;
wire n_318;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_299;
wire n_338;
wire n_256;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_271;
wire n_302;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_219;
wire n_133;
wire n_149;
wire n_214;
wire n_204;
wire n_430;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_379;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_193;
wire n_273;
wire n_390;
wire n_245;
wire n_357;
wire n_260;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_419;
wire n_396;
wire n_168;
wire n_398;
wire n_438;
wire n_134;
wire n_429;
wire n_233;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_203;
wire n_300;
wire n_158;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_418;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_371;
wire n_323;
wire n_347;
wire n_258;
wire n_253;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_176;
wire n_123;
wire n_223;
wire n_372;
wire n_194;
wire n_287;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_395;
wire n_406;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g122 ( .A(n_19), .Y(n_122) );
HB1xp67_ASAP7_75t_L g123 ( .A(n_88), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_105), .Y(n_124) );
HB1xp67_ASAP7_75t_L g125 ( .A(n_114), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_62), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_20), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_24), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_90), .Y(n_129) );
INVx1_ASAP7_75t_SL g130 ( .A(n_72), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_96), .Y(n_131) );
INVxp67_ASAP7_75t_SL g132 ( .A(n_92), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_67), .Y(n_133) );
CKINVDCx16_ASAP7_75t_R g134 ( .A(n_18), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_2), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_91), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_93), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_43), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_99), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_71), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_41), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_86), .Y(n_142) );
BUFx10_ASAP7_75t_L g143 ( .A(n_100), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_113), .Y(n_144) );
INVx1_ASAP7_75t_SL g145 ( .A(n_30), .Y(n_145) );
CKINVDCx16_ASAP7_75t_R g146 ( .A(n_109), .Y(n_146) );
NOR2xp67_ASAP7_75t_L g147 ( .A(n_117), .B(n_51), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_81), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_17), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_58), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_27), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_25), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_83), .Y(n_153) );
HB1xp67_ASAP7_75t_L g154 ( .A(n_47), .Y(n_154) );
BUFx10_ASAP7_75t_L g155 ( .A(n_8), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_115), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_26), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_31), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_107), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_50), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_52), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_108), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_77), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_56), .Y(n_164) );
CKINVDCx5p33_ASAP7_75t_R g165 ( .A(n_89), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_60), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_120), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_36), .Y(n_168) );
BUFx3_ASAP7_75t_L g169 ( .A(n_106), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_112), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_35), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_68), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g173 ( .A(n_101), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_79), .Y(n_174) );
CKINVDCx5p33_ASAP7_75t_R g175 ( .A(n_103), .Y(n_175) );
BUFx10_ASAP7_75t_L g176 ( .A(n_97), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_63), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_111), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_0), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_6), .Y(n_180) );
BUFx5_ASAP7_75t_L g181 ( .A(n_4), .Y(n_181) );
HB1xp67_ASAP7_75t_L g182 ( .A(n_37), .Y(n_182) );
CKINVDCx16_ASAP7_75t_R g183 ( .A(n_5), .Y(n_183) );
CKINVDCx5p33_ASAP7_75t_R g184 ( .A(n_23), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_121), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_82), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_2), .Y(n_187) );
INVx2_ASAP7_75t_SL g188 ( .A(n_38), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_46), .Y(n_189) );
BUFx2_ASAP7_75t_L g190 ( .A(n_87), .Y(n_190) );
CKINVDCx16_ASAP7_75t_R g191 ( .A(n_28), .Y(n_191) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_98), .Y(n_192) );
CKINVDCx16_ASAP7_75t_R g193 ( .A(n_119), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_61), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_110), .Y(n_195) );
NOR2xp67_ASAP7_75t_L g196 ( .A(n_118), .B(n_85), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_102), .Y(n_197) );
INVx2_ASAP7_75t_SL g198 ( .A(n_49), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_40), .Y(n_199) );
BUFx2_ASAP7_75t_L g200 ( .A(n_95), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_116), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_104), .Y(n_202) );
CKINVDCx16_ASAP7_75t_R g203 ( .A(n_75), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_94), .Y(n_204) );
HB1xp67_ASAP7_75t_L g205 ( .A(n_7), .Y(n_205) );
OAI22xp5_ASAP7_75t_L g206 ( .A1(n_183), .A2(n_0), .B1(n_1), .B2(n_3), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_181), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_181), .Y(n_208) );
INVx3_ASAP7_75t_L g209 ( .A(n_143), .Y(n_209) );
AND2x2_ASAP7_75t_L g210 ( .A(n_190), .B(n_1), .Y(n_210) );
AND2x4_ASAP7_75t_L g211 ( .A(n_200), .B(n_3), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_181), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_205), .B(n_4), .Y(n_213) );
CKINVDCx6p67_ASAP7_75t_R g214 ( .A(n_143), .Y(n_214) );
AND2x4_ASAP7_75t_L g215 ( .A(n_135), .B(n_5), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_181), .Y(n_216) );
AND2x4_ASAP7_75t_L g217 ( .A(n_123), .B(n_6), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_188), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_198), .Y(n_219) );
AND2x4_ASAP7_75t_L g220 ( .A(n_179), .B(n_7), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_136), .Y(n_221) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_142), .Y(n_222) );
AND2x4_ASAP7_75t_L g223 ( .A(n_125), .B(n_9), .Y(n_223) );
AND2x6_ASAP7_75t_L g224 ( .A(n_122), .B(n_10), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_154), .B(n_11), .Y(n_225) );
INVx2_ASAP7_75t_SL g226 ( .A(n_209), .Y(n_226) );
BUFx6f_ASAP7_75t_L g227 ( .A(n_222), .Y(n_227) );
INVx4_ASAP7_75t_L g228 ( .A(n_224), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_207), .Y(n_229) );
AND2x2_ASAP7_75t_L g230 ( .A(n_214), .B(n_134), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_218), .B(n_182), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_208), .Y(n_232) );
AND2x2_ASAP7_75t_L g233 ( .A(n_210), .B(n_146), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_208), .Y(n_234) );
INVx3_ASAP7_75t_L g235 ( .A(n_215), .Y(n_235) );
OAI22xp33_ASAP7_75t_L g236 ( .A1(n_213), .A2(n_187), .B1(n_180), .B2(n_191), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_212), .Y(n_237) );
CKINVDCx5p33_ASAP7_75t_R g238 ( .A(n_223), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_234), .B(n_224), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_235), .B(n_211), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_226), .B(n_217), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_228), .B(n_193), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_234), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_233), .B(n_225), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_236), .B(n_215), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_237), .B(n_220), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_237), .Y(n_247) );
INVx2_ASAP7_75t_L g248 ( .A(n_232), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_231), .B(n_220), .Y(n_249) );
INVx2_ASAP7_75t_SL g250 ( .A(n_230), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_238), .B(n_219), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_239), .A2(n_228), .B(n_229), .Y(n_252) );
BUFx3_ASAP7_75t_L g253 ( .A(n_250), .Y(n_253) );
A2O1A1Ixp33_ASAP7_75t_L g254 ( .A1(n_245), .A2(n_216), .B(n_212), .C(n_221), .Y(n_254) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_244), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_249), .B(n_203), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_246), .A2(n_247), .B(n_243), .Y(n_257) );
AOI22x1_ASAP7_75t_L g258 ( .A1(n_248), .A2(n_132), .B1(n_141), .B2(n_137), .Y(n_258) );
AOI21x1_ASAP7_75t_L g259 ( .A1(n_242), .A2(n_196), .B(n_147), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_240), .A2(n_127), .B(n_124), .Y(n_260) );
BUFx6f_ASAP7_75t_L g261 ( .A(n_251), .Y(n_261) );
AND2x4_ASAP7_75t_L g262 ( .A(n_241), .B(n_173), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_239), .A2(n_131), .B(n_128), .Y(n_263) );
OAI21xp5_ASAP7_75t_L g264 ( .A1(n_239), .A2(n_139), .B(n_133), .Y(n_264) );
OAI21x1_ASAP7_75t_L g265 ( .A1(n_257), .A2(n_144), .B(n_140), .Y(n_265) );
AOI22xp5_ASAP7_75t_L g266 ( .A1(n_262), .A2(n_206), .B1(n_148), .B2(n_149), .Y(n_266) );
AO31x2_ASAP7_75t_L g267 ( .A1(n_254), .A2(n_150), .A3(n_153), .B(n_151), .Y(n_267) );
O2A1O1Ixp5_ASAP7_75t_L g268 ( .A1(n_259), .A2(n_264), .B(n_263), .C(n_260), .Y(n_268) );
BUFx2_ASAP7_75t_L g269 ( .A(n_253), .Y(n_269) );
A2O1A1Ixp33_ASAP7_75t_L g270 ( .A1(n_256), .A2(n_158), .B(n_159), .C(n_157), .Y(n_270) );
INVx4_ASAP7_75t_L g271 ( .A(n_261), .Y(n_271) );
OAI21xp5_ASAP7_75t_L g272 ( .A1(n_258), .A2(n_163), .B(n_161), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_255), .B(n_164), .Y(n_273) );
AO31x2_ASAP7_75t_L g274 ( .A1(n_254), .A2(n_166), .A3(n_168), .B(n_167), .Y(n_274) );
NOR2x1_ASAP7_75t_SL g275 ( .A(n_261), .B(n_170), .Y(n_275) );
BUFx6f_ASAP7_75t_L g276 ( .A(n_261), .Y(n_276) );
BUFx8_ASAP7_75t_L g277 ( .A(n_253), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_255), .B(n_171), .Y(n_278) );
AOI21xp5_ASAP7_75t_L g279 ( .A1(n_252), .A2(n_177), .B(n_174), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_273), .Y(n_280) );
OAI21x1_ASAP7_75t_L g281 ( .A1(n_265), .A2(n_172), .B(n_162), .Y(n_281) );
OAI21x1_ASAP7_75t_L g282 ( .A1(n_279), .A2(n_268), .B(n_272), .Y(n_282) );
OAI21x1_ASAP7_75t_L g283 ( .A1(n_278), .A2(n_186), .B(n_185), .Y(n_283) );
OAI21xp5_ASAP7_75t_L g284 ( .A1(n_270), .A2(n_194), .B(n_189), .Y(n_284) );
OA21x2_ASAP7_75t_L g285 ( .A1(n_267), .A2(n_197), .B(n_195), .Y(n_285) );
NOR2xp67_ASAP7_75t_L g286 ( .A(n_271), .B(n_12), .Y(n_286) );
OAI21x1_ASAP7_75t_L g287 ( .A1(n_267), .A2(n_201), .B(n_199), .Y(n_287) );
OAI21x1_ASAP7_75t_L g288 ( .A1(n_274), .A2(n_204), .B(n_202), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_275), .Y(n_289) );
OAI21x1_ASAP7_75t_L g290 ( .A1(n_266), .A2(n_156), .B(n_142), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_276), .Y(n_291) );
OAI21x1_ASAP7_75t_L g292 ( .A1(n_276), .A2(n_156), .B(n_142), .Y(n_292) );
OAI21x1_ASAP7_75t_L g293 ( .A1(n_277), .A2(n_13), .B(n_14), .Y(n_293) );
AO21x2_ASAP7_75t_L g294 ( .A1(n_272), .A2(n_176), .B(n_155), .Y(n_294) );
OAI21x1_ASAP7_75t_L g295 ( .A1(n_265), .A2(n_15), .B(n_16), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_277), .Y(n_296) );
INVx4_ASAP7_75t_L g297 ( .A(n_276), .Y(n_297) );
OA21x2_ASAP7_75t_L g298 ( .A1(n_265), .A2(n_145), .B(n_130), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_273), .Y(n_299) );
BUFx2_ASAP7_75t_L g300 ( .A(n_276), .Y(n_300) );
OR2x6_ASAP7_75t_L g301 ( .A(n_269), .B(n_169), .Y(n_301) );
OAI21xp5_ASAP7_75t_L g302 ( .A1(n_270), .A2(n_129), .B(n_126), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_265), .Y(n_303) );
OAI21x1_ASAP7_75t_L g304 ( .A1(n_265), .A2(n_21), .B(n_22), .Y(n_304) );
AO21x2_ASAP7_75t_L g305 ( .A1(n_272), .A2(n_222), .B(n_227), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_299), .Y(n_306) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_289), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g308 ( .A1(n_281), .A2(n_152), .B(n_138), .Y(n_308) );
INVx2_ASAP7_75t_L g309 ( .A(n_285), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_291), .Y(n_310) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_300), .Y(n_311) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_292), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_286), .Y(n_313) );
OAI21x1_ASAP7_75t_L g314 ( .A1(n_290), .A2(n_29), .B(n_32), .Y(n_314) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_298), .Y(n_315) );
INVx2_ASAP7_75t_SL g316 ( .A(n_296), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_282), .B(n_160), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_294), .Y(n_318) );
INVx3_ASAP7_75t_L g319 ( .A(n_301), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_283), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_287), .Y(n_321) );
NAND2x1p5_ASAP7_75t_L g322 ( .A(n_293), .B(n_227), .Y(n_322) );
OAI21xp5_ASAP7_75t_L g323 ( .A1(n_288), .A2(n_175), .B(n_165), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_284), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_295), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_302), .B(n_178), .Y(n_326) );
INVx4_ASAP7_75t_L g327 ( .A(n_305), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_304), .Y(n_328) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_300), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_280), .Y(n_330) );
HB1xp67_ASAP7_75t_L g331 ( .A(n_303), .Y(n_331) );
BUFx2_ASAP7_75t_L g332 ( .A(n_297), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_280), .Y(n_333) );
AO21x2_ASAP7_75t_L g334 ( .A1(n_303), .A2(n_227), .B(n_34), .Y(n_334) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_303), .Y(n_335) );
OR2x2_ASAP7_75t_L g336 ( .A(n_307), .B(n_184), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_331), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_306), .B(n_192), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_330), .Y(n_339) );
AND2x4_ASAP7_75t_L g340 ( .A(n_307), .B(n_33), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_333), .Y(n_341) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_311), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_331), .Y(n_343) );
BUFx2_ASAP7_75t_L g344 ( .A(n_332), .Y(n_344) );
BUFx3_ASAP7_75t_L g345 ( .A(n_316), .Y(n_345) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_311), .Y(n_346) );
BUFx2_ASAP7_75t_L g347 ( .A(n_329), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_335), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_310), .Y(n_349) );
INVxp67_ASAP7_75t_SL g350 ( .A(n_335), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_318), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_315), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_319), .B(n_39), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_319), .B(n_42), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_315), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_309), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_313), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_320), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_324), .B(n_44), .Y(n_359) );
AND2x4_ASAP7_75t_L g360 ( .A(n_321), .B(n_45), .Y(n_360) );
NAND2x1p5_ASAP7_75t_L g361 ( .A(n_326), .B(n_48), .Y(n_361) );
HB1xp67_ASAP7_75t_L g362 ( .A(n_323), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_322), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_325), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_314), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_308), .A2(n_53), .B1(n_54), .B2(n_55), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_328), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_337), .B(n_317), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_344), .B(n_317), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_339), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_341), .Y(n_371) );
OR2x2_ASAP7_75t_L g372 ( .A(n_342), .B(n_327), .Y(n_372) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_346), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_357), .B(n_334), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_337), .B(n_334), .Y(n_375) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_350), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_343), .B(n_312), .Y(n_377) );
BUFx2_ASAP7_75t_L g378 ( .A(n_347), .Y(n_378) );
OR2x2_ASAP7_75t_L g379 ( .A(n_349), .B(n_312), .Y(n_379) );
OR2x2_ASAP7_75t_L g380 ( .A(n_348), .B(n_312), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_348), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_362), .B(n_57), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_351), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_364), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_356), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_367), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_340), .B(n_59), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_356), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_352), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_352), .Y(n_390) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_355), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_378), .B(n_355), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_373), .B(n_358), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_369), .B(n_345), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_376), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_385), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_370), .B(n_360), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_384), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_371), .B(n_363), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_383), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_381), .B(n_353), .Y(n_401) );
NOR2xp33_ASAP7_75t_SL g402 ( .A(n_387), .B(n_361), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_389), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_390), .B(n_354), .Y(n_404) );
AND2x4_ASAP7_75t_L g405 ( .A(n_372), .B(n_391), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_391), .B(n_336), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_400), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_405), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_393), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_398), .Y(n_410) );
NAND2x1_ASAP7_75t_L g411 ( .A(n_395), .B(n_394), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_403), .Y(n_412) );
CKINVDCx16_ASAP7_75t_R g413 ( .A(n_402), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_406), .B(n_368), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_398), .Y(n_415) );
OR2x2_ASAP7_75t_L g416 ( .A(n_392), .B(n_388), .Y(n_416) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_396), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_417), .Y(n_418) );
CKINVDCx16_ASAP7_75t_R g419 ( .A(n_413), .Y(n_419) );
INVxp67_ASAP7_75t_L g420 ( .A(n_411), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_409), .B(n_399), .Y(n_421) );
NOR2xp33_ASAP7_75t_SL g422 ( .A(n_408), .B(n_397), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_410), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_419), .B(n_414), .Y(n_424) );
OAI22xp5_ASAP7_75t_L g425 ( .A1(n_420), .A2(n_416), .B1(n_407), .B2(n_412), .Y(n_425) );
OAI22xp33_ASAP7_75t_L g426 ( .A1(n_422), .A2(n_410), .B1(n_404), .B2(n_401), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_418), .B(n_415), .Y(n_427) );
NOR3xp33_ASAP7_75t_SL g428 ( .A(n_424), .B(n_421), .C(n_338), .Y(n_428) );
NOR2x1_ASAP7_75t_SL g429 ( .A(n_425), .B(n_423), .Y(n_429) );
OAI322xp33_ASAP7_75t_L g430 ( .A1(n_429), .A2(n_426), .A3(n_427), .B1(n_380), .B2(n_386), .C1(n_377), .C2(n_379), .Y(n_430) );
NAND3xp33_ASAP7_75t_L g431 ( .A(n_428), .B(n_366), .C(n_382), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_431), .B(n_374), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_432), .B(n_430), .Y(n_433) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_432), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_434), .Y(n_435) );
OAI22x1_ASAP7_75t_L g436 ( .A1(n_435), .A2(n_433), .B1(n_434), .B2(n_359), .Y(n_436) );
AOI21xp5_ASAP7_75t_L g437 ( .A1(n_436), .A2(n_375), .B(n_365), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g438 ( .A1(n_437), .A2(n_64), .B1(n_65), .B2(n_66), .Y(n_438) );
AOI21xp5_ASAP7_75t_L g439 ( .A1(n_438), .A2(n_69), .B(n_70), .Y(n_439) );
AO21x2_ASAP7_75t_L g440 ( .A1(n_439), .A2(n_73), .B(n_74), .Y(n_440) );
AO21x2_ASAP7_75t_L g441 ( .A1(n_440), .A2(n_76), .B(n_78), .Y(n_441) );
AOI21xp33_ASAP7_75t_SL g442 ( .A1(n_441), .A2(n_80), .B(n_84), .Y(n_442) );
endmodule