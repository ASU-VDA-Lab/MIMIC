module fake_jpeg_5699_n_309 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_309);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_309;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_11),
.B(n_2),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_6),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_36),
.B(n_43),
.Y(n_94)
);

BUFx16f_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_37),
.Y(n_63)
);

NAND3xp33_ASAP7_75t_SL g38 ( 
.A(n_34),
.B(n_0),
.C(n_1),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_38),
.B(n_20),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_45),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_0),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_41),
.B(n_25),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_44),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_17),
.B(n_6),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_25),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_20),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_23),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_17),
.B(n_6),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_48),
.B(n_50),
.Y(n_66)
);

INVx2_ASAP7_75t_R g49 ( 
.A(n_31),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_49),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_20),
.B(n_7),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_52),
.B(n_90),
.Y(n_129)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_53),
.B(n_59),
.Y(n_102)
);

AOI21xp33_ASAP7_75t_SL g55 ( 
.A1(n_49),
.A2(n_23),
.B(n_16),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_55),
.B(n_76),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_49),
.A2(n_24),
.B1(n_18),
.B2(n_30),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_56),
.A2(n_67),
.B(n_83),
.Y(n_108)
);

AO22x1_ASAP7_75t_SL g58 ( 
.A1(n_49),
.A2(n_35),
.B1(n_22),
.B2(n_19),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_58),
.A2(n_19),
.B1(n_23),
.B2(n_32),
.Y(n_113)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_62),
.Y(n_126)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_64),
.A2(n_85),
.B1(n_92),
.B2(n_93),
.Y(n_119)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx3_ASAP7_75t_SL g117 ( 
.A(n_65),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_44),
.A2(n_24),
.B1(n_18),
.B2(n_30),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_68),
.B(n_70),
.Y(n_103)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_71),
.B(n_79),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_41),
.B(n_26),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_72),
.B(n_74),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_75),
.B(n_77),
.Y(n_115)
);

AND2x2_ASAP7_75t_SL g76 ( 
.A(n_42),
.B(n_16),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_36),
.B(n_26),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_38),
.Y(n_79)
);

CKINVDCx12_ASAP7_75t_R g80 ( 
.A(n_40),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_80),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_41),
.B(n_27),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_81),
.B(n_82),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_40),
.B(n_28),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_45),
.A2(n_24),
.B1(n_18),
.B2(n_30),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_84),
.B(n_88),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_46),
.A2(n_33),
.B1(n_35),
.B2(n_22),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_43),
.B(n_28),
.C(n_15),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_86),
.A2(n_94),
.B1(n_66),
.B2(n_90),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_87),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_46),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_50),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_89),
.B(n_96),
.Y(n_128)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_91),
.Y(n_123)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_37),
.Y(n_92)
);

AND2x2_ASAP7_75t_SL g93 ( 
.A(n_49),
.B(n_16),
.Y(n_93)
);

AND2x4_ASAP7_75t_SL g95 ( 
.A(n_49),
.B(n_35),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_95),
.A2(n_19),
.B1(n_29),
.B2(n_21),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_41),
.B(n_27),
.Y(n_96)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_97),
.Y(n_104)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_39),
.Y(n_98)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_98),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_41),
.B(n_15),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_33),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_58),
.A2(n_22),
.B1(n_33),
.B2(n_19),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_101),
.A2(n_85),
.B1(n_58),
.B2(n_83),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_110),
.B(n_86),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_124),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_113),
.A2(n_73),
.B1(n_79),
.B2(n_61),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_74),
.B(n_54),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_122),
.B(n_125),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_82),
.B(n_0),
.Y(n_125)
);

A2O1A1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_129),
.A2(n_55),
.B(n_95),
.C(n_93),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_130),
.B(n_141),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_76),
.C(n_93),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_132),
.B(n_156),
.C(n_163),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_112),
.B(n_95),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_133),
.A2(n_115),
.B(n_120),
.Y(n_184)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_134),
.B(n_137),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_84),
.Y(n_135)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_135),
.Y(n_168)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_138),
.A2(n_115),
.B(n_120),
.Y(n_187)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_103),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_139),
.B(n_140),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_128),
.B(n_87),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_128),
.B(n_87),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_102),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_142),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_98),
.Y(n_143)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_143),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_144),
.A2(n_161),
.B1(n_113),
.B2(n_125),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_145),
.A2(n_116),
.B1(n_129),
.B2(n_108),
.Y(n_170)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_103),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_146),
.B(n_153),
.Y(n_179)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_106),
.Y(n_147)
);

INVx11_ASAP7_75t_L g190 ( 
.A(n_147),
.Y(n_190)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_148),
.Y(n_165)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_126),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_149),
.Y(n_182)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_126),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_150),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_102),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_154),
.Y(n_167)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_106),
.Y(n_152)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_152),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_111),
.B(n_73),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_122),
.B(n_57),
.Y(n_154)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_117),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_155),
.Y(n_169)
);

MAJx2_ASAP7_75t_L g156 ( 
.A(n_114),
.B(n_76),
.C(n_69),
.Y(n_156)
);

INVx6_ASAP7_75t_L g157 ( 
.A(n_117),
.Y(n_157)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_157),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_118),
.B(n_64),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_158),
.B(n_159),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_118),
.B(n_92),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_107),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_160),
.B(n_164),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_119),
.A2(n_56),
.B1(n_67),
.B2(n_61),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g162 ( 
.A(n_106),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_100),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_108),
.B(n_63),
.C(n_91),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_110),
.B(n_97),
.Y(n_164)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_170),
.Y(n_205)
);

AND2x6_ASAP7_75t_L g171 ( 
.A(n_133),
.B(n_132),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_171),
.B(n_174),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_172),
.A2(n_127),
.B1(n_152),
.B2(n_149),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_133),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_176),
.B(n_109),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_130),
.A2(n_144),
.B1(n_145),
.B2(n_163),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_177),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_161),
.A2(n_146),
.B(n_131),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_181),
.A2(n_184),
.B(n_196),
.Y(n_211)
);

O2A1O1Ixp33_ASAP7_75t_L g183 ( 
.A1(n_153),
.A2(n_114),
.B(n_116),
.C(n_100),
.Y(n_183)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_183),
.Y(n_215)
);

NOR3xp33_ASAP7_75t_SL g210 ( 
.A(n_187),
.B(n_188),
.C(n_32),
.Y(n_210)
);

NOR3xp33_ASAP7_75t_SL g188 ( 
.A(n_156),
.B(n_60),
.C(n_105),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_131),
.A2(n_136),
.B1(n_157),
.B2(n_155),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_191),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_136),
.B(n_104),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_192),
.B(n_179),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_131),
.B(n_53),
.C(n_107),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_197),
.C(n_3),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_148),
.A2(n_104),
.B(n_147),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_162),
.B(n_105),
.C(n_70),
.Y(n_197)
);

OA21x2_ASAP7_75t_L g199 ( 
.A1(n_150),
.A2(n_71),
.B(n_109),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_199),
.A2(n_3),
.B(n_5),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_150),
.Y(n_200)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_200),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_201),
.A2(n_216),
.B(n_184),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_202),
.A2(n_212),
.B1(n_183),
.B2(n_176),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_181),
.A2(n_127),
.B1(n_29),
.B2(n_21),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_204),
.B(n_209),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_214),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_178),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_210),
.A2(n_185),
.B1(n_167),
.B2(n_176),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_172),
.A2(n_29),
.B1(n_32),
.B2(n_2),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_188),
.A2(n_32),
.B1(n_7),
.B2(n_8),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_213),
.A2(n_169),
.B(n_193),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_179),
.B(n_0),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_177),
.B(n_32),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_168),
.B(n_1),
.Y(n_217)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_217),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_189),
.B(n_1),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_225),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_168),
.B(n_2),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_219),
.B(n_220),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_3),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_221),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_224),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_223),
.B(n_175),
.C(n_195),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_197),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_189),
.B(n_174),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_227),
.C(n_238),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_225),
.B(n_175),
.C(n_171),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_229),
.A2(n_234),
.B(n_235),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_230),
.A2(n_239),
.B1(n_245),
.B2(n_222),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_211),
.A2(n_203),
.B(n_215),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_211),
.A2(n_191),
.B(n_170),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_205),
.C(n_206),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_207),
.A2(n_180),
.B1(n_187),
.B2(n_186),
.Y(n_239)
);

OAI322xp33_ASAP7_75t_L g257 ( 
.A1(n_242),
.A2(n_210),
.A3(n_213),
.B1(n_216),
.B2(n_214),
.C1(n_220),
.C2(n_209),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_186),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_243),
.A2(n_216),
.B1(n_202),
.B2(n_218),
.Y(n_249)
);

NOR3xp33_ASAP7_75t_SL g244 ( 
.A(n_210),
.B(n_167),
.C(n_198),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_246),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_215),
.A2(n_205),
.B(n_201),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_208),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_248),
.B(n_259),
.C(n_241),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_249),
.B(n_258),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_250),
.A2(n_243),
.B1(n_228),
.B2(n_230),
.Y(n_268)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_231),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_253),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_223),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_239),
.Y(n_264)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_231),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_240),
.Y(n_254)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_254),
.Y(n_265)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_243),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_261),
.Y(n_266)
);

AOI321xp33_ASAP7_75t_L g272 ( 
.A1(n_257),
.A2(n_236),
.A3(n_237),
.B1(n_241),
.B2(n_185),
.C(n_199),
.Y(n_272)
);

XOR2x1_ASAP7_75t_SL g258 ( 
.A(n_229),
.B(n_216),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_226),
.B(n_236),
.C(n_235),
.Y(n_259)
);

A2O1A1O1Ixp25_ASAP7_75t_L g260 ( 
.A1(n_233),
.A2(n_200),
.B(n_217),
.C(n_219),
.D(n_199),
.Y(n_260)
);

MAJx2_ASAP7_75t_L g263 ( 
.A(n_260),
.B(n_246),
.C(n_244),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_232),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_263),
.B(n_264),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_268),
.A2(n_270),
.B1(n_255),
.B2(n_249),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_259),
.A2(n_228),
.B(n_234),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_269),
.B(n_272),
.Y(n_279)
);

AO22x1_ASAP7_75t_SL g270 ( 
.A1(n_258),
.A2(n_245),
.B1(n_242),
.B2(n_240),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_256),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_273),
.B(n_256),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_247),
.C(n_248),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_260),
.B(n_182),
.Y(n_275)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_275),
.Y(n_284)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_276),
.Y(n_287)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_277),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_266),
.Y(n_278)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_278),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_173),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_282),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_270),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_273),
.A2(n_254),
.B1(n_262),
.B2(n_247),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_283),
.A2(n_279),
.B1(n_270),
.B2(n_278),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_254),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_285),
.B(n_286),
.C(n_274),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_291),
.C(n_294),
.Y(n_300)
);

AOI21x1_ASAP7_75t_L g292 ( 
.A1(n_281),
.A2(n_267),
.B(n_263),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_292),
.A2(n_293),
.B1(n_190),
.B2(n_165),
.Y(n_299)
);

INVx11_ASAP7_75t_L g293 ( 
.A(n_281),
.Y(n_293)
);

AOI322xp5_ASAP7_75t_L g294 ( 
.A1(n_284),
.A2(n_267),
.A3(n_252),
.B1(n_237),
.B2(n_286),
.C1(n_165),
.C2(n_169),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_194),
.Y(n_296)
);

OAI221xp5_ASAP7_75t_L g305 ( 
.A1(n_296),
.A2(n_301),
.B1(n_291),
.B2(n_292),
.C(n_190),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_289),
.B(n_194),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_297),
.B(n_298),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_290),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_287),
.C(n_289),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_173),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_303),
.A2(n_288),
.B(n_298),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_300),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_304),
.A2(n_305),
.B1(n_293),
.B2(n_302),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_306),
.B(n_307),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_308),
.B(n_8),
.Y(n_309)
);


endmodule