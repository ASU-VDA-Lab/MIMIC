module real_jpeg_17189_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_531;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_0),
.A2(n_20),
.B(n_532),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_0),
.B(n_533),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_1),
.B(n_207),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_1),
.B(n_107),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_1),
.B(n_276),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_1),
.B(n_302),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_1),
.B(n_130),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_1),
.B(n_416),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_1),
.B(n_420),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_1),
.B(n_436),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_2),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g249 ( 
.A(n_2),
.Y(n_249)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_2),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_3),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_3),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_3),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_3),
.B(n_119),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_3),
.B(n_82),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_3),
.B(n_196),
.Y(n_250)
);

NAND2x1_ASAP7_75t_L g251 ( 
.A(n_3),
.B(n_252),
.Y(n_251)
);

AOI22x1_ASAP7_75t_SL g326 ( 
.A1(n_3),
.A2(n_16),
.B1(n_130),
.B2(n_327),
.Y(n_326)
);

CKINVDCx14_ASAP7_75t_R g354 ( 
.A(n_3),
.Y(n_354)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_4),
.Y(n_68)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_4),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_4),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_4),
.Y(n_364)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_5),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_5),
.B(n_99),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_5),
.B(n_114),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_5),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_5),
.B(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_6),
.Y(n_300)
);

BUFx5_ASAP7_75t_L g311 ( 
.A(n_6),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_6),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_7),
.B(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_7),
.B(n_58),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_7),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_7),
.B(n_81),
.Y(n_136)
);

NAND2x1_ASAP7_75t_SL g208 ( 
.A(n_7),
.B(n_209),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_7),
.B(n_198),
.Y(n_278)
);

AND2x2_ASAP7_75t_SL g287 ( 
.A(n_7),
.B(n_288),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_7),
.B(n_315),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_8),
.B(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_8),
.B(n_363),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_8),
.B(n_381),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_8),
.B(n_405),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_8),
.B(n_450),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g461 ( 
.A(n_8),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_9),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_9),
.B(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_9),
.B(n_31),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_9),
.B(n_58),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_9),
.B(n_236),
.Y(n_235)
);

INVxp33_ASAP7_75t_L g282 ( 
.A(n_9),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_9),
.B(n_311),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_9),
.B(n_248),
.Y(n_360)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g198 ( 
.A(n_10),
.Y(n_198)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_10),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_10),
.Y(n_470)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_11),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_11),
.B(n_107),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_11),
.B(n_242),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_11),
.B(n_256),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_11),
.B(n_298),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_11),
.B(n_209),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_11),
.B(n_198),
.Y(n_359)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_11),
.B(n_99),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_12),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_12),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_12),
.B(n_86),
.Y(n_85)
);

NAND2x1_ASAP7_75t_SL g129 ( 
.A(n_12),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_12),
.B(n_165),
.Y(n_164)
);

AND2x4_ASAP7_75t_L g195 ( 
.A(n_12),
.B(n_196),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_12),
.B(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_13),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_13),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_13),
.Y(n_296)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_13),
.Y(n_408)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_14),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_14),
.Y(n_239)
);

BUFx5_ASAP7_75t_L g387 ( 
.A(n_14),
.Y(n_387)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_14),
.Y(n_453)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_15),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_16),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_16),
.B(n_232),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_16),
.B(n_295),
.Y(n_294)
);

AOI31xp33_ASAP7_75t_L g349 ( 
.A1(n_16),
.A2(n_326),
.A3(n_350),
.B(n_353),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_16),
.B(n_385),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_16),
.B(n_252),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_16),
.B(n_413),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_16),
.B(n_99),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_17),
.Y(n_162)
);

BUFx8_ASAP7_75t_L g82 ( 
.A(n_18),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_18),
.Y(n_108)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_18),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_172),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_170),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_143),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_23),
.B(n_143),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_110),
.C(n_124),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_24),
.B(n_176),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_78),
.C(n_95),
.Y(n_24)
);

INVxp33_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_26),
.B(n_182),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_46),
.C(n_62),
.Y(n_26)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_27),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_SL g27 ( 
.A(n_28),
.B(n_34),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_28),
.B(n_36),
.C(n_42),
.Y(n_121)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_33),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_36),
.B1(n_42),
.B2(n_43),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_35),
.A2(n_36),
.B1(n_113),
.B2(n_115),
.Y(n_112)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_SL g134 ( 
.A(n_36),
.B(n_113),
.C(n_116),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_42),
.A2(n_43),
.B1(n_98),
.B2(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_43),
.Y(n_42)
);

MAJx2_ASAP7_75t_L g97 ( 
.A(n_43),
.B(n_98),
.C(n_101),
.Y(n_97)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_45),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_46),
.B(n_62),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_52),
.C(n_56),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_47),
.B(n_57),
.Y(n_189)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_52),
.B(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_55),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_61),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_69),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_63),
.B(n_70),
.C(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_68),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_75),
.Y(n_69)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_74),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_75),
.Y(n_123)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_79),
.B(n_95),
.Y(n_182)
);

XNOR2x1_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_83),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_80),
.B(n_84),
.C(n_94),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_90),
.B2(n_94),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_89),
.Y(n_242)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_90),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

MAJx2_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_104),
.C(n_109),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_96),
.A2(n_97),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_97),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_98),
.B(n_191),
.C(n_195),
.Y(n_190)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_98),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_98),
.A2(n_195),
.B1(n_203),
.B2(n_229),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_100),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_101),
.A2(n_200),
.B1(n_201),
.B2(n_202),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_101),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_101),
.A2(n_200),
.B1(n_278),
.B2(n_279),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_104),
.B(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_105),
.B(n_109),
.Y(n_214)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_106),
.B(n_247),
.C(n_250),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g309 ( 
.A(n_108),
.Y(n_309)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_109),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_109),
.A2(n_211),
.B1(n_212),
.B2(n_262),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_110),
.A2(n_124),
.B1(n_125),
.B2(n_177),
.Y(n_176)
);

INVxp33_ASAP7_75t_SL g177 ( 
.A(n_110),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_121),
.C(n_122),
.Y(n_110)
);

XNOR2x2_ASAP7_75t_SL g183 ( 
.A(n_111),
.B(n_184),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_116),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_113),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_113),
.A2(n_115),
.B1(n_138),
.B2(n_142),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_114),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_136),
.C(n_138),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_118),
.Y(n_116)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_120),
.Y(n_167)
);

INVx3_ASAP7_75t_SL g207 ( 
.A(n_120),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_121),
.B(n_122),
.Y(n_184)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_133),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_126),
.B(n_134),
.C(n_169),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_132),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_129),
.C(n_132),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_135),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_138),
.Y(n_142)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_138),
.Y(n_163)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_141),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_142),
.A2(n_156),
.B1(n_157),
.B2(n_163),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_168),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_153),
.B2(n_154),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_150),
.B1(n_151),
.B2(n_152),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_149),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_150),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_164),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_162),
.Y(n_258)
);

BUFx5_ASAP7_75t_L g383 ( 
.A(n_162),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVxp33_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_216),
.B(n_528),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g529 ( 
.A1(n_174),
.A2(n_530),
.B(n_531),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_178),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g531 ( 
.A(n_175),
.B(n_178),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_183),
.C(n_185),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_180),
.A2(n_181),
.B1(n_183),
.B2(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_183),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_185),
.B(n_264),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_204),
.C(n_213),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XNOR2x1_ASAP7_75t_L g220 ( 
.A(n_187),
.B(n_221),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_190),
.C(n_199),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_188),
.B(n_190),
.Y(n_512)
);

XNOR2x1_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_228),
.Y(n_227)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_195),
.Y(n_229)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_198),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_199),
.B(n_512),
.Y(n_511)
);

MAJx2_ASAP7_75t_L g328 ( 
.A(n_200),
.B(n_275),
.C(n_278),
.Y(n_328)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_213),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_211),
.C(n_212),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_205),
.B(n_261),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_208),
.C(n_210),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_206),
.B(n_210),
.Y(n_244)
);

XOR2x1_ASAP7_75t_L g243 ( 
.A(n_208),
.B(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_211),
.Y(n_262)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_214),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_266),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_263),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_219),
.B(n_263),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_222),
.C(n_225),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_220),
.B(n_222),
.Y(n_521)
);

XNOR2x1_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_225),
.B(n_521),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_245),
.C(n_259),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_226),
.B(n_510),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_230),
.C(n_243),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_227),
.B(n_230),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_235),
.C(n_240),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_231),
.A2(n_240),
.B1(n_241),
.B2(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_231),
.Y(n_319)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_235),
.B(n_318),
.Y(n_317)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_238),
.Y(n_304)
);

INVx6_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_240),
.B(n_380),
.C(n_384),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_240),
.A2(n_241),
.B1(n_380),
.B2(n_430),
.Y(n_429)
);

INVx2_ASAP7_75t_SL g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_243),
.B(n_337),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_245),
.B(n_260),
.Y(n_510)
);

MAJx2_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_251),
.C(n_254),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_246),
.B(n_333),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_247),
.B(n_250),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_251),
.B(n_255),
.Y(n_333)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_254),
.A2(n_255),
.B1(n_361),
.B2(n_362),
.Y(n_487)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_255),
.B(n_358),
.C(n_361),
.Y(n_357)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_258),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

AO21x2_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_501),
.B(n_525),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_394),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_340),
.C(n_368),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_270),
.B(n_341),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_320),
.Y(n_270)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_271),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_305),
.C(n_317),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_272),
.B(n_343),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_280),
.C(n_292),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

XNOR2x1_ASAP7_75t_SL g390 ( 
.A(n_274),
.B(n_391),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_277),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_278),
.Y(n_279)
);

XNOR2x1_ASAP7_75t_L g391 ( 
.A(n_280),
.B(n_293),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_287),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_281),
.B(n_287),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx6_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx6_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_290),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g356 ( 
.A(n_290),
.Y(n_356)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_297),
.C(n_301),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_294),
.A2(n_297),
.B1(n_376),
.B2(n_377),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_294),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_297),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_297),
.A2(n_377),
.B1(n_448),
.B2(n_449),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_297),
.Y(n_478)
);

BUFx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_300),
.Y(n_439)
);

XOR2x2_ASAP7_75t_SL g374 ( 
.A(n_301),
.B(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_305),
.B(n_317),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_312),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_306),
.B(n_313),
.C(n_331),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.C(n_310),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_307),
.A2(n_310),
.B1(n_347),
.B2(n_348),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_307),
.Y(n_347)
);

XNOR2x2_ASAP7_75t_SL g402 ( 
.A(n_307),
.B(n_403),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_308),
.B(n_346),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_310),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_314),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g460 ( 
.A(n_316),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_321),
.A2(n_336),
.B1(n_338),
.B2(n_339),
.Y(n_320)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_321),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_329),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g505 ( 
.A(n_322),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_325),
.C(n_328),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_323),
.B(n_366),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_325),
.A2(n_326),
.B1(n_328),
.B2(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_328),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_330),
.A2(n_332),
.B1(n_334),
.B2(n_335),
.Y(n_329)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_330),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_330),
.Y(n_506)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_332),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_335),
.Y(n_507)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_336),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_336),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_338),
.Y(n_516)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_344),
.C(n_365),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_342),
.B(n_393),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_344),
.B(n_365),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_349),
.C(n_357),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_345),
.B(n_349),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_347),
.B(n_404),
.C(n_409),
.Y(n_427)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

BUFx2_ASAP7_75t_SL g351 ( 
.A(n_352),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_355),
.Y(n_353)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_357),
.B(n_371),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_SL g486 ( 
.A(n_358),
.B(n_487),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_360),
.Y(n_358)
);

XNOR2x1_ASAP7_75t_SL g434 ( 
.A(n_359),
.B(n_360),
.Y(n_434)
);

CKINVDCx16_ASAP7_75t_R g455 ( 
.A(n_359),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_359),
.A2(n_455),
.B1(n_456),
.B2(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

NOR2xp67_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_392),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_369),
.B(n_392),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_372),
.C(n_390),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_370),
.B(n_499),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_373),
.B(n_390),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_378),
.C(n_388),
.Y(n_373)
);

XOR2x1_ASAP7_75t_L g491 ( 
.A(n_374),
.B(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_379),
.B(n_389),
.Y(n_492)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_380),
.Y(n_430)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

XOR2x2_ASAP7_75t_L g428 ( 
.A(n_384),
.B(n_429),
.Y(n_428)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

NAND3xp33_ASAP7_75t_SL g394 ( 
.A(n_395),
.B(n_396),
.C(n_397),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_398),
.A2(n_495),
.B(n_500),
.Y(n_397)
);

AOI21x1_ASAP7_75t_L g398 ( 
.A1(n_399),
.A2(n_481),
.B(n_494),
.Y(n_398)
);

OAI21x1_ASAP7_75t_SL g399 ( 
.A1(n_400),
.A2(n_440),
.B(n_480),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_401),
.B(n_425),
.Y(n_400)
);

OR2x2_ASAP7_75t_L g480 ( 
.A(n_401),
.B(n_425),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_410),
.C(n_418),
.Y(n_401)
);

XOR2x1_ASAP7_75t_L g474 ( 
.A(n_402),
.B(n_475),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_409),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_410),
.A2(n_411),
.B1(n_418),
.B2(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_415),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_SL g445 ( 
.A(n_412),
.B(n_415),
.Y(n_445)
);

INVx3_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx4_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_418),
.Y(n_476)
);

AO22x1_ASAP7_75t_SL g418 ( 
.A1(n_419),
.A2(n_422),
.B1(n_423),
.B2(n_424),
.Y(n_418)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_419),
.Y(n_423)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g424 ( 
.A(n_422),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_422),
.B(n_423),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_424),
.B(n_465),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_431),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_428),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_427),
.B(n_428),
.C(n_431),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_433),
.Y(n_431)
);

MAJx2_ASAP7_75t_L g489 ( 
.A(n_432),
.B(n_434),
.C(n_435),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_435),
.Y(n_433)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

AOI21x1_ASAP7_75t_SL g440 ( 
.A1(n_441),
.A2(n_473),
.B(n_479),
.Y(n_440)
);

OAI21x1_ASAP7_75t_L g441 ( 
.A1(n_442),
.A2(n_457),
.B(n_472),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_454),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_443),
.B(n_454),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_444),
.A2(n_445),
.B1(n_446),
.B2(n_447),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_444),
.B(n_448),
.C(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_SL g454 ( 
.A(n_455),
.B(n_456),
.Y(n_454)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_456),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_458),
.A2(n_464),
.B(n_471),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_462),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_459),
.B(n_462),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_460),
.B(n_461),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g465 ( 
.A(n_461),
.B(n_466),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_474),
.B(n_477),
.Y(n_473)
);

NOR2xp67_ASAP7_75t_SL g479 ( 
.A(n_474),
.B(n_477),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_482),
.B(n_493),
.Y(n_481)
);

NOR2xp67_ASAP7_75t_L g494 ( 
.A(n_482),
.B(n_493),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_483),
.A2(n_484),
.B1(n_490),
.B2(n_491),
.Y(n_482)
);

INVxp33_ASAP7_75t_SL g483 ( 
.A(n_484),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_485),
.A2(n_486),
.B1(n_488),
.B2(n_489),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g497 ( 
.A(n_485),
.Y(n_497)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_489),
.B(n_490),
.C(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

NOR2xp67_ASAP7_75t_L g495 ( 
.A(n_496),
.B(n_498),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_496),
.B(n_498),
.Y(n_500)
);

NOR2xp67_ASAP7_75t_SL g501 ( 
.A(n_502),
.B(n_519),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_515),
.Y(n_502)
);

OR2x2_ASAP7_75t_L g526 ( 
.A(n_503),
.B(n_515),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_504),
.B(n_508),
.Y(n_503)
);

INVxp67_ASAP7_75t_SL g523 ( 
.A(n_504),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_506),
.C(n_507),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_509),
.A2(n_511),
.B1(n_513),
.B2(n_514),
.Y(n_508)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_509),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_511),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_511),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_513),
.B(n_523),
.C(n_524),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_516),
.B(n_517),
.C(n_518),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_L g525 ( 
.A1(n_519),
.A2(n_526),
.B(n_527),
.Y(n_525)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_520),
.B(n_522),
.Y(n_519)
);

OR2x2_ASAP7_75t_L g527 ( 
.A(n_520),
.B(n_522),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);


endmodule