module real_aes_6308_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_404;
wire n_147;
wire n_288;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_587;
wire n_546;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g103 ( .A(n_0), .Y(n_103) );
INVx1_ASAP7_75t_L g529 ( .A(n_1), .Y(n_529) );
INVx1_ASAP7_75t_L g194 ( .A(n_2), .Y(n_194) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_3), .A2(n_38), .B1(n_156), .B2(n_471), .Y(n_488) );
AOI21xp33_ASAP7_75t_L g135 ( .A1(n_4), .A2(n_136), .B(n_143), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_5), .B(n_129), .Y(n_520) );
AND2x6_ASAP7_75t_L g141 ( .A(n_6), .B(n_142), .Y(n_141) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_7), .A2(n_235), .B(n_236), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_8), .B(n_109), .Y(n_108) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_8), .B(n_39), .Y(n_445) );
INVx1_ASAP7_75t_L g153 ( .A(n_9), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_10), .B(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g134 ( .A(n_11), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_12), .B(n_166), .Y(n_466) );
INVx1_ASAP7_75t_L g241 ( .A(n_13), .Y(n_241) );
INVx1_ASAP7_75t_L g524 ( .A(n_14), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_15), .B(n_130), .Y(n_505) );
AO32x2_ASAP7_75t_L g486 ( .A1(n_16), .A2(n_129), .A3(n_163), .B1(n_487), .B2(n_491), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_17), .B(n_156), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_18), .B(n_182), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_19), .B(n_130), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g490 ( .A1(n_20), .A2(n_49), .B1(n_156), .B2(n_471), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_21), .B(n_136), .Y(n_206) );
AOI22xp33_ASAP7_75t_SL g499 ( .A1(n_22), .A2(n_74), .B1(n_156), .B2(n_166), .Y(n_499) );
NAND2xp5_ASAP7_75t_SL g482 ( .A(n_23), .B(n_156), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_24), .B(n_127), .Y(n_185) );
A2O1A1Ixp33_ASAP7_75t_L g238 ( .A1(n_25), .A2(n_239), .B(n_240), .C(n_242), .Y(n_238) );
OAI222xp33_ASAP7_75t_L g450 ( .A1(n_26), .A2(n_451), .B1(n_738), .B2(n_744), .C1(n_745), .C2(n_747), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_26), .Y(n_744) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_27), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_28), .B(n_159), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_29), .B(n_151), .Y(n_196) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_30), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g747 ( .A(n_31), .Y(n_747) );
INVx1_ASAP7_75t_L g172 ( .A(n_32), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_33), .B(n_159), .Y(n_484) );
INVx2_ASAP7_75t_L g139 ( .A(n_34), .Y(n_139) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_35), .B(n_156), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_36), .B(n_159), .Y(n_472) );
A2O1A1Ixp33_ASAP7_75t_L g207 ( .A1(n_37), .A2(n_141), .B(n_146), .C(n_208), .Y(n_207) );
INVx1_ASAP7_75t_L g109 ( .A(n_39), .Y(n_109) );
INVx1_ASAP7_75t_L g170 ( .A(n_40), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g255 ( .A(n_41), .B(n_151), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g514 ( .A(n_42), .B(n_156), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_43), .A2(n_84), .B1(n_213), .B2(n_471), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_44), .B(n_156), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_45), .B(n_156), .Y(n_525) );
CKINVDCx16_ASAP7_75t_R g173 ( .A(n_46), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_47), .B(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_48), .B(n_136), .Y(n_229) );
AOI22xp33_ASAP7_75t_SL g509 ( .A1(n_50), .A2(n_59), .B1(n_156), .B2(n_166), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g165 ( .A1(n_51), .A2(n_146), .B1(n_166), .B2(n_168), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g216 ( .A(n_52), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_53), .B(n_156), .Y(n_465) );
CKINVDCx16_ASAP7_75t_R g191 ( .A(n_54), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g542 ( .A(n_55), .B(n_156), .Y(n_542) );
A2O1A1Ixp33_ASAP7_75t_L g149 ( .A1(n_56), .A2(n_150), .B(n_152), .C(n_155), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g259 ( .A(n_57), .Y(n_259) );
INVx1_ASAP7_75t_L g144 ( .A(n_58), .Y(n_144) );
INVx1_ASAP7_75t_L g142 ( .A(n_60), .Y(n_142) );
OAI22xp5_ASAP7_75t_L g116 ( .A1(n_61), .A2(n_117), .B1(n_118), .B2(n_437), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_61), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_62), .B(n_156), .Y(n_530) );
INVx1_ASAP7_75t_L g133 ( .A(n_63), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g114 ( .A(n_64), .Y(n_114) );
AO32x2_ASAP7_75t_L g496 ( .A1(n_65), .A2(n_129), .A3(n_221), .B1(n_491), .B2(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g541 ( .A(n_66), .Y(n_541) );
INVx1_ASAP7_75t_L g479 ( .A(n_67), .Y(n_479) );
A2O1A1Ixp33_ASAP7_75t_SL g181 ( .A1(n_68), .A2(n_155), .B(n_182), .C(n_183), .Y(n_181) );
INVxp67_ASAP7_75t_L g184 ( .A(n_69), .Y(n_184) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_70), .B(n_166), .Y(n_480) );
INVx1_ASAP7_75t_L g107 ( .A(n_71), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g176 ( .A(n_72), .Y(n_176) );
INVx1_ASAP7_75t_L g252 ( .A(n_73), .Y(n_252) );
A2O1A1Ixp33_ASAP7_75t_L g253 ( .A1(n_75), .A2(n_141), .B(n_146), .C(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_76), .B(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g483 ( .A(n_77), .B(n_166), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_78), .B(n_195), .Y(n_209) );
INVx2_ASAP7_75t_L g131 ( .A(n_79), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_80), .B(n_182), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_81), .B(n_166), .Y(n_515) );
A2O1A1Ixp33_ASAP7_75t_L g192 ( .A1(n_82), .A2(n_141), .B(n_146), .C(n_193), .Y(n_192) );
INVx2_ASAP7_75t_L g104 ( .A(n_83), .Y(n_104) );
OR2x2_ASAP7_75t_L g442 ( .A(n_83), .B(n_443), .Y(n_442) );
OR2x2_ASAP7_75t_L g453 ( .A(n_83), .B(n_444), .Y(n_453) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_85), .A2(n_98), .B1(n_166), .B2(n_167), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_86), .B(n_159), .Y(n_158) );
CKINVDCx20_ASAP7_75t_R g199 ( .A(n_87), .Y(n_199) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_88), .A2(n_141), .B(n_146), .C(n_224), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g231 ( .A(n_89), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_90), .A2(n_100), .B1(n_110), .B2(n_751), .Y(n_99) );
INVx1_ASAP7_75t_L g180 ( .A(n_91), .Y(n_180) );
CKINVDCx16_ASAP7_75t_R g237 ( .A(n_92), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g225 ( .A(n_93), .B(n_195), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_94), .B(n_166), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_95), .B(n_129), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_96), .B(n_107), .Y(n_106) );
AOI21xp5_ASAP7_75t_L g178 ( .A1(n_97), .A2(n_136), .B(n_179), .Y(n_178) );
INVx1_ASAP7_75t_SL g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_L g752 ( .A(n_101), .Y(n_752) );
OR2x2_ASAP7_75t_L g101 ( .A(n_102), .B(n_108), .Y(n_101) );
NAND3xp33_ASAP7_75t_SL g102 ( .A(n_103), .B(n_104), .C(n_105), .Y(n_102) );
AND2x2_ASAP7_75t_L g444 ( .A(n_103), .B(n_445), .Y(n_444) );
OR2x2_ASAP7_75t_L g455 ( .A(n_104), .B(n_444), .Y(n_455) );
NOR2x2_ASAP7_75t_L g746 ( .A(n_104), .B(n_443), .Y(n_746) );
INVx1_ASAP7_75t_SL g105 ( .A(n_106), .Y(n_105) );
OAI21xp5_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_115), .B(n_449), .Y(n_110) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx2_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
BUFx2_ASAP7_75t_L g750 ( .A(n_113), .Y(n_750) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AOI21xp5_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_439), .B(n_446), .Y(n_115) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
AOI22xp5_ASAP7_75t_L g451 ( .A1(n_120), .A2(n_452), .B1(n_454), .B2(n_456), .Y(n_451) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
BUFx2_ASAP7_75t_L g438 ( .A(n_121), .Y(n_438) );
AND3x1_ASAP7_75t_L g121 ( .A(n_122), .B(n_359), .C(n_404), .Y(n_121) );
NOR4xp25_ASAP7_75t_L g122 ( .A(n_123), .B(n_282), .C(n_323), .D(n_340), .Y(n_122) );
A2O1A1Ixp33_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_186), .B(n_202), .C(n_244), .Y(n_123) );
OR2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_160), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_125), .B(n_187), .Y(n_186) );
NOR4xp25_ASAP7_75t_L g306 ( .A(n_125), .B(n_300), .C(n_307), .D(n_313), .Y(n_306) );
AND2x2_ASAP7_75t_L g379 ( .A(n_125), .B(n_268), .Y(n_379) );
AND2x2_ASAP7_75t_L g398 ( .A(n_125), .B(n_344), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_125), .B(n_393), .Y(n_407) );
AND2x2_ASAP7_75t_L g420 ( .A(n_125), .B(n_201), .Y(n_420) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx1_ASAP7_75t_SL g265 ( .A(n_126), .Y(n_265) );
AND2x2_ASAP7_75t_L g272 ( .A(n_126), .B(n_273), .Y(n_272) );
OR2x2_ASAP7_75t_L g322 ( .A(n_126), .B(n_161), .Y(n_322) );
AND2x2_ASAP7_75t_SL g333 ( .A(n_126), .B(n_268), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_126), .B(n_161), .Y(n_337) );
AND2x2_ASAP7_75t_L g346 ( .A(n_126), .B(n_271), .Y(n_346) );
BUFx2_ASAP7_75t_L g369 ( .A(n_126), .Y(n_369) );
AND2x2_ASAP7_75t_L g373 ( .A(n_126), .B(n_177), .Y(n_373) );
OA21x2_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_135), .B(n_158), .Y(n_126) );
INVx3_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
NOR2xp33_ASAP7_75t_SL g215 ( .A(n_128), .B(n_216), .Y(n_215) );
NAND3xp33_ASAP7_75t_L g506 ( .A(n_128), .B(n_491), .C(n_507), .Y(n_506) );
AO21x1_ASAP7_75t_L g544 ( .A1(n_128), .A2(n_507), .B(n_545), .Y(n_544) );
INVx4_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
OA21x2_ASAP7_75t_L g177 ( .A1(n_129), .A2(n_178), .B(n_185), .Y(n_177) );
OA21x2_ASAP7_75t_L g511 ( .A1(n_129), .A2(n_512), .B(n_520), .Y(n_511) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx1_ASAP7_75t_L g163 ( .A(n_130), .Y(n_163) );
AND2x2_ASAP7_75t_L g130 ( .A(n_131), .B(n_132), .Y(n_130) );
AND2x2_ASAP7_75t_SL g159 ( .A(n_131), .B(n_132), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_134), .Y(n_132) );
BUFx2_ASAP7_75t_L g235 ( .A(n_136), .Y(n_235) );
AND2x4_ASAP7_75t_L g136 ( .A(n_137), .B(n_141), .Y(n_136) );
NAND2x1p5_ASAP7_75t_L g174 ( .A(n_137), .B(n_141), .Y(n_174) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_140), .Y(n_137) );
INVx1_ASAP7_75t_L g519 ( .A(n_138), .Y(n_519) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g147 ( .A(n_139), .Y(n_147) );
INVx1_ASAP7_75t_L g167 ( .A(n_139), .Y(n_167) );
INVx1_ASAP7_75t_L g148 ( .A(n_140), .Y(n_148) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_140), .Y(n_151) );
INVx3_ASAP7_75t_L g154 ( .A(n_140), .Y(n_154) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_140), .Y(n_169) );
INVx1_ASAP7_75t_L g182 ( .A(n_140), .Y(n_182) );
INVx4_ASAP7_75t_SL g157 ( .A(n_141), .Y(n_157) );
OAI21xp5_ASAP7_75t_L g463 ( .A1(n_141), .A2(n_464), .B(n_468), .Y(n_463) );
OAI21xp5_ASAP7_75t_L g477 ( .A1(n_141), .A2(n_478), .B(n_481), .Y(n_477) );
BUFx3_ASAP7_75t_L g491 ( .A(n_141), .Y(n_491) );
OAI21xp5_ASAP7_75t_L g512 ( .A1(n_141), .A2(n_513), .B(n_516), .Y(n_512) );
OAI21xp5_ASAP7_75t_L g522 ( .A1(n_141), .A2(n_523), .B(n_527), .Y(n_522) );
O2A1O1Ixp33_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_145), .B(n_149), .C(n_157), .Y(n_143) );
O2A1O1Ixp33_ASAP7_75t_L g179 ( .A1(n_145), .A2(n_157), .B(n_180), .C(n_181), .Y(n_179) );
O2A1O1Ixp33_ASAP7_75t_L g236 ( .A1(n_145), .A2(n_157), .B(n_237), .C(n_238), .Y(n_236) );
INVx5_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
AND2x6_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_147), .Y(n_156) );
BUFx3_ASAP7_75t_L g213 ( .A(n_147), .Y(n_213) );
INVx1_ASAP7_75t_L g471 ( .A(n_147), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_150), .A2(n_469), .B(n_470), .Y(n_468) );
O2A1O1Ixp5_ASAP7_75t_L g540 ( .A1(n_150), .A2(n_528), .B(n_541), .C(n_542), .Y(n_540) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx4_ASAP7_75t_L g227 ( .A(n_151), .Y(n_227) );
OAI22xp5_ASAP7_75t_L g487 ( .A1(n_151), .A2(n_488), .B1(n_489), .B2(n_490), .Y(n_487) );
OAI22xp5_ASAP7_75t_SL g497 ( .A1(n_151), .A2(n_154), .B1(n_498), .B2(n_499), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g507 ( .A1(n_151), .A2(n_489), .B1(n_508), .B2(n_509), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_154), .B(n_184), .Y(n_183) );
INVx5_ASAP7_75t_L g195 ( .A(n_154), .Y(n_195) );
O2A1O1Ixp5_ASAP7_75t_SL g478 ( .A1(n_155), .A2(n_195), .B(n_479), .C(n_480), .Y(n_478) );
INVx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
HB1xp67_ASAP7_75t_L g228 ( .A(n_156), .Y(n_228) );
OAI22xp33_ASAP7_75t_L g164 ( .A1(n_157), .A2(n_165), .B1(n_173), .B2(n_174), .Y(n_164) );
INVx1_ASAP7_75t_L g200 ( .A(n_159), .Y(n_200) );
INVx2_ASAP7_75t_L g221 ( .A(n_159), .Y(n_221) );
OA21x2_ASAP7_75t_L g233 ( .A1(n_159), .A2(n_234), .B(n_243), .Y(n_233) );
OA21x2_ASAP7_75t_L g462 ( .A1(n_159), .A2(n_463), .B(n_472), .Y(n_462) );
OA21x2_ASAP7_75t_L g476 ( .A1(n_159), .A2(n_477), .B(n_484), .Y(n_476) );
OR2x2_ASAP7_75t_L g160 ( .A(n_161), .B(n_177), .Y(n_160) );
AND2x2_ASAP7_75t_L g201 ( .A(n_161), .B(n_177), .Y(n_201) );
BUFx2_ASAP7_75t_L g275 ( .A(n_161), .Y(n_275) );
AOI22xp33_ASAP7_75t_L g307 ( .A1(n_161), .A2(n_308), .B1(n_310), .B2(n_311), .Y(n_307) );
OR2x2_ASAP7_75t_L g329 ( .A(n_161), .B(n_189), .Y(n_329) );
AND2x2_ASAP7_75t_L g393 ( .A(n_161), .B(n_271), .Y(n_393) );
INVx3_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AND2x2_ASAP7_75t_L g261 ( .A(n_162), .B(n_189), .Y(n_261) );
AND2x2_ASAP7_75t_L g268 ( .A(n_162), .B(n_177), .Y(n_268) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_162), .Y(n_310) );
OR2x2_ASAP7_75t_L g345 ( .A(n_162), .B(n_188), .Y(n_345) );
AO21x2_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_164), .B(n_175), .Y(n_162) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_163), .B(n_176), .Y(n_175) );
AO21x2_ASAP7_75t_L g189 ( .A1(n_163), .A2(n_190), .B(n_198), .Y(n_189) );
INVx2_ASAP7_75t_L g214 ( .A(n_163), .Y(n_214) );
INVx2_ASAP7_75t_L g197 ( .A(n_166), .Y(n_197) );
INVx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
OAI22xp5_ASAP7_75t_SL g168 ( .A1(n_169), .A2(n_170), .B1(n_171), .B2(n_172), .Y(n_168) );
INVx2_ASAP7_75t_L g171 ( .A(n_169), .Y(n_171) );
INVx4_ASAP7_75t_L g239 ( .A(n_169), .Y(n_239) );
OAI21xp5_ASAP7_75t_L g190 ( .A1(n_174), .A2(n_191), .B(n_192), .Y(n_190) );
OAI21xp5_ASAP7_75t_L g251 ( .A1(n_174), .A2(n_252), .B(n_253), .Y(n_251) );
INVx1_ASAP7_75t_L g264 ( .A(n_177), .Y(n_264) );
INVx3_ASAP7_75t_L g273 ( .A(n_177), .Y(n_273) );
BUFx2_ASAP7_75t_L g297 ( .A(n_177), .Y(n_297) );
AND2x2_ASAP7_75t_L g330 ( .A(n_177), .B(n_265), .Y(n_330) );
INVx1_ASAP7_75t_L g467 ( .A(n_182), .Y(n_467) );
OAI22xp5_ASAP7_75t_L g415 ( .A1(n_186), .A2(n_416), .B1(n_417), .B2(n_418), .Y(n_415) );
AND2x2_ASAP7_75t_L g187 ( .A(n_188), .B(n_201), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_188), .B(n_273), .Y(n_277) );
INVx1_ASAP7_75t_L g305 ( .A(n_188), .Y(n_305) );
INVx3_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx3_ASAP7_75t_L g271 ( .A(n_189), .Y(n_271) );
O2A1O1Ixp33_ASAP7_75t_L g193 ( .A1(n_194), .A2(n_195), .B(n_196), .C(n_197), .Y(n_193) );
INVx2_ASAP7_75t_L g489 ( .A(n_195), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_195), .A2(n_514), .B(n_515), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_195), .A2(n_538), .B(n_539), .Y(n_537) );
O2A1O1Ixp33_ASAP7_75t_L g523 ( .A1(n_197), .A2(n_524), .B(n_525), .C(n_526), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_199), .B(n_200), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_200), .B(n_231), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_200), .B(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g283 ( .A(n_201), .Y(n_283) );
NAND2x1_ASAP7_75t_SL g202 ( .A(n_203), .B(n_217), .Y(n_202) );
AND2x2_ASAP7_75t_L g281 ( .A(n_203), .B(n_232), .Y(n_281) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_203), .Y(n_355) );
AND2x2_ASAP7_75t_L g382 ( .A(n_203), .B(n_302), .Y(n_382) );
AND2x2_ASAP7_75t_L g390 ( .A(n_203), .B(n_352), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_203), .B(n_247), .Y(n_417) );
INVx3_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g248 ( .A(n_204), .B(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g266 ( .A(n_204), .B(n_267), .Y(n_266) );
INVx2_ASAP7_75t_L g287 ( .A(n_204), .Y(n_287) );
INVx1_ASAP7_75t_L g293 ( .A(n_204), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g308 ( .A(n_204), .B(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g326 ( .A(n_204), .B(n_250), .Y(n_326) );
OR2x2_ASAP7_75t_L g364 ( .A(n_204), .B(n_319), .Y(n_364) );
AOI32xp33_ASAP7_75t_L g376 ( .A1(n_204), .A2(n_377), .A3(n_380), .B1(n_381), .B2(n_382), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_204), .B(n_352), .Y(n_416) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_204), .B(n_312), .Y(n_427) );
OR2x6_ASAP7_75t_L g204 ( .A(n_205), .B(n_215), .Y(n_204) );
AOI21xp5_ASAP7_75t_SL g205 ( .A1(n_206), .A2(n_207), .B(n_214), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_209), .A2(n_210), .B(n_211), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g254 ( .A1(n_211), .A2(n_255), .B(n_256), .Y(n_254) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g242 ( .A(n_213), .Y(n_242) );
INVx1_ASAP7_75t_L g257 ( .A(n_214), .Y(n_257) );
OA21x2_ASAP7_75t_L g521 ( .A1(n_214), .A2(n_522), .B(n_531), .Y(n_521) );
OA21x2_ASAP7_75t_L g535 ( .A1(n_214), .A2(n_536), .B(n_543), .Y(n_535) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
OR2x2_ASAP7_75t_L g338 ( .A(n_218), .B(n_339), .Y(n_338) );
OR2x2_ASAP7_75t_L g218 ( .A(n_219), .B(n_232), .Y(n_218) );
INVx1_ASAP7_75t_L g300 ( .A(n_219), .Y(n_300) );
AND2x2_ASAP7_75t_L g302 ( .A(n_219), .B(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_219), .B(n_249), .Y(n_319) );
AND2x2_ASAP7_75t_L g352 ( .A(n_219), .B(n_328), .Y(n_352) );
AND2x2_ASAP7_75t_L g389 ( .A(n_219), .B(n_250), .Y(n_389) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g247 ( .A(n_220), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_220), .B(n_249), .Y(n_279) );
AND2x2_ASAP7_75t_L g286 ( .A(n_220), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g327 ( .A(n_220), .B(n_328), .Y(n_327) );
AO21x2_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_222), .B(n_230), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_223), .B(n_229), .Y(n_222) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_226), .B(n_228), .Y(n_224) );
INVx2_ASAP7_75t_L g303 ( .A(n_232), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_232), .B(n_249), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_232), .B(n_294), .Y(n_375) );
INVx1_ASAP7_75t_L g397 ( .A(n_232), .Y(n_397) );
INVx1_ASAP7_75t_L g414 ( .A(n_232), .Y(n_414) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
AND2x2_ASAP7_75t_L g267 ( .A(n_233), .B(n_249), .Y(n_267) );
AND2x2_ASAP7_75t_L g289 ( .A(n_233), .B(n_250), .Y(n_289) );
INVx1_ASAP7_75t_L g328 ( .A(n_233), .Y(n_328) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_239), .B(n_241), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_239), .A2(n_482), .B(n_483), .Y(n_481) );
INVx1_ASAP7_75t_L g526 ( .A(n_239), .Y(n_526) );
AOI221x1_ASAP7_75t_SL g244 ( .A1(n_245), .A2(n_260), .B1(n_266), .B2(n_268), .C(n_269), .Y(n_244) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_245), .A2(n_333), .B1(n_400), .B2(n_401), .Y(n_399) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_248), .Y(n_245) );
AND2x2_ASAP7_75t_L g291 ( .A(n_246), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g386 ( .A(n_246), .B(n_266), .Y(n_386) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g342 ( .A(n_247), .B(n_267), .Y(n_342) );
INVx1_ASAP7_75t_L g354 ( .A(n_248), .Y(n_354) );
AND2x2_ASAP7_75t_L g365 ( .A(n_248), .B(n_352), .Y(n_365) );
AND2x2_ASAP7_75t_L g432 ( .A(n_248), .B(n_327), .Y(n_432) );
INVx2_ASAP7_75t_L g294 ( .A(n_249), .Y(n_294) );
INVx2_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
AO21x2_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_257), .B(n_258), .Y(n_250) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_261), .B(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g384 ( .A(n_261), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_262), .B(n_345), .Y(n_348) );
INVx3_ASAP7_75t_SL g262 ( .A(n_263), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g428 ( .A1(n_263), .A2(n_384), .B(n_429), .Y(n_428) );
AND2x4_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
NOR2xp33_ASAP7_75t_SL g406 ( .A(n_266), .B(n_292), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_267), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g358 ( .A(n_267), .B(n_286), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_267), .B(n_293), .Y(n_435) );
AND2x2_ASAP7_75t_L g304 ( .A(n_268), .B(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g371 ( .A(n_268), .Y(n_371) );
AOI21xp33_ASAP7_75t_L g269 ( .A1(n_270), .A2(n_274), .B(n_278), .Y(n_269) );
NAND2x1_ASAP7_75t_L g270 ( .A(n_271), .B(n_272), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_271), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g320 ( .A(n_271), .B(n_321), .Y(n_320) );
INVx1_ASAP7_75t_SL g332 ( .A(n_271), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g377 ( .A(n_271), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g356 ( .A(n_272), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_272), .B(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_272), .B(n_275), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
AOI211xp5_ASAP7_75t_L g343 ( .A1(n_275), .A2(n_314), .B(n_344), .C(n_346), .Y(n_343) );
AOI221xp5_ASAP7_75t_L g361 ( .A1(n_275), .A2(n_362), .B1(n_365), .B2(n_366), .C(n_370), .Y(n_361) );
AND2x2_ASAP7_75t_L g357 ( .A(n_276), .B(n_310), .Y(n_357) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g317 ( .A(n_281), .B(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g388 ( .A(n_281), .B(n_389), .Y(n_388) );
OAI211xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_284), .B(n_290), .C(n_315), .Y(n_282) );
NAND3xp33_ASAP7_75t_SL g401 ( .A(n_283), .B(n_402), .C(n_403), .Y(n_401) );
OR2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_288), .Y(n_284) );
OR2x2_ASAP7_75t_L g374 ( .A(n_285), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AOI221xp5_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_295), .B1(n_298), .B2(n_304), .C(n_306), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_292), .B(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_292), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g314 ( .A(n_297), .Y(n_314) );
OAI22xp5_ASAP7_75t_L g353 ( .A1(n_297), .A2(n_354), .B1(n_355), .B2(n_356), .Y(n_353) );
OR2x2_ASAP7_75t_L g434 ( .A(n_297), .B(n_345), .Y(n_434) );
NAND2xp5_ASAP7_75t_SL g298 ( .A(n_299), .B(n_301), .Y(n_298) );
INVxp67_ASAP7_75t_L g408 ( .A(n_300), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_302), .B(n_423), .Y(n_422) );
INVxp67_ASAP7_75t_L g309 ( .A(n_303), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_305), .B(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_305), .B(n_352), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_305), .B(n_372), .Y(n_411) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_309), .Y(n_335) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
OR2x2_ASAP7_75t_L g425 ( .A(n_314), .B(n_345), .Y(n_425) );
INVx1_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_320), .Y(n_316) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx1_ASAP7_75t_SL g403 ( .A(n_320), .Y(n_403) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
OAI322xp33_ASAP7_75t_SL g323 ( .A1(n_324), .A2(n_329), .A3(n_330), .B1(n_331), .B2(n_334), .C1(n_336), .C2(n_338), .Y(n_323) );
OAI322xp33_ASAP7_75t_L g405 ( .A1(n_324), .A2(n_406), .A3(n_407), .B1(n_408), .B2(n_409), .C1(n_410), .C2(n_412), .Y(n_405) );
CKINVDCx16_ASAP7_75t_R g324 ( .A(n_325), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
INVx4_ASAP7_75t_L g339 ( .A(n_326), .Y(n_339) );
AND2x2_ASAP7_75t_L g400 ( .A(n_326), .B(n_352), .Y(n_400) );
AND2x2_ASAP7_75t_L g413 ( .A(n_326), .B(n_414), .Y(n_413) );
CKINVDCx16_ASAP7_75t_R g424 ( .A(n_329), .Y(n_424) );
INVx1_ASAP7_75t_L g402 ( .A(n_330), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
OR2x2_ASAP7_75t_L g336 ( .A(n_332), .B(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g419 ( .A(n_332), .B(n_420), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_332), .B(n_373), .Y(n_430) );
OR2x2_ASAP7_75t_L g363 ( .A(n_335), .B(n_364), .Y(n_363) );
INVxp33_ASAP7_75t_L g380 ( .A(n_335), .Y(n_380) );
OAI221xp5_ASAP7_75t_SL g340 ( .A1(n_339), .A2(n_341), .B1(n_343), .B2(n_347), .C(n_349), .Y(n_340) );
NOR2xp67_ASAP7_75t_L g396 ( .A(n_339), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g423 ( .A(n_339), .Y(n_423) );
INVx1_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
INVx3_ASAP7_75t_SL g344 ( .A(n_345), .Y(n_344) );
AOI322xp5_ASAP7_75t_L g387 ( .A1(n_346), .A2(n_371), .A3(n_388), .B1(n_390), .B2(n_391), .C1(n_394), .C2(n_398), .Y(n_387) );
INVxp67_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AOI22xp5_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_353), .B1(n_357), .B2(n_358), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_360), .B(n_383), .Y(n_359) );
NAND2xp5_ASAP7_75t_SL g360 ( .A(n_361), .B(n_376), .Y(n_360) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_SL g394 ( .A(n_364), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
NAND2xp33_ASAP7_75t_SL g381 ( .A(n_367), .B(n_378), .Y(n_381) );
INVx1_ASAP7_75t_SL g368 ( .A(n_369), .Y(n_368) );
OAI322xp33_ASAP7_75t_L g421 ( .A1(n_369), .A2(n_422), .A3(n_424), .B1(n_425), .B2(n_426), .C1(n_428), .C2(n_431), .Y(n_421) );
AOI21xp33_ASAP7_75t_SL g370 ( .A1(n_371), .A2(n_372), .B(n_374), .Y(n_370) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_379), .B(n_427), .Y(n_436) );
OAI211xp5_ASAP7_75t_SL g383 ( .A1(n_384), .A2(n_385), .B(n_387), .C(n_399), .Y(n_383) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
NOR4xp25_ASAP7_75t_L g404 ( .A(n_405), .B(n_415), .C(n_421), .D(n_433), .Y(n_404) );
INVxp67_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_SL g418 ( .A(n_419), .Y(n_418) );
INVxp67_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
CKINVDCx14_ASAP7_75t_R g431 ( .A(n_432), .Y(n_431) );
OAI21xp5_ASAP7_75t_SL g433 ( .A1(n_434), .A2(n_435), .B(n_436), .Y(n_433) );
BUFx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g738 ( .A1(n_438), .A2(n_739), .B1(n_742), .B2(n_743), .Y(n_738) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
CKINVDCx20_ASAP7_75t_R g440 ( .A(n_441), .Y(n_440) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
BUFx2_ASAP7_75t_L g447 ( .A(n_442), .Y(n_447) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
OAI21xp5_ASAP7_75t_SL g449 ( .A1(n_446), .A2(n_450), .B(n_748), .Y(n_449) );
NOR2xp33_ASAP7_75t_SL g446 ( .A(n_447), .B(n_448), .Y(n_446) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g741 ( .A(n_453), .Y(n_741) );
INVx6_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g742 ( .A(n_455), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_456), .Y(n_743) );
OR2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_660), .Y(n_456) );
NAND5xp2_ASAP7_75t_L g457 ( .A(n_458), .B(n_579), .C(n_594), .D(n_620), .E(n_642), .Y(n_457) );
NOR2xp33_ASAP7_75t_SL g458 ( .A(n_459), .B(n_559), .Y(n_458) );
OAI221xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_500), .B1(n_532), .B2(n_548), .C(n_549), .Y(n_459) );
NOR2xp33_ASAP7_75t_SL g460 ( .A(n_461), .B(n_492), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_461), .B(n_609), .Y(n_608) );
INVx1_ASAP7_75t_SL g736 ( .A(n_461), .Y(n_736) );
AND2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_473), .Y(n_461) );
INVx1_ASAP7_75t_L g576 ( .A(n_462), .Y(n_576) );
AND2x2_ASAP7_75t_L g578 ( .A(n_462), .B(n_486), .Y(n_578) );
AND2x2_ASAP7_75t_L g588 ( .A(n_462), .B(n_485), .Y(n_588) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_462), .Y(n_606) );
INVx1_ASAP7_75t_L g616 ( .A(n_462), .Y(n_616) );
OR2x2_ASAP7_75t_L g654 ( .A(n_462), .B(n_553), .Y(n_654) );
INVx2_ASAP7_75t_L g704 ( .A(n_462), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_462), .B(n_552), .Y(n_721) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_466), .B(n_467), .Y(n_464) );
NOR2xp67_ASAP7_75t_L g473 ( .A(n_474), .B(n_485), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
HB1xp67_ASAP7_75t_L g570 ( .A(n_475), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_475), .B(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_SL g636 ( .A(n_475), .B(n_576), .Y(n_636) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
HB1xp67_ASAP7_75t_L g494 ( .A(n_476), .Y(n_494) );
INVx2_ASAP7_75t_L g553 ( .A(n_476), .Y(n_553) );
OR2x2_ASAP7_75t_L g615 ( .A(n_476), .B(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g554 ( .A(n_485), .B(n_496), .Y(n_554) );
AND2x2_ASAP7_75t_L g571 ( .A(n_485), .B(n_551), .Y(n_571) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g495 ( .A(n_486), .B(n_496), .Y(n_495) );
BUFx2_ASAP7_75t_L g574 ( .A(n_486), .Y(n_574) );
AND2x2_ASAP7_75t_L g703 ( .A(n_486), .B(n_704), .Y(n_703) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_489), .A2(n_517), .B(n_518), .Y(n_516) );
O2A1O1Ixp33_ASAP7_75t_L g527 ( .A1(n_489), .A2(n_528), .B(n_529), .C(n_530), .Y(n_527) );
OAI21xp5_ASAP7_75t_L g536 ( .A1(n_491), .A2(n_537), .B(n_540), .Y(n_536) );
INVx1_ASAP7_75t_L g548 ( .A(n_492), .Y(n_548) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_495), .Y(n_492) );
AND2x2_ASAP7_75t_L g666 ( .A(n_493), .B(n_554), .Y(n_666) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g667 ( .A(n_494), .B(n_578), .Y(n_667) );
O2A1O1Ixp33_ASAP7_75t_L g634 ( .A1(n_495), .A2(n_635), .B(n_637), .C(n_639), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_495), .B(n_635), .Y(n_644) );
AOI221xp5_ASAP7_75t_L g707 ( .A1(n_495), .A2(n_565), .B1(n_708), .B2(n_709), .C(n_711), .Y(n_707) );
INVx1_ASAP7_75t_L g551 ( .A(n_496), .Y(n_551) );
INVx1_ASAP7_75t_L g587 ( .A(n_496), .Y(n_587) );
BUFx6f_ASAP7_75t_L g596 ( .A(n_496), .Y(n_596) );
INVx1_ASAP7_75t_SL g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_502), .B(n_510), .Y(n_501) );
AND2x2_ASAP7_75t_L g613 ( .A(n_502), .B(n_558), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_502), .B(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_503), .B(n_582), .Y(n_581) );
OR2x2_ASAP7_75t_L g705 ( .A(n_503), .B(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g737 ( .A(n_503), .Y(n_737) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx3_ASAP7_75t_L g567 ( .A(n_504), .Y(n_567) );
AND2x2_ASAP7_75t_L g593 ( .A(n_504), .B(n_547), .Y(n_593) );
NOR2x1_ASAP7_75t_L g602 ( .A(n_504), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g609 ( .A(n_504), .B(n_610), .Y(n_609) );
AND2x4_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
INVx1_ASAP7_75t_L g545 ( .A(n_505), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_510), .B(n_649), .Y(n_684) );
INVx1_ASAP7_75t_SL g688 ( .A(n_510), .Y(n_688) );
AND2x2_ASAP7_75t_L g510 ( .A(n_511), .B(n_521), .Y(n_510) );
INVx3_ASAP7_75t_L g547 ( .A(n_511), .Y(n_547) );
AND2x2_ASAP7_75t_L g558 ( .A(n_511), .B(n_535), .Y(n_558) );
AND2x2_ASAP7_75t_L g580 ( .A(n_511), .B(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g625 ( .A(n_511), .B(n_619), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_511), .B(n_557), .Y(n_706) );
INVx2_ASAP7_75t_L g528 ( .A(n_519), .Y(n_528) );
AND2x2_ASAP7_75t_L g546 ( .A(n_521), .B(n_547), .Y(n_546) );
INVx2_ASAP7_75t_L g557 ( .A(n_521), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_521), .B(n_535), .Y(n_582) );
AND2x2_ASAP7_75t_L g618 ( .A(n_521), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_546), .Y(n_533) );
INVx1_ASAP7_75t_L g598 ( .A(n_534), .Y(n_598) );
AND2x2_ASAP7_75t_L g640 ( .A(n_534), .B(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_SL g646 ( .A(n_534), .B(n_561), .Y(n_646) );
AOI21xp5_ASAP7_75t_SL g720 ( .A1(n_534), .A2(n_552), .B(n_575), .Y(n_720) );
AND2x2_ASAP7_75t_L g534 ( .A(n_535), .B(n_544), .Y(n_534) );
OR2x2_ASAP7_75t_L g563 ( .A(n_535), .B(n_544), .Y(n_563) );
AND2x2_ASAP7_75t_L g610 ( .A(n_535), .B(n_547), .Y(n_610) );
INVx2_ASAP7_75t_L g619 ( .A(n_535), .Y(n_619) );
INVx1_ASAP7_75t_L g725 ( .A(n_535), .Y(n_725) );
AND2x2_ASAP7_75t_L g649 ( .A(n_544), .B(n_619), .Y(n_649) );
INVx1_ASAP7_75t_L g674 ( .A(n_544), .Y(n_674) );
AND2x2_ASAP7_75t_L g583 ( .A(n_546), .B(n_567), .Y(n_583) );
AND2x2_ASAP7_75t_L g595 ( .A(n_546), .B(n_596), .Y(n_595) );
INVx2_ASAP7_75t_SL g713 ( .A(n_546), .Y(n_713) );
INVx2_ASAP7_75t_L g603 ( .A(n_547), .Y(n_603) );
AND2x2_ASAP7_75t_L g641 ( .A(n_547), .B(n_557), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_547), .B(n_725), .Y(n_724) );
OAI21xp33_ASAP7_75t_L g549 ( .A1(n_550), .A2(n_554), .B(n_555), .Y(n_549) );
AND2x2_ASAP7_75t_L g656 ( .A(n_550), .B(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g710 ( .A(n_550), .Y(n_710) );
AND2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
INVx1_ASAP7_75t_L g630 ( .A(n_551), .Y(n_630) );
BUFx2_ASAP7_75t_L g729 ( .A(n_551), .Y(n_729) );
BUFx2_ASAP7_75t_L g600 ( .A(n_552), .Y(n_600) );
AND2x2_ASAP7_75t_L g702 ( .A(n_552), .B(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx1_ASAP7_75t_L g685 ( .A(n_553), .Y(n_685) );
AND2x4_ASAP7_75t_L g612 ( .A(n_554), .B(n_575), .Y(n_612) );
NAND2xp5_ASAP7_75t_SL g648 ( .A(n_554), .B(n_636), .Y(n_648) );
AOI32xp33_ASAP7_75t_L g572 ( .A1(n_555), .A2(n_573), .A3(n_575), .B1(n_577), .B2(n_578), .Y(n_572) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_558), .Y(n_555) );
INVx3_ASAP7_75t_L g561 ( .A(n_556), .Y(n_561) );
OR2x2_ASAP7_75t_L g697 ( .A(n_556), .B(n_653), .Y(n_697) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g566 ( .A(n_557), .B(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g673 ( .A(n_557), .B(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g565 ( .A(n_558), .B(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g577 ( .A(n_558), .B(n_567), .Y(n_577) );
INVx1_ASAP7_75t_L g698 ( .A(n_558), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_558), .B(n_673), .Y(n_731) );
A2O1A1Ixp33_ASAP7_75t_L g559 ( .A1(n_560), .A2(n_564), .B(n_568), .C(n_572), .Y(n_559) );
OAI322xp33_ASAP7_75t_L g668 ( .A1(n_560), .A2(n_605), .A3(n_669), .B1(n_671), .B2(n_675), .C1(n_676), .C2(n_680), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
INVxp67_ASAP7_75t_L g633 ( .A(n_561), .Y(n_633) );
INVx1_ASAP7_75t_SL g562 ( .A(n_563), .Y(n_562) );
OR2x2_ASAP7_75t_L g687 ( .A(n_563), .B(n_688), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g734 ( .A(n_563), .B(n_603), .Y(n_734) );
INVxp67_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g626 ( .A(n_566), .Y(n_626) );
OR2x2_ASAP7_75t_L g712 ( .A(n_567), .B(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_570), .B(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g621 ( .A(n_571), .B(n_600), .Y(n_621) );
AND2x2_ASAP7_75t_L g692 ( .A(n_571), .B(n_605), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_571), .B(n_679), .Y(n_714) );
AOI221xp5_ASAP7_75t_L g579 ( .A1(n_573), .A2(n_580), .B1(n_583), .B2(n_584), .C(n_589), .Y(n_579) );
OR2x2_ASAP7_75t_L g590 ( .A(n_573), .B(n_586), .Y(n_590) );
AND2x2_ASAP7_75t_L g678 ( .A(n_573), .B(n_679), .Y(n_678) );
AOI32xp33_ASAP7_75t_L g717 ( .A1(n_573), .A2(n_603), .A3(n_718), .B1(n_719), .B2(n_722), .Y(n_717) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NAND3xp33_ASAP7_75t_L g651 ( .A(n_574), .B(n_610), .C(n_633), .Y(n_651) );
AND2x2_ASAP7_75t_L g677 ( .A(n_574), .B(n_670), .Y(n_677) );
INVxp67_ASAP7_75t_L g657 ( .A(n_575), .Y(n_657) );
BUFx3_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_SL g686 ( .A(n_578), .B(n_630), .Y(n_686) );
INVx2_ASAP7_75t_L g696 ( .A(n_578), .Y(n_696) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_578), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g665 ( .A(n_581), .Y(n_665) );
OR2x2_ASAP7_75t_L g591 ( .A(n_582), .B(n_592), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g701 ( .A(n_584), .B(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_588), .Y(n_584) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_587), .Y(n_670) );
AND2x2_ASAP7_75t_L g629 ( .A(n_588), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g675 ( .A(n_588), .Y(n_675) );
HB1xp67_ASAP7_75t_L g700 ( .A(n_588), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
AOI21xp33_ASAP7_75t_SL g614 ( .A1(n_590), .A2(n_615), .B(n_617), .Y(n_614) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AND2x2_ASAP7_75t_L g708 ( .A(n_593), .B(n_618), .Y(n_708) );
AOI211xp5_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_597), .B(n_607), .C(n_614), .Y(n_594) );
AND2x2_ASAP7_75t_L g638 ( .A(n_596), .B(n_606), .Y(n_638) );
INVx2_ASAP7_75t_L g653 ( .A(n_596), .Y(n_653) );
OR2x2_ASAP7_75t_L g691 ( .A(n_596), .B(n_654), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_596), .B(n_734), .Y(n_733) );
AOI211xp5_ASAP7_75t_SL g597 ( .A1(n_598), .A2(n_599), .B(n_601), .C(n_604), .Y(n_597) );
INVxp67_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_600), .B(n_638), .Y(n_637) );
OAI211xp5_ASAP7_75t_L g719 ( .A1(n_601), .A2(n_696), .B(n_720), .C(n_721), .Y(n_719) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND2x1p5_ASAP7_75t_L g617 ( .A(n_602), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g659 ( .A(n_603), .B(n_649), .Y(n_659) );
INVx1_ASAP7_75t_L g664 ( .A(n_603), .Y(n_664) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_SL g607 ( .A(n_608), .B(n_611), .Y(n_607) );
INVxp33_ASAP7_75t_L g715 ( .A(n_609), .Y(n_715) );
AND2x2_ASAP7_75t_L g694 ( .A(n_610), .B(n_673), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
AOI21xp5_ASAP7_75t_L g676 ( .A1(n_615), .A2(n_677), .B(n_678), .Y(n_676) );
OAI322xp33_ASAP7_75t_L g695 ( .A1(n_617), .A2(n_696), .A3(n_697), .B1(n_698), .B2(n_699), .C1(n_701), .C2(n_705), .Y(n_695) );
AOI221xp5_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_622), .B1(n_627), .B2(n_631), .C(n_634), .Y(n_620) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OR2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_626), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g672 ( .A(n_625), .B(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g716 ( .A(n_629), .Y(n_716) );
INVxp67_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_632), .B(n_652), .Y(n_718) );
INVx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx1_ASAP7_75t_SL g639 ( .A(n_640), .Y(n_639) );
AND2x2_ASAP7_75t_L g681 ( .A(n_641), .B(n_649), .Y(n_681) );
AOI221xp5_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_645), .B1(n_647), .B2(n_649), .C(n_650), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AOI221xp5_ASAP7_75t_L g661 ( .A1(n_645), .A2(n_662), .B1(n_666), .B2(n_667), .C(n_668), .Y(n_661) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVxp67_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_649), .B(n_664), .Y(n_663) );
OAI22xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_652), .B1(n_655), .B2(n_658), .Y(n_650) );
OR2x2_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
INVx2_ASAP7_75t_SL g679 ( .A(n_654), .Y(n_679) );
INVxp67_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NAND5xp2_ASAP7_75t_L g660 ( .A(n_661), .B(n_682), .C(n_707), .D(n_717), .E(n_727), .Y(n_660) );
NAND2xp5_ASAP7_75t_SL g662 ( .A(n_663), .B(n_665), .Y(n_662) );
NOR4xp25_ASAP7_75t_L g735 ( .A(n_664), .B(n_670), .C(n_736), .D(n_737), .Y(n_735) );
AOI221xp5_ASAP7_75t_L g727 ( .A1(n_667), .A2(n_728), .B1(n_730), .B2(n_732), .C(n_735), .Y(n_727) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g726 ( .A(n_673), .Y(n_726) );
OAI322xp33_ASAP7_75t_L g683 ( .A1(n_677), .A2(n_684), .A3(n_685), .B1(n_686), .B2(n_687), .C1(n_689), .C2(n_693), .Y(n_683) );
INVx1_ASAP7_75t_SL g680 ( .A(n_681), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_683), .B(n_695), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_690), .B(n_692), .Y(n_689) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g728 ( .A(n_703), .B(n_729), .Y(n_728) );
OAI22xp33_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_714), .B1(n_715), .B2(n_716), .Y(n_711) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
OR2x2_ASAP7_75t_L g723 ( .A(n_724), .B(n_726), .Y(n_723) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVxp67_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_SL g739 ( .A(n_740), .Y(n_739) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx3_ASAP7_75t_SL g745 ( .A(n_746), .Y(n_745) );
INVxp67_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_SL g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
endmodule