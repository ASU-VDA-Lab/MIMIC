module fake_jpeg_30228_n_198 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_198);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_198;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

BUFx8_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

INVx4_ASAP7_75t_SL g35 ( 
.A(n_22),
.Y(n_35)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_21),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_41),
.B(n_43),
.Y(n_72)
);

AOI21xp33_ASAP7_75t_L g42 ( 
.A1(n_21),
.A2(n_16),
.B(n_28),
.Y(n_42)
);

NAND2x1_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_24),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_19),
.B(n_15),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_19),
.B(n_11),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_48),
.Y(n_58)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_17),
.B(n_10),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_17),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_32),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_42),
.A2(n_31),
.B1(n_23),
.B2(n_20),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_54),
.A2(n_67),
.B1(n_26),
.B2(n_2),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_46),
.A2(n_20),
.B1(n_23),
.B2(n_21),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_56),
.A2(n_60),
.B1(n_66),
.B2(n_74),
.Y(n_86)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_46),
.A2(n_18),
.B1(n_28),
.B2(n_16),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_62),
.A2(n_54),
.B(n_58),
.C(n_73),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_76),
.Y(n_78)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_47),
.A2(n_40),
.B1(n_37),
.B2(n_18),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_37),
.A2(n_33),
.B1(n_32),
.B2(n_27),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_69),
.Y(n_97)
);

AOI21xp33_ASAP7_75t_L g71 ( 
.A1(n_35),
.A2(n_25),
.B(n_27),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_71),
.B(n_73),
.Y(n_93)
);

NOR2x1_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_25),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_34),
.A2(n_33),
.B1(n_36),
.B2(n_35),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_38),
.B(n_24),
.Y(n_76)
);

AO22x1_ASAP7_75t_SL g77 ( 
.A1(n_62),
.A2(n_34),
.B1(n_24),
.B2(n_33),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_77),
.B(n_81),
.Y(n_117)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_61),
.Y(n_80)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_26),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_82),
.B(n_9),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_34),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_87),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_26),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_89),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_1),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_26),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_92),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_75),
.B(n_9),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_103),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_1),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_52),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_75),
.B(n_2),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_100),
.Y(n_112)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

AOI21xp33_ASAP7_75t_L g98 ( 
.A1(n_61),
.A2(n_3),
.B(n_4),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_98),
.B(n_50),
.Y(n_113)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_70),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_57),
.B(n_3),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_101),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_55),
.B(n_5),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_6),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_53),
.B(n_9),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_82),
.B(n_5),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_104),
.B(n_114),
.Y(n_135)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_106),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_90),
.A2(n_70),
.B1(n_50),
.B2(n_55),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_113),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_93),
.B(n_78),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_115),
.B(n_116),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_7),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_120),
.B(n_121),
.Y(n_141)
);

INVxp67_ASAP7_75t_SL g121 ( 
.A(n_80),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_123),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_92),
.A2(n_7),
.B1(n_8),
.B2(n_98),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_124),
.A2(n_92),
.B(n_87),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_116),
.B(n_91),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_126),
.B(n_131),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_83),
.C(n_97),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_111),
.C(n_109),
.Y(n_150)
);

NOR2xp67_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_77),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_123),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_105),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_103),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_133),
.B(n_140),
.Y(n_154)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

NAND2x1_ASAP7_75t_SL g137 ( 
.A(n_125),
.B(n_77),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_137),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_138),
.A2(n_124),
.B(n_88),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_111),
.A2(n_117),
.B1(n_118),
.B2(n_110),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_139),
.A2(n_144),
.B1(n_86),
.B2(n_130),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_81),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_81),
.Y(n_142)
);

A2O1A1O1Ixp25_ASAP7_75t_L g151 ( 
.A1(n_142),
.A2(n_133),
.B(n_140),
.C(n_122),
.D(n_136),
.Y(n_151)
);

OAI21xp33_ASAP7_75t_L g143 ( 
.A1(n_117),
.A2(n_97),
.B(n_79),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_143),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_111),
.A2(n_86),
.B1(n_79),
.B2(n_88),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_146),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_141),
.B(n_112),
.Y(n_146)
);

BUFx12_ASAP7_75t_L g147 ( 
.A(n_128),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_151),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_148),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_150),
.B(n_136),
.C(n_126),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_125),
.Y(n_152)
);

BUFx24_ASAP7_75t_SL g162 ( 
.A(n_152),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_105),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_128),
.C(n_101),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_129),
.A2(n_118),
.B1(n_106),
.B2(n_108),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_156),
.A2(n_139),
.B1(n_144),
.B2(n_132),
.Y(n_163)
);

AO21x1_ASAP7_75t_L g161 ( 
.A1(n_157),
.A2(n_129),
.B(n_142),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_160),
.B(n_166),
.C(n_155),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_161),
.A2(n_157),
.B(n_158),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_168),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_159),
.Y(n_164)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_164),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_129),
.C(n_131),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_156),
.A2(n_137),
.B1(n_138),
.B2(n_134),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_145),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_171),
.A2(n_172),
.B(n_176),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_169),
.A2(n_158),
.B(n_149),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_162),
.B(n_149),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_173),
.B(n_178),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_174),
.B(n_179),
.C(n_166),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_161),
.A2(n_137),
.B(n_155),
.Y(n_176)
);

OA21x2_ASAP7_75t_SL g178 ( 
.A1(n_165),
.A2(n_151),
.B(n_154),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_180),
.B(n_108),
.C(n_85),
.Y(n_190)
);

XOR2x2_ASAP7_75t_L g181 ( 
.A(n_174),
.B(n_167),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_181),
.A2(n_183),
.B1(n_147),
.B2(n_127),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_177),
.B(n_160),
.C(n_154),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_127),
.Y(n_189)
);

XOR2x1_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_147),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_185),
.A2(n_175),
.B1(n_148),
.B2(n_159),
.Y(n_187)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_184),
.B(n_147),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_186),
.B(n_187),
.Y(n_191)
);

NOR2xp67_ASAP7_75t_SL g193 ( 
.A(n_188),
.B(n_190),
.Y(n_193)
);

OAI21x1_ASAP7_75t_L g192 ( 
.A1(n_189),
.A2(n_183),
.B(n_8),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_192),
.B(n_186),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_191),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_194),
.B(n_195),
.C(n_190),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_196),
.A2(n_193),
.B1(n_80),
.B2(n_85),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_7),
.Y(n_198)
);


endmodule