module fake_aes_9921_n_31 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_0, n_31);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_0;
output n_31;
wire n_20;
wire n_23;
wire n_8;
wire n_28;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx2_ASAP7_75t_L g8 ( .A(n_6), .Y(n_8) );
HB1xp67_ASAP7_75t_L g9 ( .A(n_5), .Y(n_9) );
CKINVDCx5p33_ASAP7_75t_R g10 ( .A(n_3), .Y(n_10) );
INVx2_ASAP7_75t_L g11 ( .A(n_4), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_1), .Y(n_12) );
HB1xp67_ASAP7_75t_L g13 ( .A(n_7), .Y(n_13) );
AND2x4_ASAP7_75t_L g14 ( .A(n_9), .B(n_0), .Y(n_14) );
NAND2xp5_ASAP7_75t_L g15 ( .A(n_13), .B(n_0), .Y(n_15) );
AND2x4_ASAP7_75t_L g16 ( .A(n_8), .B(n_1), .Y(n_16) );
INVxp67_ASAP7_75t_L g17 ( .A(n_12), .Y(n_17) );
AOI22xp33_ASAP7_75t_L g18 ( .A1(n_16), .A2(n_11), .B1(n_10), .B2(n_2), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_17), .B(n_2), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
AND2x4_ASAP7_75t_L g21 ( .A(n_18), .B(n_14), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_21), .Y(n_22) );
INVx2_ASAP7_75t_L g23 ( .A(n_20), .Y(n_23) );
AOI22xp33_ASAP7_75t_L g24 ( .A1(n_22), .A2(n_21), .B1(n_14), .B2(n_15), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_23), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
AND2x2_ASAP7_75t_L g27 ( .A(n_24), .B(n_23), .Y(n_27) );
BUFx6f_ASAP7_75t_L g28 ( .A(n_25), .Y(n_28) );
NOR2xp33_ASAP7_75t_L g29 ( .A(n_26), .B(n_27), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_29), .Y(n_30) );
AOI22xp33_ASAP7_75t_R g31 ( .A1(n_30), .A2(n_28), .B1(n_13), .B2(n_9), .Y(n_31) );
endmodule