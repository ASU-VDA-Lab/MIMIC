module fake_jpeg_27262_n_114 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_114);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_114;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_6),
.Y(n_10)
);

INVx11_ASAP7_75t_SL g11 ( 
.A(n_2),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx24_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_2),
.B(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_25),
.Y(n_33)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_27),
.A2(n_13),
.B1(n_17),
.B2(n_12),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_30),
.A2(n_31),
.B1(n_35),
.B2(n_23),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_27),
.A2(n_23),
.B1(n_26),
.B2(n_25),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_27),
.A2(n_23),
.B1(n_26),
.B2(n_25),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_14),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_37),
.B(n_39),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_SL g57 ( 
.A1(n_38),
.A2(n_44),
.B(n_40),
.C(n_39),
.Y(n_57)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_40),
.B(n_41),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_28),
.B(n_14),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_10),
.Y(n_42)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_24),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_21),
.B(n_24),
.C(n_17),
.Y(n_53)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_45),
.A2(n_21),
.B1(n_18),
.B2(n_17),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_12),
.B1(n_16),
.B2(n_15),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_46),
.A2(n_32),
.B1(n_15),
.B2(n_10),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_45),
.A2(n_30),
.B1(n_34),
.B2(n_32),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_47),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_38),
.A2(n_30),
.B1(n_34),
.B2(n_32),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_42),
.A2(n_34),
.B1(n_31),
.B2(n_32),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_44),
.A2(n_34),
.B1(n_32),
.B2(n_16),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_54),
.Y(n_62)
);

AO22x1_ASAP7_75t_L g68 ( 
.A1(n_57),
.A2(n_58),
.B1(n_21),
.B2(n_22),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_49),
.B(n_41),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_60),
.B(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_48),
.B(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_56),
.B(n_20),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_65),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_16),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_43),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_67),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_19),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_69),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_19),
.Y(n_69)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_69),
.B(n_57),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_SL g87 ( 
.A(n_72),
.B(n_77),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_70),
.A2(n_57),
.B1(n_53),
.B2(n_55),
.Y(n_74)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

MAJx2_ASAP7_75t_L g75 ( 
.A(n_62),
.B(n_57),
.C(n_20),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_66),
.A2(n_0),
.B(n_1),
.Y(n_76)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_59),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_62),
.A2(n_19),
.B1(n_22),
.B2(n_29),
.Y(n_80)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_62),
.C(n_68),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_68),
.A2(n_5),
.B1(n_8),
.B2(n_7),
.Y(n_82)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

AOI221xp5_ASAP7_75t_L g83 ( 
.A1(n_75),
.A2(n_64),
.B1(n_6),
.B2(n_7),
.C(n_8),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_80),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_79),
.B(n_64),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_91),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_22),
.Y(n_88)
);

AOI322xp5_ASAP7_75t_SL g91 ( 
.A1(n_73),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_22),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_84),
.A2(n_77),
.B1(n_74),
.B2(n_71),
.Y(n_92)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_89),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_84),
.A2(n_71),
.B1(n_81),
.B2(n_72),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_86),
.A2(n_0),
.B(n_1),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_95),
.A2(n_86),
.B(n_88),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_90),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_98),
.B(n_93),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_99),
.B(n_100),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_96),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_102),
.B(n_104),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_105),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_94),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_99),
.A2(n_87),
.B(n_3),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_29),
.C(n_102),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_108),
.B(n_29),
.Y(n_110)
);

MAJx2_ASAP7_75t_L g109 ( 
.A(n_107),
.B(n_29),
.C(n_106),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_109),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_110),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_111),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_106),
.Y(n_114)
);


endmodule