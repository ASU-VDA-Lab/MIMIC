module real_aes_6420_n_13 (n_4, n_0, n_3, n_5, n_2, n_7, n_8, n_6, n_9, n_12, n_1, n_10, n_11, n_13);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_8;
input n_6;
input n_9;
input n_12;
input n_1;
input n_10;
input n_11;
output n_13;
wire n_28;
wire n_17;
wire n_22;
wire n_24;
wire n_41;
wire n_34;
wire n_19;
wire n_40;
wire n_25;
wire n_32;
wire n_30;
wire n_14;
wire n_16;
wire n_37;
wire n_35;
wire n_39;
wire n_15;
wire n_27;
wire n_23;
wire n_38;
wire n_29;
wire n_20;
wire n_26;
wire n_18;
wire n_21;
wire n_31;
wire n_33;
wire n_36;
NOR2xp33_ASAP7_75t_R g17 ( .A(n_0), .B(n_18), .Y(n_17) );
NAND2xp33_ASAP7_75t_SL g36 ( .A(n_0), .B(n_37), .Y(n_36) );
CKINVDCx20_ASAP7_75t_R g14 ( .A(n_1), .Y(n_14) );
NAND2xp33_ASAP7_75t_SL g25 ( .A(n_1), .B(n_26), .Y(n_25) );
NOR2xp33_ASAP7_75t_R g41 ( .A(n_1), .B(n_12), .Y(n_41) );
CKINVDCx20_ASAP7_75t_R g23 ( .A(n_2), .Y(n_23) );
NOR3xp33_ASAP7_75t_SL g21 ( .A(n_3), .B(n_9), .C(n_22), .Y(n_21) );
INVx1_ASAP7_75t_L g32 ( .A(n_4), .Y(n_32) );
NOR2xp33_ASAP7_75t_R g15 ( .A(n_5), .B(n_16), .Y(n_15) );
CKINVDCx20_ASAP7_75t_R g27 ( .A(n_5), .Y(n_27) );
AOI322xp5_ASAP7_75t_SL g13 ( .A1(n_6), .A2(n_8), .A3(n_14), .B1(n_15), .B2(n_24), .C1(n_28), .C2(n_33), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g22 ( .A(n_7), .Y(n_22) );
CKINVDCx20_ASAP7_75t_R g19 ( .A(n_10), .Y(n_19) );
NOR2xp33_ASAP7_75t_R g33 ( .A(n_10), .B(n_34), .Y(n_33) );
CKINVDCx20_ASAP7_75t_R g18 ( .A(n_11), .Y(n_18) );
NAND4xp25_ASAP7_75t_SL g16 ( .A(n_12), .B(n_17), .C(n_19), .D(n_20), .Y(n_16) );
NOR2xp33_ASAP7_75t_R g26 ( .A(n_16), .B(n_27), .Y(n_26) );
NAND2xp33_ASAP7_75t_SL g40 ( .A(n_18), .B(n_20), .Y(n_40) );
AND2x2_ASAP7_75t_L g20 ( .A(n_21), .B(n_23), .Y(n_20) );
CKINVDCx14_ASAP7_75t_R g24 ( .A(n_25), .Y(n_24) );
NAND2xp33_ASAP7_75t_SL g38 ( .A(n_27), .B(n_39), .Y(n_38) );
BUFx3_ASAP7_75t_L g28 ( .A(n_29), .Y(n_28) );
HB1xp67_ASAP7_75t_L g29 ( .A(n_30), .Y(n_29) );
HB1xp67_ASAP7_75t_L g30 ( .A(n_31), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_32), .Y(n_31) );
NAND2xp33_ASAP7_75t_SL g34 ( .A(n_35), .B(n_41), .Y(n_34) );
CKINVDCx5p33_ASAP7_75t_R g35 ( .A(n_36), .Y(n_35) );
CKINVDCx20_ASAP7_75t_R g37 ( .A(n_38), .Y(n_37) );
CKINVDCx20_ASAP7_75t_R g39 ( .A(n_40), .Y(n_39) );
endmodule