module fake_jpeg_11001_n_304 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_304);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_304;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_265;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx4f_ASAP7_75t_SL g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_43),
.Y(n_103)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_34),
.Y(n_44)
);

INVx4_ASAP7_75t_SL g116 ( 
.A(n_44),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_45),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_20),
.B(n_6),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_46),
.B(n_47),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_20),
.B(n_5),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_23),
.B(n_7),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_49),
.B(n_65),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_30),
.Y(n_52)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_53),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_54),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

BUFx4f_ASAP7_75t_SL g122 ( 
.A(n_56),
.Y(n_122)
);

INVx6_ASAP7_75t_SL g57 ( 
.A(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_58),
.Y(n_86)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_28),
.B(n_21),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_59),
.B(n_67),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_60),
.Y(n_118)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_61),
.Y(n_119)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_64),
.Y(n_88)
);

INVxp67_ASAP7_75t_SL g63 ( 
.A(n_17),
.Y(n_63)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_23),
.B(n_4),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_25),
.B(n_8),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_25),
.B(n_11),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_27),
.B(n_1),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_70),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_27),
.B(n_10),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_69),
.B(n_35),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_29),
.B(n_2),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_29),
.B(n_2),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_71),
.B(n_74),
.Y(n_105)
);

CKINVDCx9p33_ASAP7_75t_R g72 ( 
.A(n_38),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_78),
.Y(n_106)
);

BUFx4f_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

INVx6_ASAP7_75t_SL g74 ( 
.A(n_38),
.Y(n_74)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_17),
.Y(n_75)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_76),
.B(n_79),
.Y(n_107)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_81),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_31),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_35),
.B(n_2),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_83),
.Y(n_111)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_32),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_84),
.B(n_101),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_63),
.A2(n_16),
.B1(n_38),
.B2(n_22),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_95),
.A2(n_100),
.B1(n_104),
.B2(n_118),
.Y(n_158)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_44),
.A2(n_26),
.B(n_41),
.C(n_40),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_96),
.A2(n_106),
.B(n_130),
.C(n_108),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_43),
.A2(n_66),
.B1(n_55),
.B2(n_16),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_97),
.A2(n_127),
.B1(n_10),
.B2(n_60),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_45),
.A2(n_22),
.B1(n_36),
.B2(n_40),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_54),
.B(n_26),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_51),
.B(n_32),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_108),
.B(n_115),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_79),
.A2(n_22),
.B1(n_24),
.B2(n_41),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_112),
.A2(n_125),
.B1(n_106),
.B2(n_97),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_51),
.B(n_39),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_114),
.B(n_117),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_24),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_39),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_121),
.B(n_123),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_81),
.B(n_42),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_50),
.B(n_18),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_128),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_52),
.A2(n_42),
.B1(n_36),
.B2(n_18),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_53),
.A2(n_33),
.B1(n_3),
.B2(n_9),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_56),
.B(n_33),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_73),
.A2(n_0),
.B(n_3),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_130),
.B(n_115),
.C(n_101),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_107),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_131),
.B(n_155),
.Y(n_173)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_134),
.Y(n_179)
);

OAI21xp33_ASAP7_75t_L g135 ( 
.A1(n_84),
.A2(n_10),
.B(n_0),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_135),
.B(n_141),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_89),
.A2(n_75),
.B1(n_61),
.B2(n_60),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_136),
.A2(n_152),
.B1(n_160),
.B2(n_144),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_111),
.B(n_56),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_137),
.B(n_146),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_138),
.A2(n_145),
.B1(n_154),
.B2(n_158),
.Y(n_178)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_139),
.Y(n_172)
);

INVx13_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g183 ( 
.A(n_140),
.Y(n_183)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_90),
.Y(n_143)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_143),
.Y(n_185)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_90),
.Y(n_144)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_144),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_88),
.B(n_102),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_92),
.B(n_93),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_147),
.B(n_149),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_148),
.A2(n_133),
.B(n_162),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_93),
.B(n_98),
.Y(n_149)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_99),
.Y(n_151)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_89),
.A2(n_99),
.B1(n_96),
.B2(n_85),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_85),
.B(n_116),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_153),
.B(n_163),
.C(n_87),
.Y(n_175)
);

OA22x2_ASAP7_75t_L g154 ( 
.A1(n_103),
.A2(n_120),
.B1(n_119),
.B2(n_129),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_86),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_103),
.Y(n_156)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_156),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_105),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_157),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_104),
.Y(n_159)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_159),
.Y(n_195)
);

INVx3_ASAP7_75t_SL g160 ( 
.A(n_126),
.Y(n_160)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_160),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_110),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_166),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_120),
.A2(n_124),
.B(n_91),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_126),
.A2(n_113),
.B1(n_129),
.B2(n_118),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_164),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_122),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_165),
.A2(n_169),
.B1(n_160),
.B2(n_159),
.Y(n_182)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_94),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_94),
.B(n_122),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_167),
.Y(n_194)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_91),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_143),
.Y(n_191)
);

OA22x2_ASAP7_75t_L g169 ( 
.A1(n_119),
.A2(n_113),
.B1(n_122),
.B2(n_87),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_153),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_170),
.B(n_142),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_171),
.B(n_187),
.C(n_201),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_175),
.A2(n_169),
.B(n_154),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_176),
.A2(n_140),
.B1(n_199),
.B2(n_186),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_182),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_148),
.B(n_162),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_188),
.B(n_197),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_191),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_150),
.B(n_131),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_192),
.B(n_196),
.Y(n_213)
);

OAI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_141),
.A2(n_163),
.B1(n_145),
.B2(n_133),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_193),
.A2(n_200),
.B1(n_140),
.B2(n_176),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_150),
.B(n_155),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_161),
.B(n_132),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_153),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_198),
.B(n_201),
.Y(n_205)
);

OAI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_154),
.A2(n_138),
.B1(n_169),
.B2(n_156),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_142),
.B(n_134),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g202 ( 
.A1(n_187),
.A2(n_175),
.B(n_188),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_202),
.B(n_208),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_191),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_203),
.B(n_215),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_204),
.B(n_173),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_171),
.B(n_154),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_225),
.C(n_194),
.Y(n_231)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_190),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_209),
.Y(n_238)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_185),
.Y(n_210)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_210),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_178),
.A2(n_151),
.B1(n_169),
.B2(n_139),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_211),
.B(n_226),
.Y(n_239)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_185),
.Y(n_212)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_212),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g214 ( 
.A(n_170),
.B(n_165),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_214),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_177),
.B(n_165),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_177),
.B(n_166),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_216),
.B(n_217),
.Y(n_242)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_179),
.Y(n_217)
);

OA22x2_ASAP7_75t_L g233 ( 
.A1(n_218),
.A2(n_220),
.B1(n_199),
.B2(n_224),
.Y(n_233)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_186),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_221),
.B(n_223),
.Y(n_245)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_179),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_189),
.A2(n_198),
.B1(n_197),
.B2(n_184),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_224),
.A2(n_187),
.B1(n_192),
.B2(n_196),
.Y(n_228)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_190),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g252 ( 
.A(n_228),
.B(n_230),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_231),
.B(n_202),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_233),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_220),
.A2(n_174),
.B1(n_173),
.B2(n_181),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_240),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_206),
.A2(n_183),
.B1(n_195),
.B2(n_181),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_235),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_214),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_237),
.B(n_243),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_206),
.A2(n_174),
.B1(n_195),
.B2(n_180),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_172),
.C(n_180),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_241),
.B(n_214),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_183),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_246),
.B(n_250),
.C(n_253),
.Y(n_263)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_245),
.Y(n_247)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_247),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_236),
.A2(n_207),
.B(n_208),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_248),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_225),
.Y(n_253)
);

OAI322xp33_ASAP7_75t_L g254 ( 
.A1(n_230),
.A2(n_213),
.A3(n_205),
.B1(n_219),
.B2(n_221),
.C1(n_210),
.C2(n_212),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_254),
.A2(n_228),
.B1(n_234),
.B2(n_231),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_219),
.Y(n_255)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_255),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_238),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_256),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_239),
.A2(n_229),
.B(n_237),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_248),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_227),
.B(n_205),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_258),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_242),
.B(n_183),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_261),
.A2(n_229),
.B1(n_244),
.B2(n_232),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_266),
.A2(n_252),
.B1(n_249),
.B2(n_255),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_267),
.B(n_252),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_268),
.A2(n_247),
.B1(n_249),
.B2(n_251),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_246),
.B(n_241),
.C(n_239),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_270),
.B(n_250),
.C(n_259),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_240),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_270),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_282),
.C(n_281),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_281),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_258),
.Y(n_275)
);

MAJx2_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_276),
.C(n_280),
.Y(n_283)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_264),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_277),
.B(n_279),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_272),
.Y(n_278)
);

OAI31xp33_ASAP7_75t_L g288 ( 
.A1(n_278),
.A2(n_265),
.A3(n_244),
.B(n_232),
.Y(n_288)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_269),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_263),
.B(n_257),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_285),
.B(n_286),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_275),
.B(n_266),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_288),
.A2(n_251),
.B1(n_279),
.B2(n_223),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_271),
.C(n_267),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_289),
.B(n_280),
.C(n_262),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_294),
.C(n_287),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_292),
.B(n_293),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_287),
.A2(n_260),
.B1(n_269),
.B2(n_211),
.Y(n_293)
);

AOI21x1_ASAP7_75t_L g294 ( 
.A1(n_284),
.A2(n_260),
.B(n_282),
.Y(n_294)
);

INVx6_ASAP7_75t_L g296 ( 
.A(n_290),
.Y(n_296)
);

OAI21xp33_ASAP7_75t_L g298 ( 
.A1(n_296),
.A2(n_297),
.B(n_283),
.Y(n_298)
);

OR2x2_ASAP7_75t_L g300 ( 
.A(n_298),
.B(n_299),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_296),
.A2(n_291),
.B(n_293),
.Y(n_299)
);

A2O1A1Ixp33_ASAP7_75t_L g301 ( 
.A1(n_299),
.A2(n_297),
.B(n_295),
.C(n_283),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_295),
.Y(n_302)
);

OAI321xp33_ASAP7_75t_L g303 ( 
.A1(n_302),
.A2(n_300),
.A3(n_226),
.B1(n_233),
.B2(n_209),
.C(n_172),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_303),
.B(n_233),
.Y(n_304)
);


endmodule