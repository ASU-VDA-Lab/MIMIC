module fake_jpeg_23048_n_339 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_46),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_15),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_44),
.B(n_30),
.Y(n_57)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_27),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_55),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_46),
.A2(n_39),
.B1(n_20),
.B2(n_29),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_51),
.A2(n_62),
.B1(n_31),
.B2(n_24),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_27),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_57),
.B(n_21),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_47),
.A2(n_33),
.B1(n_29),
.B2(n_22),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_63),
.B(n_65),
.Y(n_72)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_64),
.B(n_66),
.Y(n_102)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_45),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_54),
.C(n_65),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_71),
.B(n_38),
.C(n_19),
.Y(n_129)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_73),
.B(n_74),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_75),
.Y(n_125)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_76),
.A2(n_77),
.B1(n_83),
.B2(n_88),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_59),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_78),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_79),
.B(n_99),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_57),
.A2(n_33),
.B1(n_49),
.B2(n_47),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_80),
.A2(n_107),
.B1(n_109),
.B2(n_25),
.Y(n_116)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_81),
.Y(n_137)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

INVx4_ASAP7_75t_SL g83 ( 
.A(n_50),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

INVx4_ASAP7_75t_SL g88 ( 
.A(n_61),
.Y(n_88)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_91),
.Y(n_130)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_92),
.Y(n_134)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_52),
.Y(n_93)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_93),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_52),
.A2(n_22),
.B1(n_29),
.B2(n_36),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_94),
.A2(n_104),
.B1(n_106),
.B2(n_83),
.Y(n_132)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_95),
.Y(n_139)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

AO21x2_ASAP7_75t_L g127 ( 
.A1(n_96),
.A2(n_98),
.B(n_101),
.Y(n_127)
);

AOI32xp33_ASAP7_75t_L g97 ( 
.A1(n_67),
.A2(n_41),
.A3(n_22),
.B1(n_43),
.B2(n_42),
.Y(n_97)
);

AOI32xp33_ASAP7_75t_L g126 ( 
.A1(n_97),
.A2(n_48),
.A3(n_38),
.B1(n_19),
.B2(n_34),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_100),
.B(n_103),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

CKINVDCx6p67_ASAP7_75t_R g103 ( 
.A(n_66),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_56),
.A2(n_43),
.B1(n_42),
.B2(n_37),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_63),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_105),
.A2(n_108),
.B(n_110),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_55),
.A2(n_41),
.B1(n_26),
.B2(n_30),
.Y(n_106)
);

O2A1O1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_55),
.A2(n_31),
.B(n_21),
.C(n_24),
.Y(n_107)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_104),
.A2(n_48),
.B1(n_37),
.B2(n_38),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_113),
.A2(n_132),
.B1(n_133),
.B2(n_110),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_116),
.A2(n_123),
.B1(n_74),
.B2(n_87),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_72),
.A2(n_25),
.B(n_32),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_122),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_107),
.A2(n_48),
.B1(n_16),
.B2(n_34),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_89),
.A2(n_32),
.B(n_34),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_138),
.C(n_103),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_126),
.A2(n_90),
.B1(n_92),
.B2(n_105),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_129),
.B(n_0),
.C(n_1),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_94),
.A2(n_34),
.B1(n_28),
.B2(n_19),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_89),
.A2(n_28),
.B(n_19),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_140),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_102),
.B(n_28),
.Y(n_138)
);

OAI32xp33_ASAP7_75t_L g140 ( 
.A1(n_103),
.A2(n_28),
.A3(n_18),
.B1(n_16),
.B2(n_35),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_141),
.Y(n_199)
);

A2O1A1Ixp33_ASAP7_75t_SL g142 ( 
.A1(n_127),
.A2(n_133),
.B(n_140),
.C(n_126),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_142),
.A2(n_139),
.B(n_6),
.Y(n_204)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_127),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_143),
.B(n_147),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_88),
.Y(n_144)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_144),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_100),
.Y(n_145)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_145),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_127),
.A2(n_76),
.B1(n_90),
.B2(n_93),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_146),
.Y(n_178)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_127),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_148),
.B(n_125),
.Y(n_188)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_131),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_149),
.B(n_152),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_150),
.A2(n_153),
.B1(n_163),
.B2(n_168),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_111),
.B(n_73),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_131),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_154),
.Y(n_173)
);

INVx3_ASAP7_75t_SL g155 ( 
.A(n_112),
.Y(n_155)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_155),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_156),
.A2(n_164),
.B1(n_167),
.B2(n_117),
.Y(n_177)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_158),
.Y(n_189)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_119),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_159),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_84),
.C(n_85),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_160),
.B(n_172),
.C(n_135),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_111),
.B(n_15),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_161),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_14),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_162),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_113),
.A2(n_18),
.B1(n_35),
.B2(n_2),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_116),
.A2(n_18),
.B1(n_35),
.B2(n_3),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_125),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_165),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_18),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_170),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_123),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_136),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_168)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_112),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_169),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_128),
.B(n_124),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_115),
.Y(n_171)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_171),
.Y(n_195)
);

AO22x1_ASAP7_75t_SL g174 ( 
.A1(n_141),
.A2(n_118),
.B1(n_122),
.B2(n_128),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_174),
.A2(n_194),
.B1(n_200),
.B2(n_155),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_118),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_175),
.B(n_180),
.C(n_183),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_177),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_235)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_141),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_182),
.B(n_184),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_117),
.C(n_137),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_141),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_130),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_185),
.B(n_139),
.C(n_159),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_137),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_186),
.B(n_167),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_188),
.B(n_165),
.Y(n_228)
);

AO21x2_ASAP7_75t_L g194 ( 
.A1(n_143),
.A2(n_114),
.B(n_121),
.Y(n_194)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_168),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_205),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_151),
.A2(n_114),
.B1(n_135),
.B2(n_121),
.Y(n_200)
);

OAI21xp33_ASAP7_75t_L g201 ( 
.A1(n_151),
.A2(n_157),
.B(n_149),
.Y(n_201)
);

OAI21xp33_ASAP7_75t_L g233 ( 
.A1(n_201),
.A2(n_14),
.B(n_6),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_157),
.B(n_130),
.Y(n_203)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_203),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_204),
.A2(n_158),
.B(n_155),
.Y(n_231)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_153),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_194),
.Y(n_207)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_207),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_178),
.A2(n_171),
.B1(n_147),
.B2(n_142),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_208),
.A2(n_225),
.B1(n_178),
.B2(n_182),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_189),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_209),
.B(n_211),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_175),
.B(n_188),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_210),
.B(n_215),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_198),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_186),
.B(n_164),
.Y(n_213)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_213),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_185),
.B(n_150),
.Y(n_215)
);

NOR2x1_ASAP7_75t_L g216 ( 
.A(n_174),
.B(n_142),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_216),
.A2(n_227),
.B(n_231),
.Y(n_249)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_190),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_224),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_173),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_220),
.B(n_226),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_187),
.B(n_156),
.Y(n_221)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_221),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_180),
.B(n_172),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_228),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_194),
.Y(n_223)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_223),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_187),
.B(n_142),
.Y(n_226)
);

FAx1_ASAP7_75t_L g227 ( 
.A(n_174),
.B(n_142),
.CI(n_163),
.CON(n_227),
.SN(n_227)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_233),
.Y(n_244)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_194),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_230),
.B(n_234),
.Y(n_237)
);

NAND2x1_ASAP7_75t_L g232 ( 
.A(n_194),
.B(n_169),
.Y(n_232)
);

XNOR2x1_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_5),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_181),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_235),
.A2(n_197),
.B1(n_191),
.B2(n_202),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_236),
.A2(n_251),
.B1(n_7),
.B2(n_8),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_225),
.A2(n_205),
.B1(n_184),
.B2(n_177),
.Y(n_239)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_239),
.Y(n_267)
);

OAI22x1_ASAP7_75t_SL g240 ( 
.A1(n_232),
.A2(n_204),
.B1(n_199),
.B2(n_200),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_240),
.A2(n_247),
.B1(n_255),
.B2(n_208),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_210),
.B(n_183),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_217),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_230),
.A2(n_203),
.B1(n_199),
.B2(n_195),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_232),
.A2(n_191),
.B1(n_195),
.B2(n_179),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_252),
.A2(n_257),
.B1(n_227),
.B2(n_7),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_211),
.B(n_196),
.Y(n_254)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_254),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_212),
.A2(n_193),
.B1(n_192),
.B2(n_206),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_219),
.B(n_179),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_256),
.B(n_216),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_212),
.A2(n_181),
.B1(n_176),
.B2(n_8),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_259),
.A2(n_231),
.B(n_218),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_260),
.B(n_261),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_240),
.A2(n_226),
.B(n_213),
.Y(n_261)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_262),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_249),
.A2(n_214),
.B(n_218),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_263),
.A2(n_279),
.B1(n_247),
.B2(n_246),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_257),
.B(n_221),
.Y(n_264)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_264),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_229),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_270),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_266),
.B(n_269),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_217),
.C(n_222),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_272),
.C(n_278),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_215),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_237),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_274),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_243),
.B(n_228),
.C(n_227),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_238),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_273),
.A2(n_275),
.B1(n_244),
.B2(n_8),
.Y(n_288)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_242),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_243),
.B(n_241),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_276),
.B(n_241),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_248),
.B(n_5),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_263),
.A2(n_245),
.B1(n_258),
.B2(n_253),
.Y(n_281)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_281),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_283),
.B(n_291),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_267),
.A2(n_245),
.B1(n_252),
.B2(n_249),
.Y(n_285)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_285),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_246),
.C(n_251),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_289),
.C(n_293),
.Y(n_299)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_287),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_288),
.B(n_271),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_260),
.B(n_272),
.C(n_265),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_244),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_261),
.B(n_7),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_R g296 ( 
.A(n_262),
.B(n_9),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_296),
.Y(n_308)
);

FAx1_ASAP7_75t_SL g300 ( 
.A(n_284),
.B(n_278),
.CI(n_274),
.CON(n_300),
.SN(n_300)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_300),
.B(n_285),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_282),
.B(n_279),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_301),
.B(n_309),
.C(n_270),
.Y(n_319)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_302),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_296),
.Y(n_303)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_303),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_294),
.B(n_273),
.Y(n_305)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_305),
.Y(n_317)
);

INVxp67_ASAP7_75t_SL g306 ( 
.A(n_293),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_270),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_286),
.B(n_275),
.C(n_277),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_290),
.A2(n_295),
.B(n_284),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_310),
.A2(n_292),
.B(n_281),
.Y(n_311)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_311),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_313),
.B(n_315),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_302),
.A2(n_282),
.B(n_289),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_310),
.A2(n_280),
.B(n_291),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_316),
.B(n_318),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_309),
.A2(n_280),
.B(n_283),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_299),
.C(n_304),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_320),
.B(n_308),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_322),
.A2(n_300),
.B(n_304),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_307),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_301),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_314),
.A2(n_297),
.B1(n_298),
.B2(n_300),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_326),
.B(n_327),
.C(n_299),
.Y(n_328)
);

OAI21x1_ASAP7_75t_L g333 ( 
.A1(n_328),
.A2(n_329),
.B(n_330),
.Y(n_333)
);

AOI21xp33_ASAP7_75t_L g329 ( 
.A1(n_321),
.A2(n_312),
.B(n_313),
.Y(n_329)
);

A2O1A1O1Ixp25_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_324),
.B(n_327),
.C(n_321),
.D(n_323),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_332),
.A2(n_326),
.B(n_10),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_333),
.B(n_10),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_336)
);

BUFx24_ASAP7_75t_SL g337 ( 
.A(n_336),
.Y(n_337)
);

OAI321xp33_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_11),
.A3(n_12),
.B1(n_13),
.B2(n_335),
.C(n_333),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_11),
.Y(n_339)
);


endmodule