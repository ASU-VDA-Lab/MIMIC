module fake_jpeg_16627_n_78 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_78);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_78;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx1_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_6),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_1),
.B(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_21),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_17),
.B(n_0),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_22),
.Y(n_29)
);

CKINVDCx9p33_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

INVx3_ASAP7_75t_SL g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx4f_ASAP7_75t_SL g24 ( 
.A(n_18),
.Y(n_24)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_26),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_17),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_27),
.B(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_25),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_33),
.B(n_38),
.Y(n_50)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_19),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_37),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_20),
.B(n_19),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_27),
.B(n_11),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_14),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_43),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_27),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_48),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_32),
.A2(n_22),
.B1(n_12),
.B2(n_14),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_12),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_47),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_39),
.A2(n_24),
.B1(n_10),
.B2(n_16),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_24),
.B1(n_15),
.B2(n_13),
.Y(n_48)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_2),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_41),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_45),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_53),
.Y(n_60)
);

NOR3xp33_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_15),
.C(n_13),
.Y(n_52)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_42),
.Y(n_63)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_58),
.Y(n_64)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_57),
.B(n_50),
.Y(n_59)
);

A2O1A1O1Ixp25_ASAP7_75t_L g68 ( 
.A1(n_59),
.A2(n_61),
.B(n_54),
.C(n_29),
.D(n_42),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_57),
.A2(n_50),
.B(n_49),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_58),
.A2(n_29),
.B1(n_50),
.B2(n_36),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_62),
.A2(n_53),
.B1(n_55),
.B2(n_57),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_62),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_66),
.Y(n_71)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_68),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_68),
.A2(n_64),
.B1(n_61),
.B2(n_59),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_36),
.C(n_29),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_70),
.A2(n_65),
.B(n_63),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_71),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_69),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_74),
.A2(n_75),
.B(n_70),
.Y(n_76)
);

AOI322xp5_ASAP7_75t_L g77 ( 
.A1(n_76),
.A2(n_5),
.A3(n_7),
.B1(n_4),
.B2(n_2),
.C1(n_3),
.C2(n_36),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_5),
.Y(n_78)
);


endmodule