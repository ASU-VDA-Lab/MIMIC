module fake_jpeg_16571_n_122 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_122);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_122;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_6),
.B(n_26),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_6),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_43),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_52),
.B(n_55),
.Y(n_64)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_0),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_49),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_59),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_0),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_53),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_61),
.B(n_66),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

NAND2xp33_ASAP7_75t_SL g67 ( 
.A(n_54),
.B(n_45),
.Y(n_67)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_46),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_70),
.B(n_72),
.Y(n_75)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_85),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_48),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_84),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_41),
.B1(n_38),
.B2(n_50),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_78),
.A2(n_83),
.B1(n_1),
.B2(n_2),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_49),
.Y(n_79)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_81),
.Y(n_88)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_63),
.A2(n_46),
.B1(n_39),
.B2(n_22),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_1),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_80),
.B(n_71),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_92),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_94),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_L g92 ( 
.A1(n_77),
.A2(n_62),
.B1(n_69),
.B2(n_23),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_73),
.B(n_2),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_3),
.Y(n_100)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_75),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_SL g95 ( 
.A(n_81),
.B(n_3),
.C(n_4),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_95),
.A2(n_7),
.B(n_8),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_87),
.C(n_94),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_97),
.B(n_103),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_101),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_96),
.Y(n_101)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_102),
.Y(n_108)
);

A2O1A1O1Ixp25_ASAP7_75t_L g103 ( 
.A1(n_90),
.A2(n_83),
.B(n_9),
.C(n_12),
.D(n_13),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_98),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_104),
.B(n_106),
.Y(n_110)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_107),
.B(n_74),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_105),
.B(n_99),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_111),
.C(n_112),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_110),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_108),
.A2(n_92),
.B1(n_86),
.B2(n_7),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_105),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_113),
.C(n_17),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_16),
.C(n_18),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_117),
.A2(n_19),
.B1(n_20),
.B2(n_27),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_118),
.B(n_29),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_119),
.A2(n_31),
.B(n_32),
.Y(n_120)
);

AOI221xp5_ASAP7_75t_L g121 ( 
.A1(n_120),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.C(n_36),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_37),
.Y(n_122)
);


endmodule