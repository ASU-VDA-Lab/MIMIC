module fake_jpeg_1402_n_189 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_189);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_189;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_2),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_8),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_31),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_30),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_37),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_3),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_13),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_9),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_1),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_33),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_32),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_59),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_71),
.Y(n_81)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_58),
.Y(n_82)
);

AND2x2_ASAP7_75t_SL g73 ( 
.A(n_51),
.B(n_48),
.Y(n_73)
);

NAND2x1_ASAP7_75t_SL g77 ( 
.A(n_73),
.B(n_61),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_68),
.A2(n_48),
.B1(n_47),
.B2(n_53),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_74),
.A2(n_86),
.B1(n_71),
.B2(n_63),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_69),
.A2(n_47),
.B1(n_61),
.B2(n_56),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_76),
.A2(n_63),
.B1(n_54),
.B2(n_52),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_71),
.Y(n_95)
);

NOR2x1_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_57),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_72),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_73),
.B(n_57),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_80),
.B(n_77),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_73),
.A2(n_50),
.B1(n_55),
.B2(n_62),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_85),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_68),
.A2(n_70),
.B1(n_50),
.B2(n_60),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_87),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_121)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_88),
.Y(n_122)
);

NAND2xp33_ASAP7_75t_R g104 ( 
.A(n_89),
.B(n_94),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_85),
.B(n_55),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_91),
.B(n_102),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_80),
.B(n_52),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_92),
.B(n_75),
.Y(n_114)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_103),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_65),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_97),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_65),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_74),
.A2(n_71),
.B1(n_72),
.B2(n_67),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_76),
.A2(n_54),
.B1(n_67),
.B2(n_3),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_5),
.Y(n_120)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_78),
.A2(n_0),
.B(n_4),
.C(n_5),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_46),
.C(n_45),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_90),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_116),
.Y(n_133)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_109),
.Y(n_134)
);

OAI32xp33_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_78),
.A3(n_82),
.B1(n_84),
.B2(n_83),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_113),
.Y(n_135)
);

OAI22x1_ASAP7_75t_SL g112 ( 
.A1(n_94),
.A2(n_84),
.B1(n_75),
.B2(n_83),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_112),
.A2(n_23),
.B1(n_39),
.B2(n_36),
.Y(n_140)
);

INVxp67_ASAP7_75t_SL g113 ( 
.A(n_94),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_114),
.B(n_118),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_102),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_44),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_90),
.A2(n_83),
.B(n_79),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_119),
.A2(n_123),
.B(n_6),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_116),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_98),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_119),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_124),
.B(n_129),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_121),
.A2(n_103),
.B1(n_7),
.B2(n_9),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_125),
.A2(n_137),
.B1(n_122),
.B2(n_15),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_104),
.B(n_114),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_126),
.B(n_109),
.Y(n_154)
);

NAND2xp33_ASAP7_75t_SL g155 ( 
.A(n_128),
.B(n_15),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_115),
.B(n_10),
.Y(n_129)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_130),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_42),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_142),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_110),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_141),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_112),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_111),
.A2(n_11),
.B(n_12),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_138),
.A2(n_122),
.B(n_108),
.Y(n_144)
);

INVxp33_ASAP7_75t_L g153 ( 
.A(n_140),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_118),
.B(n_13),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_41),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_143),
.Y(n_145)
);

AOI221xp5_ASAP7_75t_L g161 ( 
.A1(n_144),
.A2(n_155),
.B1(n_159),
.B2(n_138),
.C(n_125),
.Y(n_161)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

XOR2x1_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_122),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_154),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_150),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_133),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_132),
.B(n_14),
.Y(n_151)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_151),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_139),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_157)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_157),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_135),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_135),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_160),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_161),
.B(n_167),
.Y(n_171)
);

A2O1A1O1Ixp25_ASAP7_75t_L g167 ( 
.A1(n_147),
.A2(n_140),
.B(n_128),
.C(n_131),
.D(n_142),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_154),
.B(n_134),
.C(n_137),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_169),
.B(n_170),
.C(n_152),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_27),
.C(n_34),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_172),
.B(n_174),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_168),
.A2(n_144),
.B1(n_145),
.B2(n_156),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_173),
.A2(n_175),
.B(n_167),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_163),
.B(n_148),
.Y(n_174)
);

AOI322xp5_ASAP7_75t_L g175 ( 
.A1(n_165),
.A2(n_158),
.A3(n_153),
.B1(n_159),
.B2(n_149),
.C1(n_19),
.C2(n_22),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_170),
.B(n_153),
.C(n_28),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_176),
.B(n_29),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_177),
.B(n_180),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_173),
.A2(n_169),
.B(n_166),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_179),
.B(n_171),
.C(n_166),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_182),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_183),
.B(n_178),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_184),
.A2(n_181),
.B(n_164),
.Y(n_185)
);

A2O1A1Ixp33_ASAP7_75t_SL g186 ( 
.A1(n_185),
.A2(n_162),
.B(n_26),
.C(n_35),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_186),
.A2(n_20),
.B(n_21),
.Y(n_187)
);

OAI21x1_ASAP7_75t_L g188 ( 
.A1(n_187),
.A2(n_20),
.B(n_21),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_22),
.Y(n_189)
);


endmodule