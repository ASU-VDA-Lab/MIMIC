module real_aes_10830_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_1380;
wire n_501;
wire n_488;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_264;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_1404;
wire n_402;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_720;
wire n_354;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_1343;
wire n_719;
wire n_1156;
wire n_988;
wire n_1396;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_1352;
wire n_729;
wire n_1323;
wire n_1280;
wire n_703;
wire n_1369;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AO221x1_ASAP7_75t_L g1148 ( .A1(n_0), .A2(n_143), .B1(n_1121), .B2(n_1149), .C(n_1151), .Y(n_1148) );
AOI21xp33_ASAP7_75t_L g786 ( .A1(n_1), .A2(n_413), .B(n_661), .Y(n_786) );
INVx1_ASAP7_75t_L g817 ( .A(n_1), .Y(n_817) );
INVx1_ASAP7_75t_L g581 ( .A(n_2), .Y(n_581) );
OAI221xp5_ASAP7_75t_L g611 ( .A1(n_2), .A2(n_68), .B1(n_523), .B2(n_526), .C(n_529), .Y(n_611) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_3), .A2(n_244), .B1(n_413), .B2(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g620 ( .A(n_3), .Y(n_620) );
OAI221xp5_ASAP7_75t_L g903 ( .A1(n_4), .A2(n_532), .B1(n_904), .B2(n_906), .C(n_912), .Y(n_903) );
AOI21xp33_ASAP7_75t_L g936 ( .A1(n_4), .A2(n_579), .B(n_937), .Y(n_936) );
AOI22xp33_ASAP7_75t_SL g1024 ( .A1(n_5), .A2(n_71), .B1(n_1016), .B2(n_1017), .Y(n_1024) );
INVxp67_ASAP7_75t_SL g1043 ( .A(n_5), .Y(n_1043) );
INVx1_ASAP7_75t_L g1390 ( .A(n_6), .Y(n_1390) );
OAI221xp5_ASAP7_75t_L g1417 ( .A1(n_6), .A2(n_28), .B1(n_478), .B2(n_1418), .C(n_1419), .Y(n_1417) );
HB1xp67_ASAP7_75t_L g264 ( .A(n_7), .Y(n_264) );
AND2x2_ASAP7_75t_L g285 ( .A(n_7), .B(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g317 ( .A(n_7), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_7), .B(n_182), .Y(n_326) );
AOI221xp5_ASAP7_75t_L g639 ( .A1(n_8), .A2(n_140), .B1(n_588), .B2(n_640), .C(n_641), .Y(n_639) );
INVx1_ASAP7_75t_L g682 ( .A(n_8), .Y(n_682) );
INVx1_ASAP7_75t_L g874 ( .A(n_9), .Y(n_874) );
AOI22xp5_ASAP7_75t_L g1130 ( .A1(n_10), .A2(n_104), .B1(n_1121), .B2(n_1125), .Y(n_1130) );
XNOR2x2_ASAP7_75t_L g277 ( .A(n_11), .B(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g880 ( .A(n_12), .Y(n_880) );
OAI221xp5_ASAP7_75t_L g915 ( .A1(n_13), .A2(n_22), .B1(n_524), .B2(n_527), .C(n_530), .Y(n_915) );
CKINVDCx5p33_ASAP7_75t_R g944 ( .A(n_13), .Y(n_944) );
INVx1_ASAP7_75t_L g1329 ( .A(n_14), .Y(n_1329) );
AOI22xp33_ASAP7_75t_SL g1393 ( .A1(n_15), .A2(n_177), .B1(n_1394), .B2(n_1395), .Y(n_1393) );
AOI221xp5_ASAP7_75t_L g1426 ( .A1(n_15), .A2(n_63), .B1(n_465), .B2(n_586), .C(n_983), .Y(n_1426) );
AOI221xp5_ASAP7_75t_L g585 ( .A1(n_16), .A2(n_34), .B1(n_586), .B2(n_587), .C(n_588), .Y(n_585) );
INVx1_ASAP7_75t_L g621 ( .A(n_16), .Y(n_621) );
AOI221xp5_ASAP7_75t_L g463 ( .A1(n_17), .A2(n_234), .B1(n_464), .B2(n_465), .C(n_467), .Y(n_463) );
INVx1_ASAP7_75t_L g517 ( .A(n_17), .Y(n_517) );
AO22x1_ASAP7_75t_L g1159 ( .A1(n_18), .A2(n_240), .B1(n_1109), .B2(n_1117), .Y(n_1159) );
AO221x2_ASAP7_75t_L g1269 ( .A1(n_19), .A2(n_156), .B1(n_1149), .B2(n_1270), .C(n_1272), .Y(n_1269) );
AOI221xp5_ASAP7_75t_L g1062 ( .A1(n_20), .A2(n_205), .B1(n_465), .B2(n_660), .C(n_661), .Y(n_1062) );
INVx1_ASAP7_75t_L g1086 ( .A(n_20), .Y(n_1086) );
OAI221xp5_ASAP7_75t_L g764 ( .A1(n_21), .A2(n_712), .B1(n_765), .B2(n_771), .C(n_776), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g804 ( .A1(n_21), .A2(n_157), .B1(n_796), .B2(n_805), .Y(n_804) );
CKINVDCx5p33_ASAP7_75t_R g943 ( .A(n_22), .Y(n_943) );
AOI22xp33_ASAP7_75t_L g1396 ( .A1(n_23), .A2(n_63), .B1(n_1397), .B2(n_1398), .Y(n_1396) );
AOI22xp33_ASAP7_75t_L g1427 ( .A1(n_23), .A2(n_177), .B1(n_1064), .B2(n_1074), .Y(n_1427) );
INVx2_ASAP7_75t_L g373 ( .A(n_24), .Y(n_373) );
OR2x2_ASAP7_75t_L g446 ( .A(n_24), .B(n_371), .Y(n_446) );
AOI221xp5_ASAP7_75t_L g966 ( .A1(n_25), .A2(n_170), .B1(n_299), .B2(n_967), .C(n_968), .Y(n_966) );
INVx1_ASAP7_75t_L g977 ( .A(n_25), .Y(n_977) );
OAI22xp5_ASAP7_75t_L g1319 ( .A1(n_26), .A2(n_100), .B1(n_1320), .B2(n_1321), .Y(n_1319) );
OAI221xp5_ASAP7_75t_L g1365 ( .A1(n_26), .A2(n_100), .B1(n_526), .B2(n_529), .C(n_675), .Y(n_1365) );
OAI22xp5_ASAP7_75t_L g725 ( .A1(n_27), .A2(n_219), .B1(n_478), .B2(n_726), .Y(n_725) );
OAI221xp5_ASAP7_75t_L g739 ( .A1(n_27), .A2(n_219), .B1(n_526), .B2(n_529), .C(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g1389 ( .A(n_28), .Y(n_1389) );
BUFx2_ASAP7_75t_L g362 ( .A(n_29), .Y(n_362) );
BUFx2_ASAP7_75t_L g367 ( .A(n_29), .Y(n_367) );
INVx1_ASAP7_75t_L g434 ( .A(n_29), .Y(n_434) );
OR2x2_ASAP7_75t_L g505 ( .A(n_29), .B(n_326), .Y(n_505) );
INVx1_ASAP7_75t_L g700 ( .A(n_30), .Y(n_700) );
INVx1_ASAP7_75t_L g1342 ( .A(n_31), .Y(n_1342) );
INVx1_ASAP7_75t_L g952 ( .A(n_32), .Y(n_952) );
AOI22xp33_ASAP7_75t_SL g911 ( .A1(n_33), .A2(n_146), .B1(n_312), .B2(n_383), .Y(n_911) );
INVx1_ASAP7_75t_L g928 ( .A(n_33), .Y(n_928) );
INVx1_ASAP7_75t_L g614 ( .A(n_34), .Y(n_614) );
CKINVDCx5p33_ASAP7_75t_R g593 ( .A(n_35), .Y(n_593) );
OAI22xp5_ASAP7_75t_L g1065 ( .A1(n_36), .A2(n_62), .B1(n_475), .B2(n_1066), .Y(n_1065) );
OAI221xp5_ASAP7_75t_L g1088 ( .A1(n_36), .A2(n_62), .B1(n_523), .B2(n_526), .C(n_530), .Y(n_1088) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_37), .A2(n_127), .B1(n_470), .B2(n_598), .Y(n_785) );
INVx1_ASAP7_75t_L g818 ( .A(n_37), .Y(n_818) );
AOI22xp33_ASAP7_75t_SL g1015 ( .A1(n_38), .A2(n_167), .B1(n_1016), .B2(n_1017), .Y(n_1015) );
AOI221xp5_ASAP7_75t_L g1044 ( .A1(n_38), .A2(n_226), .B1(n_408), .B2(n_843), .C(n_1045), .Y(n_1044) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_39), .A2(n_82), .B1(n_295), .B2(n_616), .Y(n_913) );
OAI22xp5_ASAP7_75t_L g921 ( .A1(n_39), .A2(n_82), .B1(n_500), .B2(n_778), .Y(n_921) );
AOI22xp33_ASAP7_75t_L g717 ( .A1(n_40), .A2(n_188), .B1(n_643), .B2(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g745 ( .A(n_40), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g1401 ( .A1(n_41), .A2(n_50), .B1(n_1402), .B2(n_1404), .Y(n_1401) );
INVx1_ASAP7_75t_L g1429 ( .A(n_41), .Y(n_1429) );
INVx1_ASAP7_75t_L g959 ( .A(n_42), .Y(n_959) );
AOI22xp33_ASAP7_75t_L g292 ( .A1(n_43), .A2(n_46), .B1(n_293), .B2(n_299), .Y(n_292) );
OAI22xp5_ASAP7_75t_L g450 ( .A1(n_43), .A2(n_61), .B1(n_451), .B2(n_453), .Y(n_450) );
CKINVDCx5p33_ASAP7_75t_R g851 ( .A(n_44), .Y(n_851) );
INVx1_ASAP7_75t_L g1152 ( .A(n_45), .Y(n_1152) );
INVxp67_ASAP7_75t_SL g447 ( .A(n_46), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g1338 ( .A1(n_47), .A2(n_176), .B1(n_844), .B2(n_1339), .Y(n_1338) );
INVxp67_ASAP7_75t_SL g1350 ( .A(n_47), .Y(n_1350) );
INVx1_ASAP7_75t_L g908 ( .A(n_48), .Y(n_908) );
AOI21xp33_ASAP7_75t_L g926 ( .A1(n_48), .A2(n_483), .B(n_586), .Y(n_926) );
AOI22xp33_ASAP7_75t_SL g1023 ( .A1(n_49), .A2(n_85), .B1(n_1020), .B2(n_1021), .Y(n_1023) );
INVxp33_ASAP7_75t_SL g1053 ( .A(n_49), .Y(n_1053) );
INVx1_ASAP7_75t_L g1425 ( .A(n_50), .Y(n_1425) );
OAI22xp33_ASAP7_75t_L g787 ( .A1(n_51), .A2(n_157), .B1(n_496), .B2(n_500), .Y(n_787) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_51), .A2(n_241), .B1(n_798), .B2(n_802), .Y(n_801) );
INVx1_ASAP7_75t_L g348 ( .A(n_52), .Y(n_348) );
INVx1_ASAP7_75t_L g1335 ( .A(n_53), .Y(n_1335) );
AOI221xp5_ASAP7_75t_L g714 ( .A1(n_54), .A2(n_64), .B1(n_465), .B2(n_586), .C(n_715), .Y(n_714) );
INVxp67_ASAP7_75t_SL g746 ( .A(n_54), .Y(n_746) );
CKINVDCx5p33_ASAP7_75t_R g656 ( .A(n_55), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_56), .A2(n_181), .B1(n_843), .B2(n_844), .Y(n_842) );
OAI22xp33_ASAP7_75t_L g858 ( .A1(n_56), .A2(n_247), .B1(n_281), .B2(n_859), .Y(n_858) );
AOI221xp5_ASAP7_75t_L g1323 ( .A1(n_57), .A2(n_206), .B1(n_1324), .B2(n_1326), .C(n_1328), .Y(n_1323) );
INVxp33_ASAP7_75t_L g1371 ( .A(n_57), .Y(n_1371) );
INVx1_ASAP7_75t_L g1315 ( .A(n_58), .Y(n_1315) );
CKINVDCx5p33_ASAP7_75t_R g853 ( .A(n_59), .Y(n_853) );
INVx1_ASAP7_75t_L g1153 ( .A(n_60), .Y(n_1153) );
AOI221xp5_ASAP7_75t_L g304 ( .A1(n_61), .A2(n_169), .B1(n_305), .B2(n_310), .C(n_313), .Y(n_304) );
INVxp67_ASAP7_75t_SL g750 ( .A(n_64), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g1073 ( .A1(n_65), .A2(n_236), .B1(n_591), .B2(n_1074), .Y(n_1073) );
INVx1_ASAP7_75t_L g1091 ( .A(n_65), .Y(n_1091) );
AOI221xp5_ASAP7_75t_L g954 ( .A1(n_66), .A2(n_120), .B1(n_876), .B2(n_955), .C(n_956), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g984 ( .A1(n_66), .A2(n_83), .B1(n_985), .B2(n_986), .Y(n_984) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_67), .A2(n_216), .B1(n_418), .B2(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g519 ( .A(n_67), .Y(n_519) );
INVx1_ASAP7_75t_L g582 ( .A(n_68), .Y(n_582) );
CKINVDCx5p33_ASAP7_75t_R g910 ( .A(n_69), .Y(n_910) );
AO221x1_ASAP7_75t_L g1132 ( .A1(n_70), .A2(n_111), .B1(n_1121), .B2(n_1125), .C(n_1133), .Y(n_1132) );
INVxp33_ASAP7_75t_L g1052 ( .A(n_71), .Y(n_1052) );
INVx1_ASAP7_75t_L g958 ( .A(n_72), .Y(n_958) );
AOI221xp5_ASAP7_75t_L g979 ( .A1(n_72), .A2(n_120), .B1(n_980), .B2(n_981), .C(n_983), .Y(n_979) );
INVx1_ASAP7_75t_L g1275 ( .A(n_73), .Y(n_1275) );
AO221x1_ASAP7_75t_L g1138 ( .A1(n_74), .A2(n_150), .B1(n_1121), .B2(n_1125), .C(n_1139), .Y(n_1138) );
INVx1_ASAP7_75t_L g1140 ( .A(n_75), .Y(n_1140) );
INVx1_ASAP7_75t_L g371 ( .A(n_76), .Y(n_371) );
INVx1_ASAP7_75t_L g406 ( .A(n_76), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_77), .A2(n_228), .B1(n_643), .B2(n_645), .Y(n_642) );
INVx1_ASAP7_75t_L g691 ( .A(n_77), .Y(n_691) );
INVx1_ASAP7_75t_L g709 ( .A(n_78), .Y(n_709) );
INVx1_ASAP7_75t_L g969 ( .A(n_79), .Y(n_969) );
OAI221xp5_ASAP7_75t_L g973 ( .A1(n_79), .A2(n_170), .B1(n_398), .B2(n_974), .C(n_976), .Y(n_973) );
INVx1_ASAP7_75t_L g772 ( .A(n_80), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g794 ( .A1(n_80), .A2(n_142), .B1(n_795), .B2(n_796), .Y(n_794) );
NAND2xp33_ASAP7_75t_SL g576 ( .A(n_81), .B(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g606 ( .A(n_81), .Y(n_606) );
INVxp67_ASAP7_75t_SL g957 ( .A(n_83), .Y(n_957) );
INVxp67_ASAP7_75t_SL g1001 ( .A(n_84), .Y(n_1001) );
OAI22xp33_ASAP7_75t_L g1030 ( .A1(n_84), .A2(n_203), .B1(n_1031), .B2(n_1032), .Y(n_1030) );
INVxp67_ASAP7_75t_SL g1029 ( .A(n_85), .Y(n_1029) );
OAI22xp33_ASAP7_75t_L g919 ( .A1(n_86), .A2(n_136), .B1(n_504), .B2(n_820), .Y(n_919) );
AOI22xp33_ASAP7_75t_L g935 ( .A1(n_86), .A2(n_192), .B1(n_396), .B2(n_591), .Y(n_935) );
INVx1_ASAP7_75t_L g964 ( .A(n_87), .Y(n_964) );
AOI221xp5_ASAP7_75t_L g988 ( .A1(n_87), .A2(n_131), .B1(n_392), .B2(n_579), .C(n_640), .Y(n_988) );
INVx1_ASAP7_75t_L g354 ( .A(n_88), .Y(n_354) );
AOI221xp5_ASAP7_75t_L g385 ( .A1(n_88), .A2(n_238), .B1(n_386), .B2(n_391), .C(n_394), .Y(n_385) );
OAI22xp5_ASAP7_75t_L g917 ( .A1(n_89), .A2(n_192), .B1(n_821), .B2(n_918), .Y(n_917) );
INVx1_ASAP7_75t_L g933 ( .A(n_89), .Y(n_933) );
AOI22xp5_ASAP7_75t_L g1382 ( .A1(n_90), .A2(n_1383), .B1(n_1384), .B2(n_1385), .Y(n_1382) );
CKINVDCx5p33_ASAP7_75t_R g1383 ( .A(n_90), .Y(n_1383) );
CKINVDCx5p33_ASAP7_75t_R g494 ( .A(n_91), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g760 ( .A1(n_92), .A2(n_761), .B1(n_822), .B2(n_823), .Y(n_760) );
INVxp67_ASAP7_75t_SL g822 ( .A(n_92), .Y(n_822) );
CKINVDCx20_ASAP7_75t_R g568 ( .A(n_93), .Y(n_568) );
OAI21xp33_ASAP7_75t_L g948 ( .A1(n_94), .A2(n_949), .B(n_971), .Y(n_948) );
INVx1_ASAP7_75t_L g995 ( .A(n_94), .Y(n_995) );
INVx1_ASAP7_75t_L g970 ( .A(n_95), .Y(n_970) );
AOI22xp33_ASAP7_75t_L g1164 ( .A1(n_96), .A2(n_220), .B1(n_1121), .B2(n_1125), .Y(n_1164) );
AOI221xp5_ASAP7_75t_L g481 ( .A1(n_97), .A2(n_199), .B1(n_465), .B2(n_482), .C(n_483), .Y(n_481) );
INVx1_ASAP7_75t_L g545 ( .A(n_97), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_98), .A2(n_211), .B1(n_723), .B2(n_724), .Y(n_722) );
INVx1_ASAP7_75t_L g738 ( .A(n_98), .Y(n_738) );
CKINVDCx5p33_ASAP7_75t_R g596 ( .A(n_99), .Y(n_596) );
AOI221xp5_ASAP7_75t_L g721 ( .A1(n_101), .A2(n_193), .B1(n_413), .B2(n_465), .C(n_661), .Y(n_721) );
INVx1_ASAP7_75t_L g737 ( .A(n_101), .Y(n_737) );
INVx1_ASAP7_75t_L g1136 ( .A(n_102), .Y(n_1136) );
INVx1_ASAP7_75t_L g256 ( .A(n_103), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g501 ( .A(n_105), .Y(n_501) );
INVx1_ASAP7_75t_L g600 ( .A(n_106), .Y(n_600) );
CKINVDCx5p33_ASAP7_75t_R g1077 ( .A(n_107), .Y(n_1077) );
OA22x2_ASAP7_75t_L g458 ( .A1(n_108), .A2(n_459), .B1(n_558), .B2(n_559), .Y(n_458) );
INVx1_ASAP7_75t_L g559 ( .A(n_108), .Y(n_559) );
INVx1_ASAP7_75t_L g1098 ( .A(n_109), .Y(n_1098) );
AOI22xp5_ASAP7_75t_L g1108 ( .A1(n_110), .A2(n_184), .B1(n_1109), .B2(n_1117), .Y(n_1108) );
OAI221xp5_ASAP7_75t_SL g962 ( .A1(n_112), .A2(n_217), .B1(n_346), .B2(n_686), .C(n_963), .Y(n_962) );
AOI22xp33_ASAP7_75t_L g989 ( .A1(n_112), .A2(n_217), .B1(n_641), .B2(n_645), .Y(n_989) );
AOI22xp33_ASAP7_75t_L g1063 ( .A1(n_113), .A2(n_173), .B1(n_655), .B2(n_1064), .Y(n_1063) );
INVx1_ASAP7_75t_L g1083 ( .A(n_113), .Y(n_1083) );
AOI22xp33_ASAP7_75t_L g1399 ( .A1(n_114), .A2(n_171), .B1(n_293), .B2(n_1400), .Y(n_1399) );
INVx1_ASAP7_75t_L g1430 ( .A(n_114), .Y(n_1430) );
AOI22xp33_ASAP7_75t_SL g573 ( .A1(n_115), .A2(n_195), .B1(n_574), .B2(n_575), .Y(n_573) );
INVx1_ASAP7_75t_L g609 ( .A(n_115), .Y(n_609) );
XOR2xp5_ASAP7_75t_L g900 ( .A(n_116), .B(n_901), .Y(n_900) );
AOI22xp5_ASAP7_75t_L g1120 ( .A1(n_117), .A2(n_162), .B1(n_1121), .B2(n_1125), .Y(n_1120) );
AOI22xp5_ASAP7_75t_L g1165 ( .A1(n_118), .A2(n_248), .B1(n_1109), .B2(n_1117), .Y(n_1165) );
INVx1_ASAP7_75t_L g364 ( .A(n_119), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g663 ( .A(n_121), .Y(n_663) );
CKINVDCx5p33_ASAP7_75t_R g1407 ( .A(n_122), .Y(n_1407) );
CKINVDCx5p33_ASAP7_75t_R g498 ( .A(n_123), .Y(n_498) );
AOI221xp5_ASAP7_75t_L g659 ( .A1(n_124), .A2(n_245), .B1(n_640), .B2(n_660), .C(n_661), .Y(n_659) );
INVx1_ASAP7_75t_L g670 ( .A(n_124), .Y(n_670) );
CKINVDCx5p33_ASAP7_75t_R g781 ( .A(n_125), .Y(n_781) );
CKINVDCx5p33_ASAP7_75t_R g584 ( .A(n_126), .Y(n_584) );
OAI22xp5_ASAP7_75t_L g819 ( .A1(n_127), .A2(n_230), .B1(n_820), .B2(n_821), .Y(n_819) );
INVx1_ASAP7_75t_L g1273 ( .A(n_128), .Y(n_1273) );
AOI22xp33_ASAP7_75t_L g835 ( .A1(n_129), .A2(n_231), .B1(n_836), .B2(n_837), .Y(n_835) );
INVx1_ASAP7_75t_L g863 ( .A(n_129), .Y(n_863) );
INVx1_ASAP7_75t_L g650 ( .A(n_130), .Y(n_650) );
OAI221xp5_ASAP7_75t_L g674 ( .A1(n_130), .A2(n_212), .B1(n_527), .B2(n_675), .C(n_677), .Y(n_674) );
INVx1_ASAP7_75t_L g965 ( .A(n_131), .Y(n_965) );
CKINVDCx5p33_ASAP7_75t_R g1076 ( .A(n_132), .Y(n_1076) );
INVx1_ASAP7_75t_L g1406 ( .A(n_133), .Y(n_1406) );
AOI22xp33_ASAP7_75t_L g1420 ( .A1(n_133), .A2(n_208), .B1(n_396), .B2(n_399), .Y(n_1420) );
OAI22xp5_ASAP7_75t_L g318 ( .A1(n_134), .A2(n_153), .B1(n_319), .B2(n_327), .Y(n_318) );
OAI221xp5_ASAP7_75t_L g424 ( .A1(n_134), .A2(n_153), .B1(n_425), .B2(n_435), .C(n_439), .Y(n_424) );
CKINVDCx5p33_ASAP7_75t_R g1069 ( .A(n_135), .Y(n_1069) );
INVx1_ASAP7_75t_L g939 ( .A(n_136), .Y(n_939) );
CKINVDCx5p33_ASAP7_75t_R g638 ( .A(n_137), .Y(n_638) );
CKINVDCx5p33_ASAP7_75t_R g1026 ( .A(n_138), .Y(n_1026) );
INVx1_ASAP7_75t_L g713 ( .A(n_139), .Y(n_713) );
INVx1_ASAP7_75t_L g688 ( .A(n_140), .Y(n_688) );
CKINVDCx5p33_ASAP7_75t_R g883 ( .A(n_141), .Y(n_883) );
INVx1_ASAP7_75t_L g768 ( .A(n_142), .Y(n_768) );
XOR2x2_ASAP7_75t_L g996 ( .A(n_144), .B(n_997), .Y(n_996) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_145), .A2(n_247), .B1(n_412), .B2(n_839), .Y(n_841) );
OAI22xp33_ASAP7_75t_L g891 ( .A1(n_145), .A2(n_181), .B1(n_337), .B2(n_892), .Y(n_891) );
INVx1_ASAP7_75t_L g925 ( .A(n_146), .Y(n_925) );
AOI221xp5_ASAP7_75t_L g1070 ( .A1(n_147), .A2(n_209), .B1(n_417), .B2(n_715), .C(n_1071), .Y(n_1070) );
INVx1_ASAP7_75t_L g1094 ( .A(n_147), .Y(n_1094) );
AOI21xp33_ASAP7_75t_L g775 ( .A1(n_148), .A2(n_483), .B(n_641), .Y(n_775) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_148), .A2(n_229), .B1(n_798), .B2(n_800), .Y(n_797) );
AOI221xp5_ASAP7_75t_L g1336 ( .A1(n_149), .A2(n_235), .B1(n_655), .B2(n_715), .C(n_1337), .Y(n_1336) );
INVxp33_ASAP7_75t_SL g1355 ( .A(n_149), .Y(n_1355) );
INVx1_ASAP7_75t_L g1318 ( .A(n_151), .Y(n_1318) );
HB1xp67_ASAP7_75t_L g258 ( .A(n_152), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g1116 ( .A(n_152), .B(n_256), .Y(n_1116) );
AND3x2_ASAP7_75t_L g1124 ( .A(n_152), .B(n_256), .C(n_1113), .Y(n_1124) );
INVx2_ASAP7_75t_L g269 ( .A(n_154), .Y(n_269) );
INVx1_ASAP7_75t_L g727 ( .A(n_155), .Y(n_727) );
XOR2xp5_ASAP7_75t_L g1312 ( .A(n_156), .B(n_1313), .Y(n_1312) );
AOI22xp33_ASAP7_75t_L g1376 ( .A1(n_156), .A2(n_1377), .B1(n_1381), .B2(n_1432), .Y(n_1376) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_158), .A2(n_223), .B1(n_464), .B2(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g537 ( .A(n_158), .Y(n_537) );
INVx1_ASAP7_75t_L g1330 ( .A(n_159), .Y(n_1330) );
CKINVDCx5p33_ASAP7_75t_R g490 ( .A(n_160), .Y(n_490) );
CKINVDCx5p33_ASAP7_75t_R g1009 ( .A(n_161), .Y(n_1009) );
INVx1_ASAP7_75t_L g951 ( .A(n_163), .Y(n_951) );
INVxp33_ASAP7_75t_SL g1010 ( .A(n_164), .Y(n_1010) );
AOI221xp5_ASAP7_75t_L g1034 ( .A1(n_164), .A2(n_210), .B1(n_1035), .B2(n_1037), .C(n_1038), .Y(n_1034) );
CKINVDCx5p33_ASAP7_75t_R g780 ( .A(n_165), .Y(n_780) );
INVx1_ASAP7_75t_L g345 ( .A(n_166), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g1047 ( .A1(n_167), .A2(n_191), .B1(n_645), .B2(n_1048), .Y(n_1047) );
INVx1_ASAP7_75t_L g1113 ( .A(n_168), .Y(n_1113) );
INVxp67_ASAP7_75t_SL g449 ( .A(n_169), .Y(n_449) );
INVx1_ASAP7_75t_L g1416 ( .A(n_171), .Y(n_1416) );
AOI22xp33_ASAP7_75t_L g914 ( .A1(n_172), .A2(n_239), .B1(n_312), .B2(n_383), .Y(n_914) );
OAI22xp5_ASAP7_75t_L g922 ( .A1(n_172), .A2(n_239), .B1(n_496), .B2(n_712), .Y(n_922) );
INVx1_ASAP7_75t_L g1087 ( .A(n_173), .Y(n_1087) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_174), .A2(n_221), .B1(n_412), .B2(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g869 ( .A(n_174), .Y(n_869) );
CKINVDCx5p33_ASAP7_75t_R g1431 ( .A(n_175), .Y(n_1431) );
INVxp33_ASAP7_75t_L g1353 ( .A(n_176), .Y(n_1353) );
OAI211xp5_ASAP7_75t_L g280 ( .A1(n_178), .A2(n_281), .B(n_291), .C(n_329), .Y(n_280) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_178), .A2(n_187), .B1(n_408), .B2(n_412), .C(n_415), .Y(n_407) );
INVx1_ASAP7_75t_L g1343 ( .A(n_179), .Y(n_1343) );
CKINVDCx5p33_ASAP7_75t_R g1061 ( .A(n_180), .Y(n_1061) );
INVx1_ASAP7_75t_L g271 ( .A(n_182), .Y(n_271) );
INVx2_ASAP7_75t_L g286 ( .A(n_182), .Y(n_286) );
INVx1_ASAP7_75t_L g330 ( .A(n_183), .Y(n_330) );
AOI22xp5_ASAP7_75t_L g1129 ( .A1(n_185), .A2(n_201), .B1(n_1109), .B2(n_1117), .Y(n_1129) );
OR2x2_ASAP7_75t_L g762 ( .A(n_186), .B(n_503), .Y(n_762) );
OAI221xp5_ASAP7_75t_L g336 ( .A1(n_187), .A2(n_337), .B1(n_340), .B2(n_349), .C(n_358), .Y(n_336) );
INVx1_ASAP7_75t_L g751 ( .A(n_188), .Y(n_751) );
OAI22xp5_ASAP7_75t_L g703 ( .A1(n_189), .A2(n_704), .B1(n_758), .B2(n_759), .Y(n_703) );
INVx1_ASAP7_75t_L g759 ( .A(n_189), .Y(n_759) );
INVx1_ASAP7_75t_L g1409 ( .A(n_190), .Y(n_1409) );
AOI21xp33_ASAP7_75t_L g1421 ( .A1(n_190), .A2(n_579), .B(n_1422), .Y(n_1421) );
AOI22xp33_ASAP7_75t_SL g1019 ( .A1(n_191), .A2(n_226), .B1(n_1020), .B2(n_1021), .Y(n_1019) );
INVx1_ASAP7_75t_L g733 ( .A(n_193), .Y(n_733) );
CKINVDCx5p33_ASAP7_75t_R g647 ( .A(n_194), .Y(n_647) );
INVx1_ASAP7_75t_L g604 ( .A(n_195), .Y(n_604) );
CKINVDCx5p33_ASAP7_75t_R g648 ( .A(n_196), .Y(n_648) );
INVx1_ASAP7_75t_L g887 ( .A(n_197), .Y(n_887) );
CKINVDCx5p33_ASAP7_75t_R g594 ( .A(n_198), .Y(n_594) );
INVx1_ASAP7_75t_L g541 ( .A(n_199), .Y(n_541) );
CKINVDCx5p33_ASAP7_75t_R g473 ( .A(n_200), .Y(n_473) );
XOR2xp5_ASAP7_75t_L g830 ( .A(n_201), .B(n_831), .Y(n_830) );
INVx1_ASAP7_75t_L g878 ( .A(n_202), .Y(n_878) );
INVxp67_ASAP7_75t_SL g1004 ( .A(n_203), .Y(n_1004) );
INVx1_ASAP7_75t_L g1007 ( .A(n_204), .Y(n_1007) );
INVx1_ASAP7_75t_L g1084 ( .A(n_205), .Y(n_1084) );
INVxp33_ASAP7_75t_L g1368 ( .A(n_206), .Y(n_1368) );
OAI22xp5_ASAP7_75t_L g474 ( .A1(n_207), .A2(n_214), .B1(n_475), .B2(n_478), .Y(n_474) );
OAI221xp5_ASAP7_75t_L g522 ( .A1(n_207), .A2(n_214), .B1(n_523), .B2(n_526), .C(n_529), .Y(n_522) );
INVx1_ASAP7_75t_L g1410 ( .A(n_208), .Y(n_1410) );
INVx1_ASAP7_75t_L g1092 ( .A(n_209), .Y(n_1092) );
INVxp33_ASAP7_75t_SL g1006 ( .A(n_210), .Y(n_1006) );
INVx1_ASAP7_75t_L g731 ( .A(n_211), .Y(n_731) );
INVx1_ASAP7_75t_L g651 ( .A(n_212), .Y(n_651) );
INVx1_ASAP7_75t_L g664 ( .A(n_213), .Y(n_664) );
INVx1_ASAP7_75t_L g720 ( .A(n_215), .Y(n_720) );
INVx1_ASAP7_75t_L g510 ( .A(n_216), .Y(n_510) );
INVx1_ASAP7_75t_L g1114 ( .A(n_218), .Y(n_1114) );
NAND2xp5_ASAP7_75t_L g1119 ( .A(n_218), .B(n_1112), .Y(n_1119) );
INVx1_ASAP7_75t_L g867 ( .A(n_221), .Y(n_867) );
AO22x1_ASAP7_75t_L g1157 ( .A1(n_222), .A2(n_232), .B1(n_1125), .B2(n_1158), .Y(n_1157) );
INVx1_ASAP7_75t_L g547 ( .A(n_223), .Y(n_547) );
INVx2_ASAP7_75t_L g268 ( .A(n_224), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g658 ( .A(n_225), .Y(n_658) );
AOI21xp33_ASAP7_75t_L g578 ( .A1(n_227), .A2(n_413), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g608 ( .A(n_227), .Y(n_608) );
INVx1_ASAP7_75t_L g680 ( .A(n_228), .Y(n_680) );
INVx1_ASAP7_75t_L g770 ( .A(n_229), .Y(n_770) );
INVx1_ASAP7_75t_L g783 ( .A(n_230), .Y(n_783) );
INVx1_ASAP7_75t_L g862 ( .A(n_231), .Y(n_862) );
INVx1_ASAP7_75t_L g332 ( .A(n_233), .Y(n_332) );
INVx1_ASAP7_75t_L g513 ( .A(n_234), .Y(n_513) );
INVxp67_ASAP7_75t_L g1348 ( .A(n_235), .Y(n_1348) );
INVx1_ASAP7_75t_L g1095 ( .A(n_236), .Y(n_1095) );
INVx1_ASAP7_75t_L g1078 ( .A(n_237), .Y(n_1078) );
AOI21xp33_ASAP7_75t_L g355 ( .A1(n_238), .A2(n_305), .B(n_356), .Y(n_355) );
OAI211xp5_ASAP7_75t_SL g777 ( .A1(n_241), .A2(n_778), .B(n_779), .C(n_782), .Y(n_777) );
BUFx3_ASAP7_75t_L g376 ( .A(n_242), .Y(n_376) );
INVx1_ASAP7_75t_L g401 ( .A(n_242), .Y(n_401) );
BUFx3_ASAP7_75t_L g378 ( .A(n_243), .Y(n_378) );
INVx1_ASAP7_75t_L g397 ( .A(n_243), .Y(n_397) );
INVx1_ASAP7_75t_L g617 ( .A(n_244), .Y(n_617) );
INVx1_ASAP7_75t_L g672 ( .A(n_245), .Y(n_672) );
INVx1_ASAP7_75t_L g708 ( .A(n_246), .Y(n_708) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_272), .B(n_1100), .Y(n_249) );
BUFx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
INVx3_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
INVx1_ASAP7_75t_SL g252 ( .A(n_253), .Y(n_252) );
AND2x4_ASAP7_75t_L g253 ( .A(n_254), .B(n_259), .Y(n_253) );
AND2x4_ASAP7_75t_L g1375 ( .A(n_254), .B(n_260), .Y(n_1375) );
NOR2xp33_ASAP7_75t_SL g254 ( .A(n_255), .B(n_257), .Y(n_254) );
INVx1_ASAP7_75t_SL g1380 ( .A(n_255), .Y(n_1380) );
NAND2xp5_ASAP7_75t_L g1437 ( .A(n_255), .B(n_257), .Y(n_1437) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g1379 ( .A(n_257), .B(n_1380), .Y(n_1379) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_261), .B(n_265), .Y(n_260) );
INVxp67_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x2_ASAP7_75t_L g793 ( .A(n_263), .B(n_271), .Y(n_793) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g356 ( .A(n_264), .B(n_357), .Y(n_356) );
OR2x6_ASAP7_75t_L g265 ( .A(n_266), .B(n_270), .Y(n_265) );
OR2x2_ASAP7_75t_L g504 ( .A(n_266), .B(n_505), .Y(n_504) );
BUFx2_ASAP7_75t_L g536 ( .A(n_266), .Y(n_536) );
BUFx6f_ASAP7_75t_L g697 ( .A(n_266), .Y(n_697) );
INVx2_ASAP7_75t_SL g744 ( .A(n_266), .Y(n_744) );
INVx1_ASAP7_75t_L g882 ( .A(n_266), .Y(n_882) );
OAI22xp33_ASAP7_75t_L g956 ( .A1(n_266), .A2(n_539), .B1(n_957), .B2(n_958), .Y(n_956) );
OAI22xp33_ASAP7_75t_L g968 ( .A1(n_266), .A2(n_539), .B1(n_969), .B2(n_970), .Y(n_968) );
INVx2_ASAP7_75t_SL g1363 ( .A(n_266), .Y(n_1363) );
BUFx6f_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
INVx1_ASAP7_75t_L g289 ( .A(n_268), .Y(n_289) );
INVx2_ASAP7_75t_L g296 ( .A(n_268), .Y(n_296) );
AND2x4_ASAP7_75t_L g303 ( .A(n_268), .B(n_290), .Y(n_303) );
AND2x2_ASAP7_75t_L g309 ( .A(n_268), .B(n_269), .Y(n_309) );
INVx1_ASAP7_75t_L g353 ( .A(n_268), .Y(n_353) );
INVx2_ASAP7_75t_L g290 ( .A(n_269), .Y(n_290) );
INVx1_ASAP7_75t_L g298 ( .A(n_269), .Y(n_298) );
INVx1_ASAP7_75t_L g322 ( .A(n_269), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_269), .B(n_296), .Y(n_344) );
INVx1_ASAP7_75t_L g352 ( .A(n_269), .Y(n_352) );
INVx2_ASAP7_75t_SL g270 ( .A(n_271), .Y(n_270) );
OAI22xp33_ASAP7_75t_L g272 ( .A1(n_273), .A2(n_274), .B1(n_825), .B2(n_826), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AOI22xp5_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_276), .B1(n_562), .B2(n_824), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AOI22xp5_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_458), .B1(n_560), .B2(n_561), .Y(n_276) );
INVx1_ASAP7_75t_L g560 ( .A(n_277), .Y(n_560) );
NAND4xp25_ASAP7_75t_L g278 ( .A(n_279), .B(n_363), .C(n_384), .D(n_441), .Y(n_278) );
OAI21xp5_ASAP7_75t_SL g279 ( .A1(n_280), .A2(n_336), .B(n_360), .Y(n_279) );
INVx8_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x4_ASAP7_75t_L g282 ( .A(n_283), .B(n_287), .Y(n_282) );
AND2x4_ASAP7_75t_L g333 ( .A(n_283), .B(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g331 ( .A(n_285), .B(n_295), .Y(n_331) );
AND2x4_ASAP7_75t_L g338 ( .A(n_285), .B(n_339), .Y(n_338) );
AND2x4_ASAP7_75t_L g512 ( .A(n_285), .B(n_434), .Y(n_512) );
INVx1_ASAP7_75t_L g316 ( .A(n_286), .Y(n_316) );
INVx1_ASAP7_75t_L g357 ( .A(n_286), .Y(n_357) );
BUFx6f_ASAP7_75t_L g796 ( .A(n_287), .Y(n_796) );
BUFx3_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_288), .Y(n_312) );
BUFx3_ASAP7_75t_L g515 ( .A(n_288), .Y(n_515) );
BUFx6f_ASAP7_75t_L g735 ( .A(n_288), .Y(n_735) );
BUFx2_ASAP7_75t_L g815 ( .A(n_288), .Y(n_815) );
AND2x4_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_304), .B(n_318), .Y(n_291) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
BUFx6f_ASAP7_75t_L g521 ( .A(n_295), .Y(n_521) );
INVx1_ASAP7_75t_L g799 ( .A(n_295), .Y(n_799) );
BUFx6f_ASAP7_75t_L g955 ( .A(n_295), .Y(n_955) );
BUFx6f_ASAP7_75t_L g967 ( .A(n_295), .Y(n_967) );
AND2x4_ASAP7_75t_L g295 ( .A(n_296), .B(n_297), .Y(n_295) );
INVx1_ASAP7_75t_L g328 ( .A(n_296), .Y(n_328) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx2_ASAP7_75t_L g546 ( .A(n_301), .Y(n_546) );
INVx2_ASAP7_75t_L g551 ( .A(n_301), .Y(n_551) );
AND2x2_ASAP7_75t_L g732 ( .A(n_301), .B(n_512), .Y(n_732) );
INVx3_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx3_ASAP7_75t_L g347 ( .A(n_302), .Y(n_347) );
BUFx6f_ASAP7_75t_L g877 ( .A(n_302), .Y(n_877) );
INVx3_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g335 ( .A(n_303), .Y(n_335) );
BUFx6f_ASAP7_75t_L g865 ( .A(n_303), .Y(n_865) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x4_ASAP7_75t_L g518 ( .A(n_307), .B(n_512), .Y(n_518) );
BUFx2_ASAP7_75t_L g795 ( .A(n_307), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g963 ( .A1(n_307), .A2(n_815), .B1(n_964), .B2(n_965), .Y(n_963) );
BUFx3_ASAP7_75t_L g1016 ( .A(n_307), .Y(n_1016) );
INVx1_ASAP7_75t_L g1403 ( .A(n_307), .Y(n_1403) );
INVx2_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
INVx2_ASAP7_75t_SL g383 ( .A(n_308), .Y(n_383) );
INVx2_ASAP7_75t_L g1394 ( .A(n_308), .Y(n_1394) );
INVx3_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
BUFx6f_ASAP7_75t_L g339 ( .A(n_309), .Y(n_339) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx2_ASAP7_75t_SL g311 ( .A(n_312), .Y(n_311) );
BUFx2_ASAP7_75t_L g1404 ( .A(n_312), .Y(n_1404) );
INVx1_ASAP7_75t_L g884 ( .A(n_313), .Y(n_884) );
INVx2_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g807 ( .A(n_314), .B(n_361), .Y(n_807) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
OR2x6_ASAP7_75t_L g557 ( .A(n_315), .B(n_433), .Y(n_557) );
NAND2x1p5_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
NAND2x1p5_ASAP7_75t_L g319 ( .A(n_320), .B(n_323), .Y(n_319) );
NAND2x1_ASAP7_75t_SL g524 ( .A(n_320), .B(n_525), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g890 ( .A1(n_320), .A2(n_528), .B1(n_851), .B2(n_853), .Y(n_890) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
HB1xp67_ASAP7_75t_L g810 ( .A(n_322), .Y(n_810) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OR2x6_ASAP7_75t_L g327 ( .A(n_324), .B(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g358 ( .A(n_324), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g382 ( .A(n_324), .Y(n_382) );
AOI21xp33_ASAP7_75t_L g888 ( .A1(n_324), .A2(n_889), .B(n_890), .Y(n_888) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g528 ( .A(n_328), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_331), .B1(n_332), .B2(n_333), .Y(n_329) );
OAI22xp5_ASAP7_75t_L g415 ( .A1(n_330), .A2(n_332), .B1(n_416), .B2(n_419), .Y(n_415) );
INVx3_ASAP7_75t_L g892 ( .A(n_331), .Y(n_892) );
INVx3_ASAP7_75t_L g859 ( .A(n_333), .Y(n_859) );
INVx1_ASAP7_75t_L g803 ( .A(n_334), .Y(n_803) );
INVx2_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g616 ( .A(n_335), .Y(n_616) );
CKINVDCx6p67_ASAP7_75t_R g337 ( .A(n_338), .Y(n_337) );
INVx3_ASAP7_75t_L g806 ( .A(n_339), .Y(n_806) );
OAI22xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_345), .B1(n_346), .B2(n_348), .Y(n_340) );
OAI22xp5_ASAP7_75t_L g752 ( .A1(n_341), .A2(n_709), .B1(n_720), .B2(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g544 ( .A(n_343), .Y(n_544) );
INVx1_ASAP7_75t_L g907 ( .A(n_343), .Y(n_907) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g687 ( .A(n_344), .Y(n_687) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_345), .A2(n_348), .B1(n_395), .B2(n_398), .Y(n_394) );
OAI22xp5_ASAP7_75t_L g747 ( .A1(n_346), .A2(n_748), .B1(n_750), .B2(n_751), .Y(n_747) );
INVx1_ASAP7_75t_L g1400 ( .A(n_346), .Y(n_1400) );
INVx2_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
AND2x4_ASAP7_75t_L g511 ( .A(n_347), .B(n_512), .Y(n_511) );
BUFx3_ASAP7_75t_L g627 ( .A(n_347), .Y(n_627) );
INVx1_ASAP7_75t_SL g909 ( .A(n_347), .Y(n_909) );
INVx1_ASAP7_75t_L g1360 ( .A(n_347), .Y(n_1360) );
OAI21xp5_ASAP7_75t_SL g349 ( .A1(n_350), .A2(n_354), .B(n_355), .Y(n_349) );
OAI221xp5_ASAP7_75t_L g866 ( .A1(n_350), .A2(n_867), .B1(n_868), .B2(n_869), .C(n_870), .Y(n_866) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g359 ( .A(n_351), .Y(n_359) );
BUFx2_ASAP7_75t_L g624 ( .A(n_351), .Y(n_624) );
INVx3_ASAP7_75t_L g889 ( .A(n_351), .Y(n_889) );
AND2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_352), .B(n_353), .Y(n_540) );
INVx1_ASAP7_75t_L g813 ( .A(n_353), .Y(n_813) );
OR2x6_ASAP7_75t_L g532 ( .A(n_356), .B(n_362), .Y(n_532) );
INVx1_ASAP7_75t_L g554 ( .A(n_359), .Y(n_554) );
OAI22xp33_ASAP7_75t_L g1097 ( .A1(n_359), .A2(n_534), .B1(n_1069), .B2(n_1076), .Y(n_1097) );
CKINVDCx8_ASAP7_75t_R g599 ( .A(n_360), .Y(n_599) );
BUFx2_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx2_ASAP7_75t_L g380 ( .A(n_361), .Y(n_380) );
OR2x6_ASAP7_75t_L g403 ( .A(n_361), .B(n_404), .Y(n_403) );
AND2x4_ASAP7_75t_L g792 ( .A(n_361), .B(n_793), .Y(n_792) );
AND2x4_ASAP7_75t_L g1014 ( .A(n_361), .B(n_793), .Y(n_1014) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx2_ASAP7_75t_L g635 ( .A(n_362), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
OR2x6_ASAP7_75t_L g365 ( .A(n_366), .B(n_379), .Y(n_365) );
INVx2_ASAP7_75t_L g506 ( .A(n_366), .Y(n_506) );
AOI222xp33_ASAP7_75t_L g894 ( .A1(n_366), .A2(n_448), .B1(n_878), .B2(n_883), .C1(n_887), .C2(n_895), .Y(n_894) );
AND2x4_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
AND2x4_ASAP7_75t_L g422 ( .A(n_367), .B(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g991 ( .A(n_368), .Y(n_991) );
AND2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_374), .Y(n_368) );
NAND2x1p5_ASAP7_75t_L g432 ( .A(n_369), .B(n_433), .Y(n_432) );
AND2x4_ASAP7_75t_L g476 ( .A(n_369), .B(n_477), .Y(n_476) );
AND2x4_ASAP7_75t_L g479 ( .A(n_369), .B(n_437), .Y(n_479) );
BUFx2_ASAP7_75t_L g492 ( .A(n_369), .Y(n_492) );
AND2x4_ASAP7_75t_L g580 ( .A(n_369), .B(n_477), .Y(n_580) );
AND2x2_ASAP7_75t_L g652 ( .A(n_369), .B(n_437), .Y(n_652) );
INVx1_ASAP7_75t_L g1033 ( .A(n_369), .Y(n_1033) );
AND2x2_ASAP7_75t_L g1322 ( .A(n_369), .B(n_437), .Y(n_1322) );
AND2x4_ASAP7_75t_L g369 ( .A(n_370), .B(n_372), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AND2x4_ASAP7_75t_L g423 ( .A(n_372), .B(n_406), .Y(n_423) );
INVx2_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g405 ( .A(n_373), .B(n_406), .Y(n_405) );
INVx6_ASAP7_75t_L g393 ( .A(n_374), .Y(n_393) );
INVx2_ASAP7_75t_L g414 ( .A(n_374), .Y(n_414) );
BUFx2_ASAP7_75t_L g1074 ( .A(n_374), .Y(n_1074) );
AND2x4_ASAP7_75t_L g374 ( .A(n_375), .B(n_377), .Y(n_374) );
INVx1_ASAP7_75t_L g438 ( .A(n_375), .Y(n_438) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g390 ( .A(n_376), .B(n_378), .Y(n_390) );
AND2x4_ASAP7_75t_L g396 ( .A(n_376), .B(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g430 ( .A(n_377), .Y(n_430) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
AND2x4_ASAP7_75t_L g400 ( .A(n_378), .B(n_401), .Y(n_400) );
NOR2xp67_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g460 ( .A1(n_380), .A2(n_461), .B1(n_501), .B2(n_502), .Y(n_460) );
INVx2_ASAP7_75t_L g789 ( .A(n_380), .Y(n_789) );
INVx1_ASAP7_75t_L g886 ( .A(n_381), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
AND2x2_ASAP7_75t_L g905 ( .A(n_383), .B(n_512), .Y(n_905) );
AOI221xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_402), .B1(n_407), .B2(n_422), .C(n_424), .Y(n_384) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g840 ( .A(n_388), .Y(n_840) );
AND2x4_ASAP7_75t_L g1049 ( .A(n_388), .B(n_1050), .Y(n_1049) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g466 ( .A(n_389), .Y(n_466) );
BUFx6f_ASAP7_75t_L g640 ( .A(n_389), .Y(n_640) );
INVx1_ASAP7_75t_L g856 ( .A(n_389), .Y(n_856) );
BUFx6f_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
BUFx6f_ASAP7_75t_L g411 ( .A(n_390), .Y(n_411) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g464 ( .A(n_393), .Y(n_464) );
BUFx6f_ASAP7_75t_L g644 ( .A(n_393), .Y(n_644) );
INVx2_ASAP7_75t_L g937 ( .A(n_393), .Y(n_937) );
INVx2_ASAP7_75t_SL g1422 ( .A(n_393), .Y(n_1422) );
INVx2_ASAP7_75t_L g443 ( .A(n_395), .Y(n_443) );
INVx1_ASAP7_75t_L g980 ( .A(n_395), .Y(n_980) );
INVx2_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_396), .Y(n_418) );
BUFx2_ASAP7_75t_L g482 ( .A(n_396), .Y(n_482) );
BUFx3_ASAP7_75t_L g574 ( .A(n_396), .Y(n_574) );
BUFx6f_ASAP7_75t_L g586 ( .A(n_396), .Y(n_586) );
BUFx6f_ASAP7_75t_L g598 ( .A(n_396), .Y(n_598) );
BUFx6f_ASAP7_75t_L g641 ( .A(n_396), .Y(n_641) );
BUFx2_ASAP7_75t_L g655 ( .A(n_396), .Y(n_655) );
HB1xp67_ASAP7_75t_L g723 ( .A(n_396), .Y(n_723) );
INVx1_ASAP7_75t_L g457 ( .A(n_397), .Y(n_457) );
INVx1_ASAP7_75t_L g724 ( .A(n_398), .Y(n_724) );
INVx1_ASAP7_75t_L g986 ( .A(n_398), .Y(n_986) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g421 ( .A(n_399), .Y(n_421) );
BUFx6f_ASAP7_75t_L g645 ( .A(n_399), .Y(n_645) );
HB1xp67_ASAP7_75t_L g718 ( .A(n_399), .Y(n_718) );
INVx2_ASAP7_75t_L g845 ( .A(n_399), .Y(n_845) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g452 ( .A(n_400), .Y(n_452) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_400), .Y(n_470) );
INVx2_ASAP7_75t_L g488 ( .A(n_400), .Y(n_488) );
INVx1_ASAP7_75t_L g1325 ( .A(n_400), .Y(n_1325) );
INVx1_ASAP7_75t_L g456 ( .A(n_401), .Y(n_456) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
CKINVDCx5p33_ASAP7_75t_R g834 ( .A(n_403), .Y(n_834) );
INVx1_ASAP7_75t_L g589 ( .A(n_404), .Y(n_589) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx2_ASAP7_75t_SL g483 ( .A(n_405), .Y(n_483) );
BUFx3_ASAP7_75t_L g716 ( .A(n_405), .Y(n_716) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_410), .B(n_440), .Y(n_439) );
BUFx6f_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AND2x4_ASAP7_75t_L g489 ( .A(n_411), .B(n_472), .Y(n_489) );
AND2x4_ASAP7_75t_L g491 ( .A(n_411), .B(n_492), .Y(n_491) );
BUFx4f_ASAP7_75t_L g587 ( .A(n_411), .Y(n_587) );
AOI22xp5_ASAP7_75t_L g976 ( .A1(n_411), .A2(n_418), .B1(n_970), .B2(n_977), .Y(n_976) );
INVx2_ASAP7_75t_SL g982 ( .A(n_411), .Y(n_982) );
INVx1_ASAP7_75t_L g1072 ( .A(n_411), .Y(n_1072) );
BUFx3_ASAP7_75t_L g1337 ( .A(n_411), .Y(n_1337) );
BUFx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g448 ( .A(n_413), .B(n_444), .Y(n_448) );
A2O1A1Ixp33_ASAP7_75t_L g938 ( .A1(n_413), .A2(n_939), .B(n_940), .C(n_945), .Y(n_938) );
INVx2_ASAP7_75t_SL g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g1048 ( .A(n_414), .Y(n_1048) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
BUFx4f_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g471 ( .A(n_418), .B(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx4_ASAP7_75t_L g847 ( .A(n_422), .Y(n_847) );
INVx1_ASAP7_75t_L g467 ( .A(n_423), .Y(n_467) );
CKINVDCx5p33_ASAP7_75t_R g579 ( .A(n_423), .Y(n_579) );
INVx2_ASAP7_75t_SL g661 ( .A(n_423), .Y(n_661) );
HB1xp67_ASAP7_75t_L g1040 ( .A(n_423), .Y(n_1040) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g852 ( .A(n_427), .Y(n_852) );
NAND2x1p5_ASAP7_75t_L g427 ( .A(n_428), .B(n_431), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g477 ( .A(n_429), .Y(n_477) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_SL g431 ( .A(n_432), .Y(n_431) );
OR2x2_ASAP7_75t_L g435 ( .A(n_432), .B(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g440 ( .A(n_432), .Y(n_440) );
OR2x6_ASAP7_75t_L g850 ( .A(n_432), .B(n_436), .Y(n_850) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
OR2x2_ASAP7_75t_L g445 ( .A(n_434), .B(n_446), .Y(n_445) );
OR2x2_ASAP7_75t_L g1032 ( .A(n_436), .B(n_1033), .Y(n_1032) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AOI22xp5_ASAP7_75t_L g942 ( .A1(n_437), .A2(n_477), .B1(n_943), .B2(n_944), .Y(n_942) );
BUFx3_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g854 ( .A(n_440), .B(n_855), .Y(n_854) );
AOI221xp5_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_447), .B1(n_448), .B2(n_449), .C(n_450), .Y(n_441) );
AOI22xp5_ASAP7_75t_L g897 ( .A1(n_442), .A2(n_874), .B1(n_880), .B2(n_898), .Y(n_897) );
AND2x2_ASAP7_75t_L g442 ( .A(n_443), .B(n_444), .Y(n_442) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
OR2x2_ASAP7_75t_L g451 ( .A(n_445), .B(n_452), .Y(n_451) );
OR2x6_ASAP7_75t_L g453 ( .A(n_445), .B(n_454), .Y(n_453) );
OR2x6_ASAP7_75t_L g896 ( .A(n_445), .B(n_452), .Y(n_896) );
INVx2_ASAP7_75t_L g472 ( .A(n_446), .Y(n_472) );
OR2x2_ASAP7_75t_L g496 ( .A(n_446), .B(n_497), .Y(n_496) );
OR2x2_ASAP7_75t_L g500 ( .A(n_446), .B(n_488), .Y(n_500) );
INVx2_ASAP7_75t_L g575 ( .A(n_452), .Y(n_575) );
CKINVDCx6p67_ASAP7_75t_R g898 ( .A(n_453), .Y(n_898) );
OAI21xp33_ASAP7_75t_L g924 ( .A1(n_454), .A2(n_925), .B(n_926), .Y(n_924) );
OAI221xp5_ASAP7_75t_L g1038 ( .A1(n_454), .A2(n_1007), .B1(n_1009), .B2(n_1039), .C(n_1040), .Y(n_1038) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
BUFx4f_ASAP7_75t_L g774 ( .A(n_455), .Y(n_774) );
INVx1_ASAP7_75t_L g934 ( .A(n_455), .Y(n_934) );
INVx1_ASAP7_75t_L g941 ( .A(n_455), .Y(n_941) );
AND2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_457), .Y(n_455) );
OR2x2_ASAP7_75t_L g497 ( .A(n_456), .B(n_457), .Y(n_497) );
INVx3_ASAP7_75t_L g561 ( .A(n_458), .Y(n_561) );
INVx1_ASAP7_75t_L g558 ( .A(n_459), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_460), .B(n_507), .Y(n_459) );
NAND3xp33_ASAP7_75t_L g461 ( .A(n_462), .B(n_480), .C(n_493), .Y(n_461) );
AOI221xp5_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_468), .B1(n_471), .B2(n_473), .C(n_474), .Y(n_462) );
INVx3_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g577 ( .A(n_466), .Y(n_577) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g769 ( .A(n_470), .Y(n_769) );
BUFx3_ASAP7_75t_L g1037 ( .A(n_470), .Y(n_1037) );
AOI221xp5_ASAP7_75t_L g719 ( .A1(n_471), .A2(n_720), .B1(n_721), .B2(n_722), .C(n_725), .Y(n_719) );
INVx1_ASAP7_75t_L g778 ( .A(n_471), .Y(n_778) );
AND2x4_ASAP7_75t_L g597 ( .A(n_472), .B(n_598), .Y(n_597) );
AOI222xp33_ASAP7_75t_L g972 ( .A1(n_472), .A2(n_476), .B1(n_479), .B2(n_951), .C1(n_952), .C2(n_973), .Y(n_972) );
OAI22xp5_ASAP7_75t_L g548 ( .A1(n_473), .A2(n_498), .B1(n_543), .B2(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_SL g726 ( .A(n_476), .Y(n_726) );
AOI22xp5_ASAP7_75t_L g779 ( .A1(n_476), .A2(n_479), .B1(n_780), .B2(n_781), .Y(n_779) );
INVx4_ASAP7_75t_L g1418 ( .A(n_476), .Y(n_1418) );
INVx2_ASAP7_75t_SL g478 ( .A(n_479), .Y(n_478) );
AOI322xp5_ASAP7_75t_L g572 ( .A1(n_479), .A2(n_573), .A3(n_576), .B1(n_578), .B2(n_580), .C1(n_581), .C2(n_582), .Y(n_572) );
INVx2_ASAP7_75t_L g1066 ( .A(n_479), .Y(n_1066) );
AOI221xp5_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_484), .B1(n_489), .B2(n_490), .C(n_491), .Y(n_480) );
INVx1_ASAP7_75t_L g1046 ( .A(n_483), .Y(n_1046) );
INVx2_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g1064 ( .A(n_486), .Y(n_1064) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g591 ( .A(n_488), .Y(n_591) );
AOI221xp5_ASAP7_75t_L g583 ( .A1(n_489), .A2(n_491), .B1(n_584), .B2(n_585), .C(n_590), .Y(n_583) );
AOI221xp5_ASAP7_75t_L g637 ( .A1(n_489), .A2(n_491), .B1(n_638), .B2(n_639), .C(n_642), .Y(n_637) );
INVx2_ASAP7_75t_SL g712 ( .A(n_489), .Y(n_712) );
BUFx6f_ASAP7_75t_L g1042 ( .A(n_489), .Y(n_1042) );
HB1xp67_ASAP7_75t_L g1068 ( .A(n_489), .Y(n_1068) );
INVx1_ASAP7_75t_L g1334 ( .A(n_489), .Y(n_1334) );
HB1xp67_ASAP7_75t_L g1424 ( .A(n_489), .Y(n_1424) );
OAI22xp33_ASAP7_75t_L g552 ( .A1(n_490), .A2(n_494), .B1(n_534), .B2(n_553), .Y(n_552) );
AOI221xp5_ASAP7_75t_L g710 ( .A1(n_491), .A2(n_711), .B1(n_713), .B2(n_714), .C(n_717), .Y(n_710) );
INVx1_ASAP7_75t_L g776 ( .A(n_491), .Y(n_776) );
AOI21xp5_ASAP7_75t_L g978 ( .A1(n_491), .A2(n_979), .B(n_984), .Y(n_978) );
AOI221xp5_ASAP7_75t_L g1067 ( .A1(n_491), .A2(n_1068), .B1(n_1069), .B2(n_1070), .C(n_1073), .Y(n_1067) );
AOI221xp5_ASAP7_75t_L g1423 ( .A1(n_491), .A2(n_1424), .B1(n_1425), .B2(n_1426), .C(n_1427), .Y(n_1423) );
BUFx3_ASAP7_75t_L g945 ( .A(n_492), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_495), .B1(n_498), .B2(n_499), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_495), .A2(n_499), .B1(n_593), .B2(n_594), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_495), .A2(n_499), .B1(n_647), .B2(n_648), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g707 ( .A1(n_495), .A2(n_499), .B1(n_708), .B2(n_709), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g1051 ( .A1(n_495), .A2(n_499), .B1(n_1052), .B2(n_1053), .Y(n_1051) );
AOI22xp33_ASAP7_75t_L g1075 ( .A1(n_495), .A2(n_499), .B1(n_1076), .B2(n_1077), .Y(n_1075) );
AOI22xp33_ASAP7_75t_SL g1341 ( .A1(n_495), .A2(n_499), .B1(n_1342), .B2(n_1343), .Y(n_1341) );
AOI22xp33_ASAP7_75t_L g1428 ( .A1(n_495), .A2(n_499), .B1(n_1429), .B2(n_1430), .Y(n_1428) );
INVx6_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx2_ASAP7_75t_L g767 ( .A(n_497), .Y(n_767) );
INVx1_ASAP7_75t_L g930 ( .A(n_497), .Y(n_930) );
INVx1_ASAP7_75t_L g975 ( .A(n_497), .Y(n_975) );
INVx4_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AOI22xp5_ASAP7_75t_L g570 ( .A1(n_502), .A2(n_571), .B1(n_599), .B2(n_600), .Y(n_570) );
AOI22xp5_ASAP7_75t_L g705 ( .A1(n_502), .A2(n_599), .B1(n_706), .B2(n_727), .Y(n_705) );
INVx2_ASAP7_75t_SL g502 ( .A(n_503), .Y(n_502) );
INVx5_ASAP7_75t_L g665 ( .A(n_503), .Y(n_665) );
INVx2_ASAP7_75t_L g1079 ( .A(n_503), .Y(n_1079) );
AND2x4_ASAP7_75t_L g503 ( .A(n_504), .B(n_506), .Y(n_503) );
INVx2_ASAP7_75t_L g960 ( .A(n_504), .Y(n_960) );
INVx3_ASAP7_75t_L g525 ( .A(n_505), .Y(n_525) );
NOR3xp33_ASAP7_75t_L g507 ( .A(n_508), .B(n_522), .C(n_531), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_509), .B(n_516), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_511), .B1(n_513), .B2(n_514), .Y(n_509) );
BUFx2_ASAP7_75t_L g605 ( .A(n_511), .Y(n_605) );
BUFx2_ASAP7_75t_L g669 ( .A(n_511), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g1082 ( .A1(n_511), .A2(n_514), .B1(n_1083), .B2(n_1084), .Y(n_1082) );
BUFx2_ASAP7_75t_L g1369 ( .A(n_511), .Y(n_1369) );
AND2x6_ASAP7_75t_L g514 ( .A(n_512), .B(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g520 ( .A(n_512), .B(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g610 ( .A(n_512), .B(n_521), .Y(n_610) );
AND2x2_ASAP7_75t_L g673 ( .A(n_512), .B(n_521), .Y(n_673) );
AND2x2_ASAP7_75t_L g734 ( .A(n_512), .B(n_735), .Y(n_734) );
AOI22xp5_ASAP7_75t_L g961 ( .A1(n_512), .A2(n_807), .B1(n_962), .B2(n_966), .Y(n_961) );
AND2x2_ASAP7_75t_L g1411 ( .A(n_512), .B(n_521), .Y(n_1411) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_514), .A2(n_604), .B1(n_605), .B2(n_606), .Y(n_603) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_514), .A2(n_658), .B1(n_669), .B2(n_670), .Y(n_668) );
AOI22xp33_ASAP7_75t_L g1005 ( .A1(n_514), .A2(n_669), .B1(n_1006), .B2(n_1007), .Y(n_1005) );
AOI22xp33_ASAP7_75t_L g1367 ( .A1(n_514), .A2(n_1329), .B1(n_1368), .B2(n_1369), .Y(n_1367) );
AOI22xp33_ASAP7_75t_L g1405 ( .A1(n_514), .A2(n_1369), .B1(n_1406), .B2(n_1407), .Y(n_1405) );
NAND2x1p5_ASAP7_75t_L g530 ( .A(n_515), .B(n_525), .Y(n_530) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_518), .B1(n_519), .B2(n_520), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_518), .A2(n_608), .B1(n_609), .B2(n_610), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_518), .A2(n_656), .B1(n_672), .B2(n_673), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_518), .A2(n_610), .B1(n_737), .B2(n_738), .Y(n_736) );
AOI221xp5_ASAP7_75t_L g816 ( .A1(n_518), .A2(n_673), .B1(n_817), .B2(n_818), .C(n_819), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g1008 ( .A1(n_518), .A2(n_520), .B1(n_1009), .B2(n_1010), .Y(n_1008) );
AOI22xp33_ASAP7_75t_L g1085 ( .A1(n_518), .A2(n_520), .B1(n_1086), .B2(n_1087), .Y(n_1085) );
AOI22xp33_ASAP7_75t_L g1370 ( .A1(n_518), .A2(n_673), .B1(n_1330), .B2(n_1371), .Y(n_1370) );
AOI22xp33_ASAP7_75t_L g1408 ( .A1(n_518), .A2(n_1409), .B1(n_1410), .B2(n_1411), .Y(n_1408) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g676 ( .A(n_524), .Y(n_676) );
NAND2x1p5_ASAP7_75t_L g527 ( .A(n_525), .B(n_528), .Y(n_527) );
AND2x4_ASAP7_75t_L g809 ( .A(n_525), .B(n_810), .Y(n_809) );
AND2x4_ASAP7_75t_L g811 ( .A(n_525), .B(n_812), .Y(n_811) );
AND2x4_ASAP7_75t_L g814 ( .A(n_525), .B(n_815), .Y(n_814) );
BUFx4f_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
BUFx3_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
BUFx2_ASAP7_75t_L g677 ( .A(n_530), .Y(n_677) );
OAI33xp33_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_533), .A3(n_542), .B1(n_548), .B2(n_552), .B3(n_555), .Y(n_531) );
OAI33xp33_ASAP7_75t_L g612 ( .A1(n_532), .A2(n_555), .A3(n_613), .B1(n_618), .B2(n_622), .B3(n_625), .Y(n_612) );
OAI33xp33_ASAP7_75t_L g678 ( .A1(n_532), .A2(n_555), .A3(n_679), .B1(n_683), .B2(n_692), .B3(n_694), .Y(n_678) );
OAI33xp33_ASAP7_75t_L g741 ( .A1(n_532), .A2(n_742), .A3(n_747), .B1(n_752), .B2(n_754), .B3(n_756), .Y(n_741) );
OAI33xp33_ASAP7_75t_L g1089 ( .A1(n_532), .A2(n_557), .A3(n_1090), .B1(n_1093), .B2(n_1096), .B3(n_1097), .Y(n_1089) );
OAI33xp33_ASAP7_75t_L g1346 ( .A1(n_532), .A2(n_555), .A3(n_1347), .B1(n_1352), .B2(n_1358), .B3(n_1361), .Y(n_1346) );
OAI22xp33_ASAP7_75t_L g533 ( .A1(n_534), .A2(n_537), .B1(n_538), .B2(n_541), .Y(n_533) );
OAI22xp33_ASAP7_75t_L g622 ( .A1(n_534), .A2(n_584), .B1(n_593), .B2(n_623), .Y(n_622) );
OAI22xp33_ASAP7_75t_L g679 ( .A1(n_534), .A2(n_680), .B1(n_681), .B2(n_682), .Y(n_679) );
OAI22xp33_ASAP7_75t_L g1090 ( .A1(n_534), .A2(n_698), .B1(n_1091), .B2(n_1092), .Y(n_1090) );
INVx2_ASAP7_75t_SL g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g619 ( .A(n_535), .Y(n_619) );
INVx1_ASAP7_75t_L g868 ( .A(n_535), .Y(n_868) );
INVx2_ASAP7_75t_SL g535 ( .A(n_536), .Y(n_535) );
OAI22xp33_ASAP7_75t_L g618 ( .A1(n_538), .A2(n_619), .B1(n_620), .B2(n_621), .Y(n_618) );
BUFx3_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx2_ASAP7_75t_L g699 ( .A(n_539), .Y(n_699) );
BUFx3_ASAP7_75t_L g755 ( .A(n_539), .Y(n_755) );
OAI221xp5_ASAP7_75t_L g879 ( .A1(n_539), .A2(n_880), .B1(n_881), .B2(n_883), .C(n_884), .Y(n_879) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
OAI22xp5_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_545), .B1(n_546), .B2(n_547), .Y(n_542) );
OAI22xp5_ASAP7_75t_L g613 ( .A1(n_543), .A2(n_614), .B1(n_615), .B2(n_617), .Y(n_613) );
OAI22xp5_ASAP7_75t_L g625 ( .A1(n_543), .A2(n_594), .B1(n_596), .B2(n_626), .Y(n_625) );
BUFx2_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_SL g690 ( .A(n_546), .Y(n_690) );
OAI22xp5_ASAP7_75t_L g692 ( .A1(n_546), .A2(n_648), .B1(n_663), .B2(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g800 ( .A(n_551), .Y(n_800) );
OAI22xp33_ASAP7_75t_L g742 ( .A1(n_553), .A2(n_743), .B1(n_745), .B2(n_746), .Y(n_742) );
INVx1_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
CKINVDCx8_ASAP7_75t_R g555 ( .A(n_556), .Y(n_555) );
INVx5_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx6_ASAP7_75t_L g757 ( .A(n_557), .Y(n_757) );
OAI22xp5_ASAP7_75t_L g1133 ( .A1(n_559), .A2(n_1134), .B1(n_1136), .B2(n_1137), .Y(n_1133) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
HB1xp67_ASAP7_75t_L g824 ( .A(n_563), .Y(n_824) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_565), .B1(n_701), .B2(n_702), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AOI22xp5_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_567), .B1(n_628), .B2(n_629), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
XNOR2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_601), .Y(n_569) );
NAND4xp25_ASAP7_75t_L g571 ( .A(n_572), .B(n_583), .C(n_592), .D(n_595), .Y(n_571) );
BUFx2_ASAP7_75t_L g837 ( .A(n_575), .Y(n_837) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_580), .A2(n_650), .B1(n_651), .B2(n_652), .Y(n_649) );
INVx2_ASAP7_75t_L g1031 ( .A(n_580), .Y(n_1031) );
INVx1_ASAP7_75t_L g1320 ( .A(n_580), .Y(n_1320) );
INVx2_ASAP7_75t_L g1327 ( .A(n_586), .Y(n_1327) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g931 ( .A(n_591), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_597), .B(n_663), .Y(n_662) );
AOI211xp5_ASAP7_75t_L g1028 ( .A1(n_597), .A2(n_1029), .B(n_1030), .C(n_1034), .Y(n_1028) );
AOI221xp5_ASAP7_75t_L g1060 ( .A1(n_597), .A2(n_1061), .B1(n_1062), .B2(n_1063), .C(n_1065), .Y(n_1060) );
AOI211xp5_ASAP7_75t_L g1317 ( .A1(n_597), .A2(n_1318), .B(n_1319), .C(n_1323), .Y(n_1317) );
NOR3xp33_ASAP7_75t_SL g601 ( .A(n_602), .B(n_611), .C(n_612), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_607), .Y(n_602) );
INVx1_ASAP7_75t_L g918 ( .A(n_610), .Y(n_918) );
OAI22xp5_ASAP7_75t_L g1093 ( .A1(n_615), .A2(n_684), .B1(n_1094), .B2(n_1095), .Y(n_1093) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g753 ( .A(n_616), .Y(n_753) );
HB1xp67_ASAP7_75t_L g1398 ( .A(n_616), .Y(n_1398) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g681 ( .A(n_624), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g1096 ( .A1(n_626), .A2(n_693), .B1(n_1061), .B2(n_1077), .Y(n_1096) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
CKINVDCx5p33_ASAP7_75t_R g1351 ( .A(n_627), .Y(n_1351) );
INVx2_ASAP7_75t_SL g628 ( .A(n_629), .Y(n_628) );
XNOR2x1_ASAP7_75t_L g629 ( .A(n_630), .B(n_700), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_666), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_636), .B1(n_664), .B2(n_665), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g1058 ( .A1(n_632), .A2(n_1059), .B1(n_1078), .B2(n_1079), .Y(n_1058) );
AOI22xp5_ASAP7_75t_L g1412 ( .A1(n_632), .A2(n_1079), .B1(n_1413), .B2(n_1431), .Y(n_1412) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AOI31xp33_ASAP7_75t_L g1027 ( .A1(n_633), .A2(n_1028), .A3(n_1041), .B(n_1051), .Y(n_1027) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
BUFx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx2_ASAP7_75t_L g893 ( .A(n_635), .Y(n_893) );
NAND5xp2_ASAP7_75t_L g636 ( .A(n_637), .B(n_646), .C(n_649), .D(n_653), .E(n_662), .Y(n_636) );
OAI22xp33_ASAP7_75t_L g694 ( .A1(n_638), .A2(n_647), .B1(n_695), .B2(n_698), .Y(n_694) );
BUFx2_ASAP7_75t_L g836 ( .A(n_641), .Y(n_836) );
BUFx3_ASAP7_75t_L g843 ( .A(n_641), .Y(n_843) );
INVx1_ASAP7_75t_L g1036 ( .A(n_641), .Y(n_1036) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g660 ( .A(n_644), .Y(n_660) );
INVx1_ASAP7_75t_L g657 ( .A(n_645), .Y(n_657) );
OAI221xp5_ASAP7_75t_SL g653 ( .A1(n_654), .A2(n_656), .B1(n_657), .B2(n_658), .C(n_659), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g1331 ( .A(n_661), .Y(n_1331) );
AOI21xp5_ASAP7_75t_L g1025 ( .A1(n_665), .A2(n_1026), .B(n_1027), .Y(n_1025) );
AOI21xp33_ASAP7_75t_L g1314 ( .A1(n_665), .A2(n_1315), .B(n_1316), .Y(n_1314) );
NOR3xp33_ASAP7_75t_L g666 ( .A(n_667), .B(n_674), .C(n_678), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_668), .B(n_671), .Y(n_667) );
INVx2_ASAP7_75t_SL g675 ( .A(n_676), .Y(n_675) );
INVx2_ASAP7_75t_L g740 ( .A(n_676), .Y(n_740) );
OAI22xp5_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_688), .B1(n_689), .B2(n_691), .Y(n_683) );
INVx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g693 ( .A(n_685), .Y(n_693) );
INVx2_ASAP7_75t_L g1349 ( .A(n_685), .Y(n_1349) );
INVx2_ASAP7_75t_L g1359 ( .A(n_685), .Y(n_1359) );
INVx2_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
BUFx3_ASAP7_75t_L g749 ( .A(n_687), .Y(n_749) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
OAI22xp33_ASAP7_75t_L g754 ( .A1(n_697), .A2(n_708), .B1(n_713), .B2(n_755), .Y(n_754) );
BUFx2_ASAP7_75t_L g1354 ( .A(n_697), .Y(n_1354) );
INVx2_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx2_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
XOR2x2_ASAP7_75t_L g702 ( .A(n_703), .B(n_760), .Y(n_702) );
INVx1_ASAP7_75t_L g758 ( .A(n_704), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_705), .B(n_728), .Y(n_704) );
NAND3xp33_ASAP7_75t_L g706 ( .A(n_707), .B(n_710), .C(n_719), .Y(n_706) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx3_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVxp67_ASAP7_75t_L g983 ( .A(n_716), .Y(n_983) );
NOR3xp33_ASAP7_75t_L g728 ( .A(n_729), .B(n_739), .C(n_741), .Y(n_728) );
NAND2xp5_ASAP7_75t_SL g729 ( .A(n_730), .B(n_736), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_732), .B1(n_733), .B2(n_734), .Y(n_730) );
INVx2_ASAP7_75t_L g820 ( .A(n_732), .Y(n_820) );
INVx1_ASAP7_75t_L g821 ( .A(n_734), .Y(n_821) );
INVx2_ASAP7_75t_SL g1018 ( .A(n_735), .Y(n_1018) );
BUFx6f_ASAP7_75t_L g1395 ( .A(n_735), .Y(n_1395) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
OAI22xp5_ASAP7_75t_L g861 ( .A1(n_748), .A2(n_862), .B1(n_863), .B2(n_864), .Y(n_861) );
INVx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx2_ASAP7_75t_SL g873 ( .A(n_749), .Y(n_873) );
INVx2_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
AOI33xp33_ASAP7_75t_L g1011 ( .A1(n_757), .A2(n_1012), .A3(n_1015), .B1(n_1019), .B2(n_1023), .B3(n_1024), .Y(n_1011) );
AOI33xp33_ASAP7_75t_L g1391 ( .A1(n_757), .A2(n_1392), .A3(n_1393), .B1(n_1396), .B2(n_1399), .B3(n_1401), .Y(n_1391) );
OAI22xp33_ASAP7_75t_L g1139 ( .A1(n_759), .A2(n_1134), .B1(n_1137), .B2(n_1140), .Y(n_1139) );
INVx1_ASAP7_75t_L g823 ( .A(n_761), .Y(n_823) );
NAND4xp75_ASAP7_75t_L g761 ( .A(n_762), .B(n_763), .C(n_790), .D(n_816), .Y(n_761) );
OAI31xp33_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_777), .A3(n_787), .B(n_788), .Y(n_763) );
OAI22xp5_ASAP7_75t_L g765 ( .A1(n_766), .A2(n_768), .B1(n_769), .B2(n_770), .Y(n_765) );
INVx2_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx2_ASAP7_75t_L g1039 ( .A(n_767), .Y(n_1039) );
OAI21xp33_ASAP7_75t_L g771 ( .A1(n_772), .A2(n_773), .B(n_775), .Y(n_771) );
INVx2_ASAP7_75t_SL g773 ( .A(n_774), .Y(n_773) );
INVx1_ASAP7_75t_L g784 ( .A(n_774), .Y(n_784) );
INVx1_ASAP7_75t_L g1415 ( .A(n_778), .Y(n_1415) );
AOI221xp5_ASAP7_75t_L g808 ( .A1(n_780), .A2(n_781), .B1(n_809), .B2(n_811), .C(n_814), .Y(n_808) );
OAI211xp5_ASAP7_75t_L g782 ( .A1(n_783), .A2(n_784), .B(n_785), .C(n_786), .Y(n_782) );
INVx1_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
AOI31xp33_ASAP7_75t_SL g971 ( .A1(n_789), .A2(n_972), .A3(n_978), .B(n_987), .Y(n_971) );
AND2x2_ASAP7_75t_SL g790 ( .A(n_791), .B(n_808), .Y(n_790) );
AOI33xp33_ASAP7_75t_L g791 ( .A1(n_792), .A2(n_794), .A3(n_797), .B1(n_801), .B2(n_804), .B3(n_807), .Y(n_791) );
AOI22xp5_ASAP7_75t_L g953 ( .A1(n_792), .A2(n_954), .B1(n_959), .B2(n_960), .Y(n_953) );
BUFx2_ASAP7_75t_L g1392 ( .A(n_792), .Y(n_1392) );
INVx1_ASAP7_75t_L g871 ( .A(n_793), .Y(n_871) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g1397 ( .A(n_799), .Y(n_1397) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
INVx2_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
NAND3xp33_ASAP7_75t_L g912 ( .A(n_807), .B(n_913), .C(n_914), .Y(n_912) );
AOI221xp5_ASAP7_75t_L g950 ( .A1(n_809), .A2(n_811), .B1(n_814), .B2(n_951), .C(n_952), .Y(n_950) );
INVx1_ASAP7_75t_L g1003 ( .A(n_809), .Y(n_1003) );
AOI221xp5_ASAP7_75t_L g1388 ( .A1(n_809), .A2(n_811), .B1(n_814), .B2(n_1389), .C(n_1390), .Y(n_1388) );
HB1xp67_ASAP7_75t_L g1000 ( .A(n_811), .Y(n_1000) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
AOI221xp5_ASAP7_75t_L g999 ( .A1(n_814), .A2(n_1000), .B1(n_1001), .B2(n_1002), .C(n_1004), .Y(n_999) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
AOI22xp5_ASAP7_75t_L g826 ( .A1(n_827), .A2(n_828), .B1(n_1056), .B2(n_1099), .Y(n_826) );
INVxp67_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
AO22x2_ASAP7_75t_L g828 ( .A1(n_829), .A2(n_996), .B1(n_1054), .B2(n_1055), .Y(n_828) );
INVx1_ASAP7_75t_L g1054 ( .A(n_829), .Y(n_1054) );
XNOR2xp5_ASAP7_75t_L g829 ( .A(n_830), .B(n_899), .Y(n_829) );
NAND4xp75_ASAP7_75t_L g831 ( .A(n_832), .B(n_857), .C(n_894), .D(n_897), .Y(n_831) );
AND2x2_ASAP7_75t_SL g832 ( .A(n_833), .B(n_848), .Y(n_832) );
AOI33xp33_ASAP7_75t_L g833 ( .A1(n_834), .A2(n_835), .A3(n_838), .B1(n_841), .B2(n_842), .B3(n_846), .Y(n_833) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx1_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
AOI221xp5_ASAP7_75t_L g848 ( .A1(n_849), .A2(n_851), .B1(n_852), .B2(n_853), .C(n_854), .Y(n_848) );
INVx2_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
OAI31xp33_ASAP7_75t_L g857 ( .A1(n_858), .A2(n_860), .A3(n_891), .B(n_893), .Y(n_857) );
OAI221xp5_ASAP7_75t_L g860 ( .A1(n_861), .A2(n_866), .B1(n_872), .B2(n_879), .C(n_885), .Y(n_860) );
INVx2_ASAP7_75t_SL g864 ( .A(n_865), .Y(n_864) );
INVx2_ASAP7_75t_SL g1022 ( .A(n_865), .Y(n_1022) );
INVx2_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
OAI22xp5_ASAP7_75t_L g872 ( .A1(n_873), .A2(n_874), .B1(n_875), .B2(n_878), .Y(n_872) );
INVx1_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
INVx2_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
INVx2_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
AOI21xp5_ASAP7_75t_L g885 ( .A1(n_886), .A2(n_887), .B(n_888), .Y(n_885) );
INVx1_ASAP7_75t_L g1357 ( .A(n_889), .Y(n_1357) );
BUFx2_ASAP7_75t_L g1364 ( .A(n_889), .Y(n_1364) );
INVx2_ASAP7_75t_L g946 ( .A(n_893), .Y(n_946) );
BUFx8_ASAP7_75t_SL g1344 ( .A(n_893), .Y(n_1344) );
CKINVDCx6p67_ASAP7_75t_R g895 ( .A(n_896), .Y(n_895) );
XNOR2xp5_ASAP7_75t_L g899 ( .A(n_900), .B(n_947), .Y(n_899) );
NAND3xp33_ASAP7_75t_L g901 ( .A(n_902), .B(n_916), .C(n_920), .Y(n_901) );
NOR2xp33_ASAP7_75t_L g902 ( .A(n_903), .B(n_915), .Y(n_902) );
INVx1_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
OAI221xp5_ASAP7_75t_L g906 ( .A1(n_907), .A2(n_908), .B1(n_909), .B2(n_910), .C(n_911), .Y(n_906) );
OAI22xp5_ASAP7_75t_L g927 ( .A1(n_910), .A2(n_928), .B1(n_929), .B2(n_931), .Y(n_927) );
NOR2xp33_ASAP7_75t_SL g916 ( .A(n_917), .B(n_919), .Y(n_916) );
OAI31xp33_ASAP7_75t_SL g920 ( .A1(n_921), .A2(n_922), .A3(n_923), .B(n_946), .Y(n_920) );
OAI211xp5_ASAP7_75t_SL g923 ( .A1(n_924), .A2(n_927), .B(n_932), .C(n_938), .Y(n_923) );
OAI221xp5_ASAP7_75t_L g1328 ( .A1(n_929), .A2(n_934), .B1(n_1329), .B2(n_1330), .C(n_1331), .Y(n_1328) );
INVx2_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
OAI211xp5_ASAP7_75t_L g932 ( .A1(n_933), .A2(n_934), .B(n_935), .C(n_936), .Y(n_932) );
OAI211xp5_ASAP7_75t_L g1419 ( .A1(n_934), .A2(n_1407), .B(n_1420), .C(n_1421), .Y(n_1419) );
BUFx6f_ASAP7_75t_L g985 ( .A(n_937), .Y(n_985) );
INVx1_ASAP7_75t_L g1340 ( .A(n_937), .Y(n_1340) );
NAND2xp33_ASAP7_75t_L g940 ( .A(n_941), .B(n_942), .Y(n_940) );
NAND2xp5_ASAP7_75t_SL g947 ( .A(n_948), .B(n_992), .Y(n_947) );
INVx1_ASAP7_75t_L g994 ( .A(n_949), .Y(n_994) );
NAND3xp33_ASAP7_75t_SL g949 ( .A(n_950), .B(n_953), .C(n_961), .Y(n_949) );
AOI22xp5_ASAP7_75t_L g987 ( .A1(n_959), .A2(n_988), .B1(n_989), .B2(n_990), .Y(n_987) );
BUFx3_ASAP7_75t_L g1020 ( .A(n_967), .Y(n_1020) );
INVx1_ASAP7_75t_L g993 ( .A(n_971), .Y(n_993) );
INVx2_ASAP7_75t_L g974 ( .A(n_975), .Y(n_974) );
INVx1_ASAP7_75t_L g981 ( .A(n_982), .Y(n_981) );
INVx2_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
NAND3xp33_ASAP7_75t_L g992 ( .A(n_993), .B(n_994), .C(n_995), .Y(n_992) );
INVx2_ASAP7_75t_L g1055 ( .A(n_996), .Y(n_1055) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_998), .B(n_1025), .Y(n_997) );
AND4x1_ASAP7_75t_L g998 ( .A(n_999), .B(n_1005), .C(n_1008), .D(n_1011), .Y(n_998) );
INVx1_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
INVx2_ASAP7_75t_L g1012 ( .A(n_1013), .Y(n_1012) );
INVx2_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
INVx2_ASAP7_75t_L g1017 ( .A(n_1018), .Y(n_1017) );
INVx1_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
INVx1_ASAP7_75t_SL g1050 ( .A(n_1033), .Y(n_1050) );
INVx1_ASAP7_75t_L g1035 ( .A(n_1036), .Y(n_1035) );
AOI221xp5_ASAP7_75t_L g1041 ( .A1(n_1042), .A2(n_1043), .B1(n_1044), .B2(n_1047), .C(n_1049), .Y(n_1041) );
INVx1_ASAP7_75t_L g1045 ( .A(n_1046), .Y(n_1045) );
AOI221xp5_ASAP7_75t_L g1332 ( .A1(n_1049), .A2(n_1333), .B1(n_1335), .B2(n_1336), .C(n_1338), .Y(n_1332) );
INVx2_ASAP7_75t_L g1099 ( .A(n_1056), .Y(n_1099) );
XOR2x2_ASAP7_75t_L g1056 ( .A(n_1057), .B(n_1098), .Y(n_1056) );
NAND2xp5_ASAP7_75t_L g1057 ( .A(n_1058), .B(n_1080), .Y(n_1057) );
NAND3xp33_ASAP7_75t_L g1059 ( .A(n_1060), .B(n_1067), .C(n_1075), .Y(n_1059) );
INVx1_ASAP7_75t_L g1071 ( .A(n_1072), .Y(n_1071) );
NOR3xp33_ASAP7_75t_L g1080 ( .A(n_1081), .B(n_1088), .C(n_1089), .Y(n_1080) );
NAND2xp5_ASAP7_75t_L g1081 ( .A(n_1082), .B(n_1085), .Y(n_1081) );
OAI221xp5_ASAP7_75t_L g1100 ( .A1(n_1101), .A2(n_1308), .B1(n_1310), .B2(n_1372), .C(n_1376), .Y(n_1100) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_1102), .B(n_1235), .Y(n_1101) );
NOR2xp33_ASAP7_75t_L g1102 ( .A(n_1103), .B(n_1217), .Y(n_1102) );
NAND3xp33_ASAP7_75t_L g1103 ( .A(n_1104), .B(n_1174), .C(n_1203), .Y(n_1103) );
O2A1O1Ixp33_ASAP7_75t_L g1104 ( .A1(n_1105), .A2(n_1141), .B(n_1146), .C(n_1160), .Y(n_1104) );
AND2x2_ASAP7_75t_L g1105 ( .A(n_1106), .B(n_1126), .Y(n_1105) );
AND2x2_ASAP7_75t_L g1162 ( .A(n_1106), .B(n_1163), .Y(n_1162) );
AND2x2_ASAP7_75t_L g1183 ( .A(n_1106), .B(n_1184), .Y(n_1183) );
NOR2xp33_ASAP7_75t_L g1201 ( .A(n_1106), .B(n_1147), .Y(n_1201) );
AND2x2_ASAP7_75t_L g1206 ( .A(n_1106), .B(n_1127), .Y(n_1206) );
AND2x2_ASAP7_75t_L g1216 ( .A(n_1106), .B(n_1202), .Y(n_1216) );
OAI332xp33_ASAP7_75t_L g1239 ( .A1(n_1106), .A2(n_1171), .A3(n_1190), .B1(n_1191), .B2(n_1240), .B3(n_1243), .C1(n_1244), .C2(n_1246), .Y(n_1239) );
OAI32xp33_ASAP7_75t_L g1301 ( .A1(n_1106), .A2(n_1232), .A3(n_1257), .B1(n_1287), .B2(n_1302), .Y(n_1301) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1106), .Y(n_1303) );
INVx4_ASAP7_75t_L g1106 ( .A(n_1107), .Y(n_1106) );
NAND2xp5_ASAP7_75t_L g1143 ( .A(n_1107), .B(n_1144), .Y(n_1143) );
NAND2xp5_ASAP7_75t_L g1171 ( .A(n_1107), .B(n_1163), .Y(n_1171) );
INVx3_ASAP7_75t_L g1189 ( .A(n_1107), .Y(n_1189) );
AND2x2_ASAP7_75t_L g1197 ( .A(n_1107), .B(n_1191), .Y(n_1197) );
AND2x2_ASAP7_75t_L g1226 ( .A(n_1107), .B(n_1211), .Y(n_1226) );
OR2x2_ASAP7_75t_L g1255 ( .A(n_1107), .B(n_1163), .Y(n_1255) );
NOR2xp33_ASAP7_75t_L g1298 ( .A(n_1107), .B(n_1242), .Y(n_1298) );
NAND3xp33_ASAP7_75t_L g1305 ( .A(n_1107), .B(n_1288), .C(n_1299), .Y(n_1305) );
NOR3xp33_ASAP7_75t_L g1306 ( .A(n_1107), .B(n_1185), .C(n_1307), .Y(n_1306) );
AND2x4_ASAP7_75t_L g1107 ( .A(n_1108), .B(n_1120), .Y(n_1107) );
AND2x4_ASAP7_75t_L g1109 ( .A(n_1110), .B(n_1115), .Y(n_1109) );
INVx1_ASAP7_75t_L g1110 ( .A(n_1111), .Y(n_1110) );
OR2x2_ASAP7_75t_L g1135 ( .A(n_1111), .B(n_1116), .Y(n_1135) );
NAND2xp5_ASAP7_75t_L g1111 ( .A(n_1112), .B(n_1114), .Y(n_1111) );
HB1xp67_ASAP7_75t_L g1436 ( .A(n_1112), .Y(n_1436) );
INVx1_ASAP7_75t_L g1112 ( .A(n_1113), .Y(n_1112) );
INVx1_ASAP7_75t_L g1123 ( .A(n_1114), .Y(n_1123) );
AND2x4_ASAP7_75t_L g1117 ( .A(n_1115), .B(n_1118), .Y(n_1117) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1116), .Y(n_1115) );
OR2x2_ASAP7_75t_L g1137 ( .A(n_1116), .B(n_1119), .Y(n_1137) );
INVx1_ASAP7_75t_L g1118 ( .A(n_1119), .Y(n_1118) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1121), .Y(n_1271) );
AND2x4_ASAP7_75t_L g1121 ( .A(n_1122), .B(n_1124), .Y(n_1121) );
AND2x2_ASAP7_75t_L g1158 ( .A(n_1122), .B(n_1124), .Y(n_1158) );
HB1xp67_ASAP7_75t_L g1434 ( .A(n_1122), .Y(n_1434) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1123), .Y(n_1122) );
AND2x4_ASAP7_75t_L g1125 ( .A(n_1123), .B(n_1124), .Y(n_1125) );
INVx2_ASAP7_75t_L g1150 ( .A(n_1125), .Y(n_1150) );
OAI21xp5_ASAP7_75t_L g1168 ( .A1(n_1126), .A2(n_1169), .B(n_1170), .Y(n_1168) );
INVx1_ASAP7_75t_L g1225 ( .A(n_1126), .Y(n_1225) );
AND2x2_ASAP7_75t_L g1260 ( .A(n_1126), .B(n_1188), .Y(n_1260) );
AOI221xp5_ASAP7_75t_L g1296 ( .A1(n_1126), .A2(n_1194), .B1(n_1290), .B2(n_1297), .C(n_1298), .Y(n_1296) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_1127), .B(n_1131), .Y(n_1126) );
AND2x2_ASAP7_75t_L g1141 ( .A(n_1127), .B(n_1142), .Y(n_1141) );
NOR2x1_ASAP7_75t_L g1184 ( .A(n_1127), .B(n_1185), .Y(n_1184) );
NAND2xp5_ASAP7_75t_L g1199 ( .A(n_1127), .B(n_1185), .Y(n_1199) );
NAND2xp5_ASAP7_75t_L g1220 ( .A(n_1127), .B(n_1210), .Y(n_1220) );
AND2x2_ASAP7_75t_L g1245 ( .A(n_1127), .B(n_1180), .Y(n_1245) );
OR2x2_ASAP7_75t_L g1248 ( .A(n_1127), .B(n_1249), .Y(n_1248) );
INVx2_ASAP7_75t_L g1127 ( .A(n_1128), .Y(n_1127) );
AND2x2_ASAP7_75t_L g1167 ( .A(n_1128), .B(n_1131), .Y(n_1167) );
AND2x2_ASAP7_75t_L g1169 ( .A(n_1128), .B(n_1144), .Y(n_1169) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_1128), .B(n_1179), .Y(n_1178) );
BUFx3_ASAP7_75t_L g1191 ( .A(n_1128), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1128), .B(n_1185), .Y(n_1215) );
AND2x2_ASAP7_75t_L g1224 ( .A(n_1128), .B(n_1210), .Y(n_1224) );
OR2x2_ASAP7_75t_L g1285 ( .A(n_1128), .B(n_1286), .Y(n_1285) );
AND2x2_ASAP7_75t_L g1128 ( .A(n_1129), .B(n_1130), .Y(n_1128) );
AND2x2_ASAP7_75t_L g1196 ( .A(n_1131), .B(n_1197), .Y(n_1196) );
INVx1_ASAP7_75t_L g1242 ( .A(n_1131), .Y(n_1242) );
OAI21xp5_ASAP7_75t_L g1289 ( .A1(n_1131), .A2(n_1245), .B(n_1290), .Y(n_1289) );
AND2x2_ASAP7_75t_L g1131 ( .A(n_1132), .B(n_1138), .Y(n_1131) );
AND2x2_ASAP7_75t_L g1144 ( .A(n_1132), .B(n_1145), .Y(n_1144) );
INVx2_ASAP7_75t_L g1180 ( .A(n_1132), .Y(n_1180) );
OAI22xp33_ASAP7_75t_L g1151 ( .A1(n_1134), .A2(n_1152), .B1(n_1153), .B2(n_1154), .Y(n_1151) );
BUFx3_ASAP7_75t_L g1274 ( .A(n_1134), .Y(n_1274) );
BUFx6f_ASAP7_75t_L g1134 ( .A(n_1135), .Y(n_1134) );
HB1xp67_ASAP7_75t_L g1154 ( .A(n_1137), .Y(n_1154) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1137), .Y(n_1277) );
INVx1_ASAP7_75t_L g1145 ( .A(n_1138), .Y(n_1145) );
AND2x2_ASAP7_75t_L g1179 ( .A(n_1138), .B(n_1180), .Y(n_1179) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1138), .Y(n_1185) );
AOI221xp5_ASAP7_75t_L g1221 ( .A1(n_1141), .A2(n_1202), .B1(n_1222), .B2(n_1226), .C(n_1227), .Y(n_1221) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1144), .Y(n_1286) );
AND2x2_ASAP7_75t_L g1210 ( .A(n_1145), .B(n_1180), .Y(n_1210) );
NAND3xp33_ASAP7_75t_L g1195 ( .A(n_1146), .B(n_1193), .C(n_1196), .Y(n_1195) );
NAND2xp5_ASAP7_75t_L g1264 ( .A(n_1146), .B(n_1194), .Y(n_1264) );
AND2x4_ASAP7_75t_SL g1146 ( .A(n_1147), .B(n_1155), .Y(n_1146) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_1147), .B(n_1156), .Y(n_1176) );
OR2x2_ASAP7_75t_L g1232 ( .A(n_1147), .B(n_1155), .Y(n_1232) );
INVx2_ASAP7_75t_SL g1147 ( .A(n_1148), .Y(n_1147) );
AND2x2_ASAP7_75t_L g1173 ( .A(n_1148), .B(n_1155), .Y(n_1173) );
OR2x2_ASAP7_75t_L g1192 ( .A(n_1148), .B(n_1193), .Y(n_1192) );
INVx2_ASAP7_75t_L g1229 ( .A(n_1148), .Y(n_1229) );
INVx2_ASAP7_75t_L g1149 ( .A(n_1150), .Y(n_1149) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1150), .Y(n_1309) );
AND2x2_ASAP7_75t_L g1207 ( .A(n_1155), .B(n_1194), .Y(n_1207) );
AND2x2_ASAP7_75t_L g1288 ( .A(n_1155), .B(n_1163), .Y(n_1288) );
CKINVDCx6p67_ASAP7_75t_R g1155 ( .A(n_1156), .Y(n_1155) );
AND2x2_ASAP7_75t_L g1202 ( .A(n_1156), .B(n_1163), .Y(n_1202) );
AND2x2_ASAP7_75t_L g1211 ( .A(n_1156), .B(n_1212), .Y(n_1211) );
CKINVDCx5p33_ASAP7_75t_R g1246 ( .A(n_1156), .Y(n_1246) );
OR2x6_ASAP7_75t_L g1156 ( .A(n_1157), .B(n_1159), .Y(n_1156) );
O2A1O1Ixp33_ASAP7_75t_L g1160 ( .A1(n_1161), .A2(n_1166), .B(n_1168), .C(n_1172), .Y(n_1160) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1162), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1251 ( .A(n_1162), .B(n_1210), .Y(n_1251) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1163), .Y(n_1177) );
CKINVDCx5p33_ASAP7_75t_R g1194 ( .A(n_1163), .Y(n_1194) );
INVx1_ASAP7_75t_SL g1212 ( .A(n_1163), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1163 ( .A(n_1164), .B(n_1165), .Y(n_1163) );
AOI21xp33_ASAP7_75t_SL g1198 ( .A1(n_1166), .A2(n_1199), .B(n_1200), .Y(n_1198) );
NOR2xp33_ASAP7_75t_L g1283 ( .A(n_1166), .B(n_1194), .Y(n_1283) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1167), .Y(n_1166) );
AOI21xp5_ASAP7_75t_L g1261 ( .A1(n_1167), .A2(n_1262), .B(n_1263), .Y(n_1261) );
NAND2xp5_ASAP7_75t_L g1282 ( .A(n_1167), .B(n_1238), .Y(n_1282) );
AND2x2_ASAP7_75t_L g1227 ( .A(n_1169), .B(n_1228), .Y(n_1227) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1171), .Y(n_1170) );
INVx1_ASAP7_75t_L g1172 ( .A(n_1173), .Y(n_1172) );
NAND2xp5_ASAP7_75t_L g1218 ( .A(n_1173), .B(n_1212), .Y(n_1218) );
NAND2xp5_ASAP7_75t_L g1250 ( .A(n_1173), .B(n_1251), .Y(n_1250) );
NAND2xp5_ASAP7_75t_L g1281 ( .A(n_1173), .B(n_1189), .Y(n_1281) );
AOI211xp5_ASAP7_75t_SL g1174 ( .A1(n_1175), .A2(n_1178), .B(n_1181), .C(n_1198), .Y(n_1174) );
AND2x2_ASAP7_75t_L g1175 ( .A(n_1176), .B(n_1177), .Y(n_1175) );
INVx2_ASAP7_75t_L g1186 ( .A(n_1176), .Y(n_1186) );
NAND3xp33_ASAP7_75t_L g1302 ( .A(n_1177), .B(n_1297), .C(n_1303), .Y(n_1302) );
NAND2xp5_ASAP7_75t_L g1205 ( .A(n_1179), .B(n_1206), .Y(n_1205) );
NAND2xp5_ASAP7_75t_L g1249 ( .A(n_1179), .B(n_1189), .Y(n_1249) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1179), .Y(n_1266) );
INVx2_ASAP7_75t_L g1297 ( .A(n_1180), .Y(n_1297) );
OAI221xp5_ASAP7_75t_L g1181 ( .A1(n_1182), .A2(n_1186), .B1(n_1187), .B2(n_1192), .C(n_1195), .Y(n_1181) );
INVx1_ASAP7_75t_L g1182 ( .A(n_1183), .Y(n_1182) );
OR2x2_ASAP7_75t_L g1190 ( .A(n_1185), .B(n_1191), .Y(n_1190) );
AOI222xp33_ASAP7_75t_L g1300 ( .A1(n_1185), .A2(n_1207), .B1(n_1269), .B2(n_1301), .C1(n_1304), .C2(n_1306), .Y(n_1300) );
OR2x2_ASAP7_75t_L g1187 ( .A(n_1188), .B(n_1190), .Y(n_1187) );
NAND2xp5_ASAP7_75t_L g1256 ( .A(n_1188), .B(n_1207), .Y(n_1256) );
INVx2_ASAP7_75t_L g1188 ( .A(n_1189), .Y(n_1188) );
OR2x2_ASAP7_75t_L g1219 ( .A(n_1189), .B(n_1220), .Y(n_1219) );
NAND2xp5_ASAP7_75t_L g1234 ( .A(n_1189), .B(n_1224), .Y(n_1234) );
NAND2xp5_ASAP7_75t_L g1294 ( .A(n_1189), .B(n_1245), .Y(n_1294) );
OR2x2_ASAP7_75t_L g1265 ( .A(n_1191), .B(n_1266), .Y(n_1265) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1192), .Y(n_1262) );
INVx3_ASAP7_75t_L g1193 ( .A(n_1194), .Y(n_1193) );
NOR2xp33_ASAP7_75t_L g1292 ( .A(n_1194), .B(n_1234), .Y(n_1292) );
NAND2xp5_ASAP7_75t_L g1200 ( .A(n_1201), .B(n_1202), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1228 ( .A(n_1202), .B(n_1229), .Y(n_1228) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1202), .Y(n_1243) );
AOI221xp5_ASAP7_75t_L g1203 ( .A1(n_1204), .A2(n_1207), .B1(n_1208), .B2(n_1211), .C(n_1213), .Y(n_1203) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1205), .Y(n_1204) );
NAND2xp5_ASAP7_75t_L g1209 ( .A(n_1206), .B(n_1210), .Y(n_1209) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1209), .Y(n_1208) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1210), .Y(n_1241) );
INVx1_ASAP7_75t_L g1295 ( .A(n_1211), .Y(n_1295) );
INVxp67_ASAP7_75t_SL g1213 ( .A(n_1214), .Y(n_1213) );
NAND2xp5_ASAP7_75t_L g1214 ( .A(n_1215), .B(n_1216), .Y(n_1214) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1215), .Y(n_1257) );
OAI211xp5_ASAP7_75t_L g1217 ( .A1(n_1218), .A2(n_1219), .B(n_1221), .C(n_1230), .Y(n_1217) );
OAI221xp5_ASAP7_75t_L g1280 ( .A1(n_1218), .A2(n_1244), .B1(n_1265), .B2(n_1281), .C(n_1282), .Y(n_1280) );
NAND2xp5_ASAP7_75t_L g1222 ( .A(n_1223), .B(n_1225), .Y(n_1222) );
OAI221xp5_ASAP7_75t_L g1247 ( .A1(n_1223), .A2(n_1232), .B1(n_1246), .B2(n_1248), .C(n_1250), .Y(n_1247) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1224), .Y(n_1223) );
INVx2_ASAP7_75t_L g1238 ( .A(n_1229), .Y(n_1238) );
NOR2xp33_ASAP7_75t_L g1254 ( .A(n_1229), .B(n_1255), .Y(n_1254) );
INVx2_ASAP7_75t_L g1259 ( .A(n_1229), .Y(n_1259) );
OAI31xp33_ASAP7_75t_L g1284 ( .A1(n_1229), .A2(n_1285), .A3(n_1287), .B(n_1289), .Y(n_1284) );
AND2x2_ASAP7_75t_L g1299 ( .A(n_1229), .B(n_1269), .Y(n_1299) );
NAND2xp5_ASAP7_75t_L g1230 ( .A(n_1231), .B(n_1233), .Y(n_1230) );
INVx1_ASAP7_75t_L g1231 ( .A(n_1232), .Y(n_1231) );
INVx1_ASAP7_75t_L g1233 ( .A(n_1234), .Y(n_1233) );
AOI21xp5_ASAP7_75t_L g1235 ( .A1(n_1236), .A2(n_1267), .B(n_1278), .Y(n_1235) );
NAND3xp33_ASAP7_75t_L g1236 ( .A(n_1237), .B(n_1258), .C(n_1261), .Y(n_1236) );
AOI211xp5_ASAP7_75t_L g1237 ( .A1(n_1238), .A2(n_1239), .B(n_1247), .C(n_1252), .Y(n_1237) );
NAND2xp5_ASAP7_75t_L g1240 ( .A(n_1241), .B(n_1242), .Y(n_1240) );
INVx1_ASAP7_75t_L g1244 ( .A(n_1245), .Y(n_1244) );
OAI221xp5_ASAP7_75t_SL g1293 ( .A1(n_1246), .A2(n_1266), .B1(n_1294), .B2(n_1295), .C(n_1296), .Y(n_1293) );
AOI21xp33_ASAP7_75t_SL g1252 ( .A1(n_1253), .A2(n_1256), .B(n_1257), .Y(n_1252) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1254), .Y(n_1253) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1255), .Y(n_1290) );
NAND2xp5_ASAP7_75t_L g1258 ( .A(n_1259), .B(n_1260), .Y(n_1258) );
NOR2xp33_ASAP7_75t_L g1263 ( .A(n_1264), .B(n_1265), .Y(n_1263) );
INVx2_ASAP7_75t_L g1267 ( .A(n_1268), .Y(n_1267) );
OAI31xp33_ASAP7_75t_L g1279 ( .A1(n_1268), .A2(n_1280), .A3(n_1283), .B(n_1284), .Y(n_1279) );
BUFx3_ASAP7_75t_L g1268 ( .A(n_1269), .Y(n_1268) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1269), .Y(n_1307) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1271), .Y(n_1270) );
OAI22xp33_ASAP7_75t_L g1272 ( .A1(n_1273), .A2(n_1274), .B1(n_1275), .B2(n_1276), .Y(n_1272) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1277), .Y(n_1276) );
NAND3xp33_ASAP7_75t_L g1278 ( .A(n_1279), .B(n_1291), .C(n_1300), .Y(n_1278) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1288), .Y(n_1287) );
OAI21xp33_ASAP7_75t_L g1291 ( .A1(n_1292), .A2(n_1293), .B(n_1299), .Y(n_1291) );
INVx1_ASAP7_75t_L g1304 ( .A(n_1305), .Y(n_1304) );
INVx1_ASAP7_75t_L g1308 ( .A(n_1309), .Y(n_1308) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1311), .Y(n_1310) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1312), .Y(n_1311) );
NAND2xp5_ASAP7_75t_L g1313 ( .A(n_1314), .B(n_1345), .Y(n_1313) );
AOI31xp33_ASAP7_75t_L g1316 ( .A1(n_1317), .A2(n_1332), .A3(n_1341), .B(n_1344), .Y(n_1316) );
OAI22xp5_ASAP7_75t_L g1358 ( .A1(n_1318), .A2(n_1343), .B1(n_1359), .B2(n_1360), .Y(n_1358) );
INVx3_ASAP7_75t_L g1321 ( .A(n_1322), .Y(n_1321) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1325), .Y(n_1324) );
INVx2_ASAP7_75t_SL g1326 ( .A(n_1327), .Y(n_1326) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1334), .Y(n_1333) );
OAI22xp33_ASAP7_75t_L g1361 ( .A1(n_1335), .A2(n_1342), .B1(n_1362), .B2(n_1364), .Y(n_1361) );
INVx2_ASAP7_75t_L g1339 ( .A(n_1340), .Y(n_1339) );
NOR3xp33_ASAP7_75t_L g1345 ( .A(n_1346), .B(n_1365), .C(n_1366), .Y(n_1345) );
OAI22xp5_ASAP7_75t_L g1347 ( .A1(n_1348), .A2(n_1349), .B1(n_1350), .B2(n_1351), .Y(n_1347) );
OAI22xp33_ASAP7_75t_L g1352 ( .A1(n_1353), .A2(n_1354), .B1(n_1355), .B2(n_1356), .Y(n_1352) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1357), .Y(n_1356) );
INVx3_ASAP7_75t_L g1362 ( .A(n_1363), .Y(n_1362) );
NAND2xp5_ASAP7_75t_L g1366 ( .A(n_1367), .B(n_1370), .Y(n_1366) );
INVx4_ASAP7_75t_SL g1372 ( .A(n_1373), .Y(n_1372) );
BUFx3_ASAP7_75t_L g1373 ( .A(n_1374), .Y(n_1373) );
BUFx2_ASAP7_75t_L g1374 ( .A(n_1375), .Y(n_1374) );
INVx1_ASAP7_75t_L g1377 ( .A(n_1378), .Y(n_1377) );
CKINVDCx5p33_ASAP7_75t_R g1378 ( .A(n_1379), .Y(n_1378) );
A2O1A1Ixp33_ASAP7_75t_L g1432 ( .A1(n_1380), .A2(n_1433), .B(n_1435), .C(n_1437), .Y(n_1432) );
INVxp33_ASAP7_75t_SL g1381 ( .A(n_1382), .Y(n_1381) );
INVx1_ASAP7_75t_L g1384 ( .A(n_1385), .Y(n_1384) );
HB1xp67_ASAP7_75t_L g1385 ( .A(n_1386), .Y(n_1385) );
NAND2x1_ASAP7_75t_L g1386 ( .A(n_1387), .B(n_1412), .Y(n_1386) );
AND4x1_ASAP7_75t_L g1387 ( .A(n_1388), .B(n_1391), .C(n_1405), .D(n_1408), .Y(n_1387) );
INVx1_ASAP7_75t_L g1402 ( .A(n_1403), .Y(n_1402) );
NAND3xp33_ASAP7_75t_L g1413 ( .A(n_1414), .B(n_1423), .C(n_1428), .Y(n_1413) );
AOI21xp5_ASAP7_75t_SL g1414 ( .A1(n_1415), .A2(n_1416), .B(n_1417), .Y(n_1414) );
INVx1_ASAP7_75t_L g1433 ( .A(n_1434), .Y(n_1433) );
INVx1_ASAP7_75t_L g1435 ( .A(n_1436), .Y(n_1435) );
endmodule