module fake_jpeg_29595_n_538 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_538);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_538;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_387;
wire n_270;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_412;
wire n_249;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_1),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_14),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_55),
.Y(n_125)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_57),
.Y(n_126)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_59),
.Y(n_150)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_61),
.Y(n_153)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_62),
.Y(n_129)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_64),
.Y(n_139)
);

INVx6_ASAP7_75t_SL g65 ( 
.A(n_22),
.Y(n_65)
);

INVx6_ASAP7_75t_SL g141 ( 
.A(n_65),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_66),
.Y(n_146)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_22),
.Y(n_67)
);

INVx5_ASAP7_75t_SL g169 ( 
.A(n_67),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_68),
.Y(n_151)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_69),
.Y(n_140)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_70),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_71),
.Y(n_174)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_72),
.Y(n_144)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_73),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_74),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_46),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_75),
.B(n_78),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_76),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_21),
.B(n_0),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_77),
.B(n_91),
.Y(n_167)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_17),
.B(n_2),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_79),
.B(n_82),
.Y(n_115)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_80),
.Y(n_166)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

INVx11_ASAP7_75t_L g134 ( 
.A(n_81),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_43),
.B(n_2),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_30),
.Y(n_83)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_83),
.Y(n_154)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_84),
.Y(n_145)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_85),
.Y(n_164)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g135 ( 
.A(n_86),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_17),
.B(n_2),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_87),
.B(n_105),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_31),
.Y(n_88)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_88),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_89),
.Y(n_127)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_34),
.Y(n_90)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_90),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_52),
.B(n_4),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_46),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_92),
.B(n_97),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_31),
.Y(n_93)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_93),
.Y(n_148)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_94),
.Y(n_149)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_95),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_96),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_39),
.Y(n_97)
);

BUFx12_ASAP7_75t_L g98 ( 
.A(n_34),
.Y(n_98)
);

BUFx24_ASAP7_75t_L g171 ( 
.A(n_98),
.Y(n_171)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_47),
.Y(n_99)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_99),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_101),
.Y(n_173)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

AND2x2_ASAP7_75t_SL g103 ( 
.A(n_25),
.B(n_5),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_107),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

BUFx8_ASAP7_75t_L g159 ( 
.A(n_104),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_36),
.B(n_54),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_36),
.B(n_5),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_106),
.B(n_108),
.Y(n_147)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_25),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_26),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_26),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_109),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_40),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_18),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_50),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_111),
.B(n_54),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_118),
.B(n_124),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_101),
.A2(n_53),
.B1(n_45),
.B2(n_40),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_119),
.A2(n_136),
.B1(n_170),
.B2(n_74),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_122),
.B(n_138),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_86),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_86),
.B(n_50),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_128),
.B(n_142),
.Y(n_206)
);

BUFx12f_ASAP7_75t_SL g131 ( 
.A(n_67),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g189 ( 
.A(n_131),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_55),
.A2(n_53),
.B1(n_45),
.B2(n_35),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_133),
.A2(n_168),
.B1(n_175),
.B2(n_68),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_104),
.A2(n_32),
.B1(n_28),
.B2(n_35),
.Y(n_136)
);

INVx6_ASAP7_75t_SL g138 ( 
.A(n_81),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g210 ( 
.A(n_138),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_110),
.B(n_24),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_98),
.B(n_24),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_155),
.B(n_157),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_98),
.B(n_32),
.Y(n_157)
);

BUFx12f_ASAP7_75t_L g158 ( 
.A(n_90),
.Y(n_158)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_158),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_99),
.A2(n_32),
.B1(n_28),
.B2(n_7),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_80),
.A2(n_28),
.B1(n_6),
.B2(n_7),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_95),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_177),
.A2(n_213),
.B1(n_228),
.B2(n_229),
.Y(n_264)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_112),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_178),
.Y(n_259)
);

NAND2x1_ASAP7_75t_L g179 ( 
.A(n_121),
.B(n_102),
.Y(n_179)
);

OAI21xp33_ASAP7_75t_L g236 ( 
.A1(n_179),
.A2(n_132),
.B(n_153),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_181),
.A2(n_215),
.B1(n_162),
.B2(n_174),
.Y(n_257)
);

BUFx12f_ASAP7_75t_L g182 ( 
.A(n_131),
.Y(n_182)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_182),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_117),
.B(n_85),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_183),
.B(n_192),
.Y(n_237)
);

BUFx12f_ASAP7_75t_L g184 ( 
.A(n_150),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_184),
.Y(n_241)
);

CKINVDCx12_ASAP7_75t_R g185 ( 
.A(n_141),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_185),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_120),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_186),
.B(n_205),
.Y(n_246)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_114),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_187),
.Y(n_275)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_113),
.Y(n_188)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_188),
.Y(n_238)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_129),
.Y(n_190)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_190),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g191 ( 
.A1(n_162),
.A2(n_66),
.B1(n_57),
.B2(n_100),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_191),
.A2(n_126),
.B1(n_125),
.B2(n_146),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_109),
.Y(n_192)
);

BUFx10_ASAP7_75t_L g193 ( 
.A(n_171),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_193),
.Y(n_252)
);

INVx8_ASAP7_75t_L g194 ( 
.A(n_159),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_194),
.Y(n_249)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_135),
.Y(n_195)
);

INVx5_ASAP7_75t_L g234 ( 
.A(n_195),
.Y(n_234)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_137),
.Y(n_196)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_196),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_147),
.B(n_96),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_198),
.B(n_218),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_107),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_199),
.B(n_207),
.Y(n_239)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_130),
.Y(n_200)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_200),
.Y(n_242)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_135),
.Y(n_201)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_201),
.Y(n_253)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_139),
.Y(n_202)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_202),
.Y(n_244)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_140),
.Y(n_203)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_203),
.Y(n_255)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_144),
.Y(n_204)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_204),
.Y(n_263)
);

A2O1A1Ixp33_ASAP7_75t_L g205 ( 
.A1(n_143),
.A2(n_89),
.B(n_61),
.C(n_9),
.Y(n_205)
);

CKINVDCx12_ASAP7_75t_R g207 ( 
.A(n_171),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_152),
.Y(n_208)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_208),
.Y(n_270)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_145),
.Y(n_209)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_209),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_115),
.B(n_5),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_211),
.B(n_221),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_161),
.B(n_93),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_212),
.B(n_226),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_119),
.A2(n_88),
.B1(n_83),
.B2(n_76),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_166),
.A2(n_71),
.B1(n_9),
.B2(n_10),
.Y(n_215)
);

OR2x2_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_227),
.Y(n_235)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_169),
.Y(n_217)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_217),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_149),
.B(n_6),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_164),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_219),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_166),
.B(n_148),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_220),
.B(n_230),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_159),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_116),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_222),
.B(n_223),
.Y(n_260)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_153),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_159),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_224),
.B(n_225),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_171),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_160),
.B(n_6),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_169),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_164),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_125),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_176),
.Y(n_230)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_134),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_232),
.Y(n_254)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_134),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_136),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_233),
.B(n_202),
.C(n_190),
.Y(n_286)
);

OAI21xp33_ASAP7_75t_L g289 ( 
.A1(n_236),
.A2(n_217),
.B(n_184),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_216),
.A2(n_175),
.B1(n_173),
.B2(n_170),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_245),
.B(n_257),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_220),
.B(n_163),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_256),
.B(n_267),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_205),
.A2(n_173),
.B(n_127),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_261),
.A2(n_127),
.B(n_223),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_181),
.A2(n_215),
.B1(n_206),
.B2(n_151),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_265),
.A2(n_268),
.B1(n_274),
.B2(n_154),
.Y(n_303)
);

AO22x1_ASAP7_75t_SL g267 ( 
.A1(n_179),
.A2(n_146),
.B1(n_174),
.B2(n_151),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_216),
.B(n_126),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_269),
.B(n_123),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_214),
.A2(n_154),
.B1(n_172),
.B2(n_165),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_266),
.B(n_180),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_276),
.B(n_287),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_250),
.B(n_182),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_277),
.B(n_282),
.Y(n_333)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_248),
.Y(n_278)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_278),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_243),
.B(n_189),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_279),
.B(n_286),
.C(n_288),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_272),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_280),
.B(n_289),
.Y(n_335)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_248),
.Y(n_281)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_281),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_182),
.Y(n_282)
);

INVx13_ASAP7_75t_L g283 ( 
.A(n_272),
.Y(n_283)
);

CKINVDCx14_ASAP7_75t_R g336 ( 
.A(n_283),
.Y(n_336)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_242),
.Y(n_284)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_284),
.Y(n_320)
);

INVx5_ASAP7_75t_SL g285 ( 
.A(n_252),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_285),
.B(n_290),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_246),
.B(n_210),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_233),
.B(n_204),
.C(n_188),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_239),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_253),
.Y(n_292)
);

INVx8_ASAP7_75t_L g314 ( 
.A(n_292),
.Y(n_314)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_242),
.Y(n_293)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_293),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_262),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_294),
.B(n_295),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_235),
.Y(n_295)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_253),
.Y(n_296)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_296),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_269),
.A2(n_210),
.B(n_230),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_297),
.A2(n_301),
.B(n_156),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_237),
.B(n_243),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_298),
.B(n_302),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_235),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_299),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_235),
.B(n_203),
.C(n_200),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_303),
.A2(n_172),
.B1(n_240),
.B2(n_259),
.Y(n_332)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_234),
.Y(n_304)
);

INVxp33_ASAP7_75t_L g319 ( 
.A(n_304),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_305),
.Y(n_310)
);

INVx8_ASAP7_75t_L g306 ( 
.A(n_252),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_306),
.Y(n_315)
);

INVx11_ASAP7_75t_L g307 ( 
.A(n_234),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_307),
.Y(n_322)
);

INVx13_ASAP7_75t_L g308 ( 
.A(n_241),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_308),
.Y(n_326)
);

AND2x6_ASAP7_75t_L g309 ( 
.A(n_261),
.B(n_193),
.Y(n_309)
);

OAI32xp33_ASAP7_75t_L g329 ( 
.A1(n_309),
.A2(n_274),
.A3(n_267),
.B1(n_254),
.B2(n_260),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_291),
.A2(n_264),
.B1(n_245),
.B2(n_265),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_312),
.A2(n_321),
.B1(n_339),
.B2(n_303),
.Y(n_359)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_299),
.B(n_256),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_317),
.B(n_298),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_291),
.A2(n_257),
.B1(n_268),
.B2(n_267),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_301),
.A2(n_254),
.B(n_273),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_328),
.A2(n_330),
.B(n_331),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_SL g358 ( 
.A(n_329),
.B(n_300),
.C(n_297),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_309),
.A2(n_273),
.B(n_275),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_309),
.A2(n_258),
.B(n_267),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_332),
.A2(n_300),
.B1(n_281),
.B2(n_306),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_300),
.A2(n_258),
.B(n_240),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g351 ( 
.A1(n_337),
.A2(n_338),
.B(n_305),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_278),
.A2(n_259),
.B1(n_209),
.B2(n_208),
.Y(n_339)
);

NOR2x1_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_287),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_341),
.B(n_349),
.Y(n_397)
);

INVx13_ASAP7_75t_L g342 ( 
.A(n_314),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_342),
.B(n_350),
.Y(n_372)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_320),
.Y(n_343)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_343),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_325),
.B(n_279),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_344),
.B(n_347),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_340),
.B(n_276),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_345),
.B(n_352),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_325),
.B(n_288),
.C(n_286),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_320),
.Y(n_348)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_348),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_325),
.B(n_302),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_351),
.B(n_335),
.Y(n_388)
);

INVxp67_ASAP7_75t_SL g352 ( 
.A(n_333),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_323),
.B(n_282),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_353),
.B(n_357),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g354 ( 
.A1(n_338),
.A2(n_335),
.B(n_337),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_354),
.A2(n_335),
.B(n_337),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_355),
.B(n_370),
.Y(n_399)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_327),
.Y(n_356)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_356),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_323),
.B(n_277),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_358),
.A2(n_364),
.B(n_335),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_359),
.A2(n_365),
.B1(n_366),
.B2(n_332),
.Y(n_371)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_327),
.Y(n_360)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_360),
.Y(n_386)
);

CKINVDCx14_ASAP7_75t_R g361 ( 
.A(n_313),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_361),
.B(n_363),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_332),
.A2(n_306),
.B1(n_285),
.B2(n_280),
.Y(n_362)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_362),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_333),
.B(n_251),
.Y(n_363)
);

AND2x6_ASAP7_75t_L g364 ( 
.A(n_330),
.B(n_283),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g365 ( 
.A1(n_312),
.A2(n_285),
.B1(n_296),
.B2(n_284),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_321),
.A2(n_293),
.B1(n_292),
.B2(n_304),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_313),
.B(n_283),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_367),
.B(n_368),
.Y(n_400)
);

AOI322xp5_ASAP7_75t_L g368 ( 
.A1(n_311),
.A2(n_308),
.A3(n_292),
.B1(n_123),
.B2(n_251),
.C1(n_229),
.C2(n_184),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_316),
.Y(n_369)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_369),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_311),
.B(n_263),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_371),
.B(n_373),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_357),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_359),
.A2(n_331),
.B1(n_330),
.B2(n_316),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_374),
.B(n_382),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_369),
.Y(n_376)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_376),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_341),
.B(n_317),
.Y(n_379)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_379),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_355),
.B(n_353),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_380),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_343),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_348),
.Y(n_383)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_383),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_SL g429 ( 
.A(n_385),
.B(n_390),
.C(n_326),
.Y(n_429)
);

CKINVDCx16_ASAP7_75t_R g424 ( 
.A(n_388),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_356),
.B(n_317),
.Y(n_389)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_389),
.Y(n_420)
);

CKINVDCx16_ASAP7_75t_R g391 ( 
.A(n_360),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_391),
.B(n_315),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_354),
.B(n_351),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_393),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_358),
.A2(n_331),
.B1(n_318),
.B2(n_328),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_395),
.B(n_398),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_342),
.Y(n_398)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_366),
.Y(n_401)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_401),
.Y(n_425)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_402),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_394),
.B(n_347),
.C(n_350),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_403),
.B(n_405),
.C(n_410),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_378),
.B(n_324),
.Y(n_404)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_404),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_394),
.B(n_344),
.C(n_370),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_372),
.B(n_393),
.C(n_399),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_395),
.B(n_346),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_411),
.B(n_396),
.Y(n_445)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_397),
.B(n_346),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_414),
.B(n_417),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_393),
.B(n_328),
.C(n_365),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_415),
.B(n_418),
.C(n_422),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_397),
.B(n_329),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_399),
.B(n_324),
.C(n_310),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_373),
.A2(n_318),
.B1(n_329),
.B2(n_364),
.Y(n_419)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_419),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_385),
.B(n_315),
.C(n_322),
.Y(n_422)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_379),
.B(n_339),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_423),
.B(n_430),
.C(n_375),
.Y(n_452)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_378),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_426),
.B(n_428),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_387),
.A2(n_322),
.B1(n_336),
.B2(n_334),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_427),
.A2(n_401),
.B1(n_387),
.B2(n_371),
.Y(n_431)
);

INVxp67_ASAP7_75t_SL g428 ( 
.A(n_384),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_SL g436 ( 
.A(n_429),
.B(n_388),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_389),
.B(n_334),
.C(n_336),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g465 ( 
.A(n_431),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_409),
.A2(n_400),
.B1(n_392),
.B2(n_374),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_432),
.A2(n_450),
.B1(n_453),
.B2(n_427),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_416),
.B(n_380),
.Y(n_433)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_433),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_436),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_417),
.A2(n_388),
.B1(n_392),
.B2(n_390),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_437),
.B(n_441),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_420),
.B(n_382),
.Y(n_439)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_439),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_SL g441 ( 
.A(n_407),
.B(n_398),
.Y(n_441)
);

INVxp33_ASAP7_75t_SL g443 ( 
.A(n_429),
.Y(n_443)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_443),
.Y(n_466)
);

NAND3xp33_ASAP7_75t_L g444 ( 
.A(n_421),
.B(n_396),
.C(n_375),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_444),
.B(n_448),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_445),
.B(n_452),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_425),
.A2(n_386),
.B1(n_381),
.B2(n_377),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_408),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_449),
.B(n_308),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_408),
.A2(n_391),
.B1(n_386),
.B2(n_381),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_405),
.B(n_377),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_451),
.B(n_406),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_409),
.A2(n_383),
.B1(n_314),
.B2(n_307),
.Y(n_453)
);

OAI322xp33_ASAP7_75t_L g454 ( 
.A1(n_433),
.A2(n_412),
.A3(n_403),
.B1(n_418),
.B2(n_422),
.C1(n_410),
.C2(n_414),
.Y(n_454)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_454),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_434),
.B(n_430),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_455),
.B(n_468),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_432),
.A2(n_424),
.B1(n_411),
.B2(n_415),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_457),
.B(n_459),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_447),
.B(n_412),
.C(n_423),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_458),
.B(n_461),
.C(n_440),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_460),
.B(n_472),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_447),
.B(n_451),
.C(n_452),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_435),
.A2(n_413),
.B(n_319),
.Y(n_467)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_467),
.Y(n_482)
);

BUFx24_ASAP7_75t_SL g468 ( 
.A(n_438),
.Y(n_468)
);

OR2x2_ASAP7_75t_L g479 ( 
.A(n_470),
.B(n_463),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_442),
.B(n_271),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_471),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_474),
.B(n_478),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_476),
.B(n_469),
.Y(n_494)
);

CKINVDCx16_ASAP7_75t_R g478 ( 
.A(n_466),
.Y(n_478)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_479),
.Y(n_502)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_469),
.B(n_442),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_480),
.B(n_484),
.C(n_487),
.Y(n_492)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_464),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_483),
.B(n_486),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_461),
.B(n_440),
.C(n_445),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_456),
.A2(n_446),
.B(n_439),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_485),
.A2(n_489),
.B(n_255),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_465),
.A2(n_431),
.B1(n_437),
.B2(n_436),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_458),
.B(n_448),
.C(n_314),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g488 ( 
.A1(n_465),
.A2(n_307),
.B1(n_249),
.B2(n_244),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_488),
.B(n_249),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_456),
.A2(n_271),
.B(n_244),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g490 ( 
.A1(n_485),
.A2(n_462),
.B(n_457),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g516 ( 
.A1(n_490),
.A2(n_197),
.B(n_195),
.Y(n_516)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_491),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_494),
.B(n_497),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_482),
.A2(n_472),
.B1(n_249),
.B2(n_263),
.Y(n_496)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_496),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_477),
.A2(n_255),
.B1(n_231),
.B2(n_232),
.Y(n_498)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_498),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_475),
.B(n_270),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_499),
.B(n_501),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_476),
.B(n_270),
.C(n_247),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_500),
.B(n_480),
.C(n_481),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_479),
.B(n_247),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_473),
.B(n_238),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_503),
.B(n_504),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_487),
.B(n_238),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_SL g507 ( 
.A(n_493),
.B(n_484),
.Y(n_507)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_507),
.Y(n_519)
);

NAND2x1_ASAP7_75t_SL g508 ( 
.A(n_490),
.B(n_489),
.Y(n_508)
);

AOI322xp5_ASAP7_75t_L g518 ( 
.A1(n_508),
.A2(n_509),
.A3(n_515),
.B1(n_491),
.B2(n_502),
.C1(n_505),
.C2(n_512),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_492),
.B(n_477),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_514),
.B(n_492),
.C(n_500),
.Y(n_517)
);

OAI31xp33_ASAP7_75t_L g515 ( 
.A1(n_495),
.A2(n_486),
.A3(n_488),
.B(n_481),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_516),
.Y(n_523)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_517),
.Y(n_528)
);

AO21x1_ASAP7_75t_L g526 ( 
.A1(n_518),
.A2(n_520),
.B(n_522),
.Y(n_526)
);

AOI322xp5_ASAP7_75t_L g520 ( 
.A1(n_510),
.A2(n_498),
.A3(n_496),
.B1(n_150),
.B2(n_197),
.C1(n_123),
.C2(n_158),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_514),
.B(n_176),
.C(n_219),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_521),
.A2(n_524),
.B(n_511),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_SL g522 ( 
.A1(n_506),
.A2(n_201),
.B(n_156),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_513),
.B(n_194),
.C(n_158),
.Y(n_524)
);

AOI21x1_ASAP7_75t_L g525 ( 
.A1(n_519),
.A2(n_516),
.B(n_508),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_525),
.B(n_527),
.Y(n_532)
);

AOI21x1_ASAP7_75t_L g529 ( 
.A1(n_523),
.A2(n_515),
.B(n_193),
.Y(n_529)
);

AOI322xp5_ASAP7_75t_L g531 ( 
.A1(n_529),
.A2(n_132),
.A3(n_193),
.B1(n_12),
.B2(n_14),
.C1(n_9),
.C2(n_16),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_528),
.B(n_526),
.Y(n_530)
);

OA21x2_ASAP7_75t_L g534 ( 
.A1(n_530),
.A2(n_531),
.B(n_11),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_532),
.B(n_132),
.C(n_12),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_533),
.B(n_534),
.C(n_11),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_535),
.B(n_14),
.C(n_15),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_536),
.B(n_14),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_537),
.B(n_15),
.Y(n_538)
);


endmodule