module fake_jpeg_20611_n_304 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_304);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_304;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_181;
wire n_26;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_155;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx6_ASAP7_75t_SL g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_5),
.Y(n_24)
);

OR2x2_ASAP7_75t_L g25 ( 
.A(n_0),
.B(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_20),
.Y(n_53)
);

AOI21xp33_ASAP7_75t_SL g39 ( 
.A1(n_25),
.A2(n_0),
.B(n_1),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_39),
.B(n_24),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx5_ASAP7_75t_SL g54 ( 
.A(n_41),
.Y(n_54)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_35),
.A2(n_24),
.B1(n_18),
.B2(n_17),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_45),
.A2(n_28),
.B1(n_34),
.B2(n_33),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_46),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_50),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_25),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_51),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_25),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_42),
.B(n_29),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_52),
.B(n_65),
.Y(n_84)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_56),
.B(n_59),
.Y(n_85)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_42),
.Y(n_59)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_38),
.A2(n_17),
.B1(n_18),
.B2(n_32),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_64),
.A2(n_32),
.B1(n_29),
.B2(n_30),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_38),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_72),
.A2(n_78),
.B1(n_81),
.B2(n_87),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_63),
.A2(n_30),
.B1(n_27),
.B2(n_19),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g103 ( 
.A(n_73),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_48),
.A2(n_19),
.B(n_27),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_82),
.C(n_33),
.Y(n_106)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_77),
.B(n_88),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_52),
.A2(n_33),
.B1(n_41),
.B2(n_37),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_80),
.B(n_83),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_64),
.A2(n_43),
.B1(n_41),
.B2(n_37),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_43),
.Y(n_82)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_44),
.Y(n_86)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_56),
.A2(n_61),
.B1(n_60),
.B2(n_58),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_47),
.Y(n_89)
);

BUFx24_ASAP7_75t_SL g114 ( 
.A(n_89),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_57),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_90),
.B(n_49),
.Y(n_119)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_92),
.A2(n_54),
.B1(n_69),
.B2(n_57),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_50),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_93),
.B(n_100),
.Y(n_145)
);

OA22x2_ASAP7_75t_L g94 ( 
.A1(n_87),
.A2(n_65),
.B1(n_60),
.B2(n_44),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_94),
.A2(n_98),
.B(n_71),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_85),
.B(n_16),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_97),
.B(n_105),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_85),
.B(n_62),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_66),
.B(n_55),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_70),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_106),
.A2(n_112),
.B1(n_54),
.B2(n_79),
.Y(n_128)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_82),
.B(n_84),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_108),
.B(n_113),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_76),
.B(n_15),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_118),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_55),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_86),
.Y(n_115)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_115),
.Y(n_127)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_75),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_55),
.Y(n_117)
);

AND2x2_ASAP7_75t_SL g139 ( 
.A(n_117),
.B(n_49),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_76),
.B(n_14),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g134 ( 
.A(n_119),
.Y(n_134)
);

NAND3xp33_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_74),
.C(n_1),
.Y(n_120)
);

NAND3xp33_ASAP7_75t_L g155 ( 
.A(n_120),
.B(n_146),
.C(n_113),
.Y(n_155)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_101),
.A2(n_103),
.B1(n_107),
.B2(n_105),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_124),
.A2(n_94),
.B1(n_115),
.B2(n_96),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_104),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_125),
.B(n_132),
.Y(n_177)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_126),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_128),
.A2(n_143),
.B(n_144),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_94),
.A2(n_72),
.B1(n_54),
.B2(n_79),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_129),
.A2(n_136),
.B1(n_147),
.B2(n_139),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_90),
.C(n_75),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_139),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_104),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_95),
.Y(n_133)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_133),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_91),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_135),
.B(n_141),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_101),
.A2(n_79),
.B1(n_68),
.B2(n_69),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_94),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_91),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_97),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_131),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_98),
.A2(n_71),
.B(n_34),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_98),
.A2(n_69),
.B(n_88),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_94),
.A2(n_77),
.B(n_28),
.Y(n_146)
);

OAI32xp33_ASAP7_75t_L g147 ( 
.A1(n_93),
.A2(n_83),
.A3(n_43),
.B1(n_41),
.B2(n_37),
.Y(n_147)
);

NOR3xp33_ASAP7_75t_SL g149 ( 
.A(n_140),
.B(n_119),
.C(n_106),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_149),
.B(n_150),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_127),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_152),
.B(n_154),
.Y(n_197)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_127),
.Y(n_153)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_153),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_121),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_L g191 ( 
.A1(n_155),
.A2(n_12),
.B(n_1),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_99),
.Y(n_156)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_156),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_158),
.A2(n_128),
.B1(n_134),
.B2(n_147),
.Y(n_181)
);

INVx2_ASAP7_75t_SL g159 ( 
.A(n_137),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_159),
.B(n_171),
.Y(n_196)
);

AOI21xp33_ASAP7_75t_L g162 ( 
.A1(n_143),
.A2(n_100),
.B(n_95),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_162),
.A2(n_165),
.B(n_43),
.Y(n_201)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_163),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_122),
.B(n_117),
.Y(n_164)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_164),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_124),
.B(n_102),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_167),
.B(n_169),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_168),
.A2(n_165),
.B1(n_172),
.B2(n_177),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_125),
.B(n_102),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_170),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_132),
.B(n_96),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_139),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_176),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_134),
.B(n_109),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_173),
.Y(n_180)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_126),
.Y(n_174)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_137),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_137),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_109),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_123),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_179),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_181),
.A2(n_182),
.B1(n_190),
.B2(n_159),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_158),
.A2(n_145),
.B1(n_148),
.B2(n_146),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_130),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_183),
.B(n_184),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_160),
.B(n_148),
.Y(n_184)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_187),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_145),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_193),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_168),
.A2(n_138),
.B1(n_144),
.B2(n_49),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_191),
.B(n_195),
.Y(n_212)
);

MAJx2_ASAP7_75t_L g193 ( 
.A(n_161),
.B(n_31),
.C(n_26),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_153),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_200),
.A2(n_159),
.B1(n_176),
.B2(n_157),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_201),
.A2(n_178),
.B(n_157),
.Y(n_214)
);

NAND2xp33_ASAP7_75t_SL g204 ( 
.A(n_165),
.B(n_41),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_36),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_205),
.A2(n_175),
.B1(n_152),
.B2(n_154),
.Y(n_206)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_206),
.Y(n_230)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_198),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_207),
.B(n_218),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_197),
.B(n_163),
.Y(n_210)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_210),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_189),
.A2(n_149),
.B1(n_151),
.B2(n_170),
.Y(n_211)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_211),
.Y(n_234)
);

AND2x2_ASAP7_75t_SL g213 ( 
.A(n_190),
.B(n_151),
.Y(n_213)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_213),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_214),
.B(n_227),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_215),
.B(n_221),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_183),
.B(n_174),
.C(n_166),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_216),
.B(n_223),
.C(n_224),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_199),
.B(n_192),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_180),
.B(n_179),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_219),
.B(n_222),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_220),
.A2(n_229),
.B1(n_187),
.B2(n_203),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_166),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_194),
.B(n_12),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_184),
.B(n_37),
.C(n_36),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_188),
.B(n_36),
.C(n_26),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_11),
.Y(n_225)
);

INVxp33_ASAP7_75t_L g245 ( 
.A(n_225),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_185),
.B(n_11),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_226),
.A2(n_228),
.B1(n_212),
.B2(n_221),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_202),
.B(n_10),
.Y(n_228)
);

AO22x1_ASAP7_75t_L g229 ( 
.A1(n_186),
.A2(n_31),
.B1(n_26),
.B2(n_23),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_208),
.B(n_182),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_227),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_248),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_216),
.B(n_201),
.C(n_200),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_209),
.C(n_215),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_220),
.A2(n_181),
.B1(n_186),
.B2(n_204),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_239),
.A2(n_241),
.B1(n_246),
.B2(n_213),
.Y(n_250)
);

XOR2x2_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_193),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_242),
.A2(n_214),
.B1(n_224),
.B2(n_223),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_210),
.A2(n_180),
.B1(n_203),
.B2(n_198),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_209),
.B(n_31),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_247),
.B(n_229),
.Y(n_254)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_207),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_249),
.B(n_259),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_250),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_233),
.B(n_213),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_255),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_254),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_217),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_234),
.A2(n_227),
.B1(n_23),
.B2(n_3),
.Y(n_256)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_256),
.Y(n_271)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_244),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_257),
.Y(n_268)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_231),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_258),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_230),
.B(n_8),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_261),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_9),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_243),
.B(n_9),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_262),
.A2(n_248),
.B1(n_245),
.B2(n_232),
.Y(n_273)
);

BUFx24_ASAP7_75t_SL g266 ( 
.A(n_251),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_270),
.Y(n_284)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_255),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_249),
.A2(n_240),
.B(n_242),
.Y(n_272)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_272),
.Y(n_275)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_273),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_253),
.C(n_232),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_276),
.A2(n_278),
.B(n_283),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_271),
.A2(n_235),
.B1(n_239),
.B2(n_254),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_277),
.A2(n_281),
.B1(n_13),
.B2(n_4),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_268),
.A2(n_237),
.B(n_247),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_263),
.B(n_259),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_9),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_265),
.A2(n_237),
.B1(n_23),
.B2(n_3),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_274),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_13),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_264),
.A2(n_7),
.B(n_2),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_275),
.A2(n_272),
.B(n_269),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_285),
.B(n_288),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_279),
.A2(n_269),
.B1(n_2),
.B2(n_3),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_289),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_291),
.Y(n_297)
);

NOR2xp67_ASAP7_75t_L g291 ( 
.A(n_282),
.B(n_4),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_284),
.A2(n_16),
.B1(n_4),
.B2(n_5),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_292),
.B(n_7),
.Y(n_294)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_294),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_280),
.C(n_14),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_296),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_293),
.A2(n_290),
.B(n_288),
.Y(n_298)
);

OAI211xp5_ASAP7_75t_L g301 ( 
.A1(n_298),
.A2(n_297),
.B(n_295),
.C(n_15),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_301),
.Y(n_302)
);

OAI21x1_ASAP7_75t_L g303 ( 
.A1(n_302),
.A2(n_299),
.B(n_300),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_303),
.B(n_0),
.Y(n_304)
);


endmodule