module real_aes_11660_n_344 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_1934, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_1935, n_63, n_1, n_237, n_91, n_344);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_1934;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_1935;
input n_63;
input n_1;
input n_237;
input n_91;
output n_344;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1929;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1888;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_549;
wire n_571;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_1920;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_595;
wire n_1893;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_1883;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_1872;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1890;
wire n_1675;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1250;
wire n_1095;
wire n_1284;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_1906;
wire n_351;
wire n_898;
wire n_1926;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_1301;
wire n_728;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_346;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1813;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_1921;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_1914;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_1499;
wire n_700;
wire n_399;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_1930;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_1856;
wire n_658;
wire n_676;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_1569;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_1907;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1580;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_1915;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_1633;
wire n_442;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1910;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1908;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1811;
wire n_1066;
wire n_1917;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_1928;
wire n_977;
wire n_943;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1932;
wire n_1707;
wire n_856;
wire n_594;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1913;
wire n_1470;
wire n_816;
wire n_1899;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1923;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1927;
wire n_1411;
wire n_1263;
wire n_1922;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1802;
wire n_1605;
wire n_1855;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1785;
wire n_1774;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1496;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_1226;
wire n_525;
wire n_1617;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_1176;
wire n_640;
wire n_1721;
wire n_1691;
wire n_1931;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1292;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_1911;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1912;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_1919;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_578;
wire n_372;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_1584;
wire n_559;
wire n_1277;
wire n_1049;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_1916;
wire n_1025;
wire n_532;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_1909;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1891;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1925;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1894;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_1481;
wire n_907;
wire n_1430;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1877;
wire n_1697;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_1573;
wire n_1130;
wire n_1918;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1924;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_1280;
wire n_729;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
OAI221xp5_ASAP7_75t_L g1843 ( .A1(n_0), .A2(n_653), .B1(n_1505), .B2(n_1844), .C(n_1850), .Y(n_1843) );
AOI21xp33_ASAP7_75t_L g1872 ( .A1(n_0), .A2(n_575), .B(n_784), .Y(n_1872) );
INVx1_ASAP7_75t_L g1564 ( .A(n_1), .Y(n_1564) );
OA22x2_ASAP7_75t_L g1482 ( .A1(n_2), .A2(n_1483), .B1(n_1536), .B2(n_1537), .Y(n_1482) );
INVxp67_ASAP7_75t_SL g1537 ( .A(n_2), .Y(n_1537) );
CKINVDCx5p33_ASAP7_75t_R g1304 ( .A(n_3), .Y(n_1304) );
INVx1_ASAP7_75t_L g374 ( .A(n_4), .Y(n_374) );
INVx1_ASAP7_75t_L g1305 ( .A(n_5), .Y(n_1305) );
OAI221xp5_ASAP7_75t_L g1853 ( .A1(n_6), .A2(n_185), .B1(n_643), .B2(n_648), .C(n_651), .Y(n_1853) );
CKINVDCx5p33_ASAP7_75t_R g1877 ( .A(n_6), .Y(n_1877) );
INVx1_ASAP7_75t_L g602 ( .A(n_7), .Y(n_602) );
OAI221xp5_ASAP7_75t_L g1552 ( .A1(n_8), .A2(n_318), .B1(n_641), .B2(n_648), .C(n_650), .Y(n_1552) );
OAI22xp33_ASAP7_75t_SL g1573 ( .A1(n_8), .A2(n_318), .B1(n_841), .B2(n_1134), .Y(n_1573) );
INVx1_ASAP7_75t_L g1636 ( .A(n_9), .Y(n_1636) );
INVxp33_ASAP7_75t_L g1398 ( .A(n_10), .Y(n_1398) );
AOI22xp33_ASAP7_75t_L g1479 ( .A1(n_10), .A2(n_107), .B1(n_1195), .B2(n_1470), .Y(n_1479) );
INVxp33_ASAP7_75t_L g1548 ( .A(n_11), .Y(n_1548) );
AOI221xp5_ASAP7_75t_L g1569 ( .A1(n_11), .A2(n_105), .B1(n_736), .B2(n_783), .C(n_1570), .Y(n_1569) );
AOI221xp5_ASAP7_75t_L g1293 ( .A1(n_12), .A2(n_102), .B1(n_736), .B2(n_1294), .C(n_1295), .Y(n_1293) );
INVx1_ASAP7_75t_L g1312 ( .A(n_12), .Y(n_1312) );
AOI22xp33_ASAP7_75t_SL g1193 ( .A1(n_13), .A2(n_162), .B1(n_1194), .B2(n_1195), .Y(n_1193) );
AOI22xp33_ASAP7_75t_L g1220 ( .A1(n_13), .A2(n_59), .B1(n_732), .B2(n_1129), .Y(n_1220) );
INVx1_ASAP7_75t_L g1562 ( .A(n_14), .Y(n_1562) );
AOI221xp5_ASAP7_75t_L g1046 ( .A1(n_15), .A2(n_268), .B1(n_791), .B2(n_1047), .C(n_1048), .Y(n_1046) );
INVx1_ASAP7_75t_L g1084 ( .A(n_15), .Y(n_1084) );
INVx1_ASAP7_75t_L g995 ( .A(n_16), .Y(n_995) );
XNOR2x2_ASAP7_75t_L g1186 ( .A(n_17), .B(n_1187), .Y(n_1186) );
CKINVDCx5p33_ASAP7_75t_R g1360 ( .A(n_18), .Y(n_1360) );
AOI22xp33_ASAP7_75t_SL g1197 ( .A1(n_19), .A2(n_59), .B1(n_1025), .B2(n_1198), .Y(n_1197) );
AOI21xp33_ASAP7_75t_L g1221 ( .A1(n_19), .A2(n_439), .B(n_861), .Y(n_1221) );
OAI22xp5_ASAP7_75t_L g1485 ( .A1(n_20), .A2(n_244), .B1(n_1002), .B2(n_1486), .Y(n_1485) );
CKINVDCx5p33_ASAP7_75t_R g1532 ( .A(n_20), .Y(n_1532) );
CKINVDCx5p33_ASAP7_75t_R g1898 ( .A(n_21), .Y(n_1898) );
AOI22xp5_ASAP7_75t_L g1661 ( .A1(n_22), .A2(n_133), .B1(n_1622), .B2(n_1625), .Y(n_1661) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_23), .A2(n_293), .B1(n_456), .B2(n_458), .Y(n_985) );
INVxp67_ASAP7_75t_SL g1029 ( .A(n_23), .Y(n_1029) );
INVxp33_ASAP7_75t_L g1404 ( .A(n_24), .Y(n_1404) );
AOI22xp33_ASAP7_75t_L g1477 ( .A1(n_24), .A2(n_210), .B1(n_1472), .B2(n_1478), .Y(n_1477) );
INVxp33_ASAP7_75t_L g394 ( .A(n_25), .Y(n_394) );
AOI221xp5_ASAP7_75t_L g504 ( .A1(n_25), .A2(n_82), .B1(n_505), .B2(n_507), .C(n_510), .Y(n_504) );
OAI221xp5_ASAP7_75t_L g769 ( .A1(n_26), .A2(n_73), .B1(n_770), .B2(n_772), .C(n_773), .Y(n_769) );
INVx1_ASAP7_75t_L g814 ( .A(n_26), .Y(n_814) );
CKINVDCx5p33_ASAP7_75t_R g1848 ( .A(n_27), .Y(n_1848) );
INVx1_ASAP7_75t_L g1212 ( .A(n_28), .Y(n_1212) );
AOI22xp33_ASAP7_75t_L g1224 ( .A1(n_28), .A2(n_301), .B1(n_439), .B2(n_732), .Y(n_1224) );
OAI22xp5_ASAP7_75t_L g1044 ( .A1(n_29), .A2(n_343), .B1(n_584), .B2(n_1045), .Y(n_1044) );
INVx1_ASAP7_75t_L g1070 ( .A(n_29), .Y(n_1070) );
INVx1_ASAP7_75t_L g698 ( .A(n_30), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_30), .A2(n_57), .B1(n_753), .B2(n_755), .Y(n_752) );
INVxp67_ASAP7_75t_SL g1106 ( .A(n_31), .Y(n_1106) );
AOI221xp5_ASAP7_75t_L g1125 ( .A1(n_31), .A2(n_327), .B1(n_595), .B2(n_775), .C(n_788), .Y(n_1125) );
OAI22xp5_ASAP7_75t_L g1855 ( .A1(n_32), .A2(n_69), .B1(n_1856), .B2(n_1857), .Y(n_1855) );
INVx1_ASAP7_75t_L g1869 ( .A(n_32), .Y(n_1869) );
INVxp33_ASAP7_75t_L g685 ( .A(n_33), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_33), .A2(n_85), .B1(n_731), .B2(n_732), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_34), .A2(n_330), .B1(n_445), .B2(n_448), .Y(n_444) );
INVxp67_ASAP7_75t_SL g536 ( .A(n_34), .Y(n_536) );
AOI221xp5_ASAP7_75t_L g1300 ( .A1(n_35), .A2(n_234), .B1(n_595), .B2(n_954), .C(n_1301), .Y(n_1300) );
INVx1_ASAP7_75t_L g1323 ( .A(n_35), .Y(n_1323) );
OAI211xp5_ASAP7_75t_SL g979 ( .A1(n_36), .A2(n_613), .B(n_980), .C(n_988), .Y(n_979) );
AOI221xp5_ASAP7_75t_L g1022 ( .A1(n_36), .A2(n_195), .B1(n_1023), .B2(n_1025), .C(n_1026), .Y(n_1022) );
CKINVDCx5p33_ASAP7_75t_R g1339 ( .A(n_37), .Y(n_1339) );
INVx1_ASAP7_75t_L g794 ( .A(n_38), .Y(n_794) );
INVx1_ASAP7_75t_L g349 ( .A(n_39), .Y(n_349) );
AOI22xp5_ASAP7_75t_L g1656 ( .A1(n_40), .A2(n_125), .B1(n_1622), .B2(n_1625), .Y(n_1656) );
INVx1_ASAP7_75t_L g1603 ( .A(n_41), .Y(n_1603) );
INVx1_ASAP7_75t_L g1055 ( .A(n_42), .Y(n_1055) );
AOI22xp33_ASAP7_75t_L g1078 ( .A1(n_42), .A2(n_315), .B1(n_505), .B2(n_1079), .Y(n_1078) );
OAI221xp5_ASAP7_75t_L g692 ( .A1(n_43), .A2(n_199), .B1(n_651), .B2(n_693), .C(n_694), .Y(n_692) );
OAI33xp33_ASAP7_75t_L g741 ( .A1(n_43), .A2(n_199), .A3(n_426), .B1(n_605), .B2(n_742), .B3(n_1934), .Y(n_741) );
INVx1_ASAP7_75t_L g1342 ( .A(n_44), .Y(n_1342) );
AOI221xp5_ASAP7_75t_L g1367 ( .A1(n_44), .A2(n_191), .B1(n_599), .B2(n_1368), .C(n_1370), .Y(n_1367) );
AOI22xp5_ASAP7_75t_L g1889 ( .A1(n_45), .A2(n_1890), .B1(n_1928), .B2(n_1929), .Y(n_1889) );
CKINVDCx5p33_ASAP7_75t_R g1928 ( .A(n_45), .Y(n_1928) );
OAI221xp5_ASAP7_75t_L g1490 ( .A1(n_46), .A2(n_74), .B1(n_650), .B2(n_693), .C(n_694), .Y(n_1490) );
OAI222xp33_ASAP7_75t_L g1516 ( .A1(n_46), .A2(n_74), .B1(n_230), .B2(n_793), .C1(n_1517), .C2(n_1518), .Y(n_1516) );
OAI22xp5_ASAP7_75t_L g583 ( .A1(n_47), .A2(n_64), .B1(n_584), .B2(n_587), .Y(n_583) );
OAI221xp5_ASAP7_75t_L g640 ( .A1(n_47), .A2(n_64), .B1(n_641), .B2(n_647), .C(n_650), .Y(n_640) );
AOI21xp33_ASAP7_75t_L g1905 ( .A1(n_48), .A2(n_750), .B(n_1375), .Y(n_1905) );
AOI221xp5_ASAP7_75t_L g1923 ( .A1(n_48), .A2(n_94), .B1(n_502), .B2(n_639), .C(n_1924), .Y(n_1923) );
INVx1_ASAP7_75t_L g410 ( .A(n_49), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g932 ( .A1(n_50), .A2(n_329), .B1(n_636), .B2(n_933), .Y(n_932) );
OAI22xp5_ASAP7_75t_L g961 ( .A1(n_50), .A2(n_252), .B1(n_962), .B2(n_963), .Y(n_961) );
AOI22xp33_ASAP7_75t_SL g981 ( .A1(n_51), .A2(n_116), .B1(n_458), .B2(n_574), .Y(n_981) );
AOI22xp33_ASAP7_75t_SL g1004 ( .A1(n_51), .A2(n_184), .B1(n_1005), .B2(n_1006), .Y(n_1004) );
AOI221xp5_ASAP7_75t_L g986 ( .A1(n_52), .A2(n_205), .B1(n_574), .B2(n_575), .C(n_987), .Y(n_986) );
OAI21xp33_ASAP7_75t_SL g1001 ( .A1(n_52), .A2(n_1002), .B(n_1003), .Y(n_1001) );
INVx1_ASAP7_75t_L g1065 ( .A(n_53), .Y(n_1065) );
AOI22xp33_ASAP7_75t_L g1075 ( .A1(n_53), .A2(n_321), .B1(n_1005), .B2(n_1076), .Y(n_1075) );
OAI222xp33_ASAP7_75t_L g1154 ( .A1(n_54), .A2(n_181), .B1(n_273), .B2(n_1155), .C1(n_1157), .C2(n_1158), .Y(n_1154) );
AOI221xp5_ASAP7_75t_L g1180 ( .A1(n_54), .A2(n_181), .B1(n_1181), .B2(n_1182), .C(n_1184), .Y(n_1180) );
CKINVDCx5p33_ASAP7_75t_R g1191 ( .A(n_55), .Y(n_1191) );
AOI22xp33_ASAP7_75t_L g1662 ( .A1(n_56), .A2(n_79), .B1(n_1593), .B2(n_1601), .Y(n_1662) );
INVx1_ASAP7_75t_L g705 ( .A(n_57), .Y(n_705) );
INVxp67_ASAP7_75t_SL g1105 ( .A(n_58), .Y(n_1105) );
AOI22xp33_ASAP7_75t_L g1126 ( .A1(n_58), .A2(n_216), .B1(n_579), .B2(n_1127), .Y(n_1126) );
INVx1_ASAP7_75t_L g714 ( .A(n_60), .Y(n_714) );
CKINVDCx5p33_ASAP7_75t_R g1500 ( .A(n_61), .Y(n_1500) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_62), .A2(n_206), .B1(n_456), .B2(n_458), .Y(n_455) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_62), .A2(n_206), .B1(n_555), .B2(n_560), .Y(n_554) );
INVxp67_ASAP7_75t_L g1236 ( .A(n_63), .Y(n_1236) );
INVx1_ASAP7_75t_L g922 ( .A(n_65), .Y(n_922) );
AOI22xp33_ASAP7_75t_L g1852 ( .A1(n_66), .A2(n_176), .B1(n_480), .B2(n_806), .Y(n_1852) );
OAI22xp5_ASAP7_75t_L g1861 ( .A1(n_66), .A2(n_176), .B1(n_609), .B2(n_1054), .Y(n_1861) );
AOI22xp33_ASAP7_75t_L g927 ( .A1(n_67), .A2(n_161), .B1(n_804), .B2(n_928), .Y(n_927) );
AOI221xp5_ASAP7_75t_L g935 ( .A1(n_67), .A2(n_219), .B1(n_936), .B2(n_937), .C(n_939), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g1640 ( .A1(n_68), .A2(n_212), .B1(n_1622), .B2(n_1625), .Y(n_1640) );
AOI22xp33_ASAP7_75t_L g1871 ( .A1(n_69), .A2(n_124), .B1(n_378), .B2(n_964), .Y(n_1871) );
OAI221xp5_ASAP7_75t_L g1900 ( .A1(n_70), .A2(n_152), .B1(n_742), .B2(n_967), .C(n_1901), .Y(n_1900) );
INVx1_ASAP7_75t_L g1927 ( .A(n_70), .Y(n_1927) );
INVxp67_ASAP7_75t_L g1256 ( .A(n_71), .Y(n_1256) );
AOI22xp33_ASAP7_75t_L g1280 ( .A1(n_71), .A2(n_113), .B1(n_735), .B2(n_936), .Y(n_1280) );
AO22x1_ASAP7_75t_SL g1649 ( .A1(n_72), .A2(n_134), .B1(n_1622), .B2(n_1625), .Y(n_1649) );
AOI221xp5_ASAP7_75t_L g807 ( .A1(n_73), .A2(n_211), .B1(n_808), .B2(n_810), .C(n_813), .Y(n_807) );
INVx1_ASAP7_75t_L g680 ( .A(n_75), .Y(n_680) );
CKINVDCx5p33_ASAP7_75t_R g1357 ( .A(n_76), .Y(n_1357) );
CKINVDCx5p33_ASAP7_75t_R g1498 ( .A(n_77), .Y(n_1498) );
AOI21xp33_ASAP7_75t_L g848 ( .A1(n_78), .A2(n_575), .B(n_849), .Y(n_848) );
INVxp33_ASAP7_75t_L g876 ( .A(n_78), .Y(n_876) );
XOR2x2_ASAP7_75t_L g369 ( .A(n_79), .B(n_370), .Y(n_369) );
OAI22xp33_ASAP7_75t_L g1298 ( .A1(n_80), .A2(n_217), .B1(n_1134), .B2(n_1274), .Y(n_1298) );
OAI221xp5_ASAP7_75t_L g1317 ( .A1(n_80), .A2(n_217), .B1(n_694), .B2(n_1099), .C(n_1318), .Y(n_1317) );
INVxp33_ASAP7_75t_L g689 ( .A(n_81), .Y(n_689) );
AOI21xp33_ASAP7_75t_L g734 ( .A1(n_81), .A2(n_735), .B(n_736), .Y(n_734) );
INVxp33_ASAP7_75t_L g401 ( .A(n_82), .Y(n_401) );
INVx1_ASAP7_75t_L g1261 ( .A(n_83), .Y(n_1261) );
AOI22x1_ASAP7_75t_L g976 ( .A1(n_84), .A2(n_977), .B1(n_1030), .B2(n_1031), .Y(n_976) );
INVxp67_ASAP7_75t_L g1030 ( .A(n_84), .Y(n_1030) );
INVxp33_ASAP7_75t_L g690 ( .A(n_85), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g1641 ( .A1(n_86), .A2(n_229), .B1(n_1601), .B2(n_1628), .Y(n_1641) );
INVxp33_ASAP7_75t_L g1547 ( .A(n_87), .Y(n_1547) );
AOI22xp33_ASAP7_75t_L g1572 ( .A1(n_87), .A2(n_276), .B1(n_983), .B2(n_1463), .Y(n_1572) );
AOI22xp33_ASAP7_75t_L g1457 ( .A1(n_88), .A2(n_269), .B1(n_445), .B2(n_1458), .Y(n_1457) );
AOI22xp33_ASAP7_75t_L g1469 ( .A1(n_88), .A2(n_269), .B1(n_1195), .B2(n_1470), .Y(n_1469) );
INVx1_ASAP7_75t_L g914 ( .A(n_89), .Y(n_914) );
CKINVDCx20_ASAP7_75t_R g839 ( .A(n_90), .Y(n_839) );
CKINVDCx5p33_ASAP7_75t_R g1209 ( .A(n_91), .Y(n_1209) );
AOI221xp5_ASAP7_75t_L g572 ( .A1(n_92), .A2(n_333), .B1(n_573), .B2(n_574), .C(n_575), .Y(n_572) );
INVxp33_ASAP7_75t_L g630 ( .A(n_92), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g1199 ( .A1(n_93), .A2(n_187), .B1(n_502), .B2(n_1200), .Y(n_1199) );
OAI22xp5_ASAP7_75t_L g1231 ( .A1(n_93), .A2(n_187), .B1(n_947), .B2(n_1232), .Y(n_1231) );
AOI22xp33_ASAP7_75t_L g1904 ( .A1(n_94), .A2(n_237), .B1(n_732), .B2(n_754), .Y(n_1904) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_95), .A2(n_186), .B1(n_446), .B2(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g823 ( .A(n_95), .Y(n_823) );
OAI221xp5_ASAP7_75t_L g1343 ( .A1(n_96), .A2(n_167), .B1(n_647), .B2(n_693), .C(n_879), .Y(n_1343) );
OAI22xp33_ASAP7_75t_L g1365 ( .A1(n_96), .A2(n_167), .B1(n_1045), .B2(n_1366), .Y(n_1365) );
AOI22xp5_ASAP7_75t_L g1627 ( .A1(n_97), .A2(n_118), .B1(n_1601), .B2(n_1628), .Y(n_1627) );
AOI22xp33_ASAP7_75t_L g597 ( .A1(n_98), .A2(n_297), .B1(n_598), .B2(n_599), .Y(n_597) );
INVxp67_ASAP7_75t_SL g667 ( .A(n_98), .Y(n_667) );
INVx1_ASAP7_75t_L g1136 ( .A(n_99), .Y(n_1136) );
AOI22xp33_ASAP7_75t_SL g576 ( .A1(n_100), .A2(n_227), .B1(n_577), .B2(n_579), .Y(n_576) );
INVxp33_ASAP7_75t_SL g637 ( .A(n_100), .Y(n_637) );
INVx1_ASAP7_75t_L g385 ( .A(n_101), .Y(n_385) );
BUFx2_ASAP7_75t_L g436 ( .A(n_101), .Y(n_436) );
BUFx2_ASAP7_75t_L g462 ( .A(n_101), .Y(n_462) );
OR2x2_ASAP7_75t_L g619 ( .A(n_101), .B(n_479), .Y(n_619) );
INVx1_ASAP7_75t_L g1314 ( .A(n_102), .Y(n_1314) );
AOI22xp33_ASAP7_75t_SL g1849 ( .A1(n_103), .A2(n_148), .B1(n_480), .B2(n_806), .Y(n_1849) );
INVx1_ASAP7_75t_L g1867 ( .A(n_103), .Y(n_1867) );
AOI22xp33_ASAP7_75t_SL g1201 ( .A1(n_104), .A2(n_120), .B1(n_1194), .B2(n_1195), .Y(n_1201) );
INVx1_ASAP7_75t_L g1230 ( .A(n_104), .Y(n_1230) );
INVxp33_ASAP7_75t_L g1550 ( .A(n_105), .Y(n_1550) );
INVx1_ASAP7_75t_L g1610 ( .A(n_106), .Y(n_1610) );
INVxp67_ASAP7_75t_L g1416 ( .A(n_107), .Y(n_1416) );
CKINVDCx5p33_ASAP7_75t_R g836 ( .A(n_108), .Y(n_836) );
AOI221xp5_ASAP7_75t_L g853 ( .A1(n_109), .A2(n_231), .B1(n_854), .B2(n_856), .C(n_859), .Y(n_853) );
INVxp67_ASAP7_75t_SL g888 ( .A(n_109), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g1644 ( .A1(n_110), .A2(n_294), .B1(n_1622), .B2(n_1625), .Y(n_1644) );
AOI221xp5_ASAP7_75t_SL g780 ( .A1(n_111), .A2(n_117), .B1(n_575), .B2(n_781), .C(n_783), .Y(n_780) );
INVx1_ASAP7_75t_L g803 ( .A(n_111), .Y(n_803) );
INVxp33_ASAP7_75t_L g1450 ( .A(n_112), .Y(n_1450) );
AOI22xp33_ASAP7_75t_L g1464 ( .A1(n_112), .A2(n_304), .B1(n_445), .B2(n_573), .Y(n_1464) );
INVxp33_ASAP7_75t_L g1250 ( .A(n_113), .Y(n_1250) );
INVx1_ASAP7_75t_L g776 ( .A(n_114), .Y(n_776) );
AOI22xp5_ASAP7_75t_L g1333 ( .A1(n_115), .A2(n_1334), .B1(n_1383), .B2(n_1384), .Y(n_1333) );
INVx1_ASAP7_75t_L g1383 ( .A(n_115), .Y(n_1383) );
AOI22xp33_ASAP7_75t_L g1657 ( .A1(n_115), .A2(n_259), .B1(n_1593), .B2(n_1601), .Y(n_1657) );
AOI22xp33_ASAP7_75t_L g1008 ( .A1(n_116), .A2(n_129), .B1(n_1009), .B2(n_1010), .Y(n_1008) );
INVx1_ASAP7_75t_L g801 ( .A(n_117), .Y(n_801) );
INVxp67_ASAP7_75t_SL g709 ( .A(n_119), .Y(n_709) );
AOI221xp5_ASAP7_75t_L g746 ( .A1(n_119), .A2(n_303), .B1(n_747), .B2(n_749), .C(n_750), .Y(n_746) );
NOR2xp33_ASAP7_75t_L g1215 ( .A(n_120), .B(n_609), .Y(n_1215) );
OAI22xp5_ASAP7_75t_L g1487 ( .A1(n_121), .A2(n_230), .B1(n_618), .B2(n_1488), .Y(n_1487) );
CKINVDCx5p33_ASAP7_75t_R g1530 ( .A(n_121), .Y(n_1530) );
INVxp33_ASAP7_75t_L g1443 ( .A(n_122), .Y(n_1443) );
AOI22xp33_ASAP7_75t_L g1465 ( .A1(n_122), .A2(n_283), .B1(n_755), .B2(n_1147), .Y(n_1465) );
INVx1_ASAP7_75t_L g1267 ( .A(n_123), .Y(n_1267) );
OAI22xp33_ASAP7_75t_L g1858 ( .A1(n_124), .A2(n_142), .B1(n_618), .B2(n_1488), .Y(n_1858) );
INVxp67_ASAP7_75t_L g1246 ( .A(n_126), .Y(n_1246) );
AOI22xp33_ASAP7_75t_L g1272 ( .A1(n_126), .A2(n_158), .B1(n_731), .B2(n_791), .Y(n_1272) );
INVx1_ASAP7_75t_L g1652 ( .A(n_127), .Y(n_1652) );
AOI22xp33_ASAP7_75t_L g1910 ( .A1(n_128), .A2(n_261), .B1(n_439), .B2(n_460), .Y(n_1910) );
OAI211xp5_ASAP7_75t_L g1912 ( .A1(n_128), .A2(n_1913), .B(n_1914), .C(n_1916), .Y(n_1912) );
AOI221xp5_ASAP7_75t_L g982 ( .A1(n_129), .A2(n_184), .B1(n_788), .B2(n_983), .C(n_984), .Y(n_982) );
INVx1_ASAP7_75t_L g1283 ( .A(n_130), .Y(n_1283) );
CKINVDCx5p33_ASAP7_75t_R g1292 ( .A(n_131), .Y(n_1292) );
INVx1_ASAP7_75t_L g1561 ( .A(n_132), .Y(n_1561) );
AOI221xp5_ASAP7_75t_L g787 ( .A1(n_135), .A2(n_193), .B1(n_595), .B2(n_788), .C(n_789), .Y(n_787) );
AOI221xp5_ASAP7_75t_L g818 ( .A1(n_135), .A2(n_186), .B1(n_819), .B2(n_821), .C(n_822), .Y(n_818) );
INVx1_ASAP7_75t_L g959 ( .A(n_136), .Y(n_959) );
CKINVDCx5p33_ASAP7_75t_R g1359 ( .A(n_137), .Y(n_1359) );
OAI222xp33_ASAP7_75t_L g1159 ( .A1(n_138), .A2(n_202), .B1(n_328), .B2(n_793), .C1(n_1134), .C2(n_1160), .Y(n_1159) );
INVx1_ASAP7_75t_L g1171 ( .A(n_138), .Y(n_1171) );
AOI221xp5_ASAP7_75t_L g1056 ( .A1(n_139), .A2(n_307), .B1(n_861), .B2(n_983), .C(n_1057), .Y(n_1056) );
AOI22xp33_ASAP7_75t_L g1074 ( .A1(n_139), .A2(n_224), .B1(n_671), .B2(n_1005), .Y(n_1074) );
OAI22xp33_ASAP7_75t_L g1896 ( .A1(n_140), .A2(n_310), .B1(n_967), .B2(n_1062), .Y(n_1896) );
AOI22xp33_ASAP7_75t_L g1922 ( .A1(n_140), .A2(n_192), .B1(n_506), .B2(n_802), .Y(n_1922) );
INVxp67_ASAP7_75t_L g1245 ( .A(n_141), .Y(n_1245) );
AOI221xp5_ASAP7_75t_L g1271 ( .A1(n_141), .A2(n_196), .B1(n_573), .B2(n_575), .C(n_849), .Y(n_1271) );
INVx1_ASAP7_75t_L g1874 ( .A(n_142), .Y(n_1874) );
AOI21xp5_ASAP7_75t_L g1911 ( .A1(n_143), .A2(n_735), .B(n_736), .Y(n_1911) );
INVx1_ASAP7_75t_L g1917 ( .A(n_143), .Y(n_1917) );
OAI22xp5_ASAP7_75t_L g1894 ( .A1(n_144), .A2(n_192), .B1(n_962), .B2(n_1895), .Y(n_1894) );
AOI22xp5_ASAP7_75t_L g1921 ( .A1(n_144), .A2(n_310), .B1(n_627), .B2(n_1198), .Y(n_1921) );
CKINVDCx5p33_ASAP7_75t_R g1289 ( .A(n_145), .Y(n_1289) );
OAI221xp5_ASAP7_75t_L g1098 ( .A1(n_146), .A2(n_179), .B1(n_641), .B2(n_648), .C(n_1099), .Y(n_1098) );
OAI22xp33_ASAP7_75t_L g1133 ( .A1(n_146), .A2(n_179), .B1(n_841), .B2(n_1134), .Y(n_1133) );
INVx1_ASAP7_75t_L g916 ( .A(n_147), .Y(n_916) );
INVx1_ASAP7_75t_L g1864 ( .A(n_148), .Y(n_1864) );
XNOR2xp5_ASAP7_75t_L g1542 ( .A(n_149), .B(n_1543), .Y(n_1542) );
CKINVDCx5p33_ASAP7_75t_R g1903 ( .A(n_150), .Y(n_1903) );
OAI221xp5_ASAP7_75t_L g1247 ( .A1(n_151), .A2(n_190), .B1(n_650), .B2(n_693), .C(n_694), .Y(n_1247) );
OAI22xp5_ASAP7_75t_L g1273 ( .A1(n_151), .A2(n_190), .B1(n_1274), .B2(n_1275), .Y(n_1273) );
INVx1_ASAP7_75t_L g1915 ( .A(n_152), .Y(n_1915) );
INVx1_ASAP7_75t_L g778 ( .A(n_153), .Y(n_778) );
AOI221xp5_ASAP7_75t_L g1146 ( .A1(n_154), .A2(n_302), .B1(n_861), .B2(n_954), .C(n_1147), .Y(n_1146) );
INVx1_ASAP7_75t_L g1179 ( .A(n_154), .Y(n_1179) );
CKINVDCx5p33_ASAP7_75t_R g1503 ( .A(n_155), .Y(n_1503) );
INVx1_ASAP7_75t_L g1418 ( .A(n_156), .Y(n_1418) );
OAI22xp5_ASAP7_75t_L g1436 ( .A1(n_156), .A2(n_288), .B1(n_1437), .B2(n_1439), .Y(n_1436) );
CKINVDCx5p33_ASAP7_75t_R g1362 ( .A(n_157), .Y(n_1362) );
INVxp67_ASAP7_75t_L g1241 ( .A(n_158), .Y(n_1241) );
INVx1_ASAP7_75t_L g1598 ( .A(n_159), .Y(n_1598) );
CKINVDCx5p33_ASAP7_75t_R g723 ( .A(n_160), .Y(n_723) );
INVx1_ASAP7_75t_L g942 ( .A(n_161), .Y(n_942) );
INVx1_ASAP7_75t_L g1218 ( .A(n_162), .Y(n_1218) );
AOI221xp5_ASAP7_75t_L g1591 ( .A1(n_163), .A2(n_247), .B1(n_1592), .B2(n_1599), .C(n_1602), .Y(n_1591) );
INVx1_ASAP7_75t_L g687 ( .A(n_164), .Y(n_687) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_164), .B(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g423 ( .A(n_165), .Y(n_423) );
INVxp67_ASAP7_75t_L g1559 ( .A(n_166), .Y(n_1559) );
AOI22xp33_ASAP7_75t_L g1579 ( .A1(n_166), .A2(n_207), .B1(n_1127), .B2(n_1580), .Y(n_1579) );
INVx1_ASAP7_75t_L g1596 ( .A(n_168), .Y(n_1596) );
NAND2xp5_ASAP7_75t_L g1614 ( .A(n_168), .B(n_1609), .Y(n_1614) );
AOI22xp33_ASAP7_75t_L g785 ( .A1(n_169), .A2(n_248), .B1(n_577), .B2(n_599), .Y(n_785) );
OAI221xp5_ASAP7_75t_L g798 ( .A1(n_169), .A2(n_248), .B1(n_496), .B2(n_799), .C(n_800), .Y(n_798) );
AOI22xp33_ASAP7_75t_SL g437 ( .A1(n_170), .A2(n_197), .B1(n_438), .B2(n_440), .Y(n_437) );
INVxp67_ASAP7_75t_SL g533 ( .A(n_170), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g1058 ( .A1(n_171), .A2(n_224), .B1(n_1059), .B2(n_1061), .Y(n_1058) );
AOI22xp33_ASAP7_75t_SL g1072 ( .A1(n_171), .A2(n_307), .B1(n_802), .B2(n_1073), .Y(n_1072) );
AOI21xp5_ASAP7_75t_L g1050 ( .A1(n_172), .A2(n_849), .B(n_1051), .Y(n_1050) );
INVx1_ASAP7_75t_L g1083 ( .A(n_172), .Y(n_1083) );
INVx1_ASAP7_75t_L g1565 ( .A(n_173), .Y(n_1565) );
INVx2_ASAP7_75t_L g361 ( .A(n_174), .Y(n_361) );
OAI22x1_ASAP7_75t_SL g1392 ( .A1(n_175), .A2(n_1393), .B1(n_1480), .B2(n_1481), .Y(n_1392) );
INVx1_ASAP7_75t_L g1480 ( .A(n_175), .Y(n_1480) );
AO221x2_ASAP7_75t_L g1632 ( .A1(n_175), .A2(n_221), .B1(n_1593), .B2(n_1633), .C(n_1634), .Y(n_1632) );
AOI221xp5_ASAP7_75t_L g590 ( .A1(n_177), .A2(n_322), .B1(n_578), .B2(n_591), .C(n_595), .Y(n_590) );
INVxp33_ASAP7_75t_SL g660 ( .A(n_177), .Y(n_660) );
BUFx3_ASAP7_75t_L g380 ( .A(n_178), .Y(n_380) );
INVx1_ASAP7_75t_L g392 ( .A(n_178), .Y(n_392) );
INVx1_ASAP7_75t_L g989 ( .A(n_180), .Y(n_989) );
INVx1_ASAP7_75t_L g1346 ( .A(n_182), .Y(n_1346) );
AOI22xp33_ASAP7_75t_L g1380 ( .A1(n_182), .A2(n_286), .B1(n_448), .B2(n_753), .Y(n_1380) );
INVx1_ASAP7_75t_L g386 ( .A(n_183), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g1878 ( .A(n_185), .Y(n_1878) );
INVx1_ASAP7_75t_L g716 ( .A(n_188), .Y(n_716) );
INVxp33_ASAP7_75t_L g1096 ( .A(n_189), .Y(n_1096) );
AOI221xp5_ASAP7_75t_L g1131 ( .A1(n_189), .A2(n_228), .B1(n_735), .B2(n_736), .C(n_954), .Y(n_1131) );
INVx1_ASAP7_75t_L g1338 ( .A(n_191), .Y(n_1338) );
INVx1_ASAP7_75t_L g824 ( .A(n_193), .Y(n_824) );
OAI221xp5_ASAP7_75t_SL g840 ( .A1(n_194), .A2(n_332), .B1(n_587), .B2(n_841), .C(n_843), .Y(n_840) );
OAI221xp5_ASAP7_75t_L g878 ( .A1(n_194), .A2(n_332), .B1(n_648), .B2(n_693), .C(n_879), .Y(n_878) );
INVxp67_ASAP7_75t_SL g990 ( .A(n_195), .Y(n_990) );
INVxp67_ASAP7_75t_L g1242 ( .A(n_196), .Y(n_1242) );
INVxp67_ASAP7_75t_SL g544 ( .A(n_197), .Y(n_544) );
INVx1_ASAP7_75t_L g777 ( .A(n_198), .Y(n_777) );
CKINVDCx5p33_ASAP7_75t_R g1501 ( .A(n_200), .Y(n_1501) );
CKINVDCx5p33_ASAP7_75t_R g469 ( .A(n_201), .Y(n_469) );
INVx1_ASAP7_75t_L g1164 ( .A(n_202), .Y(n_1164) );
INVxp33_ASAP7_75t_SL g909 ( .A(n_203), .Y(n_909) );
AOI221xp5_ASAP7_75t_L g945 ( .A1(n_203), .A2(n_254), .B1(n_936), .B2(n_946), .C(n_948), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g1145 ( .A1(n_204), .A2(n_291), .B1(n_456), .B2(n_1061), .Y(n_1145) );
INVx1_ASAP7_75t_L g1169 ( .A(n_204), .Y(n_1169) );
INVxp33_ASAP7_75t_SL g1019 ( .A(n_205), .Y(n_1019) );
INVxp33_ASAP7_75t_L g1555 ( .A(n_207), .Y(n_1555) );
INVx1_ASAP7_75t_L g867 ( .A(n_208), .Y(n_867) );
INVx1_ASAP7_75t_L g384 ( .A(n_209), .Y(n_384) );
INVx1_ASAP7_75t_L g434 ( .A(n_209), .Y(n_434) );
INVxp33_ASAP7_75t_L g1413 ( .A(n_210), .Y(n_1413) );
INVx1_ASAP7_75t_L g774 ( .A(n_211), .Y(n_774) );
INVxp33_ASAP7_75t_SL g1093 ( .A(n_213), .Y(n_1093) );
AOI22xp33_ASAP7_75t_L g1132 ( .A1(n_213), .A2(n_218), .B1(n_789), .B2(n_964), .Y(n_1132) );
INVx1_ASAP7_75t_L g713 ( .A(n_214), .Y(n_713) );
INVx1_ASAP7_75t_L g582 ( .A(n_215), .Y(n_582) );
INVx1_ASAP7_75t_L g1110 ( .A(n_216), .Y(n_1110) );
INVxp33_ASAP7_75t_SL g1097 ( .A(n_218), .Y(n_1097) );
INVx1_ASAP7_75t_L g926 ( .A(n_219), .Y(n_926) );
CKINVDCx5p33_ASAP7_75t_R g1907 ( .A(n_220), .Y(n_1907) );
AOI22xp33_ASAP7_75t_SL g451 ( .A1(n_222), .A2(n_282), .B1(n_440), .B2(n_452), .Y(n_451) );
OAI211xp5_ASAP7_75t_SL g484 ( .A1(n_222), .A2(n_485), .B(n_495), .C(n_515), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g1621 ( .A1(n_223), .A2(n_267), .B1(n_1622), .B2(n_1625), .Y(n_1621) );
XOR2xp5_ASAP7_75t_L g1840 ( .A(n_223), .B(n_1841), .Y(n_1840) );
AOI22xp33_ASAP7_75t_L g1883 ( .A1(n_223), .A2(n_1884), .B1(n_1888), .B2(n_1930), .Y(n_1883) );
INVx1_ASAP7_75t_L g1086 ( .A(n_225), .Y(n_1086) );
AOI22xp5_ASAP7_75t_L g1645 ( .A1(n_225), .A2(n_295), .B1(n_1601), .B2(n_1628), .Y(n_1645) );
AOI221xp5_ASAP7_75t_L g1144 ( .A1(n_226), .A2(n_308), .B1(n_575), .B2(n_781), .C(n_783), .Y(n_1144) );
INVx1_ASAP7_75t_L g1167 ( .A(n_226), .Y(n_1167) );
INVxp33_ASAP7_75t_L g624 ( .A(n_227), .Y(n_624) );
INVxp33_ASAP7_75t_L g1094 ( .A(n_228), .Y(n_1094) );
INVx1_ASAP7_75t_L g885 ( .A(n_231), .Y(n_885) );
CKINVDCx5p33_ASAP7_75t_R g1190 ( .A(n_232), .Y(n_1190) );
AOI22xp33_ASAP7_75t_L g1296 ( .A1(n_233), .A2(n_239), .B1(n_983), .B2(n_1297), .Y(n_1296) );
INVx1_ASAP7_75t_L g1310 ( .A(n_233), .Y(n_1310) );
INVx1_ASAP7_75t_L g1325 ( .A(n_234), .Y(n_1325) );
INVxp67_ASAP7_75t_L g1253 ( .A(n_235), .Y(n_1253) );
AOI221xp5_ASAP7_75t_L g1277 ( .A1(n_235), .A2(n_249), .B1(n_457), .B2(n_1278), .C(n_1279), .Y(n_1277) );
AOI22xp33_ASAP7_75t_L g862 ( .A1(n_236), .A2(n_298), .B1(n_863), .B2(n_864), .Y(n_862) );
INVx1_ASAP7_75t_L g884 ( .A(n_236), .Y(n_884) );
INVx1_ASAP7_75t_L g1925 ( .A(n_237), .Y(n_1925) );
INVxp67_ASAP7_75t_L g1558 ( .A(n_238), .Y(n_1558) );
AOI221xp5_ASAP7_75t_L g1577 ( .A1(n_238), .A2(n_338), .B1(n_595), .B2(n_788), .C(n_1578), .Y(n_1577) );
INVx1_ASAP7_75t_L g1315 ( .A(n_239), .Y(n_1315) );
INVx1_ASAP7_75t_L g1653 ( .A(n_240), .Y(n_1653) );
XNOR2xp5_ASAP7_75t_L g1284 ( .A(n_241), .B(n_1285), .Y(n_1284) );
OAI211xp5_ASAP7_75t_SL g991 ( .A1(n_242), .A2(n_992), .B(n_993), .C(n_998), .Y(n_991) );
INVx1_ASAP7_75t_L g1027 ( .A(n_242), .Y(n_1027) );
INVx1_ASAP7_75t_L g1213 ( .A(n_243), .Y(n_1213) );
OAI211xp5_ASAP7_75t_L g1228 ( .A1(n_243), .A2(n_793), .B(n_1229), .C(n_1233), .Y(n_1228) );
CKINVDCx5p33_ASAP7_75t_R g1528 ( .A(n_244), .Y(n_1528) );
CKINVDCx5p33_ASAP7_75t_R g1504 ( .A(n_245), .Y(n_1504) );
CKINVDCx20_ASAP7_75t_R g1635 ( .A(n_246), .Y(n_1635) );
INVxp33_ASAP7_75t_L g1251 ( .A(n_249), .Y(n_1251) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_250), .A2(n_257), .B1(n_457), .B2(n_460), .Y(n_847) );
INVxp33_ASAP7_75t_L g877 ( .A(n_250), .Y(n_877) );
INVx1_ASAP7_75t_L g1351 ( .A(n_251), .Y(n_1351) );
AOI221xp5_ASAP7_75t_L g1374 ( .A1(n_251), .A2(n_263), .B1(n_1279), .B2(n_1375), .C(n_1376), .Y(n_1374) );
INVxp67_ASAP7_75t_SL g931 ( .A(n_252), .Y(n_931) );
XNOR2x1_ASAP7_75t_L g1140 ( .A(n_253), .B(n_1141), .Y(n_1140) );
INVxp33_ASAP7_75t_SL g913 ( .A(n_254), .Y(n_913) );
INVx1_ASAP7_75t_L g379 ( .A(n_255), .Y(n_379) );
BUFx3_ASAP7_75t_L g391 ( .A(n_255), .Y(n_391) );
CKINVDCx5p33_ASAP7_75t_R g1496 ( .A(n_256), .Y(n_1496) );
INVxp33_ASAP7_75t_L g873 ( .A(n_257), .Y(n_873) );
INVx1_ASAP7_75t_L g899 ( .A(n_258), .Y(n_899) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_260), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_260), .B(n_326), .Y(n_479) );
AND2x2_ASAP7_75t_L g489 ( .A(n_260), .B(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g514 ( .A(n_260), .Y(n_514) );
INVx1_ASAP7_75t_L g1918 ( .A(n_261), .Y(n_1918) );
OAI332xp33_ASAP7_75t_L g1491 ( .A1(n_262), .A2(n_653), .A3(n_677), .B1(n_1492), .B2(n_1495), .B3(n_1499), .C1(n_1502), .C2(n_1505), .Y(n_1491) );
INVx1_ASAP7_75t_L g1534 ( .A(n_262), .Y(n_1534) );
INVx1_ASAP7_75t_L g1349 ( .A(n_263), .Y(n_1349) );
INVx1_ASAP7_75t_L g607 ( .A(n_264), .Y(n_607) );
INVx1_ASAP7_75t_L g958 ( .A(n_265), .Y(n_958) );
OR2x2_ASAP7_75t_L g383 ( .A(n_266), .B(n_384), .Y(n_383) );
INVx2_ASAP7_75t_L g421 ( .A(n_266), .Y(n_421) );
INVx1_ASAP7_75t_L g1081 ( .A(n_268), .Y(n_1081) );
CKINVDCx5p33_ASAP7_75t_R g1494 ( .A(n_270), .Y(n_1494) );
INVx1_ASAP7_75t_L g1259 ( .A(n_271), .Y(n_1259) );
AOI22xp33_ASAP7_75t_L g1851 ( .A1(n_272), .A2(n_289), .B1(n_557), .B2(n_1264), .Y(n_1851) );
OAI22xp5_ASAP7_75t_L g1860 ( .A1(n_272), .A2(n_289), .B1(n_613), .B2(n_1122), .Y(n_1860) );
INVx1_ASAP7_75t_L g1185 ( .A(n_273), .Y(n_1185) );
CKINVDCx16_ASAP7_75t_R g765 ( .A(n_274), .Y(n_765) );
INVx1_ASAP7_75t_L g1113 ( .A(n_275), .Y(n_1113) );
INVxp33_ASAP7_75t_SL g1551 ( .A(n_276), .Y(n_1551) );
INVx1_ASAP7_75t_L g1066 ( .A(n_277), .Y(n_1066) );
INVx1_ASAP7_75t_L g611 ( .A(n_278), .Y(n_611) );
INVx1_ASAP7_75t_L g1846 ( .A(n_279), .Y(n_1846) );
AOI21xp33_ASAP7_75t_L g1865 ( .A1(n_279), .A2(n_861), .B(n_944), .Y(n_1865) );
INVxp67_ASAP7_75t_SL g994 ( .A(n_280), .Y(n_994) );
OAI211xp5_ASAP7_75t_SL g1012 ( .A1(n_280), .A2(n_700), .B(n_1013), .C(n_1016), .Y(n_1012) );
INVx1_ASAP7_75t_L g852 ( .A(n_281), .Y(n_852) );
OAI221xp5_ASAP7_75t_L g523 ( .A1(n_282), .A2(n_524), .B1(n_526), .B2(n_540), .C(n_551), .Y(n_523) );
INVxp67_ASAP7_75t_L g1447 ( .A(n_283), .Y(n_1447) );
INVx1_ASAP7_75t_L g1409 ( .A(n_284), .Y(n_1409) );
AOI22xp33_ASAP7_75t_L g1148 ( .A1(n_285), .A2(n_305), .B1(n_579), .B2(n_1149), .Y(n_1148) );
INVx1_ASAP7_75t_L g1178 ( .A(n_285), .Y(n_1178) );
INVx1_ASAP7_75t_L g1354 ( .A(n_286), .Y(n_1354) );
INVx1_ASAP7_75t_L g678 ( .A(n_287), .Y(n_678) );
INVx1_ASAP7_75t_L g1423 ( .A(n_288), .Y(n_1423) );
INVx1_ASAP7_75t_L g1204 ( .A(n_290), .Y(n_1204) );
AOI21xp5_ASAP7_75t_L g1225 ( .A1(n_290), .A2(n_754), .B(n_1226), .Y(n_1225) );
INVx1_ASAP7_75t_L g1166 ( .A(n_291), .Y(n_1166) );
CKINVDCx5p33_ASAP7_75t_R g1341 ( .A(n_292), .Y(n_1341) );
INVxp33_ASAP7_75t_L g1020 ( .A(n_293), .Y(n_1020) );
AOI22xp33_ASAP7_75t_L g1461 ( .A1(n_296), .A2(n_313), .B1(n_1462), .B2(n_1463), .Y(n_1461) );
AOI22xp33_ASAP7_75t_L g1471 ( .A1(n_296), .A2(n_313), .B1(n_1472), .B2(n_1473), .Y(n_1471) );
INVxp33_ASAP7_75t_L g657 ( .A(n_297), .Y(n_657) );
INVx1_ASAP7_75t_L g891 ( .A(n_298), .Y(n_891) );
INVx1_ASAP7_75t_L g718 ( .A(n_299), .Y(n_718) );
CKINVDCx5p33_ASAP7_75t_R g1356 ( .A(n_300), .Y(n_1356) );
INVx1_ASAP7_75t_L g1208 ( .A(n_301), .Y(n_1208) );
AOI221xp5_ASAP7_75t_L g1175 ( .A1(n_302), .A2(n_305), .B1(n_808), .B2(n_1176), .C(n_1177), .Y(n_1175) );
INVxp33_ASAP7_75t_L g699 ( .A(n_303), .Y(n_699) );
INVxp67_ASAP7_75t_L g1430 ( .A(n_304), .Y(n_1430) );
AOI22xp33_ASAP7_75t_L g1302 ( .A1(n_306), .A2(n_334), .B1(n_574), .B2(n_964), .Y(n_1302) );
INVx1_ASAP7_75t_L g1327 ( .A(n_306), .Y(n_1327) );
INVx1_ASAP7_75t_L g1174 ( .A(n_308), .Y(n_1174) );
CKINVDCx5p33_ASAP7_75t_R g1153 ( .A(n_309), .Y(n_1153) );
INVx1_ASAP7_75t_L g1266 ( .A(n_311), .Y(n_1266) );
INVx1_ASAP7_75t_L g615 ( .A(n_312), .Y(n_615) );
INVx1_ASAP7_75t_L g844 ( .A(n_314), .Y(n_844) );
INVx1_ASAP7_75t_L g1064 ( .A(n_315), .Y(n_1064) );
INVx1_ASAP7_75t_L g1088 ( .A(n_316), .Y(n_1088) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_317), .Y(n_351) );
AND3x2_ASAP7_75t_L g1597 ( .A(n_317), .B(n_349), .C(n_1598), .Y(n_1597) );
NAND2xp5_ASAP7_75t_L g1607 ( .A(n_317), .B(n_349), .Y(n_1607) );
INVx2_ASAP7_75t_L g362 ( .A(n_319), .Y(n_362) );
XNOR2x2_ASAP7_75t_L g905 ( .A(n_320), .B(n_906), .Y(n_905) );
INVx1_ASAP7_75t_L g1043 ( .A(n_321), .Y(n_1043) );
INVxp67_ASAP7_75t_SL g663 ( .A(n_322), .Y(n_663) );
INVx1_ASAP7_75t_L g911 ( .A(n_323), .Y(n_911) );
CKINVDCx5p33_ASAP7_75t_R g1493 ( .A(n_324), .Y(n_1493) );
INVx1_ASAP7_75t_L g1116 ( .A(n_325), .Y(n_1116) );
INVx1_ASAP7_75t_L g364 ( .A(n_326), .Y(n_364) );
INVx2_ASAP7_75t_L g490 ( .A(n_326), .Y(n_490) );
INVxp67_ASAP7_75t_SL g1109 ( .A(n_327), .Y(n_1109) );
INVx1_ASAP7_75t_L g1163 ( .A(n_328), .Y(n_1163) );
OAI22xp33_ASAP7_75t_L g965 ( .A1(n_329), .A2(n_339), .B1(n_966), .B2(n_967), .Y(n_965) );
INVxp67_ASAP7_75t_SL g550 ( .A(n_330), .Y(n_550) );
INVx1_ASAP7_75t_L g1114 ( .A(n_331), .Y(n_1114) );
INVxp33_ASAP7_75t_L g634 ( .A(n_333), .Y(n_634) );
INVx1_ASAP7_75t_L g1322 ( .A(n_334), .Y(n_1322) );
INVx1_ASAP7_75t_L g996 ( .A(n_335), .Y(n_996) );
INVx1_ASAP7_75t_L g1582 ( .A(n_336), .Y(n_1582) );
CKINVDCx5p33_ASAP7_75t_R g1290 ( .A(n_337), .Y(n_1290) );
INVxp33_ASAP7_75t_L g1556 ( .A(n_338), .Y(n_1556) );
INVxp67_ASAP7_75t_SL g930 ( .A(n_339), .Y(n_930) );
INVx1_ASAP7_75t_L g866 ( .A(n_340), .Y(n_866) );
INVx1_ASAP7_75t_L g1117 ( .A(n_341), .Y(n_1117) );
CKINVDCx5p33_ASAP7_75t_R g1049 ( .A(n_342), .Y(n_1049) );
INVx1_ASAP7_75t_L g1069 ( .A(n_343), .Y(n_1069) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_365), .B(n_1584), .Y(n_344) );
BUFx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x4_ASAP7_75t_L g346 ( .A(n_347), .B(n_352), .Y(n_346) );
AND2x4_ASAP7_75t_L g1882 ( .A(n_347), .B(n_353), .Y(n_1882) );
NOR2xp33_ASAP7_75t_SL g347 ( .A(n_348), .B(n_350), .Y(n_347) );
INVx1_ASAP7_75t_SL g1887 ( .A(n_348), .Y(n_1887) );
NAND2xp5_ASAP7_75t_L g1932 ( .A(n_348), .B(n_350), .Y(n_1932) );
HB1xp67_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g1886 ( .A(n_350), .B(n_1887), .Y(n_1886) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_354), .B(n_358), .Y(n_353) );
INVxp67_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OR2x2_ASAP7_75t_L g1453 ( .A(n_355), .B(n_462), .Y(n_1453) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g539 ( .A(n_356), .B(n_364), .Y(n_539) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
OR2x2_ASAP7_75t_L g654 ( .A(n_357), .B(n_655), .Y(n_654) );
INVx8_ASAP7_75t_L g1449 ( .A(n_358), .Y(n_1449) );
OR2x6_ASAP7_75t_L g358 ( .A(n_359), .B(n_363), .Y(n_358) );
INVx2_ASAP7_75t_SL g535 ( .A(n_359), .Y(n_535) );
OR2x2_ASAP7_75t_L g618 ( .A(n_359), .B(n_619), .Y(n_618) );
BUFx6f_ASAP7_75t_L g659 ( .A(n_359), .Y(n_659) );
INVx2_ASAP7_75t_SL g704 ( .A(n_359), .Y(n_704) );
INVx1_ASAP7_75t_L g883 ( .A(n_359), .Y(n_883) );
BUFx2_ASAP7_75t_L g1015 ( .A(n_359), .Y(n_1015) );
OAI22xp33_ASAP7_75t_L g1184 ( .A1(n_359), .A2(n_529), .B1(n_1153), .B2(n_1185), .Y(n_1184) );
OR2x6_ASAP7_75t_L g1452 ( .A(n_359), .B(n_1442), .Y(n_1452) );
OAI22xp5_ASAP7_75t_L g1924 ( .A1(n_359), .A2(n_529), .B1(n_1903), .B2(n_1925), .Y(n_1924) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_361), .B(n_362), .Y(n_360) );
AND2x2_ASAP7_75t_L g482 ( .A(n_361), .B(n_362), .Y(n_482) );
INVx1_ASAP7_75t_L g493 ( .A(n_361), .Y(n_493) );
INVx2_ASAP7_75t_L g500 ( .A(n_361), .Y(n_500) );
AND2x4_ASAP7_75t_L g503 ( .A(n_361), .B(n_494), .Y(n_503) );
INVx1_ASAP7_75t_L g532 ( .A(n_361), .Y(n_532) );
INVx2_ASAP7_75t_L g494 ( .A(n_362), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_362), .B(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g519 ( .A(n_362), .Y(n_519) );
INVx1_ASAP7_75t_L g531 ( .A(n_362), .Y(n_531) );
INVx1_ASAP7_75t_L g559 ( .A(n_362), .Y(n_559) );
AND2x4_ASAP7_75t_L g1438 ( .A(n_363), .B(n_519), .Y(n_1438) );
INVx2_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
OR2x2_ASAP7_75t_L g1439 ( .A(n_364), .B(n_830), .Y(n_1439) );
XNOR2xp5_ASAP7_75t_L g365 ( .A(n_366), .B(n_1387), .Y(n_365) );
AOI22xp5_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_1033), .B1(n_1034), .B2(n_1386), .Y(n_366) );
INVx1_ASAP7_75t_L g1386 ( .A(n_367), .Y(n_1386) );
XNOR2xp5_ASAP7_75t_L g367 ( .A(n_368), .B(n_760), .Y(n_367) );
XNOR2x1_ASAP7_75t_L g368 ( .A(n_369), .B(n_565), .Y(n_368) );
NAND3xp33_ASAP7_75t_L g370 ( .A(n_371), .B(n_468), .C(n_483), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_372), .B(n_408), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_393), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_375), .B1(n_386), .B2(n_387), .Y(n_373) );
OAI221xp5_ASAP7_75t_L g495 ( .A1(n_374), .A2(n_386), .B1(n_496), .B2(n_501), .C(n_504), .Y(n_495) );
AND2x2_ASAP7_75t_L g375 ( .A(n_376), .B(n_381), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g1301 ( .A(n_377), .Y(n_1301) );
INVx2_ASAP7_75t_SL g1375 ( .A(n_377), .Y(n_1375) );
INVx2_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
BUFx3_ASAP7_75t_L g439 ( .A(n_378), .Y(n_439) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_378), .Y(n_457) );
BUFx6f_ASAP7_75t_L g578 ( .A(n_378), .Y(n_578) );
BUFx2_ASAP7_75t_L g731 ( .A(n_378), .Y(n_731) );
BUFx6f_ASAP7_75t_L g775 ( .A(n_378), .Y(n_775) );
BUFx2_ASAP7_75t_L g789 ( .A(n_378), .Y(n_789) );
BUFx6f_ASAP7_75t_L g944 ( .A(n_378), .Y(n_944) );
HB1xp67_ASAP7_75t_L g1147 ( .A(n_378), .Y(n_1147) );
AND2x6_ASAP7_75t_L g1405 ( .A(n_378), .B(n_1406), .Y(n_1405) );
HB1xp67_ASAP7_75t_L g1578 ( .A(n_378), .Y(n_1578) );
AND2x4_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
INVx1_ASAP7_75t_L g407 ( .A(n_379), .Y(n_407) );
INVx2_ASAP7_75t_L g399 ( .A(n_380), .Y(n_399) );
AND2x2_ASAP7_75t_L g443 ( .A(n_380), .B(n_391), .Y(n_443) );
AND2x2_ASAP7_75t_L g395 ( .A(n_381), .B(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
OR2x6_ASAP7_75t_L g388 ( .A(n_382), .B(n_389), .Y(n_388) );
OR2x6_ASAP7_75t_L g403 ( .A(n_382), .B(n_404), .Y(n_403) );
OR2x2_ASAP7_75t_L g382 ( .A(n_383), .B(n_385), .Y(n_382) );
INVx2_ASAP7_75t_L g581 ( .A(n_383), .Y(n_581) );
OR2x2_ASAP7_75t_L g609 ( .A(n_383), .B(n_610), .Y(n_609) );
OR2x2_ASAP7_75t_L g613 ( .A(n_383), .B(n_614), .Y(n_613) );
A2O1A1Ixp33_ASAP7_75t_SL g1507 ( .A1(n_383), .A2(n_1508), .B(n_1511), .C(n_1515), .Y(n_1507) );
INVx1_ASAP7_75t_L g419 ( .A(n_384), .Y(n_419) );
INVx1_ASAP7_75t_L g422 ( .A(n_385), .Y(n_422) );
AND2x4_ASAP7_75t_L g629 ( .A(n_385), .B(n_489), .Y(n_629) );
CKINVDCx6p67_ASAP7_75t_R g387 ( .A(n_388), .Y(n_387) );
INVx2_ASAP7_75t_L g1510 ( .A(n_389), .Y(n_1510) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
BUFx6f_ASAP7_75t_L g450 ( .A(n_390), .Y(n_450) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_390), .Y(n_460) );
INVx1_ASAP7_75t_L g600 ( .A(n_390), .Y(n_600) );
INVx2_ASAP7_75t_L g614 ( .A(n_390), .Y(n_614) );
AND2x4_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .Y(n_390) );
INVx2_ASAP7_75t_L g400 ( .A(n_391), .Y(n_400) );
INVx1_ASAP7_75t_L g406 ( .A(n_392), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_395), .B1(n_401), .B2(n_402), .Y(n_393) );
A2O1A1Ixp33_ASAP7_75t_L g1873 ( .A1(n_396), .A2(n_955), .B(n_1874), .C(n_1875), .Y(n_1873) );
INVx2_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g598 ( .A(n_397), .Y(n_598) );
INVx1_ASAP7_75t_L g1294 ( .A(n_397), .Y(n_1294) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx6_ASAP7_75t_L g447 ( .A(n_398), .Y(n_447) );
AND2x2_ASAP7_75t_L g472 ( .A(n_398), .B(n_418), .Y(n_472) );
BUFx2_ASAP7_75t_L g735 ( .A(n_398), .Y(n_735) );
AND2x4_ASAP7_75t_L g1410 ( .A(n_398), .B(n_1411), .Y(n_1410) );
AND2x4_ASAP7_75t_L g398 ( .A(n_399), .B(n_400), .Y(n_398) );
INVx1_ASAP7_75t_L g428 ( .A(n_399), .Y(n_428) );
INVx1_ASAP7_75t_L g415 ( .A(n_400), .Y(n_415) );
CKINVDCx6p67_ASAP7_75t_R g402 ( .A(n_403), .Y(n_402) );
BUFx3_ASAP7_75t_L g1223 ( .A(n_404), .Y(n_1223) );
OAI21xp33_ASAP7_75t_L g1863 ( .A1(n_404), .A2(n_1864), .B(n_1865), .Y(n_1863) );
INVx1_ASAP7_75t_L g1909 ( .A(n_404), .Y(n_1909) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g740 ( .A(n_405), .Y(n_740) );
BUFx4f_ASAP7_75t_L g846 ( .A(n_405), .Y(n_846) );
BUFx2_ASAP7_75t_L g941 ( .A(n_405), .Y(n_941) );
INVx1_ASAP7_75t_L g1156 ( .A(n_405), .Y(n_1156) );
INVx1_ASAP7_75t_L g1870 ( .A(n_405), .Y(n_1870) );
AND2x2_ASAP7_75t_L g405 ( .A(n_406), .B(n_407), .Y(n_405) );
OR2x2_ASAP7_75t_L g610 ( .A(n_406), .B(n_407), .Y(n_610) );
NAND3xp33_ASAP7_75t_SL g408 ( .A(n_409), .B(n_429), .C(n_464), .Y(n_408) );
AOI22xp33_ASAP7_75t_L g409 ( .A1(n_410), .A2(n_411), .B1(n_423), .B2(n_424), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_410), .A2(n_423), .B1(n_516), .B2(n_520), .Y(n_515) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
NAND2x1p5_ASAP7_75t_L g412 ( .A(n_413), .B(n_416), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx2_ASAP7_75t_L g586 ( .A(n_414), .Y(n_586) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g1422 ( .A(n_415), .Y(n_1422) );
INVx2_ASAP7_75t_SL g416 ( .A(n_417), .Y(n_416) );
OR2x6_ASAP7_75t_L g425 ( .A(n_417), .B(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g467 ( .A(n_417), .Y(n_467) );
NAND2x1p5_ASAP7_75t_L g417 ( .A(n_418), .B(n_422), .Y(n_417) );
AND2x4_ASAP7_75t_L g585 ( .A(n_418), .B(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g588 ( .A(n_418), .B(n_427), .Y(n_588) );
INVx1_ASAP7_75t_L g605 ( .A(n_418), .Y(n_605) );
AND2x4_ASAP7_75t_L g842 ( .A(n_418), .B(n_586), .Y(n_842) );
BUFx2_ASAP7_75t_L g956 ( .A(n_418), .Y(n_956) );
AND2x2_ASAP7_75t_L g997 ( .A(n_418), .B(n_427), .Y(n_997) );
AND2x4_ASAP7_75t_L g1135 ( .A(n_418), .B(n_427), .Y(n_1135) );
AND2x4_ASAP7_75t_L g418 ( .A(n_419), .B(n_420), .Y(n_418) );
AND2x4_ASAP7_75t_L g463 ( .A(n_420), .B(n_434), .Y(n_463) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g433 ( .A(n_421), .B(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g1402 ( .A(n_421), .Y(n_1402) );
INVx1_ASAP7_75t_L g1407 ( .A(n_421), .Y(n_1407) );
HB1xp67_ASAP7_75t_L g1412 ( .A(n_421), .Y(n_1412) );
OR2x6_ASAP7_75t_L g677 ( .A(n_422), .B(n_512), .Y(n_677) );
INVx2_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
OR2x2_ASAP7_75t_L g1518 ( .A(n_426), .B(n_605), .Y(n_1518) );
INVx2_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
AOI22xp5_ASAP7_75t_L g1876 ( .A1(n_427), .A2(n_586), .B1(n_1877), .B2(n_1878), .Y(n_1876) );
INVx1_ASAP7_75t_L g1901 ( .A(n_427), .Y(n_1901) );
BUFx3_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
AND2x6_ASAP7_75t_L g1424 ( .A(n_428), .B(n_1407), .Y(n_1424) );
AOI33xp33_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_437), .A3(n_444), .B1(n_451), .B2(n_455), .B3(n_461), .Y(n_429) );
CKINVDCx5p33_ASAP7_75t_R g430 ( .A(n_431), .Y(n_430) );
CKINVDCx5p33_ASAP7_75t_R g1456 ( .A(n_431), .Y(n_1456) );
OR2x6_ASAP7_75t_L g431 ( .A(n_432), .B(n_435), .Y(n_431) );
INVx1_ASAP7_75t_L g751 ( .A(n_432), .Y(n_751) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
BUFx3_ASAP7_75t_L g596 ( .A(n_433), .Y(n_596) );
INVx2_ASAP7_75t_SL g861 ( .A(n_433), .Y(n_861) );
INVx1_ASAP7_75t_L g1279 ( .A(n_433), .Y(n_1279) );
INVx1_ASAP7_75t_L g1395 ( .A(n_434), .Y(n_1395) );
INVx2_ASAP7_75t_L g474 ( .A(n_435), .Y(n_474) );
AOI31xp33_ASAP7_75t_L g724 ( .A1(n_435), .A2(n_725), .A3(n_743), .B(n_757), .Y(n_724) );
AND2x4_ASAP7_75t_L g817 ( .A(n_435), .B(n_539), .Y(n_817) );
BUFx2_ASAP7_75t_L g969 ( .A(n_435), .Y(n_969) );
AND2x4_ASAP7_75t_L g1011 ( .A(n_435), .B(n_539), .Y(n_1011) );
AND2x2_ASAP7_75t_L g1202 ( .A(n_435), .B(n_511), .Y(n_1202) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
BUFx2_ASAP7_75t_L g564 ( .A(n_436), .Y(n_564) );
OR2x6_ASAP7_75t_L g653 ( .A(n_436), .B(n_654), .Y(n_653) );
BUFx3_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_SL g1513 ( .A(n_439), .Y(n_1513) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_441), .B(n_467), .Y(n_466) );
HB1xp67_ASAP7_75t_L g1417 ( .A(n_441), .Y(n_1417) );
BUFx2_ASAP7_75t_SL g1514 ( .A(n_441), .Y(n_1514) );
BUFx6f_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
BUFx4f_ASAP7_75t_L g573 ( .A(n_442), .Y(n_573) );
AND2x4_ASAP7_75t_L g601 ( .A(n_442), .B(n_581), .Y(n_601) );
INVx2_ASAP7_75t_SL g782 ( .A(n_442), .Y(n_782) );
BUFx3_ASAP7_75t_L g788 ( .A(n_442), .Y(n_788) );
AND2x4_ASAP7_75t_L g1151 ( .A(n_442), .B(n_956), .Y(n_1151) );
INVx1_ASAP7_75t_L g1571 ( .A(n_442), .Y(n_1571) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
BUFx6f_ASAP7_75t_L g594 ( .A(n_443), .Y(n_594) );
BUFx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_447), .Y(n_454) );
INVx1_ASAP7_75t_L g754 ( .A(n_447), .Y(n_754) );
INVx2_ASAP7_75t_L g784 ( .A(n_447), .Y(n_784) );
INVx2_ASAP7_75t_L g849 ( .A(n_447), .Y(n_849) );
INVx2_ASAP7_75t_SL g1129 ( .A(n_447), .Y(n_1129) );
HB1xp67_ASAP7_75t_L g1150 ( .A(n_447), .Y(n_1150) );
INVx2_ASAP7_75t_L g1403 ( .A(n_447), .Y(n_1403) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g756 ( .A(n_450), .Y(n_756) );
BUFx6f_ASAP7_75t_L g864 ( .A(n_450), .Y(n_864) );
BUFx6f_ASAP7_75t_L g936 ( .A(n_450), .Y(n_936) );
INVx2_ASAP7_75t_L g1062 ( .A(n_450), .Y(n_1062) );
AND2x6_ASAP7_75t_L g1414 ( .A(n_450), .B(n_1401), .Y(n_1414) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx4_ASAP7_75t_L g574 ( .A(n_454), .Y(n_574) );
INVx1_ASAP7_75t_L g1899 ( .A(n_454), .Y(n_1899) );
BUFx3_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g947 ( .A(n_457), .Y(n_947) );
INVx2_ASAP7_75t_L g966 ( .A(n_457), .Y(n_966) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
BUFx6f_ASAP7_75t_L g579 ( .A(n_460), .Y(n_579) );
BUFx3_ASAP7_75t_L g1297 ( .A(n_460), .Y(n_1297) );
BUFx4f_ASAP7_75t_L g1466 ( .A(n_461), .Y(n_1466) );
AND2x4_ASAP7_75t_L g461 ( .A(n_462), .B(n_463), .Y(n_461) );
AND2x4_ASAP7_75t_L g471 ( .A(n_462), .B(n_472), .Y(n_471) );
CKINVDCx5p33_ASAP7_75t_R g575 ( .A(n_463), .Y(n_575) );
INVx1_ASAP7_75t_L g736 ( .A(n_463), .Y(n_736) );
HB1xp67_ASAP7_75t_L g951 ( .A(n_463), .Y(n_951) );
INVx2_ASAP7_75t_L g1051 ( .A(n_463), .Y(n_1051) );
INVx2_ASAP7_75t_SL g1226 ( .A(n_463), .Y(n_1226) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
OR2x6_ASAP7_75t_L g470 ( .A(n_471), .B(n_473), .Y(n_470) );
INVx2_ASAP7_75t_L g620 ( .A(n_471), .Y(n_620) );
INVx2_ASAP7_75t_L g793 ( .A(n_472), .Y(n_793) );
NOR2xp67_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
INVx2_ASAP7_75t_L g795 ( .A(n_474), .Y(n_795) );
AOI211xp5_ASAP7_75t_L g1891 ( .A1(n_474), .A2(n_1892), .B(n_1912), .C(n_1919), .Y(n_1891) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_480), .Y(n_475) );
AND2x2_ASAP7_75t_L g517 ( .A(n_476), .B(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
OR2x6_ASAP7_75t_L g521 ( .A(n_477), .B(n_522), .Y(n_521) );
OR2x2_ASAP7_75t_L g551 ( .A(n_477), .B(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
AND2x2_ASAP7_75t_L g1173 ( .A(n_480), .B(n_629), .Y(n_1173) );
INVx2_ASAP7_75t_SL g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_SL g636 ( .A(n_481), .Y(n_636) );
INVx2_ASAP7_75t_L g1009 ( .A(n_481), .Y(n_1009) );
INVx3_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
BUFx6f_ASAP7_75t_L g509 ( .A(n_482), .Y(n_509) );
OAI31xp33_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_523), .A3(n_554), .B(n_562), .Y(n_483) );
INVx8_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AND2x4_ASAP7_75t_L g486 ( .A(n_487), .B(n_491), .Y(n_486) );
AND2x4_ASAP7_75t_L g561 ( .A(n_487), .B(n_548), .Y(n_561) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AND2x4_ASAP7_75t_L g525 ( .A(n_489), .B(n_509), .Y(n_525) );
AND2x2_ASAP7_75t_L g556 ( .A(n_489), .B(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g513 ( .A(n_490), .Y(n_513) );
INVx1_ASAP7_75t_L g655 ( .A(n_490), .Y(n_655) );
BUFx6f_ASAP7_75t_L g933 ( .A(n_491), .Y(n_933) );
BUFx3_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_492), .Y(n_506) );
BUFx3_ASAP7_75t_L g632 ( .A(n_492), .Y(n_632) );
BUFx6f_ASAP7_75t_L g806 ( .A(n_492), .Y(n_806) );
BUFx2_ASAP7_75t_L g832 ( .A(n_492), .Y(n_832) );
INVx1_ASAP7_75t_L g1196 ( .A(n_492), .Y(n_1196) );
AND2x4_ASAP7_75t_L g1433 ( .A(n_492), .B(n_1434), .Y(n_1433) );
AND2x4_ASAP7_75t_L g492 ( .A(n_493), .B(n_494), .Y(n_492) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx2_ASAP7_75t_L g708 ( .A(n_497), .Y(n_708) );
INVx2_ASAP7_75t_SL g712 ( .A(n_497), .Y(n_712) );
INVx2_ASAP7_75t_L g1260 ( .A(n_497), .Y(n_1260) );
BUFx3_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g666 ( .A(n_498), .Y(n_666) );
INVx1_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g543 ( .A(n_499), .Y(n_543) );
BUFx2_ASAP7_75t_L g921 ( .A(n_499), .Y(n_921) );
INVx1_ASAP7_75t_L g522 ( .A(n_500), .Y(n_522) );
AND2x4_ASAP7_75t_L g557 ( .A(n_500), .B(n_558), .Y(n_557) );
OAI22xp33_ASAP7_75t_L g697 ( .A1(n_501), .A2(n_698), .B1(n_699), .B2(n_700), .Y(n_697) );
INVxp67_ASAP7_75t_L g821 ( .A(n_501), .Y(n_821) );
INVx2_ASAP7_75t_SL g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_SL g668 ( .A(n_502), .Y(n_668) );
INVx2_ASAP7_75t_SL g799 ( .A(n_502), .Y(n_799) );
BUFx3_ASAP7_75t_L g890 ( .A(n_502), .Y(n_890) );
INVx4_ASAP7_75t_L g1007 ( .A(n_502), .Y(n_1007) );
BUFx6f_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g549 ( .A(n_503), .Y(n_549) );
INVx3_ASAP7_75t_L g628 ( .A(n_503), .Y(n_628) );
INVx1_ASAP7_75t_L g1446 ( .A(n_503), .Y(n_1446) );
BUFx6f_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AND2x2_ASAP7_75t_L g1243 ( .A(n_506), .B(n_629), .Y(n_1243) );
INVx2_ASAP7_75t_SL g507 ( .A(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g928 ( .A(n_508), .Y(n_928) );
INVx2_ASAP7_75t_L g1194 ( .A(n_508), .Y(n_1194) );
INVx3_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
BUFx6f_ASAP7_75t_L g802 ( .A(n_509), .Y(n_802) );
BUFx2_ASAP7_75t_L g1470 ( .A(n_509), .Y(n_1470) );
INVx2_ASAP7_75t_SL g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
NAND2x1p5_ASAP7_75t_L g512 ( .A(n_513), .B(n_514), .Y(n_512) );
INVx1_ASAP7_75t_L g1435 ( .A(n_513), .Y(n_1435) );
HB1xp67_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AND2x4_ASAP7_75t_L g827 ( .A(n_518), .B(n_646), .Y(n_827) );
HB1xp67_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
INVx1_ASAP7_75t_L g645 ( .A(n_519), .Y(n_645) );
CKINVDCx11_ASAP7_75t_R g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g649 ( .A(n_522), .Y(n_649) );
CKINVDCx6p67_ASAP7_75t_R g524 ( .A(n_525), .Y(n_524) );
OAI221xp5_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_533), .B1(n_534), .B2(n_536), .C(n_537), .Y(n_526) );
BUFx3_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
OAI22xp5_ASAP7_75t_L g1495 ( .A1(n_528), .A2(n_1496), .B1(n_1497), .B2(n_1498), .Y(n_1495) );
BUFx3_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g701 ( .A(n_529), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g1177 ( .A1(n_529), .A2(n_1015), .B1(n_1178), .B2(n_1179), .Y(n_1177) );
BUFx6f_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_532), .Y(n_530) );
AND2x2_ASAP7_75t_L g553 ( .A(n_531), .B(n_532), .Y(n_553) );
INVx1_ASAP7_75t_L g830 ( .A(n_532), .Y(n_830) );
OAI22xp5_ASAP7_75t_SL g1265 ( .A1(n_534), .A2(n_700), .B1(n_1266), .B2(n_1267), .Y(n_1265) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_544), .B1(n_545), .B2(n_550), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g887 ( .A(n_543), .Y(n_887) );
INVx1_ASAP7_75t_L g1255 ( .A(n_543), .Y(n_1255) );
INVx1_ASAP7_75t_L g1845 ( .A(n_543), .Y(n_1845) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g1264 ( .A(n_549), .Y(n_1264) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_552), .Y(n_717) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
INVx2_ASAP7_75t_L g661 ( .A(n_553), .Y(n_661) );
BUFx2_ASAP7_75t_L g674 ( .A(n_553), .Y(n_674) );
INVx3_ASAP7_75t_L g815 ( .A(n_553), .Y(n_815) );
INVx3_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
BUFx6f_ASAP7_75t_L g639 ( .A(n_557), .Y(n_639) );
INVx1_ASAP7_75t_L g809 ( .A(n_557), .Y(n_809) );
INVx1_ASAP7_75t_L g820 ( .A(n_557), .Y(n_820) );
BUFx2_ASAP7_75t_L g1005 ( .A(n_557), .Y(n_1005) );
BUFx6f_ASAP7_75t_L g1198 ( .A(n_557), .Y(n_1198) );
BUFx6f_ASAP7_75t_L g1200 ( .A(n_557), .Y(n_1200) );
AND2x4_ASAP7_75t_L g1441 ( .A(n_557), .B(n_1442), .Y(n_1441) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx3_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx5_ASAP7_75t_L g999 ( .A(n_562), .Y(n_999) );
BUFx8_ASAP7_75t_SL g562 ( .A(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g569 ( .A(n_563), .Y(n_569) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
BUFx2_ASAP7_75t_L g869 ( .A(n_564), .Y(n_869) );
AND2x4_ASAP7_75t_L g1394 ( .A(n_564), .B(n_1395), .Y(n_1394) );
AO22x2_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_679), .B1(n_758), .B2(n_759), .Y(n_565) );
INVx1_ASAP7_75t_L g759 ( .A(n_566), .Y(n_759) );
XOR2x2_ASAP7_75t_L g566 ( .A(n_567), .B(n_678), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_621), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_570), .B1(n_615), .B2(n_616), .Y(n_568) );
AOI22xp5_ASAP7_75t_L g1286 ( .A1(n_569), .A2(n_1287), .B1(n_1305), .B2(n_1306), .Y(n_1286) );
OAI31xp33_ASAP7_75t_SL g1859 ( .A1(n_569), .A2(n_1860), .A3(n_1861), .B(n_1862), .Y(n_1859) );
NAND3xp33_ASAP7_75t_L g570 ( .A(n_571), .B(n_589), .C(n_606), .Y(n_570) );
AOI221xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_576), .B1(n_580), .B2(n_582), .C(n_583), .Y(n_571) );
BUFx2_ASAP7_75t_L g749 ( .A(n_573), .Y(n_749) );
A2O1A1Ixp33_ASAP7_75t_L g1229 ( .A1(n_573), .A2(n_581), .B(n_1230), .C(n_1231), .Y(n_1229) );
AOI22xp33_ASAP7_75t_L g1508 ( .A1(n_574), .A2(n_1501), .B1(n_1503), .B2(n_1509), .Y(n_1508) );
INVxp67_ASAP7_75t_L g1529 ( .A(n_577), .Y(n_1529) );
BUFx3_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x4_ASAP7_75t_L g580 ( .A(n_578), .B(n_581), .Y(n_580) );
INVx2_ASAP7_75t_SL g748 ( .A(n_578), .Y(n_748) );
INVx1_ASAP7_75t_L g1369 ( .A(n_578), .Y(n_1369) );
INVx1_ASAP7_75t_L g1523 ( .A(n_579), .Y(n_1523) );
INVx1_ASAP7_75t_L g727 ( .A(n_580), .Y(n_727) );
AOI21xp5_ASAP7_75t_L g838 ( .A1(n_580), .A2(n_839), .B(n_840), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g988 ( .A1(n_580), .A2(n_608), .B1(n_989), .B2(n_990), .Y(n_988) );
AOI22xp33_ASAP7_75t_L g1063 ( .A1(n_580), .A2(n_608), .B1(n_1064), .B2(n_1065), .Y(n_1063) );
AOI211xp5_ASAP7_75t_L g1364 ( .A1(n_580), .A2(n_1357), .B(n_1365), .C(n_1367), .Y(n_1364) );
AOI22xp33_ASAP7_75t_L g1581 ( .A1(n_580), .A2(n_608), .B1(n_1561), .B2(n_1564), .Y(n_1581) );
AOI222xp33_ASAP7_75t_L g768 ( .A1(n_581), .A2(n_585), .B1(n_588), .B2(n_769), .C1(n_777), .C2(n_778), .Y(n_768) );
OAI21xp5_ASAP7_75t_L g960 ( .A1(n_581), .A2(n_961), .B(n_965), .Y(n_960) );
AND2x2_ASAP7_75t_L g1123 ( .A(n_581), .B(n_775), .Y(n_1123) );
AOI221xp5_ASAP7_75t_L g1152 ( .A1(n_581), .A2(n_608), .B1(n_1153), .B2(n_1154), .C(n_1159), .Y(n_1152) );
OAI21xp5_ASAP7_75t_L g1893 ( .A1(n_581), .A2(n_1894), .B(n_1896), .Y(n_1893) );
OAI22xp5_ASAP7_75t_L g669 ( .A1(n_582), .A2(n_611), .B1(n_664), .B2(n_670), .Y(n_669) );
INVx2_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g957 ( .A1(n_585), .A2(n_588), .B1(n_958), .B2(n_959), .Y(n_957) );
AOI222xp33_ASAP7_75t_L g993 ( .A1(n_585), .A2(n_792), .B1(n_994), .B2(n_995), .C1(n_996), .C2(n_997), .Y(n_993) );
INVx1_ASAP7_75t_L g1366 ( .A(n_585), .Y(n_1366) );
INVx2_ASAP7_75t_SL g1517 ( .A(n_585), .Y(n_1517) );
INVxp67_ASAP7_75t_L g742 ( .A(n_586), .Y(n_742) );
INVx3_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AOI221xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_597), .B1(n_601), .B2(n_602), .C(n_603), .Y(n_589) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g1057 ( .A(n_592), .Y(n_1057) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
AND2x4_ASAP7_75t_L g603 ( .A(n_593), .B(n_604), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g773 ( .A1(n_593), .A2(n_774), .B1(n_775), .B2(n_776), .Y(n_773) );
BUFx6f_ASAP7_75t_L g954 ( .A(n_593), .Y(n_954) );
BUFx6f_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g858 ( .A(n_594), .Y(n_858) );
BUFx6f_ASAP7_75t_L g1278 ( .A(n_594), .Y(n_1278) );
INVx2_ASAP7_75t_L g1379 ( .A(n_594), .Y(n_1379) );
AND2x4_ASAP7_75t_L g1426 ( .A(n_594), .B(n_1427), .Y(n_1426) );
INVx3_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g984 ( .A(n_596), .Y(n_984) );
OAI221xp5_ASAP7_75t_L g1524 ( .A1(n_596), .A2(n_739), .B1(n_1493), .B2(n_1498), .C(n_1525), .Y(n_1524) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g791 ( .A(n_600), .Y(n_791) );
INVx1_ASAP7_75t_L g1463 ( .A(n_600), .Y(n_1463) );
INVx1_ASAP7_75t_L g745 ( .A(n_601), .Y(n_745) );
BUFx6f_ASAP7_75t_L g851 ( .A(n_601), .Y(n_851) );
INVx1_ASAP7_75t_L g992 ( .A(n_601), .Y(n_992) );
INVx2_ASAP7_75t_SL g1054 ( .A(n_601), .Y(n_1054) );
AOI221xp5_ASAP7_75t_L g1276 ( .A1(n_601), .A2(n_1151), .B1(n_1267), .B2(n_1277), .C(n_1280), .Y(n_1276) );
INVx1_ASAP7_75t_L g1576 ( .A(n_601), .Y(n_1576) );
OAI22xp33_ASAP7_75t_L g672 ( .A1(n_602), .A2(n_607), .B1(n_658), .B2(n_673), .Y(n_672) );
AOI221xp5_ASAP7_75t_L g743 ( .A1(n_603), .A2(n_718), .B1(n_744), .B2(n_746), .C(n_752), .Y(n_743) );
AOI21xp33_ASAP7_75t_L g779 ( .A1(n_603), .A2(n_780), .B(n_785), .Y(n_779) );
AOI221xp5_ASAP7_75t_L g850 ( .A1(n_603), .A2(n_851), .B1(n_852), .B2(n_853), .C(n_862), .Y(n_850) );
INVx1_ASAP7_75t_L g998 ( .A(n_603), .Y(n_998) );
AOI221xp5_ASAP7_75t_L g1052 ( .A1(n_603), .A2(n_1053), .B1(n_1055), .B2(n_1056), .C(n_1058), .Y(n_1052) );
AOI221xp5_ASAP7_75t_L g1124 ( .A1(n_603), .A2(n_1053), .B1(n_1117), .B2(n_1125), .C(n_1126), .Y(n_1124) );
AOI221xp5_ASAP7_75t_L g1373 ( .A1(n_603), .A2(n_744), .B1(n_1360), .B2(n_1374), .C(n_1380), .Y(n_1373) );
INVx1_ASAP7_75t_L g1515 ( .A(n_603), .Y(n_1515) );
AOI221xp5_ASAP7_75t_L g1574 ( .A1(n_603), .A2(n_1565), .B1(n_1575), .B2(n_1577), .C(n_1579), .Y(n_1574) );
INVx1_ASAP7_75t_SL g604 ( .A(n_605), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_608), .B1(n_611), .B2(n_612), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_608), .A2(n_612), .B1(n_714), .B2(n_716), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_608), .A2(n_612), .B1(n_866), .B2(n_867), .Y(n_865) );
AOI22xp5_ASAP7_75t_L g1120 ( .A1(n_608), .A2(n_1113), .B1(n_1116), .B2(n_1121), .Y(n_1120) );
AOI22xp5_ASAP7_75t_L g1281 ( .A1(n_608), .A2(n_612), .B1(n_1261), .B2(n_1266), .Y(n_1281) );
AOI22xp33_ASAP7_75t_L g1288 ( .A1(n_608), .A2(n_1123), .B1(n_1289), .B2(n_1290), .Y(n_1288) );
AOI22xp33_ASAP7_75t_L g1381 ( .A1(n_608), .A2(n_612), .B1(n_1356), .B2(n_1359), .Y(n_1381) );
INVx6_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g771 ( .A(n_610), .Y(n_771) );
INVx1_ASAP7_75t_L g950 ( .A(n_610), .Y(n_950) );
AOI211xp5_ASAP7_75t_L g1042 ( .A1(n_612), .A2(n_1043), .B(n_1044), .C(n_1046), .Y(n_1042) );
AOI221xp5_ASAP7_75t_L g1130 ( .A1(n_612), .A2(n_1114), .B1(n_1131), .B2(n_1132), .C(n_1133), .Y(n_1130) );
AOI221xp5_ASAP7_75t_L g1291 ( .A1(n_612), .A2(n_1292), .B1(n_1293), .B2(n_1296), .C(n_1298), .Y(n_1291) );
AOI221xp5_ASAP7_75t_L g1568 ( .A1(n_612), .A2(n_1562), .B1(n_1569), .B2(n_1572), .C(n_1573), .Y(n_1568) );
INVx4_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx2_ASAP7_75t_L g733 ( .A(n_614), .Y(n_733) );
INVx1_ASAP7_75t_L g964 ( .A(n_614), .Y(n_964) );
AOI21xp33_ASAP7_75t_SL g835 ( .A1(n_616), .A2(n_836), .B(n_837), .Y(n_835) );
AOI22xp5_ASAP7_75t_L g1040 ( .A1(n_616), .A2(n_869), .B1(n_1041), .B2(n_1066), .Y(n_1040) );
INVx5_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g722 ( .A(n_617), .Y(n_722) );
INVx1_ASAP7_75t_L g1137 ( .A(n_617), .Y(n_1137) );
INVx2_ASAP7_75t_SL g1282 ( .A(n_617), .Y(n_1282) );
INVx2_ASAP7_75t_L g1306 ( .A(n_617), .Y(n_1306) );
AND2x4_ASAP7_75t_L g617 ( .A(n_618), .B(n_620), .Y(n_617) );
INVx2_ASAP7_75t_L g825 ( .A(n_618), .Y(n_825) );
INVx3_ASAP7_75t_L g646 ( .A(n_619), .Y(n_646) );
NOR3xp33_ASAP7_75t_L g621 ( .A(n_622), .B(n_640), .C(n_652), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_623), .B(n_633), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_625), .B1(n_630), .B2(n_631), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g1021 ( .A1(n_625), .A2(n_720), .B1(n_1022), .B2(n_1029), .Y(n_1021) );
AOI22xp33_ASAP7_75t_L g1080 ( .A1(n_625), .A2(n_631), .B1(n_1049), .B2(n_1081), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g1092 ( .A1(n_625), .A2(n_631), .B1(n_1093), .B2(n_1094), .Y(n_1092) );
BUFx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
BUFx2_ASAP7_75t_L g686 ( .A(n_626), .Y(n_686) );
BUFx2_ASAP7_75t_L g874 ( .A(n_626), .Y(n_874) );
BUFx2_ASAP7_75t_L g910 ( .A(n_626), .Y(n_910) );
BUFx2_ASAP7_75t_L g1170 ( .A(n_626), .Y(n_1170) );
BUFx2_ASAP7_75t_L g1311 ( .A(n_626), .Y(n_1311) );
AND2x4_ASAP7_75t_L g626 ( .A(n_627), .B(n_629), .Y(n_626) );
BUFx3_ASAP7_75t_L g671 ( .A(n_627), .Y(n_671) );
INVx1_ASAP7_75t_SL g1847 ( .A(n_627), .Y(n_1847) );
INVx3_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx3_ASAP7_75t_L g812 ( .A(n_628), .Y(n_812) );
BUFx6f_ASAP7_75t_L g925 ( .A(n_628), .Y(n_925) );
AND2x6_ASAP7_75t_L g631 ( .A(n_629), .B(n_632), .Y(n_631) );
AND2x4_ASAP7_75t_L g635 ( .A(n_629), .B(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g638 ( .A(n_629), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g691 ( .A(n_629), .B(n_639), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_629), .A2(n_720), .B1(n_798), .B2(n_807), .Y(n_797) );
AND2x2_ASAP7_75t_L g1085 ( .A(n_629), .B(n_639), .Y(n_1085) );
AND2x2_ASAP7_75t_L g1207 ( .A(n_629), .B(n_639), .Y(n_1207) );
AND2x2_ASAP7_75t_L g1211 ( .A(n_629), .B(n_812), .Y(n_1211) );
AND2x2_ASAP7_75t_L g1316 ( .A(n_629), .B(n_639), .Y(n_1316) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_631), .A2(n_685), .B1(n_686), .B2(n_687), .Y(n_684) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_631), .A2(n_844), .B1(n_873), .B2(n_874), .Y(n_872) );
AOI22xp33_ASAP7_75t_L g908 ( .A1(n_631), .A2(n_909), .B1(n_910), .B2(n_911), .Y(n_908) );
INVx1_ASAP7_75t_SL g1002 ( .A(n_631), .Y(n_1002) );
AOI22xp5_ASAP7_75t_L g1165 ( .A1(n_631), .A2(n_1085), .B1(n_1166), .B2(n_1167), .Y(n_1165) );
AOI22xp33_ASAP7_75t_L g1206 ( .A1(n_631), .A2(n_1207), .B1(n_1208), .B2(n_1209), .Y(n_1206) );
AOI22xp33_ASAP7_75t_L g1309 ( .A1(n_631), .A2(n_1310), .B1(n_1311), .B2(n_1312), .Y(n_1309) );
AOI22xp33_ASAP7_75t_L g1337 ( .A1(n_631), .A2(n_1170), .B1(n_1338), .B2(n_1339), .Y(n_1337) );
AOI22xp33_ASAP7_75t_L g1546 ( .A1(n_631), .A2(n_874), .B1(n_1547), .B2(n_1548), .Y(n_1546) );
NAND2x1p5_ASAP7_75t_L g651 ( .A(n_632), .B(n_646), .Y(n_651) );
BUFx2_ASAP7_75t_L g1010 ( .A(n_632), .Y(n_1010) );
AOI22xp33_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_635), .B1(n_637), .B2(n_638), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_635), .A2(n_689), .B1(n_690), .B2(n_691), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_635), .A2(n_638), .B1(n_876), .B2(n_877), .Y(n_875) );
AOI21xp5_ASAP7_75t_L g915 ( .A1(n_635), .A2(n_916), .B(n_917), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g1018 ( .A1(n_635), .A2(n_638), .B1(n_1019), .B2(n_1020), .Y(n_1018) );
AOI22xp33_ASAP7_75t_L g1082 ( .A1(n_635), .A2(n_1083), .B1(n_1084), .B2(n_1085), .Y(n_1082) );
AOI22xp33_ASAP7_75t_L g1095 ( .A1(n_635), .A2(n_1085), .B1(n_1096), .B2(n_1097), .Y(n_1095) );
NAND2xp5_ASAP7_75t_L g1203 ( .A(n_635), .B(n_1204), .Y(n_1203) );
AOI22xp33_ASAP7_75t_L g1313 ( .A1(n_635), .A2(n_1314), .B1(n_1315), .B2(n_1316), .Y(n_1313) );
AOI22xp33_ASAP7_75t_L g1340 ( .A1(n_635), .A2(n_691), .B1(n_1341), .B2(n_1342), .Y(n_1340) );
AOI22xp33_ASAP7_75t_L g1549 ( .A1(n_635), .A2(n_1316), .B1(n_1550), .B2(n_1551), .Y(n_1549) );
INVx2_ASAP7_75t_SL g1024 ( .A(n_639), .Y(n_1024) );
INVx2_ASAP7_75t_SL g641 ( .A(n_642), .Y(n_641) );
INVx2_ASAP7_75t_L g693 ( .A(n_642), .Y(n_693) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
HB1xp67_ASAP7_75t_L g1318 ( .A(n_643), .Y(n_1318) );
NAND2x1_ASAP7_75t_SL g643 ( .A(n_644), .B(n_646), .Y(n_643) );
AOI22xp33_ASAP7_75t_L g1016 ( .A1(n_644), .A2(n_649), .B1(n_995), .B2(n_996), .Y(n_1016) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
NAND2x1p5_ASAP7_75t_L g648 ( .A(n_646), .B(n_649), .Y(n_648) );
AND2x4_ASAP7_75t_L g828 ( .A(n_646), .B(n_829), .Y(n_828) );
AND2x4_ASAP7_75t_L g831 ( .A(n_646), .B(n_832), .Y(n_831) );
AOI32xp33_ASAP7_75t_L g1003 ( .A1(n_646), .A2(n_1004), .A3(n_1008), .B1(n_1011), .B2(n_1012), .Y(n_1003) );
BUFx4f_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
BUFx4f_ASAP7_75t_L g694 ( .A(n_648), .Y(n_694) );
BUFx3_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
BUFx2_ASAP7_75t_L g879 ( .A(n_651), .Y(n_879) );
BUFx2_ASAP7_75t_L g1099 ( .A(n_651), .Y(n_1099) );
OAI33xp33_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_656), .A3(n_662), .B1(n_669), .B2(n_672), .B3(n_675), .Y(n_652) );
HB1xp67_ASAP7_75t_L g696 ( .A(n_653), .Y(n_696) );
OAI33xp33_ASAP7_75t_L g880 ( .A1(n_653), .A2(n_675), .A3(n_881), .B1(n_886), .B2(n_892), .B3(n_895), .Y(n_880) );
OAI22xp5_ASAP7_75t_L g917 ( .A1(n_653), .A2(n_675), .B1(n_918), .B2(n_929), .Y(n_917) );
HB1xp67_ASAP7_75t_L g1101 ( .A(n_653), .Y(n_1101) );
OAI33xp33_ASAP7_75t_L g1248 ( .A1(n_653), .A2(n_719), .A3(n_1249), .B1(n_1252), .B2(n_1258), .B3(n_1265), .Y(n_1248) );
OAI33xp33_ASAP7_75t_L g1319 ( .A1(n_653), .A2(n_675), .A3(n_1320), .B1(n_1324), .B2(n_1329), .B3(n_1330), .Y(n_1319) );
OAI33xp33_ASAP7_75t_L g1344 ( .A1(n_653), .A2(n_675), .A3(n_1345), .B1(n_1350), .B2(n_1355), .B3(n_1358), .Y(n_1344) );
INVx1_ASAP7_75t_L g1442 ( .A(n_655), .Y(n_1442) );
OAI22xp33_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_658), .B1(n_660), .B2(n_661), .Y(n_656) );
BUFx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
OAI22xp33_ASAP7_75t_L g715 ( .A1(n_659), .A2(n_716), .B1(n_717), .B2(n_718), .Y(n_715) );
OAI22xp33_ASAP7_75t_L g813 ( .A1(n_659), .A2(n_776), .B1(n_814), .B2(n_815), .Y(n_813) );
OAI22xp5_ASAP7_75t_L g822 ( .A1(n_659), .A2(n_815), .B1(n_823), .B2(n_824), .Y(n_822) );
INVx1_ASAP7_75t_L g897 ( .A(n_659), .Y(n_897) );
INVx1_ASAP7_75t_L g1104 ( .A(n_659), .Y(n_1104) );
OAI22xp33_ASAP7_75t_L g1355 ( .A1(n_659), .A2(n_1112), .B1(n_1356), .B2(n_1357), .Y(n_1355) );
OAI22xp5_ASAP7_75t_SL g1502 ( .A1(n_659), .A2(n_700), .B1(n_1503), .B2(n_1504), .Y(n_1502) );
OAI22xp33_ASAP7_75t_L g1249 ( .A1(n_661), .A2(n_1013), .B1(n_1250), .B2(n_1251), .Y(n_1249) );
OAI22xp5_ASAP7_75t_SL g662 ( .A1(n_663), .A2(n_664), .B1(n_667), .B2(n_668), .Y(n_662) );
INVx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx2_ASAP7_75t_L g1326 ( .A(n_665), .Y(n_1326) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
BUFx2_ASAP7_75t_L g1112 ( .A(n_666), .Y(n_1112) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_668), .A2(n_711), .B1(n_713), .B2(n_714), .Y(n_710) );
OAI221xp5_ASAP7_75t_L g929 ( .A1(n_668), .A2(n_712), .B1(n_930), .B2(n_931), .C(n_932), .Y(n_929) );
OAI22xp33_ASAP7_75t_L g1358 ( .A1(n_670), .A2(n_1347), .B1(n_1359), .B2(n_1360), .Y(n_1358) );
CKINVDCx5p33_ASAP7_75t_R g670 ( .A(n_671), .Y(n_670) );
OAI22xp33_ASAP7_75t_L g881 ( .A1(n_673), .A2(n_882), .B1(n_884), .B2(n_885), .Y(n_881) );
OAI22xp33_ASAP7_75t_L g1320 ( .A1(n_673), .A2(n_1321), .B1(n_1322), .B2(n_1323), .Y(n_1320) );
INVx2_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
OAI33xp33_ASAP7_75t_L g1100 ( .A1(n_675), .A2(n_1101), .A3(n_1102), .B1(n_1107), .B2(n_1111), .B3(n_1115), .Y(n_1100) );
OAI33xp33_ASAP7_75t_L g1553 ( .A1(n_675), .A2(n_1101), .A3(n_1554), .B1(n_1557), .B2(n_1560), .B3(n_1563), .Y(n_1553) );
CKINVDCx8_ASAP7_75t_R g675 ( .A(n_676), .Y(n_675) );
INVx5_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx6_ASAP7_75t_L g720 ( .A(n_677), .Y(n_720) );
INVx1_ASAP7_75t_L g758 ( .A(n_679), .Y(n_758) );
XNOR2xp5_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_682), .B(n_721), .Y(n_681) );
NOR3xp33_ASAP7_75t_SL g682 ( .A(n_683), .B(n_692), .C(n_695), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_684), .B(n_688), .Y(n_683) );
AOI22xp33_ASAP7_75t_SL g912 ( .A1(n_691), .A2(n_825), .B1(n_913), .B2(n_914), .Y(n_912) );
OAI33xp33_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_697), .A3(n_702), .B1(n_710), .B2(n_715), .B3(n_719), .Y(n_695) );
OAI22xp33_ASAP7_75t_L g1115 ( .A1(n_700), .A2(n_1103), .B1(n_1116), .B2(n_1117), .Y(n_1115) );
OAI22xp33_ASAP7_75t_L g1330 ( .A1(n_700), .A2(n_1289), .B1(n_1304), .B2(n_1321), .Y(n_1330) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx2_ASAP7_75t_L g1028 ( .A(n_701), .Y(n_1028) );
OAI22xp33_ASAP7_75t_SL g702 ( .A1(n_703), .A2(n_705), .B1(n_706), .B2(n_709), .Y(n_702) );
OAI22xp33_ASAP7_75t_L g1345 ( .A1(n_703), .A2(n_1346), .B1(n_1347), .B2(n_1349), .Y(n_1345) );
INVx3_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g892 ( .A1(n_708), .A2(n_839), .B1(n_867), .B2(n_893), .Y(n_892) );
OAI22xp5_ASAP7_75t_L g1492 ( .A1(n_708), .A2(n_1007), .B1(n_1493), .B2(n_1494), .Y(n_1492) );
OAI22xp5_ASAP7_75t_L g1560 ( .A1(n_708), .A2(n_893), .B1(n_1561), .B2(n_1562), .Y(n_1560) );
BUFx2_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
AOI21xp5_ASAP7_75t_L g725 ( .A1(n_713), .A2(n_726), .B(n_728), .Y(n_725) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
AOI33xp33_ASAP7_75t_L g1071 ( .A1(n_720), .A2(n_817), .A3(n_1072), .B1(n_1074), .B2(n_1075), .B3(n_1078), .Y(n_1071) );
AOI222xp33_ASAP7_75t_L g1172 ( .A1(n_720), .A2(n_817), .B1(n_1173), .B2(n_1174), .C1(n_1175), .C2(n_1180), .Y(n_1172) );
AOI33xp33_ASAP7_75t_L g1467 ( .A1(n_720), .A2(n_1468), .A3(n_1469), .B1(n_1471), .B2(n_1477), .B3(n_1479), .Y(n_1467) );
AOI322xp5_ASAP7_75t_L g1920 ( .A1(n_720), .A2(n_817), .A3(n_1243), .B1(n_1907), .B2(n_1921), .C1(n_1922), .C2(n_1923), .Y(n_1920) );
AOI21xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_723), .B(n_724), .Y(n_721) );
AOI21xp5_ASAP7_75t_L g1361 ( .A1(n_722), .A2(n_1362), .B(n_1363), .Y(n_1361) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
AOI31xp33_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_734), .A3(n_737), .B(n_741), .Y(n_729) );
INVx1_ASAP7_75t_L g1157 ( .A(n_731), .Y(n_1157) );
INVx1_ASAP7_75t_L g772 ( .A(n_732), .Y(n_772) );
BUFx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx2_ASAP7_75t_L g1232 ( .A(n_733), .Y(n_1232) );
A2O1A1Ixp33_ASAP7_75t_L g953 ( .A1(n_735), .A2(n_914), .B(n_954), .C(n_955), .Y(n_953) );
INVx1_ASAP7_75t_L g1535 ( .A(n_736), .Y(n_1535) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
OAI221xp5_ASAP7_75t_L g1531 ( .A1(n_739), .A2(n_1532), .B1(n_1533), .B2(n_1534), .C(n_1535), .Y(n_1531) );
BUFx2_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
HB1xp67_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g938 ( .A(n_754), .Y(n_938) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
OAI22xp5_ASAP7_75t_L g760 ( .A1(n_761), .A2(n_901), .B1(n_902), .B2(n_1032), .Y(n_760) );
INVx1_ASAP7_75t_L g1032 ( .A(n_761), .Y(n_1032) );
OAI22xp5_ASAP7_75t_L g761 ( .A1(n_762), .A2(n_763), .B1(n_833), .B2(n_900), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
XNOR2x1_ASAP7_75t_L g764 ( .A(n_765), .B(n_766), .Y(n_764) );
OR2x2_ASAP7_75t_L g766 ( .A(n_767), .B(n_796), .Y(n_766) );
AOI31xp33_ASAP7_75t_SL g767 ( .A1(n_768), .A2(n_779), .A3(n_786), .B(n_795), .Y(n_767) );
INVx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx2_ASAP7_75t_L g962 ( .A(n_771), .Y(n_962) );
HB1xp67_ASAP7_75t_L g1522 ( .A(n_771), .Y(n_1522) );
INVx2_ASAP7_75t_L g1533 ( .A(n_771), .Y(n_1533) );
INVx1_ASAP7_75t_L g855 ( .A(n_775), .Y(n_855) );
BUFx2_ASAP7_75t_L g1462 ( .A(n_775), .Y(n_1462) );
INVx1_ASAP7_75t_L g1895 ( .A(n_775), .Y(n_1895) );
AOI221xp5_ASAP7_75t_L g826 ( .A1(n_777), .A2(n_778), .B1(n_827), .B2(n_828), .C(n_831), .Y(n_826) );
INVx2_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g987 ( .A(n_782), .Y(n_987) );
INVx1_ASAP7_75t_L g1295 ( .A(n_782), .Y(n_1295) );
BUFx6f_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g1060 ( .A(n_784), .Y(n_1060) );
AOI22xp5_ASAP7_75t_L g786 ( .A1(n_787), .A2(n_790), .B1(n_792), .B2(n_794), .Y(n_786) );
INVx2_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
AOI22xp5_ASAP7_75t_L g816 ( .A1(n_794), .A2(n_817), .B1(n_818), .B2(n_825), .Y(n_816) );
NAND3xp33_ASAP7_75t_L g796 ( .A(n_797), .B(n_816), .C(n_826), .Y(n_796) );
OAI22xp5_ASAP7_75t_L g1557 ( .A1(n_799), .A2(n_1108), .B1(n_1558), .B2(n_1559), .Y(n_1557) );
AOI22xp5_ASAP7_75t_L g800 ( .A1(n_801), .A2(n_802), .B1(n_803), .B2(n_804), .Y(n_800) );
INVx2_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
INVx2_ASAP7_75t_L g1073 ( .A(n_805), .Y(n_1073) );
INVx2_ASAP7_75t_SL g805 ( .A(n_806), .Y(n_805) );
INVx2_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx1_ASAP7_75t_L g1353 ( .A(n_811), .Y(n_1353) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx2_ASAP7_75t_L g894 ( .A(n_812), .Y(n_894) );
INVx2_ASAP7_75t_L g1077 ( .A(n_812), .Y(n_1077) );
INVx2_ASAP7_75t_L g1183 ( .A(n_812), .Y(n_1183) );
BUFx2_ASAP7_75t_L g898 ( .A(n_815), .Y(n_898) );
INVx1_ASAP7_75t_L g1348 ( .A(n_815), .Y(n_1348) );
AOI33xp33_ASAP7_75t_L g1192 ( .A1(n_817), .A2(n_1193), .A3(n_1197), .B1(n_1199), .B2(n_1201), .B3(n_1202), .Y(n_1192) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
INVx1_ASAP7_75t_L g1181 ( .A(n_820), .Y(n_1181) );
AOI22xp5_ASAP7_75t_L g1168 ( .A1(n_825), .A2(n_1169), .B1(n_1170), .B2(n_1171), .Y(n_1168) );
AOI22xp33_ASAP7_75t_L g1210 ( .A1(n_825), .A2(n_1211), .B1(n_1212), .B2(n_1213), .Y(n_1210) );
AOI22xp33_ASAP7_75t_L g1914 ( .A1(n_825), .A2(n_828), .B1(n_1898), .B2(n_1915), .Y(n_1914) );
INVx1_ASAP7_75t_L g974 ( .A(n_827), .Y(n_974) );
AOI221xp5_ASAP7_75t_L g1068 ( .A1(n_827), .A2(n_828), .B1(n_831), .B2(n_1069), .C(n_1070), .Y(n_1068) );
AOI221xp5_ASAP7_75t_L g1162 ( .A1(n_827), .A2(n_828), .B1(n_831), .B2(n_1163), .C(n_1164), .Y(n_1162) );
AOI221xp5_ASAP7_75t_L g1189 ( .A1(n_827), .A2(n_828), .B1(n_831), .B2(n_1190), .C(n_1191), .Y(n_1189) );
AOI21xp5_ASAP7_75t_L g1926 ( .A1(n_827), .A2(n_831), .B(n_1927), .Y(n_1926) );
INVx1_ASAP7_75t_L g972 ( .A(n_828), .Y(n_972) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
AOI221xp5_ASAP7_75t_L g970 ( .A1(n_831), .A2(n_958), .B1(n_959), .B2(n_971), .C(n_973), .Y(n_970) );
INVx1_ASAP7_75t_L g1432 ( .A(n_832), .Y(n_1432) );
INVx1_ASAP7_75t_SL g900 ( .A(n_833), .Y(n_900) );
XNOR2x1_ASAP7_75t_L g833 ( .A(n_834), .B(n_899), .Y(n_833) );
AND2x2_ASAP7_75t_L g834 ( .A(n_835), .B(n_870), .Y(n_834) );
AOI31xp33_ASAP7_75t_L g837 ( .A1(n_838), .A2(n_850), .A3(n_865), .B(n_868), .Y(n_837) );
INVx2_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
INVx1_ASAP7_75t_SL g1160 ( .A(n_842), .Y(n_1160) );
AOI22xp33_ASAP7_75t_L g1233 ( .A1(n_842), .A2(n_1135), .B1(n_1190), .B2(n_1191), .Y(n_1233) );
INVx4_ASAP7_75t_L g1274 ( .A(n_842), .Y(n_1274) );
OAI211xp5_ASAP7_75t_L g843 ( .A1(n_844), .A2(n_845), .B(n_847), .C(n_848), .Y(n_843) );
OAI221xp5_ASAP7_75t_L g948 ( .A1(n_845), .A2(n_911), .B1(n_916), .B2(n_949), .C(n_951), .Y(n_948) );
INVx2_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx2_ASAP7_75t_SL g967 ( .A(n_846), .Y(n_967) );
INVx1_ASAP7_75t_L g1219 ( .A(n_846), .Y(n_1219) );
BUFx3_ASAP7_75t_L g863 ( .A(n_849), .Y(n_863) );
OAI22xp33_ASAP7_75t_L g895 ( .A1(n_852), .A2(n_866), .B1(n_896), .B2(n_898), .Y(n_895) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
HB1xp67_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx1_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
INVx1_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
OAI221xp5_ASAP7_75t_L g939 ( .A1(n_860), .A2(n_922), .B1(n_940), .B2(n_942), .C(n_943), .Y(n_939) );
INVx1_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
INVx2_ASAP7_75t_SL g1158 ( .A(n_864), .Y(n_1158) );
AOI21xp5_ASAP7_75t_L g1142 ( .A1(n_868), .A2(n_1143), .B(n_1152), .Y(n_1142) );
INVx2_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
OAI31xp33_ASAP7_75t_L g1214 ( .A1(n_869), .A2(n_1215), .A3(n_1216), .B(n_1228), .Y(n_1214) );
NOR3xp33_ASAP7_75t_SL g870 ( .A(n_871), .B(n_878), .C(n_880), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g871 ( .A(n_872), .B(n_875), .Y(n_871) );
OAI22xp33_ASAP7_75t_L g1026 ( .A1(n_882), .A2(n_989), .B1(n_1027), .B2(n_1028), .Y(n_1026) );
INVx1_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
INVx2_ASAP7_75t_L g1497 ( .A(n_883), .Y(n_1497) );
OAI22xp5_ASAP7_75t_L g886 ( .A1(n_887), .A2(n_888), .B1(n_889), .B2(n_891), .Y(n_886) );
BUFx2_ASAP7_75t_L g1108 ( .A(n_887), .Y(n_1108) );
INVx1_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
HB1xp67_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
INVx2_ASAP7_75t_L g1176 ( .A(n_894), .Y(n_1176) );
INVx1_ASAP7_75t_L g896 ( .A(n_897), .Y(n_896) );
OAI22xp33_ASAP7_75t_L g1102 ( .A1(n_898), .A2(n_1103), .B1(n_1105), .B2(n_1106), .Y(n_1102) );
OAI22xp33_ASAP7_75t_L g1554 ( .A1(n_898), .A2(n_1103), .B1(n_1555), .B2(n_1556), .Y(n_1554) );
OAI22xp33_ASAP7_75t_L g1563 ( .A1(n_898), .A2(n_1103), .B1(n_1564), .B2(n_1565), .Y(n_1563) );
INVx1_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
OAI22xp5_ASAP7_75t_L g902 ( .A1(n_903), .A2(n_904), .B1(n_975), .B2(n_976), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
INVx1_ASAP7_75t_L g904 ( .A(n_905), .Y(n_904) );
NAND4xp25_ASAP7_75t_L g906 ( .A(n_907), .B(n_915), .C(n_934), .D(n_970), .Y(n_906) );
AND2x2_ASAP7_75t_L g907 ( .A(n_908), .B(n_912), .Y(n_907) );
OAI221xp5_ASAP7_75t_L g918 ( .A1(n_919), .A2(n_922), .B1(n_923), .B2(n_926), .C(n_927), .Y(n_918) );
OAI22xp5_ASAP7_75t_L g1350 ( .A1(n_919), .A2(n_1351), .B1(n_1352), .B2(n_1354), .Y(n_1350) );
OAI22xp5_ASAP7_75t_L g1499 ( .A1(n_919), .A2(n_1183), .B1(n_1500), .B2(n_1501), .Y(n_1499) );
INVx2_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
INVx2_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
INVx1_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
INVx2_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
INVx2_ASAP7_75t_L g1025 ( .A(n_925), .Y(n_1025) );
INVx3_ASAP7_75t_L g1478 ( .A(n_925), .Y(n_1478) );
OAI31xp33_ASAP7_75t_SL g934 ( .A1(n_935), .A2(n_945), .A3(n_952), .B(n_968), .Y(n_934) );
INVx1_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
OAI21xp5_ASAP7_75t_SL g1048 ( .A1(n_940), .A2(n_1049), .B(n_1050), .Y(n_1048) );
INVx2_ASAP7_75t_SL g940 ( .A(n_941), .Y(n_940) );
INVx1_ASAP7_75t_L g1371 ( .A(n_941), .Y(n_1371) );
INVx1_ASAP7_75t_L g983 ( .A(n_943), .Y(n_983) );
INVx2_ASAP7_75t_SL g943 ( .A(n_944), .Y(n_943) );
BUFx3_ASAP7_75t_L g1526 ( .A(n_944), .Y(n_1526) );
INVx1_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
OAI221xp5_ASAP7_75t_L g1370 ( .A1(n_949), .A2(n_1339), .B1(n_1341), .B2(n_1371), .C(n_1372), .Y(n_1370) );
OAI22xp5_ASAP7_75t_L g1866 ( .A1(n_949), .A2(n_963), .B1(n_1848), .B2(n_1867), .Y(n_1866) );
INVx2_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
NAND3xp33_ASAP7_75t_L g952 ( .A(n_953), .B(n_957), .C(n_960), .Y(n_952) );
A2O1A1Ixp33_ASAP7_75t_L g1897 ( .A1(n_955), .A2(n_1898), .B(n_1899), .C(n_1900), .Y(n_1897) );
BUFx3_ASAP7_75t_L g955 ( .A(n_956), .Y(n_955) );
INVx1_ASAP7_75t_L g963 ( .A(n_964), .Y(n_963) );
INVx1_ASAP7_75t_L g1047 ( .A(n_966), .Y(n_1047) );
AOI22xp5_ASAP7_75t_L g1268 ( .A1(n_968), .A2(n_1269), .B1(n_1282), .B2(n_1283), .Y(n_1268) );
INVx2_ASAP7_75t_L g1382 ( .A(n_968), .Y(n_1382) );
OAI31xp33_ASAP7_75t_L g1506 ( .A1(n_968), .A2(n_1507), .A3(n_1516), .B(n_1519), .Y(n_1506) );
CKINVDCx8_ASAP7_75t_R g968 ( .A(n_969), .Y(n_968) );
INVx1_ASAP7_75t_L g971 ( .A(n_972), .Y(n_971) );
INVx1_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
INVx1_ASAP7_75t_L g975 ( .A(n_976), .Y(n_975) );
INVx2_ASAP7_75t_SL g1031 ( .A(n_977), .Y(n_1031) );
AND2x2_ASAP7_75t_L g977 ( .A(n_978), .B(n_1000), .Y(n_977) );
OAI21xp33_ASAP7_75t_L g978 ( .A1(n_979), .A2(n_991), .B(n_999), .Y(n_978) );
AOI22xp5_ASAP7_75t_L g980 ( .A1(n_981), .A2(n_982), .B1(n_985), .B2(n_986), .Y(n_980) );
INVx2_ASAP7_75t_SL g1045 ( .A(n_997), .Y(n_1045) );
AOI22xp5_ASAP7_75t_L g1118 ( .A1(n_999), .A2(n_1119), .B1(n_1136), .B2(n_1137), .Y(n_1118) );
AOI22xp5_ASAP7_75t_L g1566 ( .A1(n_999), .A2(n_1306), .B1(n_1567), .B2(n_1582), .Y(n_1566) );
NOR2xp33_ASAP7_75t_L g1000 ( .A(n_1001), .B(n_1017), .Y(n_1000) );
INVx2_ASAP7_75t_L g1006 ( .A(n_1007), .Y(n_1006) );
OAI22xp5_ASAP7_75t_L g1107 ( .A1(n_1007), .A2(n_1108), .B1(n_1109), .B2(n_1110), .Y(n_1107) );
OAI22xp5_ASAP7_75t_L g1111 ( .A1(n_1007), .A2(n_1112), .B1(n_1113), .B2(n_1114), .Y(n_1111) );
BUFx3_ASAP7_75t_L g1079 ( .A(n_1009), .Y(n_1079) );
BUFx3_ASAP7_75t_L g1468 ( .A(n_1011), .Y(n_1468) );
INVx1_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
INVx2_ASAP7_75t_SL g1321 ( .A(n_1014), .Y(n_1321) );
INVx2_ASAP7_75t_SL g1014 ( .A(n_1015), .Y(n_1014) );
NAND2xp5_ASAP7_75t_L g1017 ( .A(n_1018), .B(n_1021), .Y(n_1017) );
INVx3_ASAP7_75t_L g1023 ( .A(n_1024), .Y(n_1023) );
INVx1_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
OAI21x1_ASAP7_75t_L g1034 ( .A1(n_1035), .A2(n_1331), .B(n_1385), .Y(n_1034) );
INVx1_ASAP7_75t_L g1035 ( .A(n_1036), .Y(n_1035) );
OR2x2_ASAP7_75t_L g1385 ( .A(n_1036), .B(n_1332), .Y(n_1385) );
XNOR2xp5_ASAP7_75t_L g1036 ( .A(n_1037), .B(n_1138), .Y(n_1036) );
XOR2x2_ASAP7_75t_L g1037 ( .A(n_1038), .B(n_1087), .Y(n_1037) );
XNOR2xp5_ASAP7_75t_L g1038 ( .A(n_1039), .B(n_1086), .Y(n_1038) );
AND2x2_ASAP7_75t_L g1039 ( .A(n_1040), .B(n_1067), .Y(n_1039) );
NAND3xp33_ASAP7_75t_SL g1041 ( .A(n_1042), .B(n_1052), .C(n_1063), .Y(n_1041) );
INVx1_ASAP7_75t_L g1372 ( .A(n_1051), .Y(n_1372) );
INVx1_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1054), .Y(n_1303) );
INVx2_ASAP7_75t_L g1059 ( .A(n_1060), .Y(n_1059) );
INVx1_ASAP7_75t_L g1061 ( .A(n_1062), .Y(n_1061) );
OAI22xp5_ASAP7_75t_L g1527 ( .A1(n_1062), .A2(n_1528), .B1(n_1529), .B2(n_1530), .Y(n_1527) );
INVx1_ASAP7_75t_L g1580 ( .A(n_1062), .Y(n_1580) );
AND4x1_ASAP7_75t_L g1067 ( .A(n_1068), .B(n_1071), .C(n_1080), .D(n_1082), .Y(n_1067) );
INVx2_ASAP7_75t_L g1076 ( .A(n_1077), .Y(n_1076) );
OAI22xp5_ASAP7_75t_L g1329 ( .A1(n_1077), .A2(n_1290), .B1(n_1292), .B2(n_1326), .Y(n_1329) );
XNOR2x1_ASAP7_75t_L g1087 ( .A(n_1088), .B(n_1089), .Y(n_1087) );
AND2x2_ASAP7_75t_L g1089 ( .A(n_1090), .B(n_1118), .Y(n_1089) );
NOR3xp33_ASAP7_75t_L g1090 ( .A(n_1091), .B(n_1098), .C(n_1100), .Y(n_1090) );
NAND2xp5_ASAP7_75t_L g1091 ( .A(n_1092), .B(n_1095), .Y(n_1091) );
INVx1_ASAP7_75t_L g1103 ( .A(n_1104), .Y(n_1103) );
NAND3xp33_ASAP7_75t_L g1119 ( .A(n_1120), .B(n_1124), .C(n_1130), .Y(n_1119) );
INVx1_ASAP7_75t_L g1121 ( .A(n_1122), .Y(n_1121) );
INVx1_ASAP7_75t_L g1122 ( .A(n_1123), .Y(n_1122) );
AOI221xp5_ASAP7_75t_L g1270 ( .A1(n_1123), .A2(n_1259), .B1(n_1271), .B2(n_1272), .C(n_1273), .Y(n_1270) );
INVx2_ASAP7_75t_L g1127 ( .A(n_1128), .Y(n_1127) );
INVx1_ASAP7_75t_L g1128 ( .A(n_1129), .Y(n_1128) );
INVx2_ASAP7_75t_L g1134 ( .A(n_1135), .Y(n_1134) );
INVx2_ASAP7_75t_SL g1275 ( .A(n_1135), .Y(n_1275) );
XOR2xp5_ASAP7_75t_L g1138 ( .A(n_1139), .B(n_1234), .Y(n_1138) );
XNOR2x1_ASAP7_75t_L g1139 ( .A(n_1140), .B(n_1186), .Y(n_1139) );
NOR2x1_ASAP7_75t_L g1141 ( .A(n_1142), .B(n_1161), .Y(n_1141) );
AOI221xp5_ASAP7_75t_L g1143 ( .A1(n_1144), .A2(n_1145), .B1(n_1146), .B2(n_1148), .C(n_1151), .Y(n_1143) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1150), .Y(n_1149) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1151), .Y(n_1227) );
AOI221xp5_ASAP7_75t_L g1299 ( .A1(n_1151), .A2(n_1300), .B1(n_1302), .B2(n_1303), .C(n_1304), .Y(n_1299) );
HB1xp67_ASAP7_75t_L g1155 ( .A(n_1156), .Y(n_1155) );
NAND2xp33_ASAP7_75t_L g1875 ( .A(n_1156), .B(n_1876), .Y(n_1875) );
NAND4xp25_ASAP7_75t_L g1161 ( .A(n_1162), .B(n_1165), .C(n_1168), .D(n_1172), .Y(n_1161) );
AOI22xp5_ASAP7_75t_L g1244 ( .A1(n_1173), .A2(n_1207), .B1(n_1245), .B2(n_1246), .Y(n_1244) );
INVx1_ASAP7_75t_L g1505 ( .A(n_1173), .Y(n_1505) );
AOI22xp5_ASAP7_75t_L g1916 ( .A1(n_1173), .A2(n_1211), .B1(n_1917), .B2(n_1918), .Y(n_1916) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1176), .Y(n_1328) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1182), .Y(n_1257) );
INVx2_ASAP7_75t_L g1182 ( .A(n_1183), .Y(n_1182) );
NAND3xp33_ASAP7_75t_L g1187 ( .A(n_1188), .B(n_1205), .C(n_1214), .Y(n_1187) );
AND3x1_ASAP7_75t_L g1188 ( .A(n_1189), .B(n_1192), .C(n_1203), .Y(n_1188) );
INVx2_ASAP7_75t_L g1195 ( .A(n_1196), .Y(n_1195) );
BUFx3_ASAP7_75t_L g1472 ( .A(n_1200), .Y(n_1472) );
NAND3xp33_ASAP7_75t_L g1850 ( .A(n_1202), .B(n_1851), .C(n_1852), .Y(n_1850) );
AND2x2_ASAP7_75t_L g1205 ( .A(n_1206), .B(n_1210), .Y(n_1205) );
INVx1_ASAP7_75t_L g1486 ( .A(n_1207), .Y(n_1486) );
INVx1_ASAP7_75t_L g1856 ( .A(n_1207), .Y(n_1856) );
INVx1_ASAP7_75t_L g1913 ( .A(n_1207), .Y(n_1913) );
OAI211xp5_ASAP7_75t_L g1222 ( .A1(n_1209), .A2(n_1223), .B(n_1224), .C(n_1225), .Y(n_1222) );
AOI22xp5_ASAP7_75t_L g1240 ( .A1(n_1211), .A2(n_1241), .B1(n_1242), .B2(n_1243), .Y(n_1240) );
INVx2_ASAP7_75t_L g1488 ( .A(n_1211), .Y(n_1488) );
NAND3xp33_ASAP7_75t_L g1216 ( .A(n_1217), .B(n_1222), .C(n_1227), .Y(n_1216) );
OAI211xp5_ASAP7_75t_L g1217 ( .A1(n_1218), .A2(n_1219), .B(n_1220), .C(n_1221), .Y(n_1217) );
OAI211xp5_ASAP7_75t_L g1902 ( .A1(n_1223), .A2(n_1903), .B(n_1904), .C(n_1905), .Y(n_1902) );
XNOR2xp5_ASAP7_75t_L g1234 ( .A(n_1235), .B(n_1284), .Y(n_1234) );
XNOR2x1_ASAP7_75t_L g1235 ( .A(n_1236), .B(n_1237), .Y(n_1235) );
AND2x2_ASAP7_75t_L g1237 ( .A(n_1238), .B(n_1268), .Y(n_1237) );
NOR3xp33_ASAP7_75t_L g1238 ( .A(n_1239), .B(n_1247), .C(n_1248), .Y(n_1238) );
NAND2xp5_ASAP7_75t_L g1239 ( .A(n_1240), .B(n_1244), .Y(n_1239) );
INVx1_ASAP7_75t_L g1857 ( .A(n_1243), .Y(n_1857) );
OAI22xp5_ASAP7_75t_L g1252 ( .A1(n_1253), .A2(n_1254), .B1(n_1256), .B2(n_1257), .Y(n_1252) );
BUFx2_ASAP7_75t_L g1254 ( .A(n_1255), .Y(n_1254) );
OAI22xp5_ASAP7_75t_SL g1258 ( .A1(n_1259), .A2(n_1260), .B1(n_1261), .B2(n_1262), .Y(n_1258) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1263), .Y(n_1262) );
HB1xp67_ASAP7_75t_L g1263 ( .A(n_1264), .Y(n_1263) );
NAND3xp33_ASAP7_75t_L g1269 ( .A(n_1270), .B(n_1276), .C(n_1281), .Y(n_1269) );
NAND2xp5_ASAP7_75t_L g1285 ( .A(n_1286), .B(n_1307), .Y(n_1285) );
NAND3xp33_ASAP7_75t_SL g1287 ( .A(n_1288), .B(n_1291), .C(n_1299), .Y(n_1287) );
NOR3xp33_ASAP7_75t_L g1307 ( .A(n_1308), .B(n_1317), .C(n_1319), .Y(n_1307) );
NAND2xp5_ASAP7_75t_L g1308 ( .A(n_1309), .B(n_1313), .Y(n_1308) );
OAI22xp5_ASAP7_75t_L g1324 ( .A1(n_1325), .A2(n_1326), .B1(n_1327), .B2(n_1328), .Y(n_1324) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1332), .Y(n_1331) );
HB1xp67_ASAP7_75t_L g1332 ( .A(n_1333), .Y(n_1332) );
INVx1_ASAP7_75t_L g1384 ( .A(n_1334), .Y(n_1384) );
AND2x2_ASAP7_75t_L g1334 ( .A(n_1335), .B(n_1361), .Y(n_1334) );
NOR3xp33_ASAP7_75t_L g1335 ( .A(n_1336), .B(n_1343), .C(n_1344), .Y(n_1335) );
NAND2xp5_ASAP7_75t_L g1336 ( .A(n_1337), .B(n_1340), .Y(n_1336) );
INVx1_ASAP7_75t_L g1347 ( .A(n_1348), .Y(n_1347) );
INVx2_ASAP7_75t_SL g1352 ( .A(n_1353), .Y(n_1352) );
AOI31xp33_ASAP7_75t_L g1363 ( .A1(n_1364), .A2(n_1373), .A3(n_1381), .B(n_1382), .Y(n_1363) );
INVx1_ASAP7_75t_L g1368 ( .A(n_1369), .Y(n_1368) );
INVx1_ASAP7_75t_L g1376 ( .A(n_1377), .Y(n_1376) );
INVx1_ASAP7_75t_L g1377 ( .A(n_1378), .Y(n_1377) );
INVx2_ASAP7_75t_L g1378 ( .A(n_1379), .Y(n_1378) );
INVx3_ASAP7_75t_L g1460 ( .A(n_1379), .Y(n_1460) );
OAI22xp5_ASAP7_75t_L g1387 ( .A1(n_1388), .A2(n_1389), .B1(n_1541), .B2(n_1583), .Y(n_1387) );
INVx1_ASAP7_75t_L g1388 ( .A(n_1389), .Y(n_1388) );
AOI22xp5_ASAP7_75t_L g1389 ( .A1(n_1390), .A2(n_1482), .B1(n_1538), .B2(n_1539), .Y(n_1389) );
INVx1_ASAP7_75t_L g1538 ( .A(n_1390), .Y(n_1538) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1391), .Y(n_1390) );
INVxp67_ASAP7_75t_SL g1391 ( .A(n_1392), .Y(n_1391) );
INVx2_ASAP7_75t_L g1481 ( .A(n_1393), .Y(n_1481) );
AO211x2_ASAP7_75t_L g1393 ( .A1(n_1394), .A2(n_1396), .B(n_1428), .C(n_1454), .Y(n_1393) );
NAND4xp25_ASAP7_75t_L g1396 ( .A(n_1397), .B(n_1408), .C(n_1415), .D(n_1425), .Y(n_1396) );
AOI22xp33_ASAP7_75t_L g1397 ( .A1(n_1398), .A2(n_1399), .B1(n_1404), .B2(n_1405), .Y(n_1397) );
HB1xp67_ASAP7_75t_L g1399 ( .A(n_1400), .Y(n_1399) );
AND2x4_ASAP7_75t_L g1400 ( .A(n_1401), .B(n_1403), .Y(n_1400) );
INVx1_ASAP7_75t_SL g1401 ( .A(n_1402), .Y(n_1401) );
INVx1_ASAP7_75t_L g1427 ( .A(n_1406), .Y(n_1427) );
INVx1_ASAP7_75t_L g1406 ( .A(n_1407), .Y(n_1406) );
AOI22xp33_ASAP7_75t_L g1408 ( .A1(n_1409), .A2(n_1410), .B1(n_1413), .B2(n_1414), .Y(n_1408) );
AOI22xp33_ASAP7_75t_SL g1448 ( .A1(n_1409), .A2(n_1449), .B1(n_1450), .B2(n_1451), .Y(n_1448) );
AND2x4_ASAP7_75t_L g1420 ( .A(n_1411), .B(n_1421), .Y(n_1420) );
INVx1_ASAP7_75t_L g1411 ( .A(n_1412), .Y(n_1411) );
AOI222xp33_ASAP7_75t_L g1415 ( .A1(n_1416), .A2(n_1417), .B1(n_1418), .B2(n_1419), .C1(n_1423), .C2(n_1424), .Y(n_1415) );
BUFx4f_ASAP7_75t_L g1419 ( .A(n_1420), .Y(n_1419) );
INVx1_ASAP7_75t_L g1421 ( .A(n_1422), .Y(n_1421) );
INVx5_ASAP7_75t_L g1425 ( .A(n_1426), .Y(n_1425) );
AOI31xp33_ASAP7_75t_L g1428 ( .A1(n_1429), .A2(n_1440), .A3(n_1448), .B(n_1453), .Y(n_1428) );
AOI211xp5_ASAP7_75t_L g1429 ( .A1(n_1430), .A2(n_1431), .B(n_1433), .C(n_1436), .Y(n_1429) );
INVx1_ASAP7_75t_L g1431 ( .A(n_1432), .Y(n_1431) );
INVx1_ASAP7_75t_L g1434 ( .A(n_1435), .Y(n_1434) );
INVx2_ASAP7_75t_L g1437 ( .A(n_1438), .Y(n_1437) );
AOI22xp33_ASAP7_75t_SL g1440 ( .A1(n_1441), .A2(n_1443), .B1(n_1444), .B2(n_1447), .Y(n_1440) );
AND2x4_ASAP7_75t_L g1444 ( .A(n_1442), .B(n_1445), .Y(n_1444) );
INVx1_ASAP7_75t_L g1445 ( .A(n_1446), .Y(n_1445) );
HB1xp67_ASAP7_75t_L g1476 ( .A(n_1446), .Y(n_1476) );
INVx4_ASAP7_75t_L g1451 ( .A(n_1452), .Y(n_1451) );
NAND2xp5_ASAP7_75t_L g1454 ( .A(n_1455), .B(n_1467), .Y(n_1454) );
AOI33xp33_ASAP7_75t_L g1455 ( .A1(n_1456), .A2(n_1457), .A3(n_1461), .B1(n_1464), .B2(n_1465), .B3(n_1466), .Y(n_1455) );
INVx1_ASAP7_75t_L g1458 ( .A(n_1459), .Y(n_1458) );
INVx1_ASAP7_75t_L g1459 ( .A(n_1460), .Y(n_1459) );
INVx1_ASAP7_75t_L g1473 ( .A(n_1474), .Y(n_1473) );
INVx1_ASAP7_75t_L g1474 ( .A(n_1475), .Y(n_1474) );
INVx1_ASAP7_75t_L g1475 ( .A(n_1476), .Y(n_1475) );
INVx2_ASAP7_75t_L g1540 ( .A(n_1482), .Y(n_1540) );
INVx1_ASAP7_75t_L g1536 ( .A(n_1483), .Y(n_1536) );
NAND3xp33_ASAP7_75t_L g1483 ( .A(n_1484), .B(n_1489), .C(n_1506), .Y(n_1483) );
NOR2xp33_ASAP7_75t_L g1484 ( .A(n_1485), .B(n_1487), .Y(n_1484) );
NOR2xp33_ASAP7_75t_L g1489 ( .A(n_1490), .B(n_1491), .Y(n_1489) );
OAI22xp5_ASAP7_75t_L g1520 ( .A1(n_1494), .A2(n_1496), .B1(n_1521), .B2(n_1523), .Y(n_1520) );
AOI22xp33_ASAP7_75t_L g1511 ( .A1(n_1500), .A2(n_1504), .B1(n_1512), .B2(n_1514), .Y(n_1511) );
BUFx2_ASAP7_75t_L g1509 ( .A(n_1510), .Y(n_1509) );
INVx1_ASAP7_75t_L g1512 ( .A(n_1513), .Y(n_1512) );
OAI22xp5_ASAP7_75t_L g1519 ( .A1(n_1520), .A2(n_1524), .B1(n_1527), .B2(n_1531), .Y(n_1519) );
INVx1_ASAP7_75t_L g1521 ( .A(n_1522), .Y(n_1521) );
INVx1_ASAP7_75t_L g1525 ( .A(n_1526), .Y(n_1525) );
BUFx2_ASAP7_75t_L g1539 ( .A(n_1540), .Y(n_1539) );
INVx1_ASAP7_75t_L g1583 ( .A(n_1541), .Y(n_1583) );
HB1xp67_ASAP7_75t_L g1541 ( .A(n_1542), .Y(n_1541) );
AND2x2_ASAP7_75t_L g1543 ( .A(n_1544), .B(n_1566), .Y(n_1543) );
NOR3xp33_ASAP7_75t_SL g1544 ( .A(n_1545), .B(n_1552), .C(n_1553), .Y(n_1544) );
NAND2xp5_ASAP7_75t_L g1545 ( .A(n_1546), .B(n_1549), .Y(n_1545) );
NAND3xp33_ASAP7_75t_L g1567 ( .A(n_1568), .B(n_1574), .C(n_1581), .Y(n_1567) );
INVx1_ASAP7_75t_L g1570 ( .A(n_1571), .Y(n_1570) );
INVx1_ASAP7_75t_L g1575 ( .A(n_1576), .Y(n_1575) );
OAI221xp5_ASAP7_75t_SL g1584 ( .A1(n_1585), .A2(n_1835), .B1(n_1837), .B2(n_1879), .C(n_1883), .Y(n_1584) );
AND4x1_ASAP7_75t_L g1585 ( .A(n_1586), .B(n_1801), .C(n_1820), .D(n_1825), .Y(n_1585) );
AOI211xp5_ASAP7_75t_L g1586 ( .A1(n_1587), .A2(n_1615), .B(n_1748), .C(n_1785), .Y(n_1586) );
OAI221xp5_ASAP7_75t_L g1748 ( .A1(n_1587), .A2(n_1749), .B1(n_1764), .B2(n_1780), .C(n_1935), .Y(n_1748) );
INVx3_ASAP7_75t_L g1587 ( .A(n_1588), .Y(n_1587) );
O2A1O1Ixp33_ASAP7_75t_L g1801 ( .A1(n_1588), .A2(n_1802), .B(n_1807), .C(n_1811), .Y(n_1801) );
INVx2_ASAP7_75t_L g1588 ( .A(n_1589), .Y(n_1588) );
INVx1_ASAP7_75t_L g1589 ( .A(n_1590), .Y(n_1589) );
NAND2xp5_ASAP7_75t_L g1791 ( .A(n_1590), .B(n_1648), .Y(n_1791) );
INVx1_ASAP7_75t_L g1590 ( .A(n_1591), .Y(n_1590) );
NOR2xp33_ASAP7_75t_L g1796 ( .A(n_1591), .B(n_1758), .Y(n_1796) );
NOR3xp33_ASAP7_75t_L g1819 ( .A(n_1591), .B(n_1672), .C(n_1697), .Y(n_1819) );
BUFx3_ASAP7_75t_L g1592 ( .A(n_1593), .Y(n_1592) );
INVx1_ASAP7_75t_L g1651 ( .A(n_1593), .Y(n_1651) );
AND2x4_ASAP7_75t_L g1593 ( .A(n_1594), .B(n_1597), .Y(n_1593) );
AND2x2_ASAP7_75t_L g1628 ( .A(n_1594), .B(n_1597), .Y(n_1628) );
INVx1_ASAP7_75t_L g1594 ( .A(n_1595), .Y(n_1594) );
AND2x4_ASAP7_75t_L g1601 ( .A(n_1595), .B(n_1597), .Y(n_1601) );
INVx1_ASAP7_75t_L g1595 ( .A(n_1596), .Y(n_1595) );
NAND2xp5_ASAP7_75t_L g1608 ( .A(n_1596), .B(n_1609), .Y(n_1608) );
INVx1_ASAP7_75t_L g1609 ( .A(n_1598), .Y(n_1609) );
INVx1_ASAP7_75t_L g1599 ( .A(n_1600), .Y(n_1599) );
INVx2_ASAP7_75t_L g1633 ( .A(n_1600), .Y(n_1633) );
OAI22xp5_ASAP7_75t_SL g1650 ( .A1(n_1600), .A2(n_1651), .B1(n_1652), .B2(n_1653), .Y(n_1650) );
INVx2_ASAP7_75t_L g1600 ( .A(n_1601), .Y(n_1600) );
OAI22xp33_ASAP7_75t_L g1602 ( .A1(n_1603), .A2(n_1604), .B1(n_1610), .B2(n_1611), .Y(n_1602) );
INVx1_ASAP7_75t_L g1836 ( .A(n_1604), .Y(n_1836) );
BUFx3_ASAP7_75t_L g1604 ( .A(n_1605), .Y(n_1604) );
OAI22xp33_ASAP7_75t_L g1634 ( .A1(n_1605), .A2(n_1635), .B1(n_1636), .B2(n_1637), .Y(n_1634) );
BUFx6f_ASAP7_75t_L g1605 ( .A(n_1606), .Y(n_1605) );
OR2x2_ASAP7_75t_L g1606 ( .A(n_1607), .B(n_1608), .Y(n_1606) );
OR2x2_ASAP7_75t_L g1613 ( .A(n_1607), .B(n_1614), .Y(n_1613) );
INVx1_ASAP7_75t_L g1624 ( .A(n_1607), .Y(n_1624) );
INVx1_ASAP7_75t_L g1623 ( .A(n_1608), .Y(n_1623) );
INVx1_ASAP7_75t_L g1611 ( .A(n_1612), .Y(n_1611) );
INVx1_ASAP7_75t_L g1612 ( .A(n_1613), .Y(n_1612) );
HB1xp67_ASAP7_75t_L g1637 ( .A(n_1613), .Y(n_1637) );
INVx1_ASAP7_75t_L g1626 ( .A(n_1614), .Y(n_1626) );
NAND5xp2_ASAP7_75t_L g1615 ( .A(n_1616), .B(n_1668), .C(n_1708), .D(n_1721), .E(n_1737), .Y(n_1615) );
AOI21xp5_ASAP7_75t_L g1616 ( .A1(n_1617), .A2(n_1646), .B(n_1658), .Y(n_1616) );
INVx2_ASAP7_75t_L g1617 ( .A(n_1618), .Y(n_1617) );
OR2x2_ASAP7_75t_L g1618 ( .A(n_1619), .B(n_1629), .Y(n_1618) );
AND2x2_ASAP7_75t_L g1663 ( .A(n_1619), .B(n_1664), .Y(n_1663) );
AND2x2_ASAP7_75t_L g1706 ( .A(n_1619), .B(n_1679), .Y(n_1706) );
AND2x2_ASAP7_75t_L g1722 ( .A(n_1619), .B(n_1666), .Y(n_1722) );
AND2x2_ASAP7_75t_L g1730 ( .A(n_1619), .B(n_1632), .Y(n_1730) );
OR2x2_ASAP7_75t_L g1751 ( .A(n_1619), .B(n_1752), .Y(n_1751) );
AND2x2_ASAP7_75t_L g1756 ( .A(n_1619), .B(n_1681), .Y(n_1756) );
AND2x2_ASAP7_75t_L g1817 ( .A(n_1619), .B(n_1774), .Y(n_1817) );
CKINVDCx5p33_ASAP7_75t_R g1619 ( .A(n_1620), .Y(n_1619) );
HB1xp67_ASAP7_75t_L g1683 ( .A(n_1620), .Y(n_1683) );
AND2x2_ASAP7_75t_L g1691 ( .A(n_1620), .B(n_1631), .Y(n_1691) );
AND2x2_ASAP7_75t_L g1699 ( .A(n_1620), .B(n_1700), .Y(n_1699) );
AND2x2_ASAP7_75t_L g1712 ( .A(n_1620), .B(n_1681), .Y(n_1712) );
AND2x2_ASAP7_75t_L g1720 ( .A(n_1620), .B(n_1679), .Y(n_1720) );
OR2x2_ASAP7_75t_L g1739 ( .A(n_1620), .B(n_1740), .Y(n_1739) );
OR2x2_ASAP7_75t_L g1761 ( .A(n_1620), .B(n_1700), .Y(n_1761) );
NOR2xp33_ASAP7_75t_L g1767 ( .A(n_1620), .B(n_1768), .Y(n_1767) );
NAND2xp5_ASAP7_75t_L g1771 ( .A(n_1620), .B(n_1639), .Y(n_1771) );
NOR2xp33_ASAP7_75t_L g1779 ( .A(n_1620), .B(n_1697), .Y(n_1779) );
AND2x2_ASAP7_75t_L g1797 ( .A(n_1620), .B(n_1697), .Y(n_1797) );
AND2x2_ASAP7_75t_L g1810 ( .A(n_1620), .B(n_1666), .Y(n_1810) );
AND2x4_ASAP7_75t_SL g1620 ( .A(n_1621), .B(n_1627), .Y(n_1620) );
AND2x4_ASAP7_75t_L g1622 ( .A(n_1623), .B(n_1624), .Y(n_1622) );
OAI21xp33_ASAP7_75t_SL g1931 ( .A1(n_1623), .A2(n_1887), .B(n_1932), .Y(n_1931) );
AND2x4_ASAP7_75t_L g1625 ( .A(n_1624), .B(n_1626), .Y(n_1625) );
NAND2xp5_ASAP7_75t_L g1629 ( .A(n_1630), .B(n_1638), .Y(n_1629) );
NOR2xp33_ASAP7_75t_L g1664 ( .A(n_1630), .B(n_1665), .Y(n_1664) );
INVxp67_ASAP7_75t_L g1696 ( .A(n_1630), .Y(n_1696) );
HB1xp67_ASAP7_75t_L g1711 ( .A(n_1630), .Y(n_1711) );
NOR2x1p5_ASAP7_75t_L g1774 ( .A(n_1630), .B(n_1775), .Y(n_1774) );
AND2x2_ASAP7_75t_L g1778 ( .A(n_1630), .B(n_1779), .Y(n_1778) );
AND2x2_ASAP7_75t_L g1787 ( .A(n_1630), .B(n_1703), .Y(n_1787) );
INVx2_ASAP7_75t_SL g1630 ( .A(n_1631), .Y(n_1630) );
BUFx3_ASAP7_75t_L g1672 ( .A(n_1631), .Y(n_1672) );
BUFx2_ASAP7_75t_L g1716 ( .A(n_1631), .Y(n_1716) );
NAND2xp5_ASAP7_75t_L g1760 ( .A(n_1631), .B(n_1660), .Y(n_1760) );
NOR2xp33_ASAP7_75t_L g1772 ( .A(n_1631), .B(n_1704), .Y(n_1772) );
INVx2_ASAP7_75t_SL g1631 ( .A(n_1632), .Y(n_1631) );
INVx2_ASAP7_75t_L g1775 ( .A(n_1638), .Y(n_1775) );
AND2x2_ASAP7_75t_L g1781 ( .A(n_1638), .B(n_1691), .Y(n_1781) );
AND2x2_ASAP7_75t_L g1638 ( .A(n_1639), .B(n_1642), .Y(n_1638) );
INVxp67_ASAP7_75t_SL g1667 ( .A(n_1639), .Y(n_1667) );
AND2x2_ASAP7_75t_L g1679 ( .A(n_1639), .B(n_1643), .Y(n_1679) );
INVx1_ASAP7_75t_L g1682 ( .A(n_1639), .Y(n_1682) );
INVx1_ASAP7_75t_L g1740 ( .A(n_1639), .Y(n_1740) );
AND2x2_ASAP7_75t_L g1639 ( .A(n_1640), .B(n_1641), .Y(n_1639) );
AND2x2_ASAP7_75t_L g1681 ( .A(n_1642), .B(n_1682), .Y(n_1681) );
INVx1_ASAP7_75t_L g1697 ( .A(n_1642), .Y(n_1697) );
INVx1_ASAP7_75t_L g1642 ( .A(n_1643), .Y(n_1642) );
AND2x2_ASAP7_75t_L g1666 ( .A(n_1643), .B(n_1667), .Y(n_1666) );
AND2x2_ASAP7_75t_L g1643 ( .A(n_1644), .B(n_1645), .Y(n_1643) );
AOI221xp5_ASAP7_75t_L g1764 ( .A1(n_1646), .A2(n_1765), .B1(n_1773), .B2(n_1774), .C(n_1776), .Y(n_1764) );
AND2x2_ASAP7_75t_L g1646 ( .A(n_1647), .B(n_1654), .Y(n_1646) );
NAND2xp5_ASAP7_75t_SL g1724 ( .A(n_1647), .B(n_1703), .Y(n_1724) );
AND2x2_ASAP7_75t_L g1731 ( .A(n_1647), .B(n_1704), .Y(n_1731) );
AND2x2_ASAP7_75t_L g1747 ( .A(n_1647), .B(n_1717), .Y(n_1747) );
AND2x2_ASAP7_75t_L g1815 ( .A(n_1647), .B(n_1660), .Y(n_1815) );
O2A1O1Ixp33_ASAP7_75t_L g1833 ( .A1(n_1647), .A2(n_1705), .B(n_1761), .C(n_1834), .Y(n_1833) );
CKINVDCx6p67_ASAP7_75t_R g1647 ( .A(n_1648), .Y(n_1647) );
OR2x2_ASAP7_75t_L g1685 ( .A(n_1648), .B(n_1654), .Y(n_1685) );
NAND2xp5_ASAP7_75t_L g1695 ( .A(n_1648), .B(n_1696), .Y(n_1695) );
AND2x2_ASAP7_75t_L g1702 ( .A(n_1648), .B(n_1703), .Y(n_1702) );
NAND2xp5_ASAP7_75t_L g1718 ( .A(n_1648), .B(n_1688), .Y(n_1718) );
AND2x2_ASAP7_75t_L g1734 ( .A(n_1648), .B(n_1654), .Y(n_1734) );
AND2x2_ASAP7_75t_L g1743 ( .A(n_1648), .B(n_1655), .Y(n_1743) );
CKINVDCx5p33_ASAP7_75t_R g1773 ( .A(n_1648), .Y(n_1773) );
OR2x2_ASAP7_75t_L g1800 ( .A(n_1648), .B(n_1674), .Y(n_1800) );
OR2x6_ASAP7_75t_L g1648 ( .A(n_1649), .B(n_1650), .Y(n_1648) );
OR2x2_ASAP7_75t_L g1806 ( .A(n_1649), .B(n_1650), .Y(n_1806) );
INVx1_ASAP7_75t_L g1758 ( .A(n_1654), .Y(n_1758) );
INVx1_ASAP7_75t_L g1654 ( .A(n_1655), .Y(n_1654) );
INVx1_ASAP7_75t_L g1675 ( .A(n_1655), .Y(n_1675) );
AND2x2_ASAP7_75t_L g1694 ( .A(n_1655), .B(n_1660), .Y(n_1694) );
BUFx6f_ASAP7_75t_L g1713 ( .A(n_1655), .Y(n_1713) );
AND2x2_ASAP7_75t_L g1717 ( .A(n_1655), .B(n_1704), .Y(n_1717) );
AND2x2_ASAP7_75t_L g1655 ( .A(n_1656), .B(n_1657), .Y(n_1655) );
AND2x2_ASAP7_75t_L g1658 ( .A(n_1659), .B(n_1663), .Y(n_1658) );
NAND2xp67_ASAP7_75t_L g1827 ( .A(n_1659), .B(n_1690), .Y(n_1827) );
INVx1_ASAP7_75t_L g1659 ( .A(n_1660), .Y(n_1659) );
NAND2xp5_ASAP7_75t_L g1674 ( .A(n_1660), .B(n_1675), .Y(n_1674) );
INVx1_ASAP7_75t_L g1689 ( .A(n_1660), .Y(n_1689) );
INVx1_ASAP7_75t_L g1704 ( .A(n_1660), .Y(n_1704) );
AND2x2_ASAP7_75t_L g1660 ( .A(n_1661), .B(n_1662), .Y(n_1660) );
INVx1_ASAP7_75t_L g1830 ( .A(n_1663), .Y(n_1830) );
OR2x2_ASAP7_75t_L g1752 ( .A(n_1665), .B(n_1716), .Y(n_1752) );
INVx1_ASAP7_75t_L g1665 ( .A(n_1666), .Y(n_1665) );
AND2x2_ASAP7_75t_L g1690 ( .A(n_1666), .B(n_1691), .Y(n_1690) );
AND2x2_ASAP7_75t_L g1744 ( .A(n_1666), .B(n_1730), .Y(n_1744) );
AOI321xp33_ASAP7_75t_L g1668 ( .A1(n_1669), .A2(n_1676), .A3(n_1683), .B1(n_1684), .B2(n_1686), .C(n_1692), .Y(n_1668) );
INVx1_ASAP7_75t_L g1834 ( .A(n_1669), .Y(n_1834) );
INVx1_ASAP7_75t_L g1669 ( .A(n_1670), .Y(n_1669) );
NAND2xp5_ASAP7_75t_L g1670 ( .A(n_1671), .B(n_1673), .Y(n_1670) );
AND2x2_ASAP7_75t_L g1832 ( .A(n_1671), .B(n_1681), .Y(n_1832) );
INVx1_ASAP7_75t_L g1671 ( .A(n_1672), .Y(n_1671) );
NAND2xp5_ASAP7_75t_L g1698 ( .A(n_1672), .B(n_1699), .Y(n_1698) );
A2O1A1Ixp33_ASAP7_75t_L g1753 ( .A1(n_1672), .A2(n_1754), .B(n_1755), .C(n_1757), .Y(n_1753) );
NAND2xp5_ASAP7_75t_L g1804 ( .A(n_1672), .B(n_1703), .Y(n_1804) );
AND2x2_ASAP7_75t_L g1813 ( .A(n_1672), .B(n_1756), .Y(n_1813) );
INVx1_ASAP7_75t_L g1673 ( .A(n_1674), .Y(n_1673) );
INVx2_ASAP7_75t_L g1707 ( .A(n_1674), .Y(n_1707) );
INVx1_ASAP7_75t_L g1793 ( .A(n_1674), .Y(n_1793) );
AND2x2_ASAP7_75t_L g1703 ( .A(n_1675), .B(n_1704), .Y(n_1703) );
INVx1_ASAP7_75t_L g1676 ( .A(n_1677), .Y(n_1676) );
NAND2xp5_ASAP7_75t_L g1677 ( .A(n_1678), .B(n_1680), .Y(n_1677) );
OR2x2_ASAP7_75t_L g1728 ( .A(n_1678), .B(n_1729), .Y(n_1728) );
INVx1_ASAP7_75t_L g1678 ( .A(n_1679), .Y(n_1678) );
NAND2xp5_ASAP7_75t_L g1746 ( .A(n_1679), .B(n_1747), .Y(n_1746) );
INVx1_ASAP7_75t_L g1680 ( .A(n_1681), .Y(n_1680) );
AND2x2_ASAP7_75t_L g1727 ( .A(n_1681), .B(n_1691), .Y(n_1727) );
NAND2xp5_ASAP7_75t_L g1777 ( .A(n_1684), .B(n_1778), .Y(n_1777) );
AOI222xp33_ASAP7_75t_L g1780 ( .A1(n_1684), .A2(n_1694), .B1(n_1781), .B2(n_1782), .C1(n_1783), .C2(n_1784), .Y(n_1780) );
INVx1_ASAP7_75t_L g1684 ( .A(n_1685), .Y(n_1684) );
INVxp67_ASAP7_75t_SL g1686 ( .A(n_1687), .Y(n_1686) );
NAND2xp5_ASAP7_75t_L g1687 ( .A(n_1688), .B(n_1690), .Y(n_1687) );
INVx1_ASAP7_75t_L g1790 ( .A(n_1688), .Y(n_1790) );
INVx3_ASAP7_75t_L g1688 ( .A(n_1689), .Y(n_1688) );
NAND2xp5_ASAP7_75t_L g1742 ( .A(n_1689), .B(n_1743), .Y(n_1742) );
OAI21xp33_ASAP7_75t_L g1765 ( .A1(n_1689), .A2(n_1766), .B(n_1769), .Y(n_1765) );
AOI32xp33_ASAP7_75t_L g1788 ( .A1(n_1689), .A2(n_1726), .A3(n_1752), .B1(n_1755), .B2(n_1789), .Y(n_1788) );
AND2x2_ASAP7_75t_L g1824 ( .A(n_1689), .B(n_1813), .Y(n_1824) );
OAI321xp33_ASAP7_75t_L g1692 ( .A1(n_1693), .A2(n_1695), .A3(n_1697), .B1(n_1698), .B2(n_1701), .C(n_1705), .Y(n_1692) );
INVx1_ASAP7_75t_L g1693 ( .A(n_1694), .Y(n_1693) );
AOI221xp5_ASAP7_75t_SL g1737 ( .A1(n_1694), .A2(n_1738), .B1(n_1741), .B2(n_1744), .C(n_1745), .Y(n_1737) );
NAND2xp5_ASAP7_75t_L g1763 ( .A(n_1694), .B(n_1706), .Y(n_1763) );
INVx1_ASAP7_75t_L g1700 ( .A(n_1697), .Y(n_1700) );
INVx1_ASAP7_75t_L g1701 ( .A(n_1702), .Y(n_1701) );
NAND2xp5_ASAP7_75t_L g1705 ( .A(n_1706), .B(n_1707), .Y(n_1705) );
AOI21xp5_ASAP7_75t_L g1708 ( .A1(n_1709), .A2(n_1713), .B(n_1714), .Y(n_1708) );
INVx1_ASAP7_75t_L g1709 ( .A(n_1710), .Y(n_1709) );
NAND2xp5_ASAP7_75t_L g1710 ( .A(n_1711), .B(n_1712), .Y(n_1710) );
NAND2xp5_ASAP7_75t_L g1822 ( .A(n_1712), .B(n_1823), .Y(n_1822) );
AOI211xp5_ASAP7_75t_L g1749 ( .A1(n_1713), .A2(n_1750), .B(n_1753), .C(n_1762), .Y(n_1749) );
CKINVDCx14_ASAP7_75t_R g1828 ( .A(n_1713), .Y(n_1828) );
AOI21xp5_ASAP7_75t_L g1714 ( .A1(n_1715), .A2(n_1718), .B(n_1719), .Y(n_1714) );
NAND2xp5_ASAP7_75t_L g1715 ( .A(n_1716), .B(n_1717), .Y(n_1715) );
INVx2_ASAP7_75t_L g1736 ( .A(n_1716), .Y(n_1736) );
NOR2xp33_ASAP7_75t_L g1738 ( .A(n_1716), .B(n_1739), .Y(n_1738) );
NAND2xp5_ASAP7_75t_L g1766 ( .A(n_1716), .B(n_1767), .Y(n_1766) );
INVx1_ASAP7_75t_L g1754 ( .A(n_1717), .Y(n_1754) );
OAI21xp33_ASAP7_75t_L g1798 ( .A1(n_1717), .A2(n_1750), .B(n_1799), .Y(n_1798) );
INVx1_ASAP7_75t_L g1784 ( .A(n_1718), .Y(n_1784) );
INVx1_ASAP7_75t_L g1719 ( .A(n_1720), .Y(n_1719) );
AND2x2_ASAP7_75t_L g1735 ( .A(n_1720), .B(n_1736), .Y(n_1735) );
NOR2xp33_ASAP7_75t_L g1795 ( .A(n_1720), .B(n_1756), .Y(n_1795) );
AOI221xp5_ASAP7_75t_L g1721 ( .A1(n_1722), .A2(n_1723), .B1(n_1725), .B2(n_1731), .C(n_1732), .Y(n_1721) );
INVx1_ASAP7_75t_L g1723 ( .A(n_1724), .Y(n_1723) );
NAND2xp5_ASAP7_75t_SL g1725 ( .A(n_1726), .B(n_1728), .Y(n_1725) );
INVx1_ASAP7_75t_L g1726 ( .A(n_1727), .Y(n_1726) );
INVxp67_ASAP7_75t_SL g1783 ( .A(n_1728), .Y(n_1783) );
INVx1_ASAP7_75t_L g1729 ( .A(n_1730), .Y(n_1729) );
INVx1_ASAP7_75t_L g1808 ( .A(n_1731), .Y(n_1808) );
INVxp67_ASAP7_75t_SL g1732 ( .A(n_1733), .Y(n_1732) );
NAND2xp5_ASAP7_75t_L g1733 ( .A(n_1734), .B(n_1735), .Y(n_1733) );
OAI221xp5_ASAP7_75t_L g1785 ( .A1(n_1736), .A2(n_1786), .B1(n_1791), .B2(n_1792), .C(n_1798), .Y(n_1785) );
INVx1_ASAP7_75t_L g1768 ( .A(n_1740), .Y(n_1768) );
INVx1_ASAP7_75t_L g1741 ( .A(n_1742), .Y(n_1741) );
OAI31xp33_ASAP7_75t_L g1820 ( .A1(n_1743), .A2(n_1750), .A3(n_1821), .B(n_1824), .Y(n_1820) );
INVx1_ASAP7_75t_L g1745 ( .A(n_1746), .Y(n_1745) );
AOI221xp5_ASAP7_75t_L g1825 ( .A1(n_1747), .A2(n_1826), .B1(n_1828), .B2(n_1829), .C(n_1833), .Y(n_1825) );
INVx1_ASAP7_75t_L g1750 ( .A(n_1751), .Y(n_1750) );
INVx1_ASAP7_75t_L g1755 ( .A(n_1756), .Y(n_1755) );
OAI21xp33_ASAP7_75t_L g1818 ( .A1(n_1756), .A2(n_1799), .B(n_1819), .Y(n_1818) );
NAND2xp5_ASAP7_75t_L g1757 ( .A(n_1758), .B(n_1759), .Y(n_1757) );
NOR2xp33_ASAP7_75t_L g1759 ( .A(n_1760), .B(n_1761), .Y(n_1759) );
INVxp67_ASAP7_75t_SL g1762 ( .A(n_1763), .Y(n_1762) );
INVx1_ASAP7_75t_L g1803 ( .A(n_1768), .Y(n_1803) );
INVxp67_ASAP7_75t_SL g1782 ( .A(n_1769), .Y(n_1782) );
NAND2xp5_ASAP7_75t_L g1769 ( .A(n_1770), .B(n_1772), .Y(n_1769) );
INVx1_ASAP7_75t_L g1770 ( .A(n_1771), .Y(n_1770) );
AOI21xp33_ASAP7_75t_SL g1786 ( .A1(n_1771), .A2(n_1787), .B(n_1788), .Y(n_1786) );
INVxp67_ASAP7_75t_SL g1776 ( .A(n_1777), .Y(n_1776) );
INVx1_ASAP7_75t_L g1805 ( .A(n_1781), .Y(n_1805) );
INVx1_ASAP7_75t_L g1789 ( .A(n_1790), .Y(n_1789) );
INVx1_ASAP7_75t_L g1823 ( .A(n_1790), .Y(n_1823) );
AOI22xp33_ASAP7_75t_L g1792 ( .A1(n_1793), .A2(n_1794), .B1(n_1796), .B2(n_1797), .Y(n_1792) );
INVxp33_ASAP7_75t_L g1794 ( .A(n_1795), .Y(n_1794) );
INVx1_ASAP7_75t_L g1799 ( .A(n_1800), .Y(n_1799) );
O2A1O1Ixp33_ASAP7_75t_SL g1802 ( .A1(n_1803), .A2(n_1804), .B(n_1805), .C(n_1806), .Y(n_1802) );
NOR2xp33_ASAP7_75t_L g1807 ( .A(n_1808), .B(n_1809), .Y(n_1807) );
OAI221xp5_ASAP7_75t_L g1811 ( .A1(n_1808), .A2(n_1812), .B1(n_1814), .B2(n_1816), .C(n_1818), .Y(n_1811) );
INVx1_ASAP7_75t_L g1809 ( .A(n_1810), .Y(n_1809) );
INVx1_ASAP7_75t_L g1812 ( .A(n_1813), .Y(n_1812) );
CKINVDCx5p33_ASAP7_75t_R g1814 ( .A(n_1815), .Y(n_1814) );
INVx1_ASAP7_75t_L g1816 ( .A(n_1817), .Y(n_1816) );
INVx1_ASAP7_75t_L g1821 ( .A(n_1822), .Y(n_1821) );
INVx1_ASAP7_75t_L g1826 ( .A(n_1827), .Y(n_1826) );
NAND2xp5_ASAP7_75t_L g1829 ( .A(n_1830), .B(n_1831), .Y(n_1829) );
INVxp67_ASAP7_75t_L g1831 ( .A(n_1832), .Y(n_1831) );
CKINVDCx5p33_ASAP7_75t_R g1835 ( .A(n_1836), .Y(n_1835) );
INVxp67_ASAP7_75t_SL g1837 ( .A(n_1838), .Y(n_1837) );
INVx1_ASAP7_75t_L g1838 ( .A(n_1839), .Y(n_1838) );
HB1xp67_ASAP7_75t_L g1839 ( .A(n_1840), .Y(n_1839) );
NAND3xp33_ASAP7_75t_L g1841 ( .A(n_1842), .B(n_1854), .C(n_1859), .Y(n_1841) );
NOR2xp33_ASAP7_75t_L g1842 ( .A(n_1843), .B(n_1853), .Y(n_1842) );
OAI221xp5_ASAP7_75t_L g1844 ( .A1(n_1845), .A2(n_1846), .B1(n_1847), .B2(n_1848), .C(n_1849), .Y(n_1844) );
NOR2xp33_ASAP7_75t_SL g1854 ( .A(n_1855), .B(n_1858), .Y(n_1854) );
OAI211xp5_ASAP7_75t_SL g1862 ( .A1(n_1863), .A2(n_1866), .B(n_1868), .C(n_1873), .Y(n_1862) );
OAI211xp5_ASAP7_75t_L g1868 ( .A1(n_1869), .A2(n_1870), .B(n_1871), .C(n_1872), .Y(n_1868) );
INVx2_ASAP7_75t_L g1879 ( .A(n_1880), .Y(n_1879) );
INVx1_ASAP7_75t_L g1880 ( .A(n_1881), .Y(n_1880) );
INVx1_ASAP7_75t_L g1881 ( .A(n_1882), .Y(n_1881) );
INVx1_ASAP7_75t_L g1884 ( .A(n_1885), .Y(n_1884) );
CKINVDCx5p33_ASAP7_75t_R g1885 ( .A(n_1886), .Y(n_1885) );
INVxp33_ASAP7_75t_L g1888 ( .A(n_1889), .Y(n_1888) );
INVx1_ASAP7_75t_L g1929 ( .A(n_1890), .Y(n_1929) );
HB1xp67_ASAP7_75t_L g1890 ( .A(n_1891), .Y(n_1890) );
NAND4xp25_ASAP7_75t_L g1892 ( .A(n_1893), .B(n_1897), .C(n_1902), .D(n_1906), .Y(n_1892) );
OAI211xp5_ASAP7_75t_L g1906 ( .A1(n_1907), .A2(n_1908), .B(n_1910), .C(n_1911), .Y(n_1906) );
INVx2_ASAP7_75t_L g1908 ( .A(n_1909), .Y(n_1908) );
NAND2xp5_ASAP7_75t_L g1919 ( .A(n_1920), .B(n_1926), .Y(n_1919) );
HB1xp67_ASAP7_75t_L g1930 ( .A(n_1931), .Y(n_1930) );
endmodule