module real_jpeg_28344_n_17 (n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_340, n_11, n_14, n_7, n_3, n_5, n_4, n_339, n_1, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_340;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_339;
input n_1;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_0),
.A2(n_55),
.B1(n_57),
.B2(n_78),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_0),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_0),
.A2(n_50),
.B1(n_51),
.B2(n_78),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_0),
.A2(n_24),
.B1(n_25),
.B2(n_78),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_0),
.A2(n_28),
.B1(n_29),
.B2(n_78),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_1),
.A2(n_55),
.B1(n_57),
.B2(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_1),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_1),
.A2(n_50),
.B1(n_51),
.B2(n_66),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_1),
.A2(n_24),
.B1(n_25),
.B2(n_66),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_1),
.A2(n_28),
.B1(n_29),
.B2(n_66),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_2),
.B(n_57),
.Y(n_56)
);

A2O1A1O1Ixp25_ASAP7_75t_L g59 ( 
.A1(n_2),
.A2(n_56),
.B(n_57),
.C(n_60),
.D(n_64),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_2),
.B(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_2),
.Y(n_103)
);

OAI21xp33_ASAP7_75t_L g108 ( 
.A1(n_2),
.A2(n_82),
.B(n_86),
.Y(n_108)
);

A2O1A1O1Ixp25_ASAP7_75t_L g118 ( 
.A1(n_2),
.A2(n_25),
.B(n_119),
.C(n_120),
.D(n_123),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_2),
.B(n_25),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_2),
.B(n_21),
.Y(n_148)
);

O2A1O1Ixp33_ASAP7_75t_SL g171 ( 
.A1(n_2),
.A2(n_23),
.B(n_29),
.C(n_172),
.Y(n_171)
);

OAI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_103),
.Y(n_177)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_3),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_4),
.A2(n_50),
.B1(n_51),
.B2(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_4),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_4),
.A2(n_55),
.B1(n_57),
.B2(n_133),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_133),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_4),
.A2(n_28),
.B1(n_29),
.B2(n_133),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_5),
.A2(n_50),
.B1(n_51),
.B2(n_170),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_5),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_5),
.A2(n_55),
.B1(n_57),
.B2(n_170),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_5),
.A2(n_24),
.B1(n_25),
.B2(n_170),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_170),
.Y(n_309)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_7),
.A2(n_31),
.B1(n_50),
.B2(n_51),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_7),
.A2(n_31),
.B1(n_55),
.B2(n_57),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_7),
.A2(n_24),
.B1(n_25),
.B2(n_31),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_10),
.A2(n_50),
.B1(n_51),
.B2(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_10),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_10),
.A2(n_55),
.B1(n_57),
.B2(n_152),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_152),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_152),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_11),
.A2(n_28),
.B1(n_29),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_11),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_11),
.A2(n_35),
.B1(n_50),
.B2(n_51),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_11),
.A2(n_35),
.B1(n_55),
.B2(n_57),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_11),
.A2(n_24),
.B1(n_25),
.B2(n_35),
.Y(n_294)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_12),
.B(n_51),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_12),
.B(n_57),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_12),
.A2(n_50),
.B1(n_51),
.B2(n_54),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_13),
.A2(n_50),
.B1(n_51),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_13),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_13),
.A2(n_55),
.B1(n_57),
.B2(n_85),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_13),
.A2(n_24),
.B1(n_25),
.B2(n_85),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_85),
.Y(n_221)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_15),
.A2(n_24),
.B1(n_25),
.B2(n_122),
.Y(n_121)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_15),
.Y(n_122)
);

INVx11_ASAP7_75t_SL g53 ( 
.A(n_16),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_38),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_36),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_32),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_20),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_26),
.B(n_30),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_21),
.B(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_21),
.A2(n_26),
.B1(n_30),
.B2(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_21),
.B(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_21),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_21),
.A2(n_26),
.B1(n_203),
.B2(n_221),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_21),
.A2(n_26),
.B1(n_34),
.B2(n_330),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_22),
.A2(n_23),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

OAI21xp33_ASAP7_75t_L g172 ( 
.A1(n_22),
.A2(n_25),
.B(n_103),
.Y(n_172)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx5_ASAP7_75t_SL g25 ( 
.A(n_24),
.Y(n_25)
);

AOI32xp33_ASAP7_75t_L g134 ( 
.A1(n_24),
.A2(n_57),
.A3(n_119),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_26),
.A2(n_177),
.B(n_178),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_26),
.B(n_180),
.Y(n_205)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_26),
.Y(n_244)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_28),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_33),
.B(n_336),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_33),
.B(n_336),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_335),
.B(n_337),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_323),
.B(n_334),
.Y(n_39)
);

OAI321xp33_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_287),
.A3(n_316),
.B1(n_321),
.B2(n_322),
.C(n_339),
.Y(n_40)
);

AOI321xp33_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_237),
.A3(n_276),
.B1(n_281),
.B2(n_286),
.C(n_340),
.Y(n_41)
);

NOR3xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_190),
.C(n_233),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_161),
.B(n_189),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_138),
.B(n_160),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_114),
.B(n_137),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_92),
.B(n_113),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_68),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_48),
.B(n_68),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_49),
.B(n_59),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_49),
.B(n_59),
.Y(n_99)
);

AOI32xp33_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_54),
.A3(n_55),
.B1(n_56),
.B2(n_58),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_50),
.B(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2x1_ASAP7_75t_SL g82 ( 
.A(n_51),
.B(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_55),
.A2(n_57),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

NAND2xp33_ASAP7_75t_SL g136 ( 
.A(n_55),
.B(n_74),
.Y(n_136)
);

O2A1O1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_57),
.A2(n_61),
.B(n_62),
.C(n_63),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_60),
.B(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_60),
.A2(n_63),
.B1(n_127),
.B2(n_128),
.Y(n_126)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_60),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_60),
.A2(n_63),
.B1(n_252),
.B2(n_253),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_60),
.A2(n_63),
.B1(n_253),
.B2(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_64),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_67),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_65),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_67),
.A2(n_77),
.B(n_79),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_67),
.B(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_67),
.A2(n_79),
.B(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_67),
.A2(n_157),
.B1(n_188),
.B2(n_212),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_67),
.A2(n_157),
.B1(n_212),
.B2(n_229),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_67),
.A2(n_157),
.B(n_262),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_81),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_75),
.B2(n_76),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_70),
.B(n_76),
.C(n_81),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_72),
.B(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_72),
.A2(n_120),
.B1(n_184),
.B2(n_185),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_72),
.A2(n_120),
.B1(n_264),
.B2(n_265),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_72),
.A2(n_120),
.B1(n_265),
.B2(n_294),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_72),
.A2(n_120),
.B(n_328),
.Y(n_327)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_77),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_84),
.B(n_86),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_82),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_88),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_82),
.A2(n_132),
.B1(n_151),
.B2(n_153),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_82),
.A2(n_90),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_82),
.A2(n_153),
.B1(n_210),
.B2(n_227),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_82),
.A2(n_90),
.B(n_227),
.Y(n_255)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_83),
.A2(n_96),
.B(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_103),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_84),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_89),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_89),
.A2(n_95),
.B1(n_97),
.B2(n_98),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_89),
.A2(n_106),
.B(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx5_ASAP7_75t_SL g153 ( 
.A(n_91),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_91),
.A2(n_97),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_100),
.B(n_112),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_99),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_94),
.B(n_99),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g100 ( 
.A1(n_101),
.A2(n_107),
.B(n_111),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_104),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_102),
.B(n_104),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_115),
.B(n_116),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_129),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_126),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_126),
.C(n_129),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_120),
.B(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_120),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_123),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_124),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_125),
.A2(n_143),
.B(n_144),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_125),
.A2(n_144),
.B(n_224),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_125),
.A2(n_198),
.B1(n_224),
.B2(n_247),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_125),
.A2(n_198),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_128),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_134),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_130),
.B(n_134),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_139),
.B(n_140),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_154),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_155),
.C(n_156),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_142),
.B(n_146),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_142),
.B(n_147),
.C(n_150),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_143),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_149),
.B2(n_150),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_151),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_158),
.B(n_159),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_162),
.B(n_163),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_175),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_166),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_165),
.B(n_166),
.C(n_175),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_171),
.B1(n_173),
.B2(n_174),
.Y(n_166)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_167),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_169),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_171),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_173),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g175 ( 
.A(n_176),
.B(n_181),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_176),
.B(n_183),
.C(n_186),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_179),
.A2(n_244),
.B(n_245),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_186),
.B2(n_187),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_185),
.Y(n_199)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_191),
.A2(n_283),
.B(n_284),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_214),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_192),
.B(n_214),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_207),
.C(n_213),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_193),
.B(n_236),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_194),
.B(n_196),
.C(n_206),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_201),
.B2(n_206),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_199),
.B(n_200),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_201),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_204),
.B(n_205),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_204),
.A2(n_205),
.B(n_272),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_204),
.A2(n_244),
.B1(n_272),
.B2(n_299),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_204),
.A2(n_244),
.B1(n_299),
.B2(n_309),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_207),
.B(n_213),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_211),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_208),
.B(n_211),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_230),
.B1(n_231),
.B2(n_232),
.Y(n_214)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_215),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g215 ( 
.A(n_216),
.B(n_225),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_216),
.B(n_225),
.C(n_232),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_217),
.B(n_220),
.C(n_222),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_222),
.B2(n_223),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_221),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_228),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_228),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_229),
.Y(n_252)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_230),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_234),
.B(n_235),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_257),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_238),
.B(n_257),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_249),
.C(n_256),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_239),
.B(n_249),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_242),
.B2(n_248),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_240),
.Y(n_248)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_243),
.B(n_246),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_243),
.B(n_246),
.C(n_248),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_247),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_254),
.B2(n_255),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_255),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_254),
.A2(n_255),
.B1(n_270),
.B2(n_271),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

AOI21xp33_ASAP7_75t_L g303 ( 
.A1(n_255),
.A2(n_270),
.B(n_273),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_280),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_275),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_267),
.B1(n_268),
.B2(n_274),
.Y(n_258)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_259),
.Y(n_274)
);

OAI21xp33_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_263),
.B(n_266),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_260),
.B(n_263),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_266),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_266),
.A2(n_289),
.B1(n_290),
.B2(n_301),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_267),
.B(n_274),
.C(n_275),
.Y(n_317)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_273),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_277),
.A2(n_282),
.B(n_285),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_278),
.B(n_279),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_304),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_288),
.B(n_304),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_301),
.C(n_302),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_291),
.A2(n_292),
.B1(n_298),
.B2(n_300),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_295),
.B1(n_296),
.B2(n_297),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_293),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_293),
.B(n_297),
.C(n_298),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_294),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_295),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_295),
.A2(n_297),
.B1(n_311),
.B2(n_312),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_297),
.B(n_308),
.C(n_312),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_298),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_298),
.A2(n_300),
.B1(n_306),
.B2(n_307),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_298),
.B(n_307),
.C(n_315),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_302),
.A2(n_303),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_315),
.Y(n_304)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_310),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_309),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_312),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_314),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_317),
.B(n_318),
.Y(n_321)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_324),
.B(n_325),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_333),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_327),
.A2(n_329),
.B1(n_331),
.B2(n_332),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_327),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_329),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_329),
.B(n_332),
.C(n_333),
.Y(n_336)
);


endmodule