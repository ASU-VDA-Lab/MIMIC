module fake_jpeg_31710_n_505 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_505);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_505;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx13_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx6_ASAP7_75t_SL g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_8),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_12),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_3),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_54),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_55),
.Y(n_149)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_56),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_16),
.B(n_26),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_57),
.B(n_95),
.Y(n_163)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_60),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_61),
.Y(n_138)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_62),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_63),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g145 ( 
.A(n_64),
.Y(n_145)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_65),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_24),
.B(n_0),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_66),
.B(n_83),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_67),
.Y(n_142)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_68),
.Y(n_151)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g158 ( 
.A(n_72),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_24),
.B(n_0),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_73),
.B(n_105),
.Y(n_115)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_74),
.Y(n_156)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_50),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_77),
.Y(n_112)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_29),
.Y(n_78)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_29),
.Y(n_79)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_79),
.Y(n_140)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_80),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx8_ASAP7_75t_L g153 ( 
.A(n_81),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_82),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_35),
.B(n_3),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_19),
.Y(n_84)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_84),
.Y(n_159)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_32),
.Y(n_85)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_45),
.Y(n_86)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_86),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_87),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_20),
.Y(n_88)
);

INVx5_ASAP7_75t_SL g130 ( 
.A(n_88),
.Y(n_130)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_89),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_90),
.Y(n_148)
);

INVx13_ASAP7_75t_L g91 ( 
.A(n_20),
.Y(n_91)
);

CKINVDCx6p67_ASAP7_75t_R g117 ( 
.A(n_91),
.Y(n_117)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_93),
.Y(n_160)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_27),
.Y(n_94)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_94),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_20),
.B(n_4),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_96),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_30),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_97),
.A2(n_47),
.B1(n_44),
.B2(n_43),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_33),
.Y(n_99)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_100),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_51),
.Y(n_101)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_101),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_35),
.B(n_4),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_102),
.B(n_53),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_103),
.Y(n_152)
);

BUFx12_ASAP7_75t_L g104 ( 
.A(n_17),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_104),
.B(n_107),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_41),
.B(n_4),
.Y(n_105)
);

INVx4_ASAP7_75t_SL g106 ( 
.A(n_17),
.Y(n_106)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_106),
.Y(n_162)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_19),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_105),
.B(n_49),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_108),
.B(n_116),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_57),
.B(n_49),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_106),
.A2(n_34),
.B1(n_30),
.B2(n_31),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_123),
.A2(n_76),
.B1(n_98),
.B2(n_79),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_56),
.A2(n_34),
.B1(n_30),
.B2(n_31),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_133),
.A2(n_82),
.B1(n_103),
.B2(n_101),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_135),
.A2(n_143),
.B1(n_36),
.B2(n_42),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_47),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_137),
.B(n_141),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_83),
.B(n_41),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_61),
.A2(n_34),
.B1(n_38),
.B2(n_39),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_95),
.B(n_44),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_146),
.B(n_150),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_88),
.B(n_43),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_154),
.B(n_48),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_77),
.B(n_53),
.Y(n_155)
);

AND2x2_ASAP7_75t_SL g182 ( 
.A(n_155),
.B(n_164),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_64),
.B(n_37),
.Y(n_164)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_89),
.Y(n_167)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_167),
.Y(n_177)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_170),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_163),
.A2(n_42),
.B1(n_36),
.B2(n_33),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_171),
.B(n_184),
.Y(n_227)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_110),
.Y(n_172)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_172),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_117),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_174),
.B(n_186),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_138),
.Y(n_176)
);

INVx5_ASAP7_75t_L g243 ( 
.A(n_176),
.Y(n_243)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_169),
.Y(n_178)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_178),
.Y(n_255)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_161),
.Y(n_179)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_179),
.Y(n_235)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_114),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_180),
.Y(n_247)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_139),
.Y(n_181)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_181),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_185),
.A2(n_195),
.B1(n_210),
.B2(n_212),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_117),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_126),
.A2(n_81),
.B1(n_93),
.B2(n_67),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_187),
.B(n_86),
.Y(n_236)
);

BUFx4f_ASAP7_75t_L g188 ( 
.A(n_117),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_188),
.Y(n_220)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_118),
.Y(n_189)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_189),
.Y(n_223)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_159),
.Y(n_190)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_190),
.Y(n_225)
);

INVxp67_ASAP7_75t_SL g191 ( 
.A(n_112),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_191),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_163),
.A2(n_37),
.B(n_48),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_192),
.B(n_219),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_132),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_193),
.Y(n_231)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_159),
.Y(n_194)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_194),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_112),
.A2(n_94),
.B1(n_25),
.B2(n_21),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_138),
.Y(n_196)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_196),
.Y(n_250)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_145),
.Y(n_197)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_197),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_142),
.Y(n_198)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_198),
.Y(n_254)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_121),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_199),
.B(n_200),
.Y(n_233)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_148),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_160),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_201),
.B(n_202),
.Y(n_234)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_113),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_119),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_203),
.B(n_204),
.Y(n_237)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_122),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_130),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_205),
.B(n_207),
.Y(n_242)
);

NOR2x1_ASAP7_75t_L g256 ( 
.A(n_206),
.B(n_215),
.Y(n_256)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_113),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_208),
.B(n_209),
.Y(n_248)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_136),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_142),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_165),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_213),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_158),
.A2(n_149),
.B1(n_109),
.B2(n_165),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_127),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_118),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_214),
.A2(n_166),
.B1(n_140),
.B2(n_153),
.Y(n_229)
);

BUFx12f_ASAP7_75t_L g215 ( 
.A(n_129),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_124),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_217),
.Y(n_221)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_128),
.Y(n_217)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_127),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_109),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_115),
.B(n_104),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_222),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_229),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_182),
.B(n_125),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_232),
.B(n_239),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_236),
.A2(n_134),
.B1(n_120),
.B2(n_129),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_182),
.B(n_147),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_189),
.A2(n_134),
.B1(n_166),
.B2(n_152),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_240),
.A2(n_212),
.B1(n_195),
.B2(n_185),
.Y(n_258)
);

OR2x4_ASAP7_75t_L g241 ( 
.A(n_191),
.B(n_162),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_241),
.B(n_151),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_183),
.B(n_157),
.C(n_156),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_227),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_177),
.B(n_173),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_249),
.B(n_252),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_175),
.B(n_111),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g314 ( 
.A1(n_258),
.A2(n_215),
.B1(n_243),
.B2(n_226),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_221),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_260),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_261),
.A2(n_223),
.B1(n_247),
.B2(n_231),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_256),
.A2(n_90),
.B1(n_87),
.B2(n_133),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_262),
.A2(n_280),
.B1(n_220),
.B2(n_223),
.Y(n_292)
);

OAI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_256),
.A2(n_214),
.B1(n_193),
.B2(n_209),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_263),
.A2(n_271),
.B1(n_272),
.B2(n_274),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_242),
.B(n_174),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_264),
.B(n_266),
.Y(n_290)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_221),
.Y(n_265)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_265),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_232),
.B(n_170),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_233),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_267),
.B(n_276),
.Y(n_298)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_233),
.Y(n_268)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_268),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_269),
.B(n_285),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_238),
.A2(n_123),
.B1(n_140),
.B2(n_153),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_236),
.A2(n_157),
.B1(n_136),
.B2(n_156),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_242),
.B(n_168),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_273),
.B(n_226),
.Y(n_297)
);

OAI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_256),
.A2(n_208),
.B1(n_202),
.B2(n_179),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_227),
.A2(n_188),
.B(n_218),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_275),
.A2(n_277),
.B(n_248),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_249),
.B(n_130),
.Y(n_276)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_234),
.Y(n_279)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_279),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_227),
.A2(n_151),
.B1(n_210),
.B2(n_198),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_239),
.B(n_188),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_283),
.Y(n_302)
);

O2A1O1Ixp33_ASAP7_75t_L g283 ( 
.A1(n_241),
.A2(n_91),
.B(n_158),
.C(n_213),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_244),
.B(n_21),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_284),
.B(n_286),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_252),
.B(n_25),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_244),
.B(n_21),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_243),
.Y(n_287)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_287),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_253),
.B(n_52),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_288),
.B(n_289),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_253),
.B(n_246),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_292),
.A2(n_303),
.B1(n_308),
.B2(n_312),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_222),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_293),
.B(n_259),
.C(n_278),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_289),
.B(n_248),
.C(n_245),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_295),
.B(n_305),
.C(n_313),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_297),
.B(n_306),
.Y(n_326)
);

CKINVDCx14_ASAP7_75t_R g336 ( 
.A(n_300),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_277),
.A2(n_224),
.B(n_237),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_304),
.A2(n_302),
.B(n_283),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_259),
.C(n_278),
.Y(n_305)
);

INVxp33_ASAP7_75t_L g306 ( 
.A(n_264),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_281),
.A2(n_247),
.B1(n_234),
.B2(n_254),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_265),
.Y(n_310)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_310),
.Y(n_319)
);

BUFx24_ASAP7_75t_SL g311 ( 
.A(n_273),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_311),
.Y(n_335)
);

OAI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_268),
.A2(n_279),
.B1(n_281),
.B2(n_274),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_285),
.B(n_245),
.C(n_225),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_314),
.A2(n_271),
.B(n_277),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_262),
.A2(n_176),
.B1(n_196),
.B2(n_237),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_316),
.A2(n_282),
.B1(n_266),
.B2(n_288),
.Y(n_332)
);

INVx2_ASAP7_75t_SL g317 ( 
.A(n_287),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_317),
.B(n_307),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_300),
.A2(n_275),
.B(n_277),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_320),
.A2(n_342),
.B(n_346),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_291),
.B(n_260),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_322),
.B(n_328),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_323),
.A2(n_292),
.B1(n_296),
.B2(n_308),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_SL g356 ( 
.A(n_325),
.B(n_296),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_327),
.B(n_330),
.C(n_334),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_291),
.B(n_267),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_309),
.A2(n_258),
.B1(n_270),
.B2(n_272),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_329),
.A2(n_343),
.B(n_250),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_293),
.B(n_286),
.C(n_284),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_309),
.Y(n_331)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_331),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_332),
.A2(n_254),
.B1(n_250),
.B2(n_225),
.Y(n_359)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_301),
.Y(n_333)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_333),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_294),
.B(n_276),
.C(n_280),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_298),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_337),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_338),
.Y(n_370)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_301),
.Y(n_339)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_339),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_298),
.B(n_283),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_340),
.B(n_345),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_297),
.B(n_231),
.Y(n_341)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_341),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_302),
.A2(n_251),
.B(n_230),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_304),
.A2(n_251),
.B(n_261),
.Y(n_343)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_307),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_344),
.B(n_215),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_290),
.B(n_230),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_317),
.A2(n_287),
.B1(n_131),
.B2(n_197),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_290),
.B(n_310),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_347),
.B(n_52),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_321),
.B(n_294),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_348),
.B(n_353),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_335),
.B(n_318),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_352),
.B(n_362),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_321),
.B(n_315),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_354),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_321),
.B(n_295),
.C(n_315),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_355),
.B(n_360),
.C(n_368),
.Y(n_386)
);

CKINVDCx14_ASAP7_75t_R g387 ( 
.A(n_356),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_337),
.A2(n_299),
.B1(n_317),
.B2(n_313),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_357),
.B(n_358),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_322),
.A2(n_299),
.B1(n_305),
.B2(n_318),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_359),
.A2(n_366),
.B1(n_333),
.B2(n_331),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_327),
.B(n_235),
.C(n_228),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_330),
.B(n_235),
.Y(n_363)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_363),
.B(n_376),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_336),
.A2(n_255),
.B1(n_228),
.B2(n_257),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_334),
.B(n_255),
.C(n_257),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_369),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_372),
.B(n_341),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g373 ( 
.A(n_328),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_373),
.B(n_374),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_336),
.B(n_131),
.C(n_52),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_347),
.B(n_21),
.Y(n_376)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_375),
.Y(n_378)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_378),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_367),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_380),
.B(n_383),
.Y(n_407)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_364),
.Y(n_381)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_381),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_382),
.A2(n_396),
.B1(n_329),
.B2(n_332),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_364),
.Y(n_383)
);

INVx13_ASAP7_75t_L g384 ( 
.A(n_366),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_384),
.B(n_391),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_365),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_385),
.B(n_389),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_372),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_351),
.Y(n_390)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_390),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_350),
.A2(n_320),
.B(n_340),
.Y(n_391)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_361),
.Y(n_393)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_393),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_394),
.B(n_395),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_370),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_371),
.Y(n_396)
);

A2O1A1Ixp33_ASAP7_75t_L g398 ( 
.A1(n_362),
.A2(n_325),
.B(n_326),
.C(n_342),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_398),
.B(n_400),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_359),
.B(n_326),
.Y(n_400)
);

OR2x6_ASAP7_75t_L g402 ( 
.A(n_350),
.B(n_323),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_402),
.A2(n_354),
.B1(n_324),
.B2(n_346),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_358),
.B(n_345),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_403),
.B(n_376),
.Y(n_404)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_404),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_405),
.A2(n_391),
.B(n_402),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_386),
.B(n_348),
.C(n_353),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_409),
.B(n_410),
.C(n_411),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_386),
.B(n_349),
.C(n_355),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_377),
.B(n_349),
.C(n_363),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_392),
.B(n_368),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_413),
.B(n_400),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_377),
.B(n_360),
.C(n_357),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_415),
.B(n_424),
.C(n_401),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_399),
.A2(n_356),
.B1(n_324),
.B2(n_319),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_417),
.A2(n_419),
.B1(n_382),
.B2(n_395),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_399),
.A2(n_319),
.B1(n_339),
.B2(n_343),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_392),
.B(n_374),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_420),
.B(n_425),
.Y(n_437)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_421),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_388),
.B(n_338),
.C(n_344),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_388),
.B(n_344),
.Y(n_425)
);

XOR2x2_ASAP7_75t_L g426 ( 
.A(n_425),
.B(n_402),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_SL g452 ( 
.A(n_426),
.B(n_428),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_427),
.A2(n_426),
.B1(n_439),
.B2(n_428),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_407),
.A2(n_380),
.B1(n_397),
.B2(n_402),
.Y(n_429)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_429),
.Y(n_444)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_432),
.B(n_439),
.Y(n_453)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_418),
.Y(n_434)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_434),
.Y(n_448)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_414),
.Y(n_435)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_435),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_412),
.B(n_379),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_436),
.B(n_442),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_405),
.A2(n_402),
.B1(n_387),
.B2(n_383),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_438),
.A2(n_419),
.B1(n_408),
.B2(n_417),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_420),
.B(n_402),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_440),
.B(n_396),
.C(n_393),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_409),
.B(n_398),
.C(n_378),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_441),
.B(n_443),
.C(n_415),
.Y(n_446)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_416),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_410),
.B(n_389),
.C(n_394),
.Y(n_443)
);

OR2x2_ASAP7_75t_L g445 ( 
.A(n_438),
.B(n_381),
.Y(n_445)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_445),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_446),
.B(n_449),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_441),
.A2(n_406),
.B(n_412),
.Y(n_447)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_447),
.A2(n_457),
.B(n_458),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_451),
.B(n_7),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_431),
.A2(n_379),
.B1(n_422),
.B2(n_424),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_454),
.A2(n_437),
.B1(n_390),
.B2(n_9),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_433),
.B(n_411),
.C(n_413),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_455),
.B(n_437),
.C(n_432),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_443),
.A2(n_430),
.B(n_440),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_433),
.A2(n_384),
.B(n_423),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_459),
.B(n_452),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_460),
.B(n_467),
.C(n_468),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_461),
.B(n_463),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_450),
.B(n_39),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_462),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_446),
.B(n_39),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_444),
.A2(n_38),
.B1(n_31),
.B2(n_52),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_465),
.A2(n_473),
.B1(n_40),
.B2(n_10),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_455),
.B(n_51),
.C(n_38),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_453),
.B(n_25),
.C(n_21),
.Y(n_468)
);

XOR2x2_ASAP7_75t_L g469 ( 
.A(n_453),
.B(n_451),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_469),
.B(n_471),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_472),
.B(n_8),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_457),
.B(n_25),
.Y(n_473)
);

OAI321xp33_ASAP7_75t_L g474 ( 
.A1(n_466),
.A2(n_448),
.A3(n_456),
.B1(n_445),
.B2(n_449),
.C(n_458),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_474),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_SL g477 ( 
.A1(n_464),
.A2(n_470),
.B(n_460),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g487 ( 
.A1(n_477),
.A2(n_480),
.B(n_8),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_469),
.B(n_459),
.C(n_452),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_479),
.B(n_483),
.Y(n_485)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_467),
.A2(n_40),
.B(n_25),
.Y(n_480)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_482),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_472),
.B(n_40),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_484),
.B(n_476),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_481),
.A2(n_468),
.B1(n_10),
.B2(n_11),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_486),
.B(n_487),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_SL g488 ( 
.A(n_479),
.B(n_476),
.Y(n_488)
);

O2A1O1Ixp33_ASAP7_75t_SL g493 ( 
.A1(n_488),
.A2(n_475),
.B(n_484),
.C(n_483),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_489),
.A2(n_475),
.B(n_12),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_SL g492 ( 
.A(n_490),
.B(n_478),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_492),
.B(n_493),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_495),
.B(n_10),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_494),
.B(n_485),
.C(n_491),
.Y(n_496)
);

OAI21xp33_ASAP7_75t_L g500 ( 
.A1(n_496),
.A2(n_497),
.B(n_14),
.Y(n_500)
);

A2O1A1Ixp33_ASAP7_75t_L g499 ( 
.A1(n_498),
.A2(n_10),
.B(n_12),
.C(n_13),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_499),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_501),
.Y(n_502)
);

AOI21x1_ASAP7_75t_L g503 ( 
.A1(n_502),
.A2(n_500),
.B(n_14),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_R g504 ( 
.A(n_503),
.B(n_14),
.C(n_15),
.Y(n_504)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_504),
.B(n_14),
.Y(n_505)
);


endmodule