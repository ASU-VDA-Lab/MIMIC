module fake_jpeg_14004_n_263 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_263);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_263;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_57;
wire n_21;
wire n_187;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_6),
.B(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx2_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_10),
.B(n_0),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_47),
.Y(n_121)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_50),
.B(n_57),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

INVxp67_ASAP7_75t_SL g55 ( 
.A(n_31),
.Y(n_55)
);

CKINVDCx6p67_ASAP7_75t_R g106 ( 
.A(n_55),
.Y(n_106)
);

BUFx10_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_19),
.B(n_15),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_58),
.B(n_64),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

BUFx16f_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_60),
.B(n_61),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_31),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_19),
.B(n_7),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_63),
.B(n_79),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_15),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

CKINVDCx5p33_ASAP7_75t_R g66 ( 
.A(n_36),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_66),
.B(n_68),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_67),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_42),
.B(n_7),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_69),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_43),
.A2(n_4),
.B1(n_5),
.B2(n_8),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_71),
.A2(n_85),
.B1(n_40),
.B2(n_32),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_73),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_20),
.B(n_4),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_74),
.B(n_76),
.Y(n_120)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_78),
.B(n_86),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_21),
.B(n_14),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_25),
.B(n_5),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_80),
.B(n_83),
.Y(n_111)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_81),
.B(n_89),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_25),
.B(n_5),
.Y(n_83)
);

BUFx10_ASAP7_75t_L g84 ( 
.A(n_17),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_84),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_23),
.A2(n_1),
.B1(n_2),
.B2(n_12),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_21),
.B(n_14),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_87),
.B(n_30),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_90),
.Y(n_127)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_17),
.Y(n_89)
);

BUFx4f_ASAP7_75t_SL g90 ( 
.A(n_17),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_55),
.A2(n_23),
.B1(n_37),
.B2(n_59),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_95),
.A2(n_108),
.B1(n_117),
.B2(n_118),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_63),
.B(n_29),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_100),
.B(n_133),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_86),
.A2(n_23),
.B1(n_46),
.B2(n_33),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_56),
.A2(n_29),
.B1(n_35),
.B2(n_34),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_56),
.A2(n_28),
.B1(n_35),
.B2(n_34),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_77),
.A2(n_45),
.B1(n_33),
.B2(n_28),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_122),
.A2(n_125),
.B1(n_131),
.B2(n_132),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_51),
.A2(n_40),
.B1(n_16),
.B2(n_32),
.Y(n_125)
);

NAND3xp33_ASAP7_75t_L g141 ( 
.A(n_128),
.B(n_1),
.C(n_2),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_87),
.B(n_83),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_129),
.B(n_130),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_80),
.B(n_30),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_69),
.A2(n_26),
.B1(n_45),
.B2(n_27),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_74),
.B(n_16),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_90),
.B(n_22),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_134),
.B(n_84),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_52),
.A2(n_22),
.B1(n_27),
.B2(n_1),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_135),
.A2(n_112),
.B1(n_123),
.B2(n_101),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_111),
.A2(n_85),
.B1(n_70),
.B2(n_72),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_137),
.Y(n_199)
);

OAI32xp33_ASAP7_75t_L g138 ( 
.A1(n_98),
.A2(n_84),
.A3(n_82),
.B1(n_60),
.B2(n_17),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_138),
.B(n_141),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_139),
.B(n_144),
.Y(n_190)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_17),
.C(n_92),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_143),
.B(n_151),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_102),
.B(n_120),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_94),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_94),
.Y(n_146)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_146),
.Y(n_180)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_132),
.A2(n_104),
.B1(n_99),
.B2(n_109),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_148),
.A2(n_172),
.B1(n_137),
.B2(n_158),
.Y(n_194)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_121),
.A2(n_114),
.B1(n_113),
.B2(n_119),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_149),
.A2(n_152),
.B1(n_164),
.B2(n_169),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_96),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_150),
.B(n_154),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_124),
.B(n_110),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_104),
.A2(n_98),
.B1(n_111),
.B2(n_99),
.Y(n_152)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_91),
.Y(n_153)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_153),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_100),
.B(n_128),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_110),
.Y(n_155)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_133),
.A2(n_136),
.B(n_107),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_156),
.B(n_167),
.Y(n_193)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_115),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_105),
.B(n_127),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_163),
.Y(n_197)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_91),
.Y(n_161)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_161),
.Y(n_198)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_106),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_162),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_107),
.B(n_106),
.Y(n_163)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_93),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_168),
.Y(n_176)
);

OAI32xp33_ASAP7_75t_L g166 ( 
.A1(n_121),
.A2(n_101),
.A3(n_106),
.B1(n_119),
.B2(n_113),
.Y(n_166)
);

NOR2x1_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_175),
.Y(n_184)
);

O2A1O1Ixp33_ASAP7_75t_L g167 ( 
.A1(n_106),
.A2(n_97),
.B(n_123),
.C(n_115),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_114),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_109),
.A2(n_119),
.B1(n_93),
.B2(n_113),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_126),
.B(n_93),
.C(n_97),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_171),
.B(n_174),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_126),
.A2(n_71),
.B1(n_132),
.B2(n_104),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_103),
.B(n_129),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_140),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_103),
.B(n_102),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_116),
.B(n_92),
.C(n_110),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g177 ( 
.A1(n_152),
.A2(n_159),
.B1(n_148),
.B2(n_151),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_177),
.A2(n_166),
.B1(n_171),
.B2(n_153),
.Y(n_203)
);

OAI21xp33_ASAP7_75t_L g206 ( 
.A1(n_179),
.A2(n_167),
.B(n_162),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_175),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_181),
.B(n_182),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_140),
.B(n_151),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_173),
.B(n_143),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_192),
.Y(n_204)
);

NOR2x1_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_138),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_189),
.A2(n_193),
.B(n_185),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_155),
.B(n_170),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_194),
.A2(n_199),
.B1(n_178),
.B2(n_189),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_146),
.B(n_147),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_176),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_190),
.B(n_150),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_201),
.B(n_202),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_190),
.B(n_168),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_203),
.A2(n_209),
.B1(n_194),
.B2(n_200),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_183),
.B(n_145),
.C(n_157),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_205),
.B(n_215),
.Y(n_227)
);

OAI21xp33_ASAP7_75t_L g231 ( 
.A1(n_206),
.A2(n_211),
.B(n_214),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_142),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_208),
.B(n_186),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_199),
.A2(n_165),
.B1(n_161),
.B2(n_169),
.Y(n_209)
);

MAJx2_ASAP7_75t_L g210 ( 
.A(n_181),
.B(n_179),
.C(n_182),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_210),
.B(n_217),
.Y(n_220)
);

AND2x4_ASAP7_75t_L g211 ( 
.A(n_196),
.B(n_184),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_212),
.A2(n_193),
.B1(n_200),
.B2(n_184),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_213),
.A2(n_216),
.B(n_184),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g214 ( 
.A(n_178),
.B(n_191),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_178),
.B(n_191),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_180),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_192),
.B(n_197),
.C(n_193),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_195),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_219),
.B(n_211),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_222),
.B(n_228),
.Y(n_240)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_223),
.B(n_225),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_224),
.A2(n_228),
.B1(n_219),
.B2(n_211),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_209),
.A2(n_198),
.B1(n_187),
.B2(n_186),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_217),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_188),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_212),
.A2(n_207),
.B1(n_203),
.B2(n_218),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_229),
.B(n_204),
.Y(n_232)
);

OAI21xp33_ASAP7_75t_SL g230 ( 
.A1(n_213),
.A2(n_189),
.B(n_185),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g236 ( 
.A(n_230),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_232),
.A2(n_220),
.B1(n_227),
.B2(n_205),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_234),
.B(n_238),
.Y(n_248)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_223),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_239),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_237),
.A2(n_224),
.B(n_216),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_226),
.B(n_215),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_204),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_241),
.A2(n_211),
.B1(n_216),
.B2(n_210),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_246),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_232),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_233),
.A2(n_231),
.B(n_229),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_245),
.B(n_247),
.Y(n_249)
);

O2A1O1Ixp33_ASAP7_75t_SL g247 ( 
.A1(n_237),
.A2(n_227),
.B(n_214),
.C(n_176),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_250),
.B(n_251),
.Y(n_255)
);

OAI221xp5_ASAP7_75t_L g251 ( 
.A1(n_242),
.A2(n_235),
.B1(n_238),
.B2(n_237),
.C(n_221),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_244),
.B(n_195),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_252),
.Y(n_254)
);

XOR2x1_ASAP7_75t_SL g256 ( 
.A(n_249),
.B(n_245),
.Y(n_256)
);

AOI322xp5_ASAP7_75t_L g258 ( 
.A1(n_256),
.A2(n_257),
.A3(n_241),
.B1(n_248),
.B2(n_243),
.C1(n_247),
.C2(n_246),
.Y(n_258)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_248),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_258),
.B(n_259),
.Y(n_261)
);

AOI322xp5_ASAP7_75t_L g259 ( 
.A1(n_254),
.A2(n_233),
.A3(n_240),
.B1(n_236),
.B2(n_247),
.C1(n_253),
.C2(n_198),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_258),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_260),
.B(n_255),
.Y(n_262)
);

AOI221xp5_ASAP7_75t_L g263 ( 
.A1(n_262),
.A2(n_261),
.B1(n_253),
.B2(n_240),
.C(n_187),
.Y(n_263)
);


endmodule