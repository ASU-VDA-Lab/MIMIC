module fake_jpeg_17287_n_349 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_349);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_349;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_12),
.B(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_4),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx24_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_6),
.B(n_3),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_13),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_42),
.Y(n_101)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_43),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_15),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_46),
.B(n_54),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_30),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_47),
.A2(n_58),
.B1(n_69),
.B2(n_34),
.Y(n_124)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_50),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_29),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_56),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_52),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_14),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_27),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_27),
.B(n_0),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_57),
.B(n_61),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_30),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_21),
.Y(n_59)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_59),
.Y(n_108)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_62),
.B(n_64),
.Y(n_97)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_18),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_65),
.Y(n_117)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_67),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_68),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_37),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_69)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

INVx4_ASAP7_75t_SL g72 ( 
.A(n_38),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_72),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_36),
.B(n_3),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_74),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_36),
.B(n_4),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_35),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_72),
.A2(n_40),
.B1(n_42),
.B2(n_61),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_76),
.A2(n_80),
.B1(n_84),
.B2(n_92),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_48),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_79),
.B(n_82),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_43),
.A2(n_32),
.B1(n_24),
.B2(n_19),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_24),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_72),
.A2(n_40),
.B1(n_32),
.B2(n_31),
.Y(n_84)
);

NAND3xp33_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_28),
.C(n_31),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g145 ( 
.A1(n_85),
.A2(n_111),
.B(n_8),
.C(n_9),
.Y(n_145)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_65),
.A2(n_38),
.B1(n_28),
.B2(n_34),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_86),
.A2(n_124),
.B1(n_127),
.B2(n_8),
.Y(n_144)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_88),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_70),
.A2(n_40),
.B1(n_49),
.B2(n_60),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_22),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_96),
.B(n_103),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_63),
.A2(n_38),
.B1(n_16),
.B2(n_20),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_98),
.A2(n_34),
.B1(n_25),
.B2(n_35),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_99),
.B(n_110),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_55),
.B(n_22),
.Y(n_103)
);

INVx13_ASAP7_75t_L g110 ( 
.A(n_51),
.Y(n_110)
);

HAxp5_ASAP7_75t_SL g111 ( 
.A(n_47),
.B(n_22),
.CON(n_111),
.SN(n_111)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_66),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g153 ( 
.A(n_112),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_41),
.B(n_35),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_114),
.B(n_115),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_62),
.B(n_35),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_50),
.Y(n_116)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_64),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_118),
.B(n_128),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_44),
.B(n_22),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_122),
.B(n_126),
.Y(n_164)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_50),
.Y(n_123)
);

BUFx2_ASAP7_75t_SL g173 ( 
.A(n_123),
.Y(n_173)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_45),
.Y(n_125)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_125),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_52),
.B(n_22),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_53),
.A2(n_20),
.B1(n_33),
.B2(n_38),
.Y(n_127)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_59),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_93),
.B(n_71),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_131),
.B(n_132),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_68),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_67),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_133),
.B(n_142),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_97),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_134),
.B(n_137),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_86),
.B(n_4),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_135),
.A2(n_47),
.B(n_156),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_101),
.A2(n_20),
.B1(n_34),
.B2(n_25),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_136),
.A2(n_158),
.B1(n_154),
.B2(n_137),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g137 ( 
.A(n_77),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_138),
.A2(n_143),
.B1(n_155),
.B2(n_112),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_77),
.Y(n_139)
);

INVx11_ASAP7_75t_L g212 ( 
.A(n_139),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_91),
.Y(n_140)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_140),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_111),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_141),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_95),
.B(n_106),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_98),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_144),
.A2(n_156),
.B1(n_140),
.B2(n_159),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_145),
.Y(n_194)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_113),
.Y(n_146)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_146),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_76),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_147),
.B(n_161),
.Y(n_189)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_113),
.Y(n_150)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_150),
.Y(n_218)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_80),
.Y(n_151)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_151),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_84),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_81),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_101),
.A2(n_10),
.B1(n_125),
.B2(n_78),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_91),
.Y(n_159)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_159),
.Y(n_183)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_117),
.Y(n_161)
);

AOI32xp33_ASAP7_75t_L g162 ( 
.A1(n_81),
.A2(n_78),
.A3(n_88),
.B1(n_83),
.B2(n_118),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_145),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_109),
.B(n_110),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_169),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_86),
.B(n_92),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_165),
.B(n_116),
.C(n_129),
.Y(n_185)
);

A2O1A1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_90),
.A2(n_105),
.B(n_104),
.C(n_123),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_166),
.B(n_168),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_100),
.B(n_128),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_167),
.B(n_171),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_87),
.B(n_94),
.Y(n_168)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_102),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_105),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_172),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_100),
.B(n_104),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_119),
.Y(n_172)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_108),
.Y(n_175)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_175),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_120),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_177),
.Y(n_197)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_121),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_89),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_179),
.Y(n_199)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_119),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_144),
.A2(n_87),
.B1(n_94),
.B2(n_89),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_181),
.A2(n_190),
.B1(n_208),
.B2(n_180),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_182),
.A2(n_195),
.B1(n_203),
.B2(n_208),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_185),
.B(n_193),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_188),
.B(n_201),
.Y(n_234)
);

AO22x1_ASAP7_75t_SL g190 ( 
.A1(n_165),
.A2(n_135),
.B1(n_151),
.B2(n_147),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_132),
.B(n_133),
.C(n_148),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_135),
.A2(n_131),
.B1(n_164),
.B2(n_142),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_167),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_204),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_200),
.Y(n_224)
);

NOR2x1_ASAP7_75t_L g201 ( 
.A(n_141),
.B(n_166),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_201),
.A2(n_207),
.B(n_194),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_134),
.A2(n_171),
.B1(n_146),
.B2(n_161),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_160),
.Y(n_204)
);

INVxp33_ASAP7_75t_L g205 ( 
.A(n_173),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_205),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_156),
.B(n_130),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_206),
.A2(n_219),
.B(n_220),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_154),
.A2(n_150),
.B1(n_177),
.B2(n_169),
.Y(n_208)
);

OAI32xp33_ASAP7_75t_L g209 ( 
.A1(n_152),
.A2(n_157),
.A3(n_149),
.B1(n_130),
.B2(n_174),
.Y(n_209)
);

A2O1A1O1Ixp25_ASAP7_75t_L g228 ( 
.A1(n_209),
.A2(n_201),
.B(n_195),
.C(n_206),
.D(n_211),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_153),
.B(n_176),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_210),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_174),
.B(n_153),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_185),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_175),
.B(n_179),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_214),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_139),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_215),
.B(n_212),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_216),
.A2(n_221),
.B1(n_219),
.B2(n_202),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_132),
.A2(n_133),
.B(n_151),
.Y(n_219)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_186),
.Y(n_226)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_226),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_228),
.A2(n_234),
.B(n_239),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_198),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_229),
.B(n_243),
.Y(n_261)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_186),
.Y(n_230)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_230),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_196),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_240),
.Y(n_259)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_218),
.Y(n_232)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_232),
.Y(n_279)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_235),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_236),
.B(n_225),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_202),
.B(n_194),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_237),
.B(n_240),
.Y(n_268)
);

OAI22x1_ASAP7_75t_SL g238 ( 
.A1(n_190),
.A2(n_181),
.B1(n_216),
.B2(n_206),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_238),
.A2(n_254),
.B1(n_251),
.B2(n_222),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_211),
.B(n_217),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_241),
.A2(n_246),
.B1(n_253),
.B2(n_255),
.Y(n_264)
);

A2O1A1Ixp33_ASAP7_75t_L g242 ( 
.A1(n_207),
.A2(n_190),
.B(n_220),
.C(n_188),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_249),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_198),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_221),
.Y(n_244)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_244),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_189),
.A2(n_213),
.B(n_190),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_245),
.A2(n_252),
.B(n_215),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_184),
.A2(n_193),
.B1(n_182),
.B2(n_204),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_199),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_250),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_184),
.B(n_203),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_218),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_209),
.A2(n_191),
.B(n_187),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_197),
.A2(n_180),
.B1(n_192),
.B2(n_183),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_183),
.A2(n_185),
.B1(n_221),
.B2(n_144),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_229),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_257),
.B(n_258),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_243),
.Y(n_258)
);

AOI221xp5_ASAP7_75t_L g305 ( 
.A1(n_262),
.A2(n_273),
.B1(n_256),
.B2(n_264),
.C(n_260),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_231),
.B(n_212),
.Y(n_265)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_265),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_233),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_266),
.B(n_270),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_268),
.B(n_277),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_244),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_237),
.B(n_249),
.Y(n_271)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_271),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_272),
.A2(n_281),
.B1(n_262),
.B2(n_265),
.Y(n_299)
);

AOI322xp5_ASAP7_75t_L g273 ( 
.A1(n_234),
.A2(n_238),
.A3(n_252),
.B1(n_239),
.B2(n_242),
.C1(n_248),
.C2(n_228),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_248),
.A2(n_224),
.B(n_234),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_274),
.A2(n_280),
.B(n_260),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_225),
.B(n_236),
.C(n_245),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_276),
.C(n_278),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_222),
.B(n_251),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_246),
.B(n_255),
.C(n_254),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_223),
.A2(n_227),
.B1(n_253),
.B2(n_233),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_227),
.B(n_223),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_283),
.B(n_270),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_276),
.B(n_247),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_284),
.B(n_275),
.C(n_256),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_277),
.A2(n_250),
.B1(n_235),
.B2(n_232),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_286),
.A2(n_292),
.B1(n_272),
.B2(n_258),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_263),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_287),
.B(n_288),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_261),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_267),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_289),
.B(n_298),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_264),
.A2(n_226),
.B1(n_230),
.B2(n_278),
.Y(n_292)
);

NAND3xp33_ASAP7_75t_L g293 ( 
.A(n_261),
.B(n_267),
.C(n_257),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_293),
.B(n_304),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_274),
.A2(n_266),
.B1(n_280),
.B2(n_258),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_294),
.B(n_269),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_297),
.B(n_305),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_263),
.Y(n_298)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_282),
.Y(n_301)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_301),
.Y(n_318)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_282),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_303),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_268),
.B(n_259),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_279),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_257),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_308),
.B(n_319),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_309),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_291),
.B(n_271),
.C(n_259),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_316),
.C(n_317),
.Y(n_323)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_315),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_291),
.B(n_273),
.C(n_283),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_284),
.B(n_281),
.C(n_279),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_SL g319 ( 
.A(n_297),
.B(n_270),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_292),
.B(n_269),
.C(n_266),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_322),
.C(n_288),
.Y(n_328)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_321),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_295),
.B(n_299),
.C(n_294),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_320),
.A2(n_290),
.B1(n_286),
.B2(n_300),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_327),
.A2(n_330),
.B1(n_324),
.B2(n_328),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_328),
.B(n_327),
.C(n_334),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_314),
.B(n_285),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_329),
.B(n_331),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_311),
.B(n_296),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_313),
.B(n_296),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_333),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_312),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_321),
.A2(n_290),
.B1(n_287),
.B2(n_298),
.Y(n_334)
);

OA21x2_ASAP7_75t_SL g335 ( 
.A1(n_307),
.A2(n_301),
.B(n_302),
.Y(n_335)
);

NAND4xp25_ASAP7_75t_SL g336 ( 
.A(n_335),
.B(n_306),
.C(n_318),
.D(n_319),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_338),
.B(n_330),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_323),
.B(n_326),
.C(n_331),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_337),
.A2(n_325),
.B(n_324),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_343),
.A2(n_341),
.B(n_336),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_344),
.A2(n_341),
.B(n_342),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_344),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_346),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_347),
.B(n_339),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_348),
.B(n_340),
.Y(n_349)
);


endmodule