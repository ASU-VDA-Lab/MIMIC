module real_aes_3335_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_577;
wire n_580;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_560;
wire n_260;
wire n_594;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_92;
wire n_519;
wire n_564;
wire n_573;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_570;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_547;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_93;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_85;
wire n_605;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_87;
wire n_171;
wire n_78;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_622;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_589;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_597;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_601;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_91;
NAND2xp5_ASAP7_75t_L g301 ( .A(n_0), .B(n_281), .Y(n_301) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_1), .Y(n_317) );
O2A1O1Ixp33_ASAP7_75t_SL g353 ( .A1(n_2), .A2(n_225), .B(n_354), .C(n_355), .Y(n_353) );
OAI22xp33_ASAP7_75t_L g306 ( .A1(n_3), .A2(n_64), .B1(n_223), .B2(n_253), .Y(n_306) );
INVx1_ASAP7_75t_L g157 ( .A(n_4), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g332 ( .A(n_5), .Y(n_332) );
OAI22xp5_ASAP7_75t_L g250 ( .A1(n_6), .A2(n_54), .B1(n_251), .B2(n_253), .Y(n_250) );
CKINVDCx5p33_ASAP7_75t_R g272 ( .A(n_7), .Y(n_272) );
INVx1_ASAP7_75t_L g107 ( .A(n_8), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g152 ( .A(n_8), .B(n_56), .Y(n_152) );
INVxp67_ASAP7_75t_L g174 ( .A(n_8), .Y(n_174) );
HB1xp67_ASAP7_75t_L g185 ( .A(n_9), .Y(n_185) );
AOI22xp5_ASAP7_75t_L g248 ( .A1(n_10), .A2(n_45), .B1(n_223), .B2(n_249), .Y(n_248) );
OA21x2_ASAP7_75t_L g238 ( .A1(n_11), .A2(n_53), .B(n_239), .Y(n_238) );
OA21x2_ASAP7_75t_L g243 ( .A1(n_11), .A2(n_53), .B(n_239), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g103 ( .A(n_12), .B(n_92), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g327 ( .A(n_13), .Y(n_327) );
BUFx3_ASAP7_75t_L g195 ( .A(n_14), .Y(n_195) );
O2A1O1Ixp33_ASAP7_75t_L g359 ( .A1(n_15), .A2(n_307), .B(n_360), .C(n_361), .Y(n_359) );
INVx1_ASAP7_75t_L g164 ( .A(n_16), .Y(n_164) );
OAI22xp33_ASAP7_75t_SL g304 ( .A1(n_17), .A2(n_31), .B1(n_223), .B2(n_271), .Y(n_304) );
AOI22xp33_ASAP7_75t_L g291 ( .A1(n_18), .A2(n_23), .B1(n_271), .B2(n_276), .Y(n_291) );
BUFx6f_ASAP7_75t_L g92 ( .A(n_19), .Y(n_92) );
O2A1O1Ixp5_ASAP7_75t_L g218 ( .A1(n_20), .A2(n_219), .B(n_222), .C(n_225), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_21), .B(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g93 ( .A(n_22), .Y(n_93) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_22), .B(n_55), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_24), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_25), .B(n_297), .Y(n_296) );
AOI22xp33_ASAP7_75t_L g128 ( .A1(n_26), .A2(n_49), .B1(n_129), .B2(n_132), .Y(n_128) );
HB1xp67_ASAP7_75t_L g177 ( .A(n_27), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_28), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_29), .Y(n_179) );
XOR2xp5_ASAP7_75t_L g618 ( .A(n_30), .B(n_82), .Y(n_618) );
INVx1_ASAP7_75t_L g239 ( .A(n_32), .Y(n_239) );
HB1xp67_ASAP7_75t_L g206 ( .A(n_33), .Y(n_206) );
AND2x4_ASAP7_75t_L g235 ( .A(n_33), .B(n_204), .Y(n_235) );
AND2x4_ASAP7_75t_L g256 ( .A(n_33), .B(n_204), .Y(n_256) );
AOI22xp5_ASAP7_75t_L g180 ( .A1(n_34), .A2(n_181), .B1(n_184), .B2(n_185), .Y(n_180) );
INVx2_ASAP7_75t_L g183 ( .A(n_34), .Y(n_183) );
INVx1_ASAP7_75t_L g160 ( .A(n_35), .Y(n_160) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_36), .Y(n_226) );
CKINVDCx5p33_ASAP7_75t_R g315 ( .A(n_37), .Y(n_315) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_38), .Y(n_232) );
INVx2_ASAP7_75t_L g277 ( .A(n_39), .Y(n_277) );
O2A1O1Ixp33_ASAP7_75t_L g329 ( .A1(n_40), .A2(n_225), .B(n_330), .C(n_331), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_41), .Y(n_314) );
INVx1_ASAP7_75t_L g146 ( .A(n_42), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_43), .B(n_257), .Y(n_319) );
AOI22xp33_ASAP7_75t_L g134 ( .A1(n_44), .A2(n_69), .B1(n_135), .B2(n_136), .Y(n_134) );
AOI22xp5_ASAP7_75t_L g292 ( .A1(n_46), .A2(n_62), .B1(n_293), .B2(n_294), .Y(n_292) );
OA22x2_ASAP7_75t_L g98 ( .A1(n_47), .A2(n_56), .B1(n_92), .B2(n_96), .Y(n_98) );
INVx1_ASAP7_75t_L g124 ( .A(n_47), .Y(n_124) );
AOI21xp5_ASAP7_75t_SL g142 ( .A1(n_48), .A2(n_143), .B(n_145), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g318 ( .A(n_50), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g86 ( .A1(n_51), .A2(n_57), .B1(n_87), .B2(n_110), .Y(n_86) );
NAND2xp33_ASAP7_75t_R g258 ( .A(n_52), .B(n_243), .Y(n_258) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_52), .A2(n_76), .B1(n_297), .B2(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g109 ( .A(n_55), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_55), .B(n_122), .Y(n_155) );
HB1xp67_ASAP7_75t_L g198 ( .A(n_55), .Y(n_198) );
OAI21xp33_ASAP7_75t_L g125 ( .A1(n_56), .A2(n_63), .B(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g139 ( .A(n_58), .Y(n_139) );
AOI22xp5_ASAP7_75t_L g113 ( .A1(n_59), .A2(n_70), .B1(n_114), .B2(n_119), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_60), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_61), .Y(n_273) );
INVx1_ASAP7_75t_L g95 ( .A(n_63), .Y(n_95) );
NOR2xp33_ASAP7_75t_L g153 ( .A(n_63), .B(n_73), .Y(n_153) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_65), .Y(n_221) );
BUFx5_ASAP7_75t_L g223 ( .A(n_65), .Y(n_223) );
INVx1_ASAP7_75t_L g252 ( .A(n_65), .Y(n_252) );
INVx2_ASAP7_75t_L g365 ( .A(n_66), .Y(n_365) );
INVx2_ASAP7_75t_L g334 ( .A(n_67), .Y(n_334) );
CKINVDCx5p33_ASAP7_75t_R g362 ( .A(n_68), .Y(n_362) );
INVx2_ASAP7_75t_SL g204 ( .A(n_71), .Y(n_204) );
HB1xp67_ASAP7_75t_L g80 ( .A(n_72), .Y(n_80) );
INVx1_ASAP7_75t_L g230 ( .A(n_72), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g101 ( .A(n_73), .B(n_102), .Y(n_101) );
INVx2_ASAP7_75t_L g241 ( .A(n_74), .Y(n_241) );
OAI21xp33_ASAP7_75t_SL g325 ( .A1(n_75), .A2(n_223), .B(n_326), .Y(n_325) );
INVxp67_ASAP7_75t_SL g279 ( .A(n_76), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_76), .B(n_297), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_190), .B1(n_207), .B2(n_604), .C(n_611), .Y(n_77) );
XOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_176), .Y(n_78) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_80), .A2(n_81), .B1(n_82), .B2(n_175), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g175 ( .A(n_80), .Y(n_175) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_81), .A2(n_82), .B1(n_613), .B2(n_614), .Y(n_612) );
INVx1_ASAP7_75t_L g81 ( .A(n_82), .Y(n_81) );
INVxp33_ASAP7_75t_L g82 ( .A(n_83), .Y(n_82) );
AND2x2_ASAP7_75t_L g83 ( .A(n_84), .B(n_137), .Y(n_83) );
NOR2xp33_ASAP7_75t_L g84 ( .A(n_85), .B(n_127), .Y(n_84) );
NAND2xp5_ASAP7_75t_L g85 ( .A(n_86), .B(n_113), .Y(n_85) );
AND2x4_ASAP7_75t_L g87 ( .A(n_88), .B(n_99), .Y(n_87) );
AND2x4_ASAP7_75t_L g110 ( .A(n_88), .B(n_111), .Y(n_110) );
AND2x4_ASAP7_75t_L g129 ( .A(n_88), .B(n_130), .Y(n_129) );
AND2x4_ASAP7_75t_L g132 ( .A(n_88), .B(n_133), .Y(n_132) );
AND2x4_ASAP7_75t_L g88 ( .A(n_89), .B(n_97), .Y(n_88) );
AND2x2_ASAP7_75t_L g144 ( .A(n_89), .B(n_98), .Y(n_144) );
INVx1_ASAP7_75t_L g89 ( .A(n_90), .Y(n_89) );
AND2x2_ASAP7_75t_L g115 ( .A(n_90), .B(n_98), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g90 ( .A(n_91), .B(n_94), .Y(n_90) );
NAND2xp33_ASAP7_75t_L g91 ( .A(n_92), .B(n_93), .Y(n_91) );
INVx2_ASAP7_75t_L g96 ( .A(n_92), .Y(n_96) );
INVx3_ASAP7_75t_L g102 ( .A(n_92), .Y(n_102) );
NAND2xp33_ASAP7_75t_L g108 ( .A(n_92), .B(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g126 ( .A(n_92), .Y(n_126) );
HB1xp67_ASAP7_75t_L g150 ( .A(n_92), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_93), .B(n_124), .Y(n_123) );
INVxp67_ASAP7_75t_L g199 ( .A(n_93), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g94 ( .A(n_95), .B(n_96), .Y(n_94) );
OAI21xp5_ASAP7_75t_L g173 ( .A1(n_95), .A2(n_126), .B(n_174), .Y(n_173) );
INVx1_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
AND2x2_ASAP7_75t_L g172 ( .A(n_98), .B(n_173), .Y(n_172) );
AND2x4_ASAP7_75t_L g159 ( .A(n_99), .B(n_144), .Y(n_159) );
AND2x4_ASAP7_75t_L g166 ( .A(n_99), .B(n_115), .Y(n_166) );
AND2x4_ASAP7_75t_L g99 ( .A(n_100), .B(n_104), .Y(n_99) );
INVx2_ASAP7_75t_L g112 ( .A(n_100), .Y(n_112) );
OR2x2_ASAP7_75t_L g117 ( .A(n_100), .B(n_118), .Y(n_117) );
AND2x4_ASAP7_75t_L g130 ( .A(n_100), .B(n_131), .Y(n_130) );
AND2x2_ASAP7_75t_L g169 ( .A(n_100), .B(n_170), .Y(n_169) );
AND2x4_ASAP7_75t_L g100 ( .A(n_101), .B(n_103), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_102), .B(n_107), .Y(n_106) );
INVxp67_ASAP7_75t_L g122 ( .A(n_102), .Y(n_122) );
NAND3xp33_ASAP7_75t_L g154 ( .A(n_103), .B(n_121), .C(n_155), .Y(n_154) );
AND2x4_ASAP7_75t_L g111 ( .A(n_104), .B(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g118 ( .A(n_105), .Y(n_118) );
AND2x2_ASAP7_75t_L g105 ( .A(n_106), .B(n_108), .Y(n_105) );
AND2x2_ASAP7_75t_L g141 ( .A(n_111), .B(n_115), .Y(n_141) );
AND2x2_ASAP7_75t_L g143 ( .A(n_111), .B(n_144), .Y(n_143) );
AND2x4_ASAP7_75t_L g162 ( .A(n_111), .B(n_120), .Y(n_162) );
AND2x4_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
AND2x4_ASAP7_75t_L g135 ( .A(n_115), .B(n_130), .Y(n_135) );
AND2x4_ASAP7_75t_L g119 ( .A(n_116), .B(n_120), .Y(n_119) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g133 ( .A(n_117), .Y(n_133) );
INVx1_ASAP7_75t_L g131 ( .A(n_118), .Y(n_131) );
AND2x4_ASAP7_75t_L g136 ( .A(n_120), .B(n_130), .Y(n_136) );
AND2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_125), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g121 ( .A(n_122), .B(n_123), .Y(n_121) );
HB1xp67_ASAP7_75t_L g200 ( .A(n_124), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_134), .Y(n_127) );
NOR3xp33_ASAP7_75t_L g137 ( .A(n_138), .B(n_156), .C(n_163), .Y(n_137) );
OAI21xp33_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_140), .B(n_142), .Y(n_138) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
NOR2xp33_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
AO21x2_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_151), .B(n_154), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_150), .B(n_171), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
OAI22xp33_ASAP7_75t_L g156 ( .A1(n_157), .A2(n_158), .B1(n_160), .B2(n_161), .Y(n_156) );
INVx2_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
OAI21xp5_ASAP7_75t_SL g163 ( .A1(n_164), .A2(n_165), .B(n_167), .Y(n_163) );
INVx1_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
AND2x4_ASAP7_75t_L g168 ( .A(n_169), .B(n_172), .Y(n_168) );
HB1xp67_ASAP7_75t_L g196 ( .A(n_171), .Y(n_196) );
AOI22xp5_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_178), .B1(n_188), .B2(n_189), .Y(n_176) );
CKINVDCx5p33_ASAP7_75t_R g188 ( .A(n_177), .Y(n_188) );
CKINVDCx20_ASAP7_75t_R g189 ( .A(n_178), .Y(n_189) );
AOI22xp5_ASAP7_75t_L g178 ( .A1(n_179), .A2(n_180), .B1(n_186), .B2(n_187), .Y(n_178) );
CKINVDCx5p33_ASAP7_75t_R g186 ( .A(n_179), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_180), .Y(n_187) );
CKINVDCx5p33_ASAP7_75t_R g181 ( .A(n_182), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
BUFx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
CKINVDCx5p33_ASAP7_75t_R g191 ( .A(n_192), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_193), .B(n_201), .Y(n_192) );
INVxp67_ASAP7_75t_SL g193 ( .A(n_194), .Y(n_193) );
AND2x2_ASAP7_75t_L g616 ( .A(n_194), .B(n_201), .Y(n_616) );
AOI211xp5_ASAP7_75t_L g194 ( .A1(n_195), .A2(n_196), .B(n_197), .C(n_200), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_202), .B(n_205), .Y(n_201) );
OR2x2_ASAP7_75t_L g620 ( .A(n_202), .B(n_206), .Y(n_620) );
INVx1_ASAP7_75t_L g623 ( .A(n_202), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_202), .B(n_205), .Y(n_624) );
HB1xp67_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
HB1xp67_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
AND4x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_462), .C(n_502), .D(n_571), .Y(n_210) );
NOR2x1_ASAP7_75t_L g211 ( .A(n_212), .B(n_400), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_213), .B(n_380), .Y(n_212) );
O2A1O1Ixp33_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_259), .B(n_283), .C(n_335), .Y(n_213) );
AND2x2_ASAP7_75t_L g394 ( .A(n_214), .B(n_395), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_214), .B(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g448 ( .A(n_214), .Y(n_448) );
AND2x2_ASAP7_75t_L g468 ( .A(n_214), .B(n_337), .Y(n_468) );
AND2x2_ASAP7_75t_L g570 ( .A(n_214), .B(n_551), .Y(n_570) );
AND2x4_ASAP7_75t_L g214 ( .A(n_215), .B(n_244), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_215), .B(n_387), .Y(n_386) );
OR2x2_ASAP7_75t_L g596 ( .A(n_215), .B(n_535), .Y(n_596) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
AND2x2_ASAP7_75t_L g367 ( .A(n_216), .B(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g374 ( .A(n_216), .Y(n_374) );
BUFx2_ASAP7_75t_R g434 ( .A(n_216), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_216), .B(n_351), .Y(n_543) );
AND2x2_ASAP7_75t_L g547 ( .A(n_216), .B(n_350), .Y(n_547) );
AO21x2_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_236), .B(n_240), .Y(n_216) );
NOR3xp33_ASAP7_75t_L g217 ( .A(n_218), .B(n_227), .C(n_234), .Y(n_217) );
INVx1_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
INVx1_ASAP7_75t_L g228 ( .A(n_220), .Y(n_228) );
INVx1_ASAP7_75t_L g330 ( .A(n_220), .Y(n_330) );
INVx3_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx2_ASAP7_75t_L g249 ( .A(n_221), .Y(n_249) );
INVx2_ASAP7_75t_L g253 ( .A(n_221), .Y(n_253) );
INVx6_ASAP7_75t_L g271 ( .A(n_221), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_223), .B(n_224), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_223), .B(n_232), .Y(n_231) );
AOI22xp5_ASAP7_75t_L g270 ( .A1(n_223), .A2(n_271), .B1(n_272), .B2(n_273), .Y(n_270) );
AOI22xp33_ASAP7_75t_SL g313 ( .A1(n_223), .A2(n_271), .B1(n_314), .B2(n_315), .Y(n_313) );
AOI22xp33_ASAP7_75t_L g316 ( .A1(n_223), .A2(n_249), .B1(n_317), .B2(n_318), .Y(n_316) );
NAND2xp5_ASAP7_75t_SL g326 ( .A(n_223), .B(n_327), .Y(n_326) );
AOI22xp5_ASAP7_75t_L g247 ( .A1(n_225), .A2(n_233), .B1(n_248), .B2(n_250), .Y(n_247) );
OAI22xp33_ASAP7_75t_L g269 ( .A1(n_225), .A2(n_233), .B1(n_270), .B2(n_274), .Y(n_269) );
OAI221xp5_ASAP7_75t_L g312 ( .A1(n_225), .A2(n_256), .B1(n_307), .B2(n_313), .C(n_316), .Y(n_312) );
INVx1_ASAP7_75t_L g393 ( .A(n_225), .Y(n_393) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_226), .B(n_230), .Y(n_229) );
INVx4_ASAP7_75t_L g233 ( .A(n_226), .Y(n_233) );
BUFx6f_ASAP7_75t_L g290 ( .A(n_226), .Y(n_290) );
INVx1_ASAP7_75t_L g295 ( .A(n_226), .Y(n_295) );
NAND2xp5_ASAP7_75t_SL g303 ( .A(n_226), .B(n_304), .Y(n_303) );
INVx3_ASAP7_75t_L g307 ( .A(n_226), .Y(n_307) );
OAI22xp5_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_229), .B1(n_231), .B2(n_233), .Y(n_227) );
INVx2_ASAP7_75t_L g328 ( .A(n_233), .Y(n_328) );
NOR2xp33_ASAP7_75t_SL g363 ( .A(n_234), .B(n_281), .Y(n_363) );
AOI221xp5_ASAP7_75t_L g390 ( .A1(n_234), .A2(n_328), .B1(n_391), .B2(n_392), .C(n_393), .Y(n_390) );
INVx4_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_235), .B(n_267), .Y(n_288) );
AND2x2_ASAP7_75t_L g322 ( .A(n_235), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_SL g389 ( .A(n_236), .B(n_390), .Y(n_389) );
BUFx3_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx3_ASAP7_75t_L g257 ( .A(n_237), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_237), .B(n_334), .Y(n_333) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx4_ASAP7_75t_L g282 ( .A(n_238), .Y(n_282) );
BUFx3_ASAP7_75t_L g344 ( .A(n_238), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_241), .B(n_242), .Y(n_240) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
BUFx3_ASAP7_75t_L g268 ( .A(n_243), .Y(n_268) );
INVx1_ASAP7_75t_L g323 ( .A(n_243), .Y(n_323) );
INVx2_ASAP7_75t_L g521 ( .A(n_243), .Y(n_521) );
INVx1_ASAP7_75t_SL g261 ( .A(n_244), .Y(n_261) );
INVx1_ASAP7_75t_L g375 ( .A(n_244), .Y(n_375) );
AND2x2_ASAP7_75t_L g457 ( .A(n_244), .B(n_350), .Y(n_457) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g368 ( .A(n_245), .Y(n_368) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_245), .Y(n_384) );
AND2x2_ASAP7_75t_L g472 ( .A(n_245), .B(n_374), .Y(n_472) );
AND2x2_ASAP7_75t_L g544 ( .A(n_245), .B(n_264), .Y(n_544) );
AND2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_258), .Y(n_245) );
AND2x2_ASAP7_75t_L g518 ( .A(n_246), .B(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_247), .B(n_254), .Y(n_246) );
AOI22xp5_ASAP7_75t_L g274 ( .A1(n_249), .A2(n_275), .B1(n_276), .B2(n_277), .Y(n_274) );
INVx1_ASAP7_75t_L g360 ( .A(n_249), .Y(n_360) );
INVx2_ASAP7_75t_L g293 ( .A(n_251), .Y(n_293) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
INVx2_ASAP7_75t_L g276 ( .A(n_252), .Y(n_276) );
NOR2xp67_ASAP7_75t_L g254 ( .A(n_255), .B(n_257), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
BUFx6f_ASAP7_75t_L g266 ( .A(n_256), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_256), .B(n_282), .Y(n_308) );
INVxp67_ASAP7_75t_SL g259 ( .A(n_260), .Y(n_259) );
OR2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_262), .B(n_366), .Y(n_593) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x4_ASAP7_75t_L g459 ( .A(n_264), .B(n_351), .Y(n_459) );
OAI21x1_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_269), .B(n_278), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
AND2x2_ASAP7_75t_L g605 ( .A(n_266), .B(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g391 ( .A(n_270), .Y(n_391) );
INVx2_ASAP7_75t_SL g294 ( .A(n_271), .Y(n_294) );
INVx2_ASAP7_75t_L g356 ( .A(n_271), .Y(n_356) );
INVx1_ASAP7_75t_L g613 ( .A(n_272), .Y(n_613) );
INVx1_ASAP7_75t_L g626 ( .A(n_273), .Y(n_626) );
INVx1_ASAP7_75t_L g392 ( .A(n_274), .Y(n_392) );
NAND2xp5_ASAP7_75t_SL g331 ( .A(n_276), .B(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_276), .B(n_362), .Y(n_361) );
OR2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
INVx2_ASAP7_75t_L g311 ( .A(n_280), .Y(n_311) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g297 ( .A(n_282), .Y(n_297) );
NOR2xp33_ASAP7_75t_SL g364 ( .A(n_282), .B(n_365), .Y(n_364) );
INVxp67_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_298), .Y(n_284) );
AND2x4_ASAP7_75t_L g377 ( .A(n_285), .B(n_378), .Y(n_377) );
INVx2_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g461 ( .A(n_286), .B(n_430), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_286), .B(n_455), .Y(n_474) );
OR2x2_ASAP7_75t_L g578 ( .A(n_286), .B(n_534), .Y(n_578) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
INVx2_ASAP7_75t_L g414 ( .A(n_287), .Y(n_414) );
OAI21x1_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_289), .B(n_296), .Y(n_287) );
INVx1_ASAP7_75t_L g342 ( .A(n_289), .Y(n_342) );
OA22x2_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_291), .B1(n_292), .B2(n_295), .Y(n_289) );
INVx4_ASAP7_75t_L g610 ( .A(n_290), .Y(n_610) );
INVx1_ASAP7_75t_L g354 ( .A(n_293), .Y(n_354) );
INVx1_ASAP7_75t_L g345 ( .A(n_296), .Y(n_345) );
BUFx2_ASAP7_75t_SL g442 ( .A(n_298), .Y(n_442) );
NOR2xp67_ASAP7_75t_L g298 ( .A(n_299), .B(n_309), .Y(n_298) );
INVx1_ASAP7_75t_L g397 ( .A(n_299), .Y(n_397) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g379 ( .A(n_300), .Y(n_379) );
INVx3_ASAP7_75t_L g416 ( .A(n_300), .Y(n_416) );
AND2x2_ASAP7_75t_L g451 ( .A(n_300), .B(n_417), .Y(n_451) );
AND2x2_ASAP7_75t_L g481 ( .A(n_300), .B(n_320), .Y(n_481) );
AND2x4_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_305), .Y(n_302) );
AOI21xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_307), .B(n_308), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_320), .Y(n_309) );
INVx2_ASAP7_75t_L g346 ( .A(n_310), .Y(n_346) );
INVx2_ASAP7_75t_L g399 ( .A(n_310), .Y(n_399) );
OA21x2_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_312), .B(n_319), .Y(n_310) );
OA21x2_ASAP7_75t_L g417 ( .A1(n_311), .A2(n_312), .B(n_319), .Y(n_417) );
INVx1_ASAP7_75t_L g338 ( .A(n_320), .Y(n_338) );
AND2x2_ASAP7_75t_L g398 ( .A(n_320), .B(n_399), .Y(n_398) );
OR2x2_ASAP7_75t_L g424 ( .A(n_320), .B(n_379), .Y(n_424) );
INVx2_ASAP7_75t_L g430 ( .A(n_320), .Y(n_430) );
AND2x2_ASAP7_75t_L g455 ( .A(n_320), .B(n_416), .Y(n_455) );
BUFx2_ASAP7_75t_L g524 ( .A(n_320), .Y(n_524) );
INVx2_ASAP7_75t_L g535 ( .A(n_320), .Y(n_535) );
INVx3_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AOI21x1_ASAP7_75t_L g321 ( .A1(n_322), .A2(n_324), .B(n_333), .Y(n_321) );
AOI21xp5_ASAP7_75t_L g324 ( .A1(n_325), .A2(n_328), .B(n_329), .Y(n_324) );
OAI22xp5_ASAP7_75t_L g335 ( .A1(n_336), .A2(n_347), .B1(n_369), .B2(n_376), .Y(n_335) );
OR2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_339), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g436 ( .A(n_340), .B(n_429), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_340), .B(n_481), .Y(n_480) );
INVx2_ASAP7_75t_SL g530 ( .A(n_340), .Y(n_530) );
AND2x4_ASAP7_75t_L g340 ( .A(n_341), .B(n_346), .Y(n_340) );
OR2x2_ASAP7_75t_L g422 ( .A(n_341), .B(n_417), .Y(n_422) );
AOI21xp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_343), .B(n_345), .Y(n_341) );
INVx3_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
AND2x4_ASAP7_75t_L g378 ( .A(n_346), .B(n_379), .Y(n_378) );
NAND3xp33_ASAP7_75t_L g402 ( .A(n_347), .B(n_403), .C(n_407), .Y(n_402) );
OR2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_366), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OR2x2_ASAP7_75t_L g385 ( .A(n_349), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g395 ( .A(n_351), .B(n_387), .Y(n_395) );
INVx1_ASAP7_75t_L g406 ( .A(n_351), .Y(n_406) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_351), .Y(n_410) );
OR2x2_ASAP7_75t_L g439 ( .A(n_351), .B(n_387), .Y(n_439) );
INVx1_ASAP7_75t_L g476 ( .A(n_351), .Y(n_476) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_351), .Y(n_598) );
AO31x2_ASAP7_75t_L g351 ( .A1(n_352), .A2(n_358), .A3(n_363), .B(n_364), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_356), .B(n_357), .Y(n_355) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_360), .Y(n_608) );
OR2x2_ASAP7_75t_L g425 ( .A(n_366), .B(n_426), .Y(n_425) );
INVx2_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
AND2x4_ASAP7_75t_L g437 ( .A(n_367), .B(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g446 ( .A(n_367), .B(n_395), .Y(n_446) );
AND2x4_ASAP7_75t_L g482 ( .A(n_367), .B(n_459), .Y(n_482) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
OR2x2_ASAP7_75t_L g527 ( .A(n_372), .B(n_410), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_375), .Y(n_372) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_373), .B(n_387), .Y(n_567) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_374), .Y(n_501) );
AND2x2_ASAP7_75t_L g552 ( .A(n_374), .B(n_517), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_376), .B(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AND2x2_ASAP7_75t_L g559 ( .A(n_377), .B(n_512), .Y(n_559) );
NAND2x1p5_ASAP7_75t_L g523 ( .A(n_378), .B(n_524), .Y(n_523) );
NAND2x1p5_ASAP7_75t_L g569 ( .A(n_378), .B(n_564), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_378), .B(n_461), .Y(n_582) );
AND2x2_ASAP7_75t_L g444 ( .A(n_379), .B(n_414), .Y(n_444) );
OAI21xp5_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_394), .B(n_396), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
OR2x2_ASAP7_75t_L g382 ( .A(n_383), .B(n_385), .Y(n_382) );
AND2x2_ASAP7_75t_L g404 ( .A(n_383), .B(n_405), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_383), .B(n_459), .Y(n_458) );
OR2x2_ASAP7_75t_L g485 ( .A(n_383), .B(n_486), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_383), .B(n_538), .Y(n_537) );
INVx2_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
INVx2_ASAP7_75t_L g531 ( .A(n_385), .Y(n_531) );
INVx1_ASAP7_75t_L g602 ( .A(n_386), .Y(n_602) );
AND2x2_ASAP7_75t_L g405 ( .A(n_387), .B(n_406), .Y(n_405) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_387), .Y(n_491) );
AND2x2_ASAP7_75t_L g387 ( .A(n_388), .B(n_389), .Y(n_387) );
AND2x2_ASAP7_75t_L g517 ( .A(n_389), .B(n_518), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_395), .B(n_434), .Y(n_433) );
BUFx6f_ASAP7_75t_L g538 ( .A(n_395), .Y(n_538) );
AOI22xp5_ASAP7_75t_SL g477 ( .A1(n_396), .A2(n_478), .B1(n_479), .B2(n_482), .Y(n_477) );
AND2x4_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_401), .B(n_435), .Y(n_400) );
AOI21xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_411), .B(n_418), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g449 ( .A(n_405), .Y(n_449) );
OR2x2_ASAP7_75t_L g515 ( .A(n_406), .B(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g587 ( .A(n_406), .B(n_544), .Y(n_587) );
INVxp67_ASAP7_75t_SL g478 ( .A(n_407), .Y(n_478) );
BUFx3_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVxp67_ASAP7_75t_L g426 ( .A(n_409), .Y(n_426) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
AND2x2_ASAP7_75t_L g411 ( .A(n_412), .B(n_415), .Y(n_411) );
A2O1A1Ixp33_ASAP7_75t_L g483 ( .A1(n_412), .A2(n_481), .B(n_484), .C(n_487), .Y(n_483) );
OR2x2_ASAP7_75t_L g556 ( .A(n_412), .B(n_424), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_412), .B(n_415), .Y(n_590) );
AND2x2_ASAP7_75t_L g603 ( .A(n_412), .B(n_451), .Y(n_603) );
INVx3_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
AND2x4_ASAP7_75t_L g511 ( .A(n_413), .B(n_415), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_413), .B(n_451), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_413), .B(n_455), .Y(n_574) );
AND2x2_ASAP7_75t_L g579 ( .A(n_413), .B(n_481), .Y(n_579) );
INVx3_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g467 ( .A(n_414), .Y(n_467) );
AND2x2_ASAP7_75t_L g585 ( .A(n_414), .B(n_417), .Y(n_585) );
AND2x2_ASAP7_75t_L g492 ( .A(n_415), .B(n_461), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_415), .B(n_524), .Y(n_555) );
AND2x4_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_416), .B(n_535), .Y(n_534) );
AND2x2_ASAP7_75t_L g466 ( .A(n_417), .B(n_467), .Y(n_466) );
OAI22xp5_ASAP7_75t_SL g418 ( .A1(n_419), .A2(n_425), .B1(n_427), .B2(n_431), .Y(n_418) );
INVx2_ASAP7_75t_SL g419 ( .A(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_421), .B(n_423), .Y(n_420) );
AND2x2_ASAP7_75t_L g428 ( .A(n_421), .B(n_429), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_421), .B(n_564), .Y(n_563) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g453 ( .A(n_422), .Y(n_453) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_SL g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_L g512 ( .A(n_429), .Y(n_512) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g495 ( .A(n_430), .B(n_444), .Y(n_495) );
AND2x2_ASAP7_75t_L g497 ( .A(n_430), .B(n_451), .Y(n_497) );
INVx1_ASAP7_75t_L g565 ( .A(n_430), .Y(n_565) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_432), .A2(n_570), .B1(n_577), .B2(n_579), .Y(n_576) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g507 ( .A(n_434), .Y(n_507) );
AOI211xp5_ASAP7_75t_SL g435 ( .A1(n_436), .A2(n_437), .B(n_440), .C(n_447), .Y(n_435) );
NOR2x1_ASAP7_75t_L g575 ( .A(n_437), .B(n_541), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_438), .B(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
AOI21xp33_ASAP7_75t_L g440 ( .A1(n_441), .A2(n_443), .B(n_445), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
OAI332xp33_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_449), .A3(n_450), .B1(n_452), .B2(n_454), .B3(n_456), .C1(n_458), .C2(n_460), .Y(n_447) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g540 ( .A1(n_451), .A2(n_541), .B1(n_545), .B2(n_546), .Y(n_540) );
INVxp67_ASAP7_75t_SL g545 ( .A(n_452), .Y(n_545) );
INVx2_ASAP7_75t_SL g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_SL g600 ( .A(n_454), .Y(n_600) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
AND2x2_ASAP7_75t_L g566 ( .A(n_457), .B(n_567), .Y(n_566) );
AND2x2_ASAP7_75t_L g601 ( .A(n_457), .B(n_602), .Y(n_601) );
INVx2_ASAP7_75t_SL g486 ( .A(n_459), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_459), .B(n_472), .Y(n_487) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AND4x1_ASAP7_75t_L g462 ( .A(n_463), .B(n_477), .C(n_483), .D(n_488), .Y(n_462) );
A2O1A1Ixp33_ASAP7_75t_L g463 ( .A1(n_464), .A2(n_468), .B(n_469), .C(n_475), .Y(n_463) );
INVxp67_ASAP7_75t_SL g464 ( .A(n_465), .Y(n_464) );
OAI321xp33_ASAP7_75t_L g591 ( .A1(n_465), .A2(n_532), .A3(n_545), .B1(n_592), .B2(n_594), .C(n_599), .Y(n_591) );
INVx3_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVxp67_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_471), .B(n_473), .Y(n_470) );
BUFx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_SL g551 ( .A(n_476), .Y(n_551) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_486), .A2(n_494), .B(n_496), .Y(n_493) );
A2O1A1Ixp33_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_492), .B(n_493), .C(n_498), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVxp67_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_497), .A2(n_514), .B1(n_522), .B2(n_525), .Y(n_513) );
INVxp67_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
NOR2x1_ASAP7_75t_L g502 ( .A(n_503), .B(n_539), .Y(n_502) );
OAI211xp5_ASAP7_75t_SL g503 ( .A1(n_504), .A2(n_508), .B(n_513), .C(n_528), .Y(n_503) );
INVxp67_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_512), .Y(n_510) );
OR2x2_ASAP7_75t_L g583 ( .A(n_512), .B(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_515), .B(n_590), .Y(n_589) );
OR2x2_ASAP7_75t_L g597 ( .A(n_516), .B(n_598), .Y(n_597) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
INVx2_ASAP7_75t_L g558 ( .A(n_517), .Y(n_558) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
HB1xp67_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
AOI32xp33_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_531), .A3(n_532), .B1(n_533), .B2(n_536), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
NAND3xp33_ASAP7_75t_SL g539 ( .A(n_540), .B(n_548), .C(n_560), .Y(n_539) );
AND2x4_ASAP7_75t_L g541 ( .A(n_542), .B(n_544), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g546 ( .A(n_544), .B(n_547), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_544), .A2(n_600), .B1(n_601), .B2(n_603), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_553), .B1(n_557), .B2(n_559), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NAND2x1p5_ASAP7_75t_SL g550 ( .A(n_551), .B(n_552), .Y(n_550) );
NAND3xp33_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .C(n_556), .Y(n_553) );
A2O1A1Ixp33_ASAP7_75t_L g572 ( .A1(n_556), .A2(n_573), .B(n_575), .C(n_576), .Y(n_572) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
AOI22xp5_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_566), .B1(n_568), .B2(n_570), .Y(n_560) );
BUFx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NOR3xp33_ASAP7_75t_L g571 ( .A(n_572), .B(n_580), .C(n_591), .Y(n_571) );
BUFx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
A2O1A1Ixp33_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_583), .B(n_586), .C(n_588), .Y(n_580) );
HB1xp67_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVxp67_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
NOR2x1_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
BUFx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
OA21x2_ASAP7_75t_L g622 ( .A1(n_606), .A2(n_623), .B(n_624), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_607), .B(n_609), .Y(n_606) );
CKINVDCx16_ASAP7_75t_R g607 ( .A(n_608), .Y(n_607) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
OAI222xp33_ASAP7_75t_L g611 ( .A1(n_612), .A2(n_615), .B1(n_617), .B2(n_619), .C1(n_621), .C2(n_625), .Y(n_611) );
INVx1_ASAP7_75t_L g614 ( .A(n_613), .Y(n_614) );
INVx1_ASAP7_75t_SL g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
BUFx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
BUFx3_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
endmodule