module real_jpeg_20412_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_330, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_330;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_0),
.A2(n_25),
.B1(n_26),
.B2(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_0),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_0),
.A2(n_47),
.B1(n_48),
.B2(n_66),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g233 ( 
.A1(n_0),
.A2(n_42),
.B1(n_43),
.B2(n_66),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_0),
.A2(n_31),
.B1(n_32),
.B2(n_66),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_1),
.A2(n_25),
.B1(n_26),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_1),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_1),
.A2(n_42),
.B1(n_43),
.B2(n_63),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_1),
.A2(n_47),
.B1(n_48),
.B2(n_63),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_1),
.A2(n_31),
.B1(n_32),
.B2(n_63),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_2),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_2),
.A2(n_24),
.B1(n_31),
.B2(n_32),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_2),
.A2(n_24),
.B1(n_47),
.B2(n_48),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_2),
.A2(n_24),
.B1(n_42),
.B2(n_43),
.Y(n_266)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_4),
.A2(n_35),
.B1(n_42),
.B2(n_43),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_35),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_4),
.A2(n_35),
.B1(n_47),
.B2(n_48),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_5),
.A2(n_42),
.B1(n_43),
.B2(n_95),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_5),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_5),
.A2(n_31),
.B1(n_32),
.B2(n_95),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_5),
.A2(n_47),
.B1(n_48),
.B2(n_95),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g256 ( 
.A1(n_5),
.A2(n_25),
.B1(n_26),
.B2(n_95),
.Y(n_256)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_6),
.Y(n_83)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_6),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_7),
.A2(n_42),
.B1(n_43),
.B2(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_7),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_7),
.A2(n_47),
.B1(n_48),
.B2(n_89),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_7),
.A2(n_31),
.B1(n_32),
.B2(n_89),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_89),
.Y(n_287)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_9),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_9),
.B(n_30),
.Y(n_134)
);

AOI21xp33_ASAP7_75t_L g155 ( 
.A1(n_9),
.A2(n_44),
.B(n_47),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_9),
.A2(n_42),
.B1(n_43),
.B2(n_104),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_9),
.A2(n_82),
.B1(n_85),
.B2(n_163),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_9),
.B(n_58),
.Y(n_176)
);

AOI21xp33_ASAP7_75t_L g193 ( 
.A1(n_9),
.A2(n_32),
.B(n_194),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_10),
.A2(n_31),
.B1(n_32),
.B2(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_10),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_10),
.A2(n_47),
.B1(n_48),
.B2(n_101),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_10),
.A2(n_42),
.B1(n_43),
.B2(n_101),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_10),
.A2(n_25),
.B1(n_26),
.B2(n_101),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_11),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_106),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_11),
.A2(n_42),
.B1(n_43),
.B2(n_106),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_11),
.A2(n_47),
.B1(n_48),
.B2(n_106),
.Y(n_163)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_13),
.A2(n_31),
.B1(n_32),
.B2(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_13),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_99),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_13),
.A2(n_47),
.B1(n_48),
.B2(n_99),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_13),
.A2(n_42),
.B1(n_43),
.B2(n_99),
.Y(n_179)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_14),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_14),
.A2(n_42),
.B1(n_43),
.B2(n_54),
.Y(n_56)
);

OAI32xp33_ASAP7_75t_L g188 ( 
.A1(n_14),
.A2(n_32),
.A3(n_43),
.B1(n_189),
.B2(n_190),
.Y(n_188)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx3_ASAP7_75t_SL g43 ( 
.A(n_17),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_72),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_71),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_36),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_22),
.B(n_36),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_27),
.B1(n_30),
.B2(n_34),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_23),
.A2(n_27),
.B1(n_30),
.B2(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_25),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g27 ( 
.A1(n_25),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_28),
.Y(n_29)
);

HAxp5_ASAP7_75t_SL g103 ( 
.A(n_25),
.B(n_104),
.CON(n_103),
.SN(n_103)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_27),
.A2(n_30),
.B1(n_103),
.B2(n_105),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_27),
.A2(n_30),
.B1(n_286),
.B2(n_287),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_28),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_30)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_28),
.B(n_32),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_29),
.A2(n_31),
.B1(n_103),
.B2(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_31),
.A2(n_54),
.B(n_55),
.C(n_56),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_31),
.B(n_54),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_31),
.B(n_104),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_67),
.C(n_69),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_37),
.A2(n_38),
.B1(n_325),
.B2(n_327),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_50),
.C(n_59),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_39),
.A2(n_296),
.B1(n_297),
.B2(n_299),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_39),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_39),
.A2(n_50),
.B1(n_299),
.B2(n_312),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_46),
.B(n_49),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_40),
.A2(n_46),
.B1(n_88),
.B2(n_90),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_40),
.A2(n_46),
.B1(n_88),
.B2(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_40),
.A2(n_46),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_40),
.A2(n_46),
.B1(n_159),
.B2(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_40),
.A2(n_46),
.B1(n_179),
.B2(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_40),
.A2(n_46),
.B1(n_94),
.B2(n_197),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_40),
.A2(n_46),
.B1(n_90),
.B2(n_233),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_40),
.A2(n_46),
.B1(n_233),
.B2(n_266),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_40),
.A2(n_46),
.B1(n_49),
.B2(n_266),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_46),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_42),
.B(n_54),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g42 ( 
.A(n_43),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_43),
.A2(n_45),
.B(n_104),
.C(n_155),
.Y(n_154)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_44),
.A2(n_45),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

CKINVDCx9p33_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_46),
.B(n_104),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g48 ( 
.A(n_47),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_48),
.B(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_50),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_57),
.B2(n_58),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_51),
.A2(n_52),
.B1(n_58),
.B2(n_298),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_52),
.A2(n_57),
.B(n_58),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_52),
.A2(n_58),
.B1(n_131),
.B2(n_133),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_52),
.A2(n_58),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_53),
.A2(n_56),
.B1(n_98),
.B2(n_100),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_53),
.A2(n_56),
.B1(n_100),
.B2(n_114),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_53),
.A2(n_56),
.B1(n_132),
.B2(n_193),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_53),
.A2(n_56),
.B1(n_114),
.B2(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_53),
.A2(n_56),
.B1(n_278),
.B2(n_279),
.Y(n_277)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_59),
.A2(n_60),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_64),
.B2(n_65),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_61),
.A2(n_64),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_61),
.A2(n_64),
.B1(n_112),
.B2(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_61),
.A2(n_64),
.B1(n_240),
.B2(n_256),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_61),
.A2(n_62),
.B1(n_64),
.B2(n_301),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_65),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_67),
.A2(n_68),
.B1(n_69),
.B2(n_326),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_69),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_322),
.B(n_328),
.Y(n_72)
);

OAI321xp33_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_291),
.A3(n_314),
.B1(n_320),
.B2(n_321),
.C(n_330),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_270),
.B(n_290),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_246),
.B(n_269),
.Y(n_75)
);

O2A1O1Ixp33_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_138),
.B(n_222),
.C(n_245),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_123),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_78),
.B(n_123),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_107),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_91),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_80),
.B(n_91),
.C(n_107),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_87),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_81),
.B(n_87),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_84),
.B1(n_85),
.B2(n_86),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_82),
.A2(n_84),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_82),
.A2(n_83),
.B1(n_120),
.B2(n_137),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_82),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_82),
.A2(n_121),
.B1(n_148),
.B2(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_82),
.A2(n_85),
.B1(n_151),
.B2(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_82),
.A2(n_121),
.B1(n_137),
.B2(n_181),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_82),
.A2(n_86),
.B1(n_121),
.B2(n_231),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_82),
.A2(n_121),
.B(n_231),
.Y(n_264)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_85),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_85),
.B(n_104),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_96),
.C(n_102),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_92),
.A2(n_93),
.B1(n_96),
.B2(n_97),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_98),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_102),
.B(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_105),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g107 ( 
.A(n_108),
.B(n_116),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_113),
.B2(n_115),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_109),
.B(n_115),
.C(n_116),
.Y(n_225)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_113),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_119),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_119),
.Y(n_127)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_126),
.C(n_128),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_124),
.B(n_219),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_126),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_134),
.C(n_135),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_130),
.B(n_207),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_134),
.A2(n_135),
.B1(n_136),
.B2(n_208),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_134),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_221),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_216),
.B(n_220),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_202),
.B(n_215),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_183),
.B(n_201),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_171),
.B(n_182),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_160),
.B(n_170),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_152),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_145),
.B(n_152),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_149),
.B2(n_150),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_156),
.B2(n_157),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_154),
.B(n_156),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_165),
.B(n_169),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_162),
.B(n_164),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_168),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_172),
.B(n_173),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_180),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_175),
.B(n_178),
.C(n_180),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_185),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_191),
.B1(n_199),
.B2(n_200),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_186),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_188),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_190),
.Y(n_194)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_191),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_195),
.B1(n_196),
.B2(n_198),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_192),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_195),
.B(n_198),
.C(n_199),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_203),
.B(n_204),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_206),
.B1(n_209),
.B2(n_210),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_212),
.C(n_213),
.Y(n_217)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_213),
.B2(n_214),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_211),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_212),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_217),
.B(n_218),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_223),
.B(n_224),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_227),
.B2(n_244),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_225),
.Y(n_244)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_234),
.B2(n_235),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_228),
.B(n_235),
.C(n_244),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_232),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_230),
.B(n_232),
.Y(n_252)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_236),
.B(n_238),
.C(n_243),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_241),
.B2(n_243),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_241),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_242),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_247),
.B(n_248),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_268),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_261),
.B2(n_262),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_262),
.C(n_268),
.Y(n_271)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_252),
.B(n_254),
.C(n_258),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_255),
.B1(n_257),
.B2(n_258),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_256),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_258),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_260),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_265),
.B2(n_267),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_263),
.A2(n_264),
.B1(n_284),
.B2(n_285),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_264),
.B(n_265),
.Y(n_282)
);

AOI21xp33_ASAP7_75t_L g305 ( 
.A1(n_264),
.A2(n_282),
.B(n_285),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_265),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_271),
.B(n_272),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_288),
.B2(n_289),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_281),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_275),
.B(n_281),
.C(n_289),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_277),
.B(n_280),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_276),
.B(n_277),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_279),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_293),
.C(n_304),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_280),
.A2(n_293),
.B1(n_294),
.B2(n_319),
.Y(n_318)
);

CKINVDCx14_ASAP7_75t_R g319 ( 
.A(n_280),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_285),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_287),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_288),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_306),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_292),
.B(n_306),
.Y(n_321)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_295),
.A2(n_300),
.B1(n_302),
.B2(n_303),
.Y(n_294)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_295),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_297),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_299),
.C(n_300),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_300),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_300),
.A2(n_303),
.B1(n_308),
.B2(n_309),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_300),
.B(n_308),
.C(n_313),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_304),
.A2(n_305),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_305),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_313),
.Y(n_306)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_311),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_315),
.B(n_316),
.Y(n_320)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_324),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_325),
.Y(n_327)
);


endmodule