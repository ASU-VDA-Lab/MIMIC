module fake_jpeg_21816_n_103 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_103);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_103;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx2_ASAP7_75t_L g11 ( 
.A(n_0),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx10_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_5),
.Y(n_17)
);

INVx13_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_23),
.Y(n_24)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_23),
.Y(n_25)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_27),
.Y(n_38)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_28),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_31),
.Y(n_35)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_31),
.B(n_13),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_34),
.B(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_29),
.B(n_13),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_27),
.B(n_22),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_22),
.Y(n_48)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_29),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_42),
.A2(n_43),
.B(n_44),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_29),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_35),
.A2(n_11),
.B(n_22),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_45),
.B(n_48),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_35),
.A2(n_11),
.B1(n_30),
.B2(n_18),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_46),
.A2(n_49),
.B1(n_51),
.B2(n_12),
.Y(n_66)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_40),
.A2(n_18),
.B1(n_21),
.B2(n_20),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_53),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_40),
.A2(n_20),
.B1(n_21),
.B2(n_17),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_37),
.B(n_38),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_57),
.C(n_58),
.Y(n_64)
);

O2A1O1Ixp33_ASAP7_75t_L g55 ( 
.A1(n_33),
.A2(n_19),
.B(n_25),
.C(n_28),
.Y(n_55)
);

OAI21xp33_ASAP7_75t_L g63 ( 
.A1(n_55),
.A2(n_18),
.B(n_19),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_15),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_14),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_15),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_28),
.C(n_25),
.Y(n_61)
);

FAx1_ASAP7_75t_SL g71 ( 
.A(n_61),
.B(n_68),
.CI(n_42),
.CON(n_71),
.SN(n_71)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_14),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_43),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_63),
.B(n_66),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_36),
.C(n_24),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_51),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_71),
.A2(n_75),
.B(n_77),
.Y(n_84)
);

A2O1A1O1Ixp25_ASAP7_75t_L g82 ( 
.A1(n_72),
.A2(n_62),
.B(n_67),
.C(n_68),
.D(n_63),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_47),
.Y(n_74)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_74),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_52),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

AO221x1_ASAP7_75t_L g86 ( 
.A1(n_76),
.A2(n_79),
.B1(n_58),
.B2(n_59),
.C(n_43),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_45),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_78),
.A2(n_61),
.B(n_55),
.Y(n_85)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_SL g90 ( 
.A1(n_80),
.A2(n_86),
.B(n_26),
.C(n_16),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_85),
.C(n_17),
.Y(n_88)
);

NAND3xp33_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_78),
.C(n_71),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_83),
.A2(n_73),
.B(n_71),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_87),
.A2(n_4),
.B(n_7),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_89),
.C(n_6),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_84),
.A2(n_16),
.B(n_12),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_90),
.A2(n_91),
.B(n_2),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_81),
.A2(n_0),
.B(n_2),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_93),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_0),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_9),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_95),
.A2(n_7),
.B1(n_9),
.B2(n_2),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_3),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_3),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_100),
.C(n_97),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_98),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_26),
.Y(n_103)
);


endmodule