module fake_jpeg_5122_n_295 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_295);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_295;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx2_ASAP7_75t_SL g17 ( 
.A(n_14),
.Y(n_17)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx13_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_1),
.Y(n_35)
);

INVx11_ASAP7_75t_SL g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_17),
.B(n_8),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_38),
.B(n_46),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_17),
.B(n_7),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_42),
.B(n_45),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_17),
.B(n_9),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_24),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_50),
.A2(n_52),
.B1(n_55),
.B2(n_21),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_51),
.Y(n_64)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_53),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_57),
.B(n_70),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_59),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_63),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_40),
.B(n_24),
.Y(n_65)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_67),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_68),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_71),
.B(n_79),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_38),
.B(n_37),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_73),
.B(n_75),
.Y(n_105)
);

INVx3_ASAP7_75t_SL g74 ( 
.A(n_53),
.Y(n_74)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_74),
.B(n_95),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_42),
.B(n_37),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_45),
.B(n_26),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_76),
.B(n_91),
.Y(n_113)
);

INVx5_ASAP7_75t_SL g77 ( 
.A(n_46),
.Y(n_77)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_77),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_78),
.Y(n_108)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_80),
.B(n_83),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_47),
.B(n_24),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_82),
.B(n_85),
.Y(n_116)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_84),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_47),
.B(n_28),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_86),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_43),
.B(n_31),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_87),
.B(n_88),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_43),
.B(n_28),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_48),
.B(n_22),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_89),
.B(n_90),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_48),
.B(n_22),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_49),
.B(n_30),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_49),
.B(n_30),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_92),
.B(n_97),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_50),
.A2(n_29),
.B1(n_21),
.B2(n_17),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_94),
.A2(n_32),
.B1(n_20),
.B2(n_35),
.Y(n_120)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_41),
.B(n_23),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_50),
.A2(n_21),
.B1(n_29),
.B2(n_26),
.Y(n_98)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_98),
.A2(n_100),
.B(n_35),
.C(n_27),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_39),
.B(n_31),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_34),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_81),
.A2(n_32),
.B1(n_23),
.B2(n_20),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_110),
.A2(n_61),
.B1(n_60),
.B2(n_79),
.Y(n_144)
);

AND2x2_ASAP7_75t_SL g111 ( 
.A(n_74),
.B(n_53),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_111),
.A2(n_123),
.B(n_124),
.Y(n_156)
);

NOR2x1_ASAP7_75t_L g119 ( 
.A(n_76),
.B(n_53),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_119),
.B(n_128),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_120),
.A2(n_122),
.B1(n_96),
.B2(n_81),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_94),
.A2(n_78),
.B1(n_98),
.B2(n_93),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_27),
.Y(n_123)
);

MAJx2_ASAP7_75t_L g124 ( 
.A(n_77),
.B(n_51),
.C(n_27),
.Y(n_124)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_72),
.A2(n_27),
.B(n_51),
.C(n_33),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_L g132 ( 
.A1(n_93),
.A2(n_34),
.B1(n_19),
.B2(n_33),
.Y(n_132)
);

OAI22xp33_ASAP7_75t_L g154 ( 
.A1(n_132),
.A2(n_58),
.B1(n_62),
.B2(n_56),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_124),
.B(n_33),
.Y(n_133)
);

OAI21xp33_ASAP7_75t_L g190 ( 
.A1(n_133),
.A2(n_136),
.B(n_160),
.Y(n_190)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_135),
.B(n_139),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_105),
.B(n_96),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_141),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_70),
.Y(n_138)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_138),
.Y(n_197)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_106),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_146),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_130),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_57),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_142),
.B(n_145),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_105),
.B(n_61),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_153),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_144),
.A2(n_154),
.B1(n_104),
.B2(n_131),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_113),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_105),
.B(n_83),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_56),
.Y(n_147)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_147),
.Y(n_185)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_106),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_150),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_126),
.Y(n_149)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_149),
.Y(n_179)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_126),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_108),
.A2(n_60),
.B1(n_64),
.B2(n_99),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_151),
.A2(n_158),
.B1(n_166),
.B2(n_104),
.Y(n_181)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_111),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_159),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_51),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_113),
.B(n_34),
.Y(n_155)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_68),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_157),
.B(n_162),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_122),
.A2(n_58),
.B1(n_80),
.B2(n_71),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_113),
.B(n_11),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_124),
.B(n_33),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_112),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_161),
.B(n_165),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_130),
.B(n_0),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_34),
.Y(n_163)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_163),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_120),
.B(n_1),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_119),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_114),
.B(n_86),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_108),
.A2(n_69),
.B1(n_66),
.B2(n_3),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_156),
.B(n_111),
.C(n_116),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_169),
.B(n_176),
.C(n_196),
.Y(n_204)
);

NOR4xp25_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_119),
.C(n_116),
.D(n_128),
.Y(n_171)
);

NAND3xp33_ASAP7_75t_L g222 ( 
.A(n_171),
.B(n_12),
.C(n_14),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_175),
.B(n_180),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_156),
.B(n_141),
.C(n_153),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_177),
.B(n_182),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_128),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_178),
.B(n_191),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_181),
.A2(n_187),
.B1(n_104),
.B2(n_131),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_133),
.B(n_114),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_133),
.B(n_160),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_147),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_137),
.B(n_127),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_134),
.A2(n_102),
.B(n_112),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_192),
.A2(n_195),
.B(n_162),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_193),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_134),
.A2(n_136),
.B(n_146),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_102),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_155),
.B(n_127),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_159),
.C(n_103),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_183),
.A2(n_160),
.B(n_145),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_202),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_212),
.Y(n_227)
);

XNOR2x2_ASAP7_75t_SL g202 ( 
.A(n_190),
.B(n_135),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_172),
.A2(n_152),
.B1(n_140),
.B2(n_164),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_205),
.A2(n_206),
.B1(n_208),
.B2(n_213),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_167),
.A2(n_166),
.B1(n_158),
.B2(n_144),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_182),
.A2(n_138),
.B(n_142),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_207),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g209 ( 
.A1(n_179),
.A2(n_161),
.B1(n_148),
.B2(n_139),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_185),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_167),
.A2(n_173),
.B1(n_188),
.B2(n_189),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_184),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_214),
.B(n_217),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_218),
.C(n_220),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_168),
.A2(n_127),
.B(n_66),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_216),
.B(n_193),
.Y(n_240)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_170),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_176),
.B(n_103),
.C(n_109),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_179),
.B(n_115),
.Y(n_219)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_219),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_178),
.B(n_117),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_181),
.A2(n_115),
.B1(n_118),
.B2(n_109),
.Y(n_221)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_221),
.Y(n_233)
);

NAND3xp33_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_189),
.C(n_188),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_200),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_224),
.B(n_231),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_204),
.B(n_169),
.C(n_173),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_226),
.B(n_236),
.C(n_242),
.Y(n_245)
);

OAI321xp33_ASAP7_75t_L g229 ( 
.A1(n_207),
.A2(n_192),
.A3(n_195),
.B1(n_194),
.B2(n_177),
.C(n_191),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_230),
.Y(n_250)
);

OAI321xp33_ASAP7_75t_L g230 ( 
.A1(n_202),
.A2(n_174),
.A3(n_196),
.B1(n_198),
.B2(n_197),
.C(n_186),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_213),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_234),
.A2(n_237),
.B(n_216),
.Y(n_246)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_205),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_212),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_174),
.C(n_185),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_238),
.A2(n_203),
.B1(n_211),
.B2(n_199),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_210),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_214),
.B(n_217),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_241),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_125),
.C(n_115),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_227),
.B(n_202),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_247),
.C(n_249),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_246),
.A2(n_129),
.B(n_10),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_227),
.B(n_225),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_210),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_248),
.B(n_223),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_218),
.C(n_215),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_239),
.A2(n_206),
.B1(n_203),
.B2(n_211),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_251),
.A2(n_254),
.B1(n_118),
.B2(n_129),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_253),
.B(n_240),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_255),
.A2(n_232),
.B(n_223),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_236),
.B(n_201),
.C(n_125),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_256),
.B(n_242),
.C(n_239),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_264),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_258),
.B(n_263),
.Y(n_269)
);

NOR3xp33_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_231),
.C(n_233),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_260),
.A2(n_266),
.B(n_267),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_261),
.A2(n_245),
.B(n_10),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_118),
.C(n_131),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_244),
.B(n_228),
.Y(n_263)
);

MAJx2_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_232),
.C(n_11),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_265),
.B(n_243),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_252),
.A2(n_1),
.B(n_2),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_268),
.B(n_275),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_264),
.A2(n_247),
.B1(n_255),
.B2(n_256),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_270),
.A2(n_274),
.B(n_4),
.Y(n_283)
);

A2O1A1O1Ixp25_ASAP7_75t_L g284 ( 
.A1(n_271),
.A2(n_273),
.B(n_4),
.C(n_6),
.D(n_9),
.Y(n_284)
);

NOR2x1_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_258),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_259),
.A2(n_245),
.B(n_10),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_272),
.B(n_266),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_279),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_269),
.B(n_1),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_273),
.A2(n_2),
.B(n_3),
.Y(n_280)
);

NOR3xp33_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_282),
.C(n_284),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_268),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_281),
.B(n_283),
.Y(n_286)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_4),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_276),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_287),
.B(n_289),
.C(n_6),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_276),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_290),
.A2(n_291),
.B(n_292),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_286),
.B(n_6),
.C(n_9),
.Y(n_291)
);

FAx1_ASAP7_75t_SL g292 ( 
.A(n_285),
.B(n_14),
.CI(n_15),
.CON(n_292),
.SN(n_292)
);

AO21x1_ASAP7_75t_L g293 ( 
.A1(n_292),
.A2(n_288),
.B(n_2),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_293),
.B(n_294),
.Y(n_295)
);


endmodule