module real_jpeg_27135_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_288;
wire n_166;
wire n_176;
wire n_215;
wire n_292;
wire n_300;
wire n_221;
wire n_249;
wire n_286;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_299;
wire n_173;
wire n_255;
wire n_115;
wire n_243;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_296;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_278;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_295;
wire n_167;
wire n_179;
wire n_216;
wire n_202;
wire n_133;
wire n_213;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;
wire n_16;

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_0),
.A2(n_87),
.B(n_88),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_0),
.B(n_54),
.Y(n_87)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_0),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_0),
.B(n_124),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_0),
.B(n_232),
.Y(n_237)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_2),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_2),
.A2(n_46),
.B1(n_50),
.B2(n_70),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_2),
.A2(n_30),
.B1(n_31),
.B2(n_70),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_2),
.A2(n_52),
.B1(n_54),
.B2(n_70),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_4),
.A2(n_30),
.B1(n_31),
.B2(n_138),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_4),
.Y(n_138)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_4),
.A2(n_24),
.B1(n_25),
.B2(n_138),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_4),
.A2(n_46),
.B1(n_50),
.B2(n_138),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_4),
.A2(n_52),
.B1(n_54),
.B2(n_138),
.Y(n_232)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_6),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_29)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_6),
.A2(n_24),
.B1(n_25),
.B2(n_32),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_6),
.A2(n_32),
.B1(n_46),
.B2(n_50),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_6),
.A2(n_32),
.B1(n_52),
.B2(n_54),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g37 ( 
.A1(n_7),
.A2(n_30),
.B(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_7),
.B(n_30),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_7),
.A2(n_46),
.B1(n_50),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_7),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_7),
.A2(n_52),
.B1(n_54),
.B2(n_58),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_7),
.A2(n_24),
.B1(n_25),
.B2(n_58),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_7),
.B(n_21),
.Y(n_188)
);

AOI21xp33_ASAP7_75t_SL g198 ( 
.A1(n_7),
.A2(n_10),
.B(n_46),
.Y(n_198)
);

AOI21xp33_ASAP7_75t_L g223 ( 
.A1(n_7),
.A2(n_49),
.B(n_52),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_7),
.B(n_67),
.Y(n_227)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_10),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_10),
.A2(n_46),
.B1(n_50),
.B2(n_66),
.Y(n_67)
);

INVx11_ASAP7_75t_SL g53 ( 
.A(n_11),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_111),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_110),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_93),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_16),
.B(n_93),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_74),
.C(n_82),
.Y(n_16)
);

FAx1_ASAP7_75t_SL g144 ( 
.A(n_17),
.B(n_74),
.CI(n_82),
.CON(n_144),
.SN(n_144)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_19),
.B1(n_39),
.B2(n_40),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_18),
.A2(n_19),
.B1(n_95),
.B2(n_96),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_19),
.B(n_41),
.C(n_60),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_33),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_20),
.B(n_134),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_28),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_21),
.B(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

A2O1A1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_22),
.A2(n_23),
.B(n_30),
.C(n_36),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_22),
.A2(n_35),
.B(n_37),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_22),
.A2(n_98),
.B(n_99),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_22),
.B(n_137),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_22)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_24),
.B(n_27),
.Y(n_174)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

O2A1O1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_25),
.A2(n_62),
.B(n_63),
.C(n_67),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_25),
.B(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_25),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_L g197 ( 
.A1(n_25),
.A2(n_58),
.B(n_62),
.C(n_198),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_29),
.B(n_35),
.Y(n_100)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_34),
.B(n_159),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_35),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_36),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_37),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_38),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_59),
.B2(n_60),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_41),
.B(n_158),
.C(n_160),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_41),
.A2(n_42),
.B1(n_160),
.B2(n_161),
.Y(n_182)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_42),
.B(n_103),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_55),
.B(n_56),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_43),
.A2(n_90),
.B(n_91),
.Y(n_89)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_44),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_44),
.B(n_57),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_44),
.B(n_205),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_51),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_45)
);

INVx4_ASAP7_75t_SL g50 ( 
.A(n_46),
.Y(n_50)
);

A2O1A1Ixp33_ASAP7_75t_L g222 ( 
.A1(n_46),
.A2(n_48),
.B(n_58),
.C(n_223),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_48),
.A2(n_49),
.B1(n_52),
.B2(n_54),
.Y(n_51)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_51),
.B(n_57),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_51),
.B(n_81),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_51),
.B(n_205),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_52),
.Y(n_54)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_54),
.B(n_247),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_55),
.A2(n_80),
.B(n_90),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_55),
.B(n_58),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_58),
.B(n_178),
.Y(n_247)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_68),
.B(n_71),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_61),
.B(n_73),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_61),
.B(n_106),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_61),
.B(n_163),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_61),
.Y(n_278)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_67),
.B(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g75 ( 
.A1(n_69),
.A2(n_76),
.B(n_77),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_71),
.B(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_72),
.B(n_171),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_74),
.A2(n_75),
.B(n_78),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_105),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_76),
.A2(n_105),
.B(n_278),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_77),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_77),
.B(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_79),
.B(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_80),
.B(n_204),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_86),
.B(n_92),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_83),
.A2(n_84),
.B1(n_141),
.B2(n_142),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_89),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_85),
.A2(n_86),
.B1(n_92),
.B2(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_85),
.A2(n_86),
.B1(n_197),
.B2(n_199),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_85),
.A2(n_86),
.B1(n_89),
.B2(n_292),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_86),
.B(n_197),
.Y(n_215)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_87),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_87),
.B(n_88),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_87),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_88),
.B(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_89),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_91),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_91),
.B(n_214),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_92),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_109),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_101),
.B1(n_102),
.B2(n_108),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_97),
.Y(n_108)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_100),
.B(n_159),
.Y(n_275)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_107),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_104),
.B(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_112),
.A2(n_145),
.B(n_301),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_144),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_113),
.B(n_144),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_139),
.C(n_140),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_114),
.A2(n_115),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_127),
.C(n_130),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_116),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_126),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_117),
.B(n_126),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_121),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_118),
.B(n_231),
.Y(n_230)
);

INVx5_ASAP7_75t_SL g178 ( 
.A(n_119),
.Y(n_178)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_121),
.A2(n_153),
.B(n_178),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_122),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_122),
.B(n_236),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_125),
.Y(n_122)
);

INVxp33_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_125),
.A2(n_153),
.B(n_154),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_127),
.A2(n_130),
.B1(n_131),
.B2(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_127),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_129),
.B(n_162),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_139),
.B(n_140),
.Y(n_299)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx24_ASAP7_75t_SL g303 ( 
.A(n_144),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_295),
.B(n_300),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_282),
.B(n_294),
.Y(n_146)
);

O2A1O1Ixp33_ASAP7_75t_SL g147 ( 
.A1(n_148),
.A2(n_191),
.B(n_265),
.C(n_281),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_179),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_149),
.B(n_179),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_164),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_157),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_151),
.B(n_157),
.C(n_164),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_155),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_152),
.B(n_155),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_154),
.B(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_154),
.B(n_231),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_156),
.B(n_204),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_165),
.B(n_172),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_169),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_166),
.B(n_169),
.C(n_172),
.Y(n_279)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_177),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_177),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_183),
.C(n_185),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_180),
.A2(n_181),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_183),
.A2(n_184),
.B1(n_185),
.B2(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_185),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.C(n_189),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_209),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_189),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_190),
.B(n_237),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_192),
.B(n_264),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_257),
.B(n_263),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_216),
.B(n_256),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_206),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_195),
.B(n_206),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_200),
.C(n_202),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_196),
.B(n_254),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_197),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_200),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_254)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_211),
.B2(n_212),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_207),
.B(n_213),
.C(n_215),
.Y(n_258)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_215),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_251),
.B(n_255),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_233),
.B(n_250),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_224),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_219),
.B(n_224),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_222),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_220),
.A2(n_221),
.B1(n_222),
.B2(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_222),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_230),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_228),
.B2(n_229),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_229),
.C(n_230),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_240),
.B(n_249),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_238),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_235),
.B(n_238),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_244),
.B(n_248),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_242),
.B(n_243),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_252),
.B(n_253),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_258),
.B(n_259),
.Y(n_263)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_266),
.B(n_267),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_279),
.B2(n_280),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_270),
.B(n_271),
.C(n_280),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_272),
.B(n_275),
.C(n_276),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_276),
.B2(n_277),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_279),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_283),
.B(n_284),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_293),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_290),
.B2(n_291),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_291),
.C(n_293),
.Y(n_296)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_296),
.B(n_297),
.Y(n_300)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);


endmodule