module fake_jpeg_10420_n_239 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_239);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_239;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_171;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_36),
.Y(n_56)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_33),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_19),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_37),
.B(n_40),
.Y(n_58)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_33),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_26),
.Y(n_59)
);

AOI21xp33_ASAP7_75t_L g42 ( 
.A1(n_17),
.A2(n_0),
.B(n_1),
.Y(n_42)
);

AND2x2_ASAP7_75t_SL g53 ( 
.A(n_42),
.B(n_16),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_35),
.A2(n_20),
.B1(n_28),
.B2(n_29),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_43),
.A2(n_46),
.B1(n_51),
.B2(n_54),
.Y(n_63)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_44),
.Y(n_80)
);

BUFx4f_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_35),
.A2(n_20),
.B1(n_28),
.B2(n_29),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_41),
.A2(n_17),
.B1(n_21),
.B2(n_16),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_47),
.A2(n_50),
.B1(n_60),
.B2(n_34),
.Y(n_82)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_52),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_41),
.A2(n_38),
.B1(n_35),
.B2(n_34),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_35),
.A2(n_38),
.B1(n_36),
.B2(n_40),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_53),
.A2(n_37),
.B(n_2),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_35),
.A2(n_25),
.B1(n_21),
.B2(n_24),
.Y(n_54)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_41),
.A2(n_34),
.B1(n_36),
.B2(n_40),
.Y(n_60)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_39),
.Y(n_67)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_64),
.B(n_68),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_55),
.A2(n_36),
.B1(n_40),
.B2(n_25),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_65),
.A2(n_70),
.B1(n_84),
.B2(n_88),
.Y(n_106)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_57),
.B(n_27),
.Y(n_69)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_59),
.A2(n_41),
.B1(n_27),
.B2(n_24),
.Y(n_70)
);

FAx1_ASAP7_75t_SL g72 ( 
.A(n_53),
.B(n_36),
.CI(n_33),
.CON(n_72),
.SN(n_72)
);

NAND2xp33_ASAP7_75t_SL g107 ( 
.A(n_72),
.B(n_31),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_75),
.Y(n_97)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_31),
.Y(n_77)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

BUFx10_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_31),
.Y(n_79)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_82),
.A2(n_50),
.B1(n_44),
.B2(n_48),
.Y(n_94)
);

AND2x2_ASAP7_75t_SL g83 ( 
.A(n_53),
.B(n_34),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_89),
.C(n_0),
.Y(n_110)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_31),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_26),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_60),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_44),
.A2(n_37),
.B1(n_26),
.B2(n_32),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_93),
.B(n_66),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_94),
.A2(n_98),
.B1(n_101),
.B2(n_113),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_82),
.A2(n_52),
.B1(n_58),
.B2(n_61),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_62),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_104),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_84),
.A2(n_61),
.B1(n_39),
.B2(n_22),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_73),
.B(n_32),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_107),
.A2(n_110),
.B(n_71),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_83),
.B(n_30),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_108),
.B(n_114),
.Y(n_120)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_109),
.Y(n_124)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_112),
.Y(n_138)
);

O2A1O1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_87),
.A2(n_39),
.B(n_49),
.C(n_30),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_83),
.B(n_0),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_114),
.A2(n_78),
.B(n_39),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_92),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_115),
.B(n_118),
.Y(n_165)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_120),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_92),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_121),
.B(n_123),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_93),
.B(n_89),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_125),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_101),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_72),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_104),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_126),
.A2(n_128),
.B(n_130),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_72),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_129),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_110),
.A2(n_98),
.B(n_111),
.Y(n_130)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_131),
.A2(n_135),
.B1(n_141),
.B2(n_64),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_94),
.B(n_71),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_140),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_106),
.A2(n_63),
.B1(n_75),
.B2(n_76),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_133),
.A2(n_111),
.B1(n_91),
.B2(n_112),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_109),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_134),
.B(n_137),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_97),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_78),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_96),
.B(n_80),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_96),
.B(n_80),
.Y(n_139)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_139),
.Y(n_147)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_100),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_129),
.B(n_91),
.C(n_105),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_142),
.B(n_162),
.C(n_130),
.Y(n_170)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_143),
.B(n_145),
.Y(n_168)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_132),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_146),
.B(n_151),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_150),
.A2(n_161),
.B1(n_115),
.B2(n_121),
.Y(n_176)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_135),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_152),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_102),
.Y(n_180)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_117),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_157),
.Y(n_167)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_122),
.B(n_90),
.Y(n_159)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_136),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_140),
.A2(n_95),
.B1(n_68),
.B2(n_81),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_102),
.C(n_85),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_126),
.Y(n_163)
);

OR2x2_ASAP7_75t_SL g166 ( 
.A(n_160),
.B(n_127),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_166),
.B(n_183),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_184),
.C(n_162),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_164),
.B(n_125),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_165),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_173),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_158),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_156),
.A2(n_153),
.B(n_155),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_176),
.A2(n_153),
.B1(n_148),
.B2(n_144),
.Y(n_195)
);

BUFx12_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

INVx11_ASAP7_75t_L g198 ( 
.A(n_177),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_143),
.B(n_120),
.Y(n_178)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_178),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_180),
.B(n_182),
.Y(n_197)
);

INVx13_ASAP7_75t_L g181 ( 
.A(n_147),
.Y(n_181)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_181),
.Y(n_191)
);

AOI32xp33_ASAP7_75t_L g182 ( 
.A1(n_159),
.A2(n_131),
.A3(n_138),
.B1(n_102),
.B2(n_124),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_95),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_85),
.C(n_138),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_150),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_185),
.B(n_85),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_186),
.B(n_167),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_169),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_185),
.A2(n_146),
.B1(n_145),
.B2(n_157),
.Y(n_189)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_149),
.C(n_156),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_194),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_144),
.C(n_178),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_195),
.A2(n_23),
.B1(n_22),
.B2(n_39),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_142),
.C(n_154),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_196),
.B(n_180),
.Y(n_203)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_167),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_186),
.C(n_196),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_198),
.A2(n_174),
.B1(n_181),
.B2(n_179),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_202),
.A2(n_200),
.B1(n_191),
.B2(n_188),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_203),
.B(n_207),
.Y(n_210)
);

NOR3xp33_ASAP7_75t_SL g205 ( 
.A(n_193),
.B(n_168),
.C(n_171),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_205),
.B(n_190),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_179),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_197),
.B(n_177),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_194),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_199),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_215),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_212),
.B(n_214),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_213),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_207),
.C(n_201),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_216),
.A2(n_23),
.B1(n_39),
.B2(n_4),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_206),
.A2(n_197),
.B1(n_191),
.B2(n_188),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_217),
.B(n_14),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_208),
.B(n_189),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_218),
.B(n_14),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_222),
.A2(n_224),
.B1(n_3),
.B2(n_5),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_223),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_221),
.A2(n_210),
.B1(n_215),
.B2(n_13),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_225),
.B(n_6),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_220),
.B(n_210),
.C(n_12),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_226),
.B(n_227),
.C(n_5),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_220),
.B(n_219),
.C(n_222),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_228),
.B(n_229),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_226),
.B(n_3),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_230),
.B(n_231),
.Y(n_234)
);

AOI322xp5_ASAP7_75t_L g235 ( 
.A1(n_233),
.A2(n_6),
.A3(n_7),
.B1(n_9),
.B2(n_39),
.C1(n_224),
.C2(n_187),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_235),
.Y(n_236)
);

OAI21x1_ASAP7_75t_L g237 ( 
.A1(n_236),
.A2(n_233),
.B(n_234),
.Y(n_237)
);

BUFx24_ASAP7_75t_SL g238 ( 
.A(n_237),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_238),
.B(n_232),
.Y(n_239)
);


endmodule