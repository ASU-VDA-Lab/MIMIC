module fake_netlist_5_1947_n_2927 (n_137, n_294, n_318, n_82, n_194, n_316, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_127, n_75, n_235, n_226, n_74, n_57, n_353, n_351, n_367, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_17, n_254, n_33, n_23, n_302, n_265, n_293, n_244, n_47, n_173, n_198, n_247, n_314, n_368, n_8, n_321, n_292, n_100, n_212, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_341, n_204, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_325, n_132, n_90, n_101, n_281, n_240, n_189, n_220, n_291, n_231, n_257, n_31, n_13, n_152, n_317, n_9, n_323, n_195, n_42, n_356, n_227, n_45, n_271, n_94, n_335, n_123, n_167, n_234, n_343, n_308, n_267, n_297, n_156, n_5, n_225, n_219, n_157, n_131, n_192, n_223, n_158, n_138, n_264, n_109, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_347, n_169, n_59, n_255, n_215, n_350, n_196, n_211, n_218, n_181, n_3, n_290, n_221, n_178, n_287, n_344, n_72, n_104, n_41, n_56, n_141, n_355, n_15, n_336, n_145, n_48, n_50, n_337, n_313, n_88, n_216, n_168, n_164, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_342, n_98, n_361, n_363, n_197, n_107, n_69, n_236, n_1, n_249, n_304, n_329, n_203, n_274, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_333, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_345, n_210, n_365, n_91, n_176, n_182, n_143, n_83, n_354, n_237, n_180, n_340, n_207, n_37, n_346, n_229, n_108, n_66, n_177, n_60, n_16, n_0, n_58, n_18, n_359, n_117, n_326, n_233, n_205, n_366, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_352, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_334, n_175, n_262, n_238, n_99, n_319, n_364, n_20, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_324, n_199, n_187, n_32, n_103, n_348, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_2927);

input n_137;
input n_294;
input n_318;
input n_82;
input n_194;
input n_316;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_353;
input n_351;
input n_367;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_17;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_368;
input n_8;
input n_321;
input n_292;
input n_100;
input n_212;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_341;
input n_204;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_31;
input n_13;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_356;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_167;
input n_234;
input n_343;
input n_308;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_158;
input n_138;
input n_264;
input n_109;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_350;
input n_196;
input n_211;
input n_218;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_287;
input n_344;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_355;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_313;
input n_88;
input n_216;
input n_168;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_342;
input n_98;
input n_361;
input n_363;
input n_197;
input n_107;
input n_69;
input n_236;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_345;
input n_210;
input n_365;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_354;
input n_237;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_16;
input n_0;
input n_58;
input n_18;
input n_359;
input n_117;
input n_326;
input n_233;
input n_205;
input n_366;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_334;
input n_175;
input n_262;
input n_238;
input n_99;
input n_319;
input n_364;
input n_20;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_324;
input n_199;
input n_187;
input n_32;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_2927;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_611;
wire n_2756;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_2739;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_469;
wire n_1508;
wire n_2771;
wire n_785;
wire n_549;
wire n_2617;
wire n_2200;
wire n_532;
wire n_1161;
wire n_1859;
wire n_2746;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_667;
wire n_2899;
wire n_790;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_2395;
wire n_880;
wire n_544;
wire n_1007;
wire n_2369;
wire n_552;
wire n_1528;
wire n_2683;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_2520;
wire n_2821;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_2568;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_2391;
wire n_1021;
wire n_1960;
wire n_2843;
wire n_2185;
wire n_551;
wire n_2143;
wire n_2853;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_2487;
wire n_1353;
wire n_800;
wire n_1347;
wire n_2495;
wire n_2880;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_2389;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_447;
wire n_2001;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_2486;
wire n_1806;
wire n_516;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2538;
wire n_2024;
wire n_2530;
wire n_1696;
wire n_2483;
wire n_1118;
wire n_755;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_1860;
wire n_2543;
wire n_1359;
wire n_530;
wire n_1728;
wire n_1107;
wire n_2076;
wire n_556;
wire n_2031;
wire n_2482;
wire n_2677;
wire n_1230;
wire n_668;
wire n_375;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_2770;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_1705;
wire n_659;
wire n_2584;
wire n_1257;
wire n_2639;
wire n_1182;
wire n_1698;
wire n_579;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2193;
wire n_2052;
wire n_2058;
wire n_2458;
wire n_2478;
wire n_2761;
wire n_731;
wire n_371;
wire n_1483;
wire n_2888;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_2537;
wire n_569;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_2515;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2466;
wire n_2635;
wire n_2652;
wire n_2715;
wire n_2085;
wire n_1669;
wire n_2566;
wire n_370;
wire n_976;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_2149;
wire n_1078;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_775;
wire n_2651;
wire n_600;
wire n_1484;
wire n_2071;
wire n_2561;
wire n_1374;
wire n_1328;
wire n_2643;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_2408;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_2384;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_2663;
wire n_1394;
wire n_436;
wire n_2659;
wire n_1414;
wire n_1216;
wire n_580;
wire n_2693;
wire n_1040;
wire n_2202;
wire n_2648;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_926;
wire n_2180;
wire n_2249;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2632;
wire n_2276;
wire n_422;
wire n_1070;
wire n_777;
wire n_1547;
wire n_475;
wire n_2089;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_1801;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_2908;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_2915;
wire n_528;
wire n_2300;
wire n_2791;
wire n_1796;
wire n_2551;
wire n_680;
wire n_1587;
wire n_1473;
wire n_2682;
wire n_395;
wire n_901;
wire n_553;
wire n_2432;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_2714;
wire n_1748;
wire n_1672;
wire n_2506;
wire n_675;
wire n_2699;
wire n_888;
wire n_1880;
wire n_2769;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_637;
wire n_2615;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_468;
wire n_2753;
wire n_464;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_2859;
wire n_2842;
wire n_1075;
wire n_1836;
wire n_2868;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2863;
wire n_2072;
wire n_2738;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_2833;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_2684;
wire n_2712;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_2855;
wire n_2713;
wire n_2644;
wire n_2700;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_2730;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_488;
wire n_736;
wire n_892;
wire n_2688;
wire n_1000;
wire n_1202;
wire n_2750;
wire n_2620;
wire n_1278;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_593;
wire n_2258;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_2784;
wire n_2919;
wire n_1053;
wire n_1224;
wire n_2865;
wire n_2557;
wire n_1926;
wire n_2706;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2757;
wire n_2152;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_2590;
wire n_2776;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2862;
wire n_2175;
wire n_2921;
wire n_2720;
wire n_2324;
wire n_1854;
wire n_2674;
wire n_2606;
wire n_1565;
wire n_2828;
wire n_1809;
wire n_1856;
wire n_647;
wire n_407;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_857;
wire n_832;
wire n_2305;
wire n_2636;
wire n_2450;
wire n_1319;
wire n_561;
wire n_2379;
wire n_2616;
wire n_2911;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_2759;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_2462;
wire n_2514;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_404;
wire n_2798;
wire n_2331;
wire n_2293;
wire n_686;
wire n_2837;
wire n_847;
wire n_1393;
wire n_2319;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_2762;
wire n_558;
wire n_2808;
wire n_702;
wire n_1276;
wire n_2548;
wire n_822;
wire n_1412;
wire n_2676;
wire n_1709;
wire n_2679;
wire n_2108;
wire n_728;
wire n_1162;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_2767;
wire n_2777;
wire n_2603;
wire n_1884;
wire n_2434;
wire n_2660;
wire n_1038;
wire n_1369;
wire n_520;
wire n_409;
wire n_2611;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2553;
wire n_2581;
wire n_2195;
wire n_2529;
wire n_2698;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_2626;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_2510;
wire n_868;
wire n_2454;
wire n_639;
wire n_2804;
wire n_914;
wire n_2120;
wire n_411;
wire n_414;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_2801;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_2763;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_2813;
wire n_2825;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_2667;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_2891;
wire n_1189;
wire n_2690;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_2449;
wire n_1733;
wire n_1244;
wire n_2413;
wire n_431;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_2621;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_2491;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_2671;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_2518;
wire n_2876;
wire n_1415;
wire n_2629;
wire n_2592;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_2838;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_2563;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2517;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_2631;
wire n_1308;
wire n_2871;
wire n_2178;
wire n_1767;
wire n_2913;
wire n_2336;
wire n_1680;
wire n_1233;
wire n_2607;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_372;
wire n_677;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_2723;
wire n_604;
wire n_2007;
wire n_433;
wire n_949;
wire n_2539;
wire n_2582;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_2736;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_2718;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_2577;
wire n_1760;
wire n_2875;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_2796;
wire n_757;
wire n_2342;
wire n_633;
wire n_2856;
wire n_439;
wire n_1832;
wire n_448;
wire n_1851;
wire n_999;
wire n_758;
wire n_2046;
wire n_2848;
wire n_2741;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_2805;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_2580;
wire n_2545;
wire n_2787;
wire n_2914;
wire n_1964;
wire n_2869;
wire n_1163;
wire n_906;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_2846;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2925;
wire n_2035;
wire n_658;
wire n_2061;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_2398;
wire n_1362;
wire n_2857;
wire n_1586;
wire n_456;
wire n_959;
wire n_2459;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_2666;
wire n_1017;
wire n_2481;
wire n_2171;
wire n_978;
wire n_2768;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_2900;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_2886;
wire n_2093;
wire n_1079;
wire n_457;
wire n_514;
wire n_1045;
wire n_1208;
wire n_2339;
wire n_2038;
wire n_2320;
wire n_2473;
wire n_2137;
wire n_603;
wire n_1431;
wire n_2583;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_2299;
wire n_2540;
wire n_2873;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_750;
wire n_742;
wire n_2029;
wire n_995;
wire n_454;
wire n_2168;
wire n_2790;
wire n_1609;
wire n_374;
wire n_1989;
wire n_2359;
wire n_396;
wire n_1887;
wire n_2523;
wire n_1383;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_662;
wire n_459;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_1336;
wire n_2882;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_2737;
wire n_1574;
wire n_2399;
wire n_2812;
wire n_473;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_2721;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_2585;
wire n_486;
wire n_1800;
wire n_1548;
wire n_2725;
wire n_614;
wire n_1421;
wire n_2571;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_2565;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_2729;
wire n_2418;
wire n_829;
wire n_2519;
wire n_2724;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_2897;
wire n_2909;
wire n_1724;
wire n_2111;
wire n_2521;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_2595;
wire n_1127;
wire n_2277;
wire n_761;
wire n_2477;
wire n_1785;
wire n_1568;
wire n_2829;
wire n_1006;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2474;
wire n_2879;
wire n_2604;
wire n_2090;
wire n_1870;
wire n_512;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_2628;
wire n_1249;
wire n_2896;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_2681;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_2775;
wire n_2716;
wire n_1913;
wire n_2878;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_2464;
wire n_1101;
wire n_2831;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_2851;
wire n_987;
wire n_1846;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_2452;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_2849;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_2905;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_2220;
wire n_2455;
wire n_628;
wire n_1849;
wire n_2410;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_2922;
wire n_1430;
wire n_2645;
wire n_2467;
wire n_513;
wire n_2727;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_2696;
wire n_1044;
wire n_1205;
wire n_2436;
wire n_1209;
wire n_1552;
wire n_2508;
wire n_495;
wire n_602;
wire n_574;
wire n_2593;
wire n_1435;
wire n_879;
wire n_2416;
wire n_2405;
wire n_623;
wire n_2088;
wire n_405;
wire n_824;
wire n_1645;
wire n_2461;
wire n_490;
wire n_1327;
wire n_2858;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_2658;
wire n_1717;
wire n_572;
wire n_2895;
wire n_815;
wire n_1795;
wire n_2128;
wire n_2578;
wire n_1821;
wire n_1381;
wire n_2555;
wire n_2662;
wire n_2740;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_2656;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_2890;
wire n_2554;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_2512;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2786;
wire n_2534;
wire n_2092;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_2694;
wire n_1776;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2281;
wire n_2131;
wire n_2789;
wire n_2216;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2308;
wire n_1893;
wire n_2910;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_2647;
wire n_1311;
wire n_2191;
wire n_2864;
wire n_1519;
wire n_950;
wire n_2428;
wire n_1553;
wire n_2664;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_389;
wire n_2465;
wire n_2824;
wire n_2650;
wire n_418;
wire n_912;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_2923;
wire n_2541;
wire n_1139;
wire n_2731;
wire n_515;
wire n_2333;
wire n_885;
wire n_2916;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_2402;
wire n_1157;
wire n_2403;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_2760;
wire n_2792;
wire n_2870;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_2304;
wire n_762;
wire n_1283;
wire n_1644;
wire n_2637;
wire n_2334;
wire n_690;
wire n_1974;
wire n_2463;
wire n_583;
wire n_2086;
wire n_2289;
wire n_1343;
wire n_2701;
wire n_2783;
wire n_2263;
wire n_2881;
wire n_1203;
wire n_1631;
wire n_2472;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_621;
wire n_753;
wire n_2475;
wire n_2733;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_2785;
wire n_2556;
wire n_507;
wire n_2269;
wire n_2732;
wire n_2309;
wire n_2415;
wire n_2646;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2816;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_2685;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_2460;
wire n_2589;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_2903;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_2743;
wire n_2675;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_2827;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_2755;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_2362;
wire n_856;
wire n_2609;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_2468;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_2364;
wire n_2533;
wire n_540;
wire n_618;
wire n_896;
wire n_2310;
wire n_2780;
wire n_2287;
wire n_2860;
wire n_2291;
wire n_2596;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_2670;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_2393;
wire n_833;
wire n_2318;
wire n_2020;
wire n_1646;
wire n_2502;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2749;
wire n_2043;
wire n_2901;
wire n_1940;
wire n_814;
wire n_2707;
wire n_2751;
wire n_2793;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_2758;
wire n_1458;
wire n_472;
wire n_669;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_2471;
wire n_1807;
wire n_387;
wire n_1149;
wire n_2618;
wire n_398;
wire n_1671;
wire n_635;
wire n_2559;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2840;
wire n_2810;
wire n_2325;
wire n_2747;
wire n_2446;
wire n_1814;
wire n_1035;
wire n_2822;
wire n_783;
wire n_555;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_2893;
wire n_1188;
wire n_2588;
wire n_1722;
wire n_661;
wire n_2441;
wire n_1802;
wire n_2600;
wire n_849;
wire n_2795;
wire n_681;
wire n_584;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_2282;
wire n_510;
wire n_2800;
wire n_2371;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2619;
wire n_2340;
wire n_2444;
wire n_2068;
wire n_875;
wire n_1110;
wire n_1655;
wire n_445;
wire n_2641;
wire n_749;
wire n_1895;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_2361;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_2638;
wire n_866;
wire n_969;
wire n_1401;
wire n_2492;
wire n_1019;
wire n_1105;
wire n_1998;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_2711;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_2653;
wire n_836;
wire n_990;
wire n_2867;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_2794;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_2608;
wire n_2657;
wire n_458;
wire n_770;
wire n_1375;
wire n_2494;
wire n_2649;
wire n_1102;
wire n_2852;
wire n_2392;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_2633;
wire n_1441;
wire n_2522;
wire n_2435;
wire n_1597;
wire n_1392;
wire n_1929;
wire n_2807;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2313;
wire n_2542;
wire n_489;
wire n_1174;
wire n_2431;
wire n_2835;
wire n_2558;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2564;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_2409;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_726;
wire n_982;
wire n_2575;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_2766;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2722;
wire n_2117;
wire n_2745;
wire n_1904;
wire n_2640;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_1514;
wire n_1335;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_1168;
wire n_707;
wire n_2219;
wire n_2437;
wire n_2885;
wire n_2877;
wire n_2148;
wire n_937;
wire n_2445;
wire n_1427;
wire n_2779;
wire n_393;
wire n_487;
wire n_1584;
wire n_1726;
wire n_1835;
wire n_665;
wire n_1440;
wire n_2164;
wire n_421;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_2845;
wire n_1787;
wire n_2634;
wire n_910;
wire n_2232;
wire n_2212;
wire n_2602;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_2811;
wire n_1496;
wire n_1125;
wire n_410;
wire n_2547;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_2501;
wire n_1915;
wire n_1109;
wire n_895;
wire n_2532;
wire n_1310;
wire n_2605;
wire n_2121;
wire n_1803;
wire n_2665;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_2924;
wire n_808;
wire n_2484;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_500;
wire n_1067;
wire n_1720;
wire n_2830;
wire n_2401;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_2692;
wire n_538;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_2754;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_2866;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_2806;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_2917;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_2926;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_2814;
wire n_1170;
wire n_2023;
wire n_2213;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_855;
wire n_1178;
wire n_1461;
wire n_2697;
wire n_850;
wire n_684;
wire n_2421;
wire n_2286;
wire n_2902;
wire n_664;
wire n_1999;
wire n_503;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_2480;
wire n_1372;
wire n_2861;
wire n_605;
wire n_2630;
wire n_1273;
wire n_1822;
wire n_2363;
wire n_643;
wire n_620;
wire n_2430;
wire n_916;
wire n_1081;
wire n_2549;
wire n_493;
wire n_2705;
wire n_2332;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_2433;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_2601;
wire n_998;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_2686;
wire n_2528;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2836;
wire n_2316;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_2906;
wire n_382;
wire n_554;
wire n_1625;
wire n_2130;
wire n_2284;
wire n_2187;
wire n_898;
wire n_2817;
wire n_2773;
wire n_2598;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_2687;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_2850;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_2654;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_2884;
wire n_1268;
wire n_559;
wire n_825;
wire n_2819;
wire n_1981;
wire n_508;
wire n_2186;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_2560;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2422;
wire n_2239;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_2448;
wire n_548;
wire n_812;
wire n_2104;
wire n_2748;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_2898;
wire n_782;
wire n_2717;
wire n_2818;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_2889;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_2772;
wire n_481;
wire n_1675;
wire n_1924;
wire n_2573;
wire n_1727;
wire n_2710;
wire n_1554;
wire n_1745;
wire n_2735;
wire n_769;
wire n_2497;
wire n_2006;
wire n_2844;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_654;
wire n_1172;
wire n_2535;
wire n_379;
wire n_428;
wire n_1341;
wire n_2726;
wire n_570;
wire n_2774;
wire n_1641;
wire n_1361;
wire n_2382;
wire n_1707;
wire n_853;
wire n_377;
wire n_2317;
wire n_751;
wire n_2799;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_392;
wire n_2579;
wire n_2476;
wire n_704;
wire n_787;
wire n_1770;
wire n_2781;
wire n_2456;
wire n_961;
wire n_2250;
wire n_2678;
wire n_1756;
wire n_771;
wire n_2778;
wire n_1716;
wire n_2788;
wire n_2872;
wire n_1225;
wire n_1520;
wire n_2451;
wire n_2887;
wire n_522;
wire n_1287;
wire n_1262;
wire n_2691;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_1962;
wire n_622;
wire n_1577;
wire n_2423;
wire n_1087;
wire n_2526;
wire n_2854;
wire n_386;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_2874;
wire n_2764;
wire n_2703;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_2680;
wire n_682;
wire n_1567;
wire n_2567;
wire n_1247;
wire n_2709;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_631;
wire n_479;
wire n_1246;
wire n_1478;
wire n_1339;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2357;
wire n_2183;
wire n_2673;
wire n_2742;
wire n_2360;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_1842;
wire n_871;
wire n_2442;
wire n_685;
wire n_598;
wire n_928;
wire n_1367;
wire n_608;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_2834;
wire n_499;
wire n_2531;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_2570;
wire n_2702;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2815;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_2744;
wire n_1348;
wire n_2030;
wire n_903;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_740;
wire n_2883;
wire n_384;
wire n_2208;
wire n_1404;
wire n_2912;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_462;
wire n_2050;
wire n_2809;
wire n_1193;
wire n_2797;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2591;
wire n_2146;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_2612;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_2841;
wire n_1627;
wire n_2918;
wire n_1245;
wire n_846;
wire n_2427;
wire n_2505;
wire n_2438;
wire n_1673;
wire n_465;
wire n_2832;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_2278;
wire n_616;
wire n_2594;
wire n_2394;
wire n_1914;
wire n_2135;
wire n_2335;
wire n_2904;
wire n_745;
wire n_2381;
wire n_1654;
wire n_2569;
wire n_2349;
wire n_1103;
wire n_648;
wire n_1379;
wire n_2734;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_2823;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2404;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_2485;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_2279;
wire n_2655;
wire n_2027;
wire n_453;
wire n_403;
wire n_2642;
wire n_1130;
wire n_720;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_2513;
wire n_2525;
wire n_2695;
wire n_1764;
wire n_2892;
wire n_712;
wire n_2414;
wire n_2907;
wire n_1583;
wire n_2426;
wire n_2826;
wire n_1042;
wire n_1402;
wire n_2820;
wire n_2049;
wire n_2273;
wire n_412;
wire n_2719;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2708;
wire n_2113;
wire n_566;
wire n_565;
wire n_2586;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_1996;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2044;
wire n_2689;
wire n_2920;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_2614;
wire n_2511;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_2752;
wire n_2894;
wire n_1693;
wire n_438;
wire n_2599;
wire n_713;
wire n_2704;
wire n_904;
wire n_2839;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_2524;
wire n_1271;
wire n_2802;
wire n_533;
wire n_1542;
wire n_1251;
wire n_2728;
wire n_2268;

INVx2_ASAP7_75t_L g370 ( 
.A(n_30),
.Y(n_370)
);

BUFx10_ASAP7_75t_L g371 ( 
.A(n_175),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_37),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_68),
.Y(n_373)
);

INVx2_ASAP7_75t_SL g374 ( 
.A(n_253),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_241),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_367),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_331),
.Y(n_377)
);

INVx2_ASAP7_75t_SL g378 ( 
.A(n_180),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_138),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_307),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_328),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_150),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_109),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_297),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_314),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_287),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_70),
.Y(n_387)
);

INVx2_ASAP7_75t_SL g388 ( 
.A(n_189),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_309),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_357),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_361),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_289),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_230),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_239),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_256),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g396 ( 
.A(n_299),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_60),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_282),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_74),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_237),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_44),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_31),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_29),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_86),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_11),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_279),
.Y(n_406)
);

BUFx10_ASAP7_75t_L g407 ( 
.A(n_284),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_80),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_155),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_366),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_84),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_354),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_192),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_224),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_4),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_293),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_223),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_242),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_157),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_30),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_28),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_324),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_158),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_9),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_137),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_236),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_353),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_345),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_330),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_47),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_220),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_54),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_205),
.Y(n_433)
);

BUFx8_ASAP7_75t_SL g434 ( 
.A(n_347),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_152),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_201),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_325),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_296),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_136),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_252),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_265),
.Y(n_441)
);

BUFx10_ASAP7_75t_L g442 ( 
.A(n_213),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_222),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_311),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_318),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_327),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_343),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_120),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_303),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_51),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_45),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_160),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_302),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_336),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_306),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_118),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_126),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_84),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_245),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_17),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_356),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_276),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_208),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_227),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_89),
.Y(n_465)
);

BUFx10_ASAP7_75t_L g466 ( 
.A(n_333),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_360),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_171),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_54),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_342),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_209),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_85),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_277),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_258),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_368),
.Y(n_475)
);

INVx1_ASAP7_75t_SL g476 ( 
.A(n_123),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_275),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_66),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_113),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_169),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_39),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_183),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_288),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_298),
.Y(n_484)
);

INVx1_ASAP7_75t_SL g485 ( 
.A(n_69),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_206),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_294),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_281),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_355),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_168),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_363),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_25),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_337),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_31),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_102),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_272),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_346),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_123),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_11),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_173),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_308),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_76),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_335),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_350),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_18),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_91),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_255),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_204),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_261),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_225),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_88),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_45),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_316),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_33),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_215),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_219),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_170),
.Y(n_517)
);

CKINVDCx5p33_ASAP7_75t_R g518 ( 
.A(n_285),
.Y(n_518)
);

BUFx8_ASAP7_75t_SL g519 ( 
.A(n_233),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_246),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_76),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_69),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_72),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_141),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_36),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_100),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_200),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_283),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_148),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_125),
.Y(n_530)
);

BUFx10_ASAP7_75t_L g531 ( 
.A(n_257),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_118),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_228),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_26),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_4),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_107),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_358),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_36),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_79),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_40),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_141),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_121),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_195),
.Y(n_543)
);

CKINVDCx16_ASAP7_75t_R g544 ( 
.A(n_46),
.Y(n_544)
);

INVx1_ASAP7_75t_SL g545 ( 
.A(n_47),
.Y(n_545)
);

INVx1_ASAP7_75t_SL g546 ( 
.A(n_349),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_120),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_0),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_348),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_292),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_238),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_67),
.Y(n_552)
);

BUFx10_ASAP7_75t_L g553 ( 
.A(n_300),
.Y(n_553)
);

CKINVDCx16_ASAP7_75t_R g554 ( 
.A(n_93),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_61),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_329),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_312),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_147),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_166),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_16),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_58),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_142),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_305),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_310),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_66),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_320),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_154),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_188),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_146),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_232),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_24),
.Y(n_571)
);

INVx1_ASAP7_75t_SL g572 ( 
.A(n_210),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_63),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_67),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_341),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_17),
.Y(n_576)
);

CKINVDCx20_ASAP7_75t_R g577 ( 
.A(n_352),
.Y(n_577)
);

INVx1_ASAP7_75t_SL g578 ( 
.A(n_317),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_60),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_112),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_359),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_5),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_364),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_280),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_109),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_92),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_89),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_63),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g589 ( 
.A(n_290),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_20),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_133),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_340),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_269),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_145),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_163),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_218),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_164),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_68),
.Y(n_598)
);

INVx1_ASAP7_75t_SL g599 ( 
.A(n_49),
.Y(n_599)
);

BUFx2_ASAP7_75t_L g600 ( 
.A(n_291),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_136),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_369),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_199),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_55),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_70),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_55),
.Y(n_606)
);

INVxp67_ASAP7_75t_SL g607 ( 
.A(n_322),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_304),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_86),
.Y(n_609)
);

BUFx3_ASAP7_75t_L g610 ( 
.A(n_18),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_33),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_326),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_115),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_93),
.Y(n_614)
);

CKINVDCx14_ASAP7_75t_R g615 ( 
.A(n_295),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_338),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_42),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_319),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_216),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_362),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_117),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_64),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_159),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_144),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_5),
.Y(n_625)
);

BUFx2_ASAP7_75t_L g626 ( 
.A(n_94),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_37),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_49),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_108),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_301),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_174),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_271),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_259),
.Y(n_633)
);

CKINVDCx16_ASAP7_75t_R g634 ( 
.A(n_321),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_90),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_162),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_179),
.Y(n_637)
);

INVx1_ASAP7_75t_SL g638 ( 
.A(n_46),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_88),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_198),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_142),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_196),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_73),
.Y(n_643)
);

INVx1_ASAP7_75t_SL g644 ( 
.A(n_351),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_140),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_16),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_332),
.Y(n_647)
);

CKINVDCx20_ASAP7_75t_R g648 ( 
.A(n_178),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_151),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_181),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_107),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_323),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_135),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_1),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_365),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_146),
.Y(n_656)
);

INVxp67_ASAP7_75t_L g657 ( 
.A(n_140),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_315),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_339),
.Y(n_659)
);

INVxp33_ASAP7_75t_L g660 ( 
.A(n_187),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_80),
.Y(n_661)
);

CKINVDCx20_ASAP7_75t_R g662 ( 
.A(n_35),
.Y(n_662)
);

CKINVDCx20_ASAP7_75t_R g663 ( 
.A(n_127),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_144),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_334),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_128),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_313),
.Y(n_667)
);

BUFx6f_ASAP7_75t_L g668 ( 
.A(n_172),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_186),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_226),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_97),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_111),
.Y(n_672)
);

CKINVDCx20_ASAP7_75t_R g673 ( 
.A(n_344),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_286),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_211),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_128),
.Y(n_676)
);

CKINVDCx16_ASAP7_75t_R g677 ( 
.A(n_544),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_635),
.Y(n_678)
);

INVxp67_ASAP7_75t_SL g679 ( 
.A(n_600),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_635),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_434),
.Y(n_681)
);

CKINVDCx20_ASAP7_75t_R g682 ( 
.A(n_472),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_635),
.Y(n_683)
);

INVxp67_ASAP7_75t_L g684 ( 
.A(n_626),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_610),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_610),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_424),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_424),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_424),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_424),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_424),
.Y(n_691)
);

BUFx6f_ASAP7_75t_L g692 ( 
.A(n_461),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_548),
.Y(n_693)
);

INVxp67_ASAP7_75t_SL g694 ( 
.A(n_500),
.Y(n_694)
);

CKINVDCx20_ASAP7_75t_R g695 ( 
.A(n_536),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_548),
.Y(n_696)
);

BUFx2_ASAP7_75t_SL g697 ( 
.A(n_375),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_548),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_554),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_548),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_548),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_621),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_621),
.Y(n_703)
);

CKINVDCx20_ASAP7_75t_R g704 ( 
.A(n_552),
.Y(n_704)
);

CKINVDCx20_ASAP7_75t_R g705 ( 
.A(n_574),
.Y(n_705)
);

CKINVDCx20_ASAP7_75t_R g706 ( 
.A(n_662),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_621),
.Y(n_707)
);

INVxp67_ASAP7_75t_L g708 ( 
.A(n_415),
.Y(n_708)
);

INVx1_ASAP7_75t_SL g709 ( 
.A(n_663),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_519),
.Y(n_710)
);

INVxp67_ASAP7_75t_L g711 ( 
.A(n_506),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_621),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_500),
.Y(n_713)
);

CKINVDCx16_ASAP7_75t_R g714 ( 
.A(n_634),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_621),
.Y(n_715)
);

INVxp67_ASAP7_75t_SL g716 ( 
.A(n_535),
.Y(n_716)
);

CKINVDCx20_ASAP7_75t_R g717 ( 
.A(n_372),
.Y(n_717)
);

CKINVDCx16_ASAP7_75t_R g718 ( 
.A(n_615),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_373),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_420),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_399),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_401),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_402),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_405),
.Y(n_724)
);

INVxp67_ASAP7_75t_L g725 ( 
.A(n_448),
.Y(n_725)
);

INVxp33_ASAP7_75t_SL g726 ( 
.A(n_372),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_450),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_457),
.Y(n_728)
);

CKINVDCx5p33_ASAP7_75t_R g729 ( 
.A(n_414),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_494),
.Y(n_730)
);

INVxp33_ASAP7_75t_L g731 ( 
.A(n_370),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_498),
.Y(n_732)
);

CKINVDCx20_ASAP7_75t_R g733 ( 
.A(n_379),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_512),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_540),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_541),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_560),
.Y(n_737)
);

INVxp67_ASAP7_75t_SL g738 ( 
.A(n_660),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_565),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_571),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_586),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_601),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_613),
.Y(n_743)
);

INVxp33_ASAP7_75t_L g744 ( 
.A(n_370),
.Y(n_744)
);

INVxp33_ASAP7_75t_L g745 ( 
.A(n_451),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_617),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_421),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_622),
.Y(n_748)
);

INVxp67_ASAP7_75t_SL g749 ( 
.A(n_380),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_425),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_627),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_451),
.Y(n_752)
);

CKINVDCx16_ASAP7_75t_R g753 ( 
.A(n_429),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_639),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_643),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_645),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_651),
.Y(n_757)
);

CKINVDCx20_ASAP7_75t_R g758 ( 
.A(n_379),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_654),
.Y(n_759)
);

CKINVDCx20_ASAP7_75t_R g760 ( 
.A(n_383),
.Y(n_760)
);

INVxp67_ASAP7_75t_SL g761 ( 
.A(n_381),
.Y(n_761)
);

BUFx3_ASAP7_75t_L g762 ( 
.A(n_371),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_656),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_661),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_672),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_382),
.Y(n_766)
);

CKINVDCx20_ASAP7_75t_R g767 ( 
.A(n_383),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_430),
.Y(n_768)
);

CKINVDCx14_ASAP7_75t_R g769 ( 
.A(n_371),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_386),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_393),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_394),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_406),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_412),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_432),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_413),
.Y(n_776)
);

CKINVDCx16_ASAP7_75t_R g777 ( 
.A(n_449),
.Y(n_777)
);

INVxp67_ASAP7_75t_SL g778 ( 
.A(n_431),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_441),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_444),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_445),
.Y(n_781)
);

CKINVDCx20_ASAP7_75t_R g782 ( 
.A(n_387),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_447),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_452),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_453),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_454),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_459),
.Y(n_787)
);

CKINVDCx16_ASAP7_75t_R g788 ( 
.A(n_488),
.Y(n_788)
);

INVxp67_ASAP7_75t_L g789 ( 
.A(n_387),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_462),
.Y(n_790)
);

CKINVDCx14_ASAP7_75t_R g791 ( 
.A(n_371),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_439),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_477),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_480),
.Y(n_794)
);

INVx1_ASAP7_75t_SL g795 ( 
.A(n_476),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_482),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_487),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_416),
.Y(n_798)
);

CKINVDCx20_ASAP7_75t_R g799 ( 
.A(n_397),
.Y(n_799)
);

HB1xp67_ASAP7_75t_L g800 ( 
.A(n_397),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_491),
.Y(n_801)
);

CKINVDCx16_ASAP7_75t_R g802 ( 
.A(n_489),
.Y(n_802)
);

BUFx3_ASAP7_75t_L g803 ( 
.A(n_407),
.Y(n_803)
);

BUFx3_ASAP7_75t_L g804 ( 
.A(n_407),
.Y(n_804)
);

INVxp33_ASAP7_75t_L g805 ( 
.A(n_511),
.Y(n_805)
);

CKINVDCx16_ASAP7_75t_R g806 ( 
.A(n_504),
.Y(n_806)
);

CKINVDCx20_ASAP7_75t_R g807 ( 
.A(n_403),
.Y(n_807)
);

INVxp33_ASAP7_75t_SL g808 ( 
.A(n_403),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_497),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_503),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_507),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_417),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_510),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_529),
.Y(n_814)
);

INVxp67_ASAP7_75t_L g815 ( 
.A(n_404),
.Y(n_815)
);

CKINVDCx20_ASAP7_75t_R g816 ( 
.A(n_404),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_689),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_SL g818 ( 
.A(n_795),
.B(n_714),
.Y(n_818)
);

AND2x4_ASAP7_75t_L g819 ( 
.A(n_762),
.B(n_374),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_690),
.Y(n_820)
);

CKINVDCx20_ASAP7_75t_R g821 ( 
.A(n_682),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_691),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_738),
.B(n_407),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_687),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_693),
.Y(n_825)
);

OA21x2_ASAP7_75t_L g826 ( 
.A1(n_687),
.A2(n_437),
.B(n_400),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_729),
.B(n_798),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_800),
.Y(n_828)
);

BUFx6f_ASAP7_75t_L g829 ( 
.A(n_692),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_696),
.Y(n_830)
);

HB1xp67_ASAP7_75t_L g831 ( 
.A(n_789),
.Y(n_831)
);

OAI22xp5_ASAP7_75t_L g832 ( 
.A1(n_679),
.A2(n_657),
.B1(n_408),
.B2(n_523),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_812),
.B(n_374),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_698),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_694),
.B(n_378),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_700),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_762),
.B(n_378),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_701),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_688),
.Y(n_839)
);

BUFx8_ASAP7_75t_L g840 ( 
.A(n_803),
.Y(n_840)
);

AND2x4_ASAP7_75t_L g841 ( 
.A(n_803),
.B(n_388),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_688),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_681),
.Y(n_843)
);

BUFx8_ASAP7_75t_L g844 ( 
.A(n_804),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_749),
.B(n_388),
.Y(n_845)
);

CKINVDCx11_ASAP7_75t_R g846 ( 
.A(n_682),
.Y(n_846)
);

OAI21x1_ASAP7_75t_L g847 ( 
.A1(n_715),
.A2(n_437),
.B(n_400),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_715),
.Y(n_848)
);

INVx5_ASAP7_75t_L g849 ( 
.A(n_692),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_804),
.B(n_607),
.Y(n_850)
);

OA21x2_ASAP7_75t_L g851 ( 
.A1(n_702),
.A2(n_630),
.B(n_537),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_761),
.B(n_537),
.Y(n_852)
);

OAI22xp5_ASAP7_75t_L g853 ( 
.A1(n_684),
.A2(n_408),
.B1(n_523),
.B2(n_411),
.Y(n_853)
);

AND2x2_ASAP7_75t_SL g854 ( 
.A(n_718),
.B(n_630),
.Y(n_854)
);

BUFx6f_ASAP7_75t_L g855 ( 
.A(n_692),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_778),
.B(n_551),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_769),
.B(n_791),
.Y(n_857)
);

BUFx8_ASAP7_75t_SL g858 ( 
.A(n_695),
.Y(n_858)
);

HB1xp67_ASAP7_75t_L g859 ( 
.A(n_815),
.Y(n_859)
);

AND2x4_ASAP7_75t_L g860 ( 
.A(n_713),
.B(n_564),
.Y(n_860)
);

AOI22xp5_ASAP7_75t_L g861 ( 
.A1(n_726),
.A2(n_563),
.B1(n_577),
.B2(n_556),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_692),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_703),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_707),
.Y(n_864)
);

INVx5_ASAP7_75t_L g865 ( 
.A(n_752),
.Y(n_865)
);

INVxp33_ASAP7_75t_SL g866 ( 
.A(n_710),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_712),
.Y(n_867)
);

AOI22xp5_ASAP7_75t_L g868 ( 
.A1(n_726),
.A2(n_619),
.B1(n_648),
.B2(n_589),
.Y(n_868)
);

INVx2_ASAP7_75t_SL g869 ( 
.A(n_720),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_713),
.B(n_568),
.Y(n_870)
);

AND2x6_ASAP7_75t_L g871 ( 
.A(n_678),
.B(n_461),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_752),
.Y(n_872)
);

INVxp67_ASAP7_75t_L g873 ( 
.A(n_716),
.Y(n_873)
);

AOI22xp5_ASAP7_75t_L g874 ( 
.A1(n_808),
.A2(n_673),
.B1(n_458),
.B2(n_460),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_697),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_680),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_683),
.Y(n_877)
);

CKINVDCx16_ASAP7_75t_R g878 ( 
.A(n_753),
.Y(n_878)
);

AOI22xp5_ASAP7_75t_L g879 ( 
.A1(n_808),
.A2(n_465),
.B1(n_469),
.B2(n_456),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_766),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_770),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_771),
.B(n_570),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_772),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_773),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_774),
.Y(n_885)
);

BUFx6f_ASAP7_75t_L g886 ( 
.A(n_719),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_776),
.B(n_581),
.Y(n_887)
);

AND2x4_ASAP7_75t_L g888 ( 
.A(n_708),
.B(n_583),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_779),
.B(n_584),
.Y(n_889)
);

INVx5_ASAP7_75t_L g890 ( 
.A(n_677),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_721),
.Y(n_891)
);

AND2x4_ASAP7_75t_L g892 ( 
.A(n_711),
.B(n_596),
.Y(n_892)
);

INVx3_ASAP7_75t_L g893 ( 
.A(n_722),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_780),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_720),
.B(n_396),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_781),
.Y(n_896)
);

INVx3_ASAP7_75t_L g897 ( 
.A(n_723),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_724),
.Y(n_898)
);

OAI22x1_ASAP7_75t_L g899 ( 
.A1(n_699),
.A2(n_624),
.B1(n_625),
.B2(n_411),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_783),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_784),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_747),
.B(n_546),
.Y(n_902)
);

HB1xp67_ASAP7_75t_L g903 ( 
.A(n_699),
.Y(n_903)
);

HB1xp67_ASAP7_75t_L g904 ( 
.A(n_747),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_727),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_785),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_769),
.B(n_442),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_786),
.Y(n_908)
);

INVx2_ASAP7_75t_L g909 ( 
.A(n_787),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_790),
.Y(n_910)
);

BUFx2_ASAP7_75t_L g911 ( 
.A(n_717),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_685),
.B(n_602),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_750),
.B(n_572),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_728),
.Y(n_914)
);

INVx2_ASAP7_75t_SL g915 ( 
.A(n_750),
.Y(n_915)
);

BUFx3_ASAP7_75t_L g916 ( 
.A(n_686),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_793),
.Y(n_917)
);

INVx6_ASAP7_75t_L g918 ( 
.A(n_777),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_794),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_796),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_730),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_797),
.Y(n_922)
);

BUFx6f_ASAP7_75t_L g923 ( 
.A(n_732),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_801),
.Y(n_924)
);

AOI22xp5_ASAP7_75t_L g925 ( 
.A1(n_768),
.A2(n_479),
.B1(n_481),
.B2(n_478),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_809),
.B(n_631),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_768),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_810),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_734),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_791),
.B(n_442),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_811),
.B(n_632),
.Y(n_931)
);

INVx4_ASAP7_75t_L g932 ( 
.A(n_775),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_813),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_814),
.Y(n_934)
);

AND2x4_ASAP7_75t_L g935 ( 
.A(n_725),
.B(n_633),
.Y(n_935)
);

OA21x2_ASAP7_75t_L g936 ( 
.A1(n_735),
.A2(n_652),
.B(n_637),
.Y(n_936)
);

OAI21x1_ASAP7_75t_L g937 ( 
.A1(n_736),
.A2(n_670),
.B(n_667),
.Y(n_937)
);

AND2x4_ASAP7_75t_L g938 ( 
.A(n_737),
.B(n_578),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_739),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_731),
.B(n_442),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_740),
.Y(n_941)
);

HB1xp67_ASAP7_75t_L g942 ( 
.A(n_940),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_843),
.Y(n_943)
);

CKINVDCx20_ASAP7_75t_R g944 ( 
.A(n_821),
.Y(n_944)
);

BUFx10_ASAP7_75t_L g945 ( 
.A(n_895),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_939),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_R g947 ( 
.A(n_927),
.B(n_775),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_824),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_858),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_941),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_858),
.Y(n_951)
);

INVx3_ASAP7_75t_L g952 ( 
.A(n_829),
.Y(n_952)
);

CKINVDCx20_ASAP7_75t_R g953 ( 
.A(n_821),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_824),
.Y(n_954)
);

CKINVDCx20_ASAP7_75t_R g955 ( 
.A(n_846),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_875),
.Y(n_956)
);

BUFx2_ASAP7_75t_L g957 ( 
.A(n_903),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_866),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_883),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_894),
.Y(n_960)
);

CKINVDCx20_ASAP7_75t_R g961 ( 
.A(n_878),
.Y(n_961)
);

HB1xp67_ASAP7_75t_L g962 ( 
.A(n_828),
.Y(n_962)
);

NOR2xp67_ASAP7_75t_L g963 ( 
.A(n_890),
.B(n_792),
.Y(n_963)
);

XNOR2xp5_ASAP7_75t_L g964 ( 
.A(n_861),
.B(n_868),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_846),
.Y(n_965)
);

HB1xp67_ASAP7_75t_L g966 ( 
.A(n_828),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_840),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_840),
.Y(n_968)
);

CKINVDCx16_ASAP7_75t_R g969 ( 
.A(n_818),
.Y(n_969)
);

CKINVDCx16_ASAP7_75t_R g970 ( 
.A(n_903),
.Y(n_970)
);

BUFx2_ASAP7_75t_L g971 ( 
.A(n_904),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_844),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_900),
.Y(n_973)
);

INVx3_ASAP7_75t_L g974 ( 
.A(n_829),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_844),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_906),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_910),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_833),
.B(n_792),
.Y(n_978)
);

INVx1_ASAP7_75t_SL g979 ( 
.A(n_911),
.Y(n_979)
);

CKINVDCx20_ASAP7_75t_R g980 ( 
.A(n_904),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_922),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_890),
.Y(n_982)
);

CKINVDCx20_ASAP7_75t_R g983 ( 
.A(n_918),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_890),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_839),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_924),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_890),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_916),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_918),
.Y(n_989)
);

CKINVDCx20_ASAP7_75t_R g990 ( 
.A(n_918),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_850),
.B(n_644),
.Y(n_991)
);

CKINVDCx20_ASAP7_75t_R g992 ( 
.A(n_932),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_827),
.Y(n_993)
);

CKINVDCx20_ASAP7_75t_R g994 ( 
.A(n_932),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_R g995 ( 
.A(n_869),
.B(n_788),
.Y(n_995)
);

BUFx2_ASAP7_75t_L g996 ( 
.A(n_907),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_R g997 ( 
.A(n_915),
.B(n_802),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_895),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_902),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_902),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_913),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_913),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_874),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_831),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_916),
.Y(n_1005)
);

INVx2_ASAP7_75t_SL g1006 ( 
.A(n_819),
.Y(n_1006)
);

HB1xp67_ASAP7_75t_L g1007 ( 
.A(n_831),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_859),
.Y(n_1008)
);

CKINVDCx20_ASAP7_75t_R g1009 ( 
.A(n_857),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_859),
.Y(n_1010)
);

OAI21x1_ASAP7_75t_L g1011 ( 
.A1(n_847),
.A2(n_742),
.B(n_741),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_873),
.B(n_731),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_877),
.Y(n_1013)
);

NAND2xp33_ASAP7_75t_R g1014 ( 
.A(n_850),
.B(n_376),
.Y(n_1014)
);

HB1xp67_ASAP7_75t_L g1015 ( 
.A(n_819),
.Y(n_1015)
);

CKINVDCx20_ASAP7_75t_R g1016 ( 
.A(n_873),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_839),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_829),
.Y(n_1018)
);

CKINVDCx20_ASAP7_75t_R g1019 ( 
.A(n_879),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_829),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_886),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_925),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_854),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_854),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_837),
.B(n_461),
.Y(n_1025)
);

NOR2xp33_ASAP7_75t_R g1026 ( 
.A(n_930),
.B(n_806),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_837),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_842),
.Y(n_1028)
);

AND2x2_ASAP7_75t_L g1029 ( 
.A(n_841),
.B(n_744),
.Y(n_1029)
);

INVx3_ASAP7_75t_L g1030 ( 
.A(n_855),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_842),
.Y(n_1031)
);

BUFx10_ASAP7_75t_L g1032 ( 
.A(n_841),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_848),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_899),
.Y(n_1034)
);

HB1xp67_ASAP7_75t_L g1035 ( 
.A(n_938),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_832),
.Y(n_1036)
);

BUFx6f_ASAP7_75t_L g1037 ( 
.A(n_855),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_856),
.Y(n_1038)
);

CKINVDCx5p33_ASAP7_75t_R g1039 ( 
.A(n_823),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_886),
.Y(n_1040)
);

CKINVDCx20_ASAP7_75t_R g1041 ( 
.A(n_823),
.Y(n_1041)
);

NAND2xp33_ASAP7_75t_SL g1042 ( 
.A(n_845),
.B(n_624),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_835),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_853),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_938),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_860),
.Y(n_1046)
);

BUFx3_ASAP7_75t_L g1047 ( 
.A(n_860),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_886),
.Y(n_1048)
);

INVxp67_ASAP7_75t_L g1049 ( 
.A(n_870),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_852),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_848),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_SL g1052 ( 
.A(n_888),
.Y(n_1052)
);

INVxp67_ASAP7_75t_L g1053 ( 
.A(n_888),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_892),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_886),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_891),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_864),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_892),
.Y(n_1058)
);

AOI21x1_ASAP7_75t_L g1059 ( 
.A1(n_882),
.A2(n_746),
.B(n_743),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_935),
.Y(n_1060)
);

BUFx10_ASAP7_75t_L g1061 ( 
.A(n_935),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_891),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_891),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_864),
.Y(n_1064)
);

INVxp67_ASAP7_75t_SL g1065 ( 
.A(n_855),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_891),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_893),
.B(n_744),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_898),
.Y(n_1068)
);

CKINVDCx20_ASAP7_75t_R g1069 ( 
.A(n_887),
.Y(n_1069)
);

CKINVDCx20_ASAP7_75t_R g1070 ( 
.A(n_889),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_912),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_898),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_898),
.Y(n_1073)
);

NOR2xp67_ASAP7_75t_L g1074 ( 
.A(n_893),
.B(n_418),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_898),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_905),
.Y(n_1076)
);

CKINVDCx20_ASAP7_75t_R g1077 ( 
.A(n_926),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_905),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_905),
.Y(n_1079)
);

CKINVDCx20_ASAP7_75t_R g1080 ( 
.A(n_931),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_905),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_914),
.Y(n_1082)
);

CKINVDCx20_ASAP7_75t_R g1083 ( 
.A(n_936),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_914),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_914),
.Y(n_1085)
);

INVx3_ASAP7_75t_L g1086 ( 
.A(n_855),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_872),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_914),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_921),
.Y(n_1089)
);

INVxp67_ASAP7_75t_SL g1090 ( 
.A(n_862),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_921),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_921),
.Y(n_1092)
);

OA21x2_ASAP7_75t_L g1093 ( 
.A1(n_937),
.A2(n_820),
.B(n_817),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_921),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_923),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_923),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_R g1097 ( 
.A(n_897),
.B(n_695),
.Y(n_1097)
);

INVx2_ASAP7_75t_SL g1098 ( 
.A(n_912),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_923),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_923),
.Y(n_1100)
);

CKINVDCx20_ASAP7_75t_R g1101 ( 
.A(n_936),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_929),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_929),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_872),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_929),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_862),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_929),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_897),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_880),
.Y(n_1109)
);

BUFx10_ASAP7_75t_L g1110 ( 
.A(n_871),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_880),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_881),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_1038),
.B(n_376),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_1050),
.B(n_936),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_1011),
.Y(n_1115)
);

BUFx6f_ASAP7_75t_L g1116 ( 
.A(n_1047),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_1043),
.B(n_377),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_998),
.B(n_709),
.Y(n_1118)
);

NAND3xp33_ASAP7_75t_L g1119 ( 
.A(n_942),
.B(n_826),
.C(n_851),
.Y(n_1119)
);

INVx5_ASAP7_75t_L g1120 ( 
.A(n_1110),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_1039),
.B(n_377),
.Y(n_1121)
);

CKINVDCx6p67_ASAP7_75t_R g1122 ( 
.A(n_955),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_946),
.Y(n_1123)
);

BUFx6f_ASAP7_75t_L g1124 ( 
.A(n_1047),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_948),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1049),
.B(n_826),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1012),
.B(n_826),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_1067),
.B(n_851),
.Y(n_1128)
);

INVxp67_ASAP7_75t_L g1129 ( 
.A(n_1029),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_950),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_948),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_954),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_1032),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_1035),
.B(n_745),
.Y(n_1134)
);

NAND2xp33_ASAP7_75t_L g1135 ( 
.A(n_993),
.B(n_419),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_954),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_985),
.Y(n_1137)
);

AO22x2_ASAP7_75t_L g1138 ( 
.A1(n_964),
.A2(n_545),
.B1(n_599),
.B2(n_485),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_1087),
.Y(n_1139)
);

BUFx2_ASAP7_75t_L g1140 ( 
.A(n_1097),
.Y(n_1140)
);

INVx4_ASAP7_75t_SL g1141 ( 
.A(n_1052),
.Y(n_1141)
);

NAND2xp33_ASAP7_75t_SL g1142 ( 
.A(n_999),
.B(n_717),
.Y(n_1142)
);

OR2x2_ASAP7_75t_L g1143 ( 
.A(n_1007),
.B(n_638),
.Y(n_1143)
);

INVxp67_ASAP7_75t_SL g1144 ( 
.A(n_1083),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_985),
.Y(n_1145)
);

OAI22xp5_ASAP7_75t_SL g1146 ( 
.A1(n_1019),
.A2(n_705),
.B1(n_706),
.B2(n_704),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_959),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1083),
.B(n_851),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1017),
.Y(n_1149)
);

NAND2x1p5_ASAP7_75t_L g1150 ( 
.A(n_1006),
.B(n_461),
.Y(n_1150)
);

BUFx3_ASAP7_75t_L g1151 ( 
.A(n_983),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_960),
.Y(n_1152)
);

CKINVDCx8_ASAP7_75t_R g1153 ( 
.A(n_949),
.Y(n_1153)
);

BUFx10_ASAP7_75t_L g1154 ( 
.A(n_958),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_973),
.Y(n_1155)
);

CKINVDCx16_ASAP7_75t_R g1156 ( 
.A(n_995),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1017),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_976),
.Y(n_1158)
);

HB1xp67_ASAP7_75t_L g1159 ( 
.A(n_1045),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_977),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_1098),
.B(n_876),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1028),
.Y(n_1162)
);

BUFx3_ASAP7_75t_L g1163 ( 
.A(n_990),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_981),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_986),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1013),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_1000),
.B(n_733),
.Y(n_1167)
);

OR2x6_ASAP7_75t_L g1168 ( 
.A(n_957),
.B(n_511),
.Y(n_1168)
);

BUFx6f_ASAP7_75t_L g1169 ( 
.A(n_1032),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_988),
.Y(n_1170)
);

AND2x4_ASAP7_75t_L g1171 ( 
.A(n_1005),
.B(n_1071),
.Y(n_1171)
);

AOI22xp33_ASAP7_75t_L g1172 ( 
.A1(n_1101),
.A2(n_573),
.B1(n_576),
.B2(n_538),
.Y(n_1172)
);

INVx4_ASAP7_75t_L g1173 ( 
.A(n_1062),
.Y(n_1173)
);

HB1xp67_ASAP7_75t_L g1174 ( 
.A(n_1015),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1087),
.Y(n_1175)
);

NOR2xp33_ASAP7_75t_L g1176 ( 
.A(n_1001),
.B(n_733),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1028),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1104),
.Y(n_1178)
);

AND2x4_ASAP7_75t_L g1179 ( 
.A(n_1053),
.B(n_876),
.Y(n_1179)
);

BUFx3_ASAP7_75t_L g1180 ( 
.A(n_989),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1101),
.B(n_822),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_L g1182 ( 
.A(n_1002),
.B(n_758),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_1031),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1031),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1033),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1104),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1057),
.Y(n_1187)
);

INVx4_ASAP7_75t_L g1188 ( 
.A(n_1063),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1033),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1051),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1057),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1051),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_978),
.B(n_758),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1064),
.Y(n_1194)
);

BUFx3_ASAP7_75t_L g1195 ( 
.A(n_961),
.Y(n_1195)
);

BUFx6f_ASAP7_75t_L g1196 ( 
.A(n_1032),
.Y(n_1196)
);

INVx4_ASAP7_75t_L g1197 ( 
.A(n_1073),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1064),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1093),
.Y(n_1199)
);

BUFx4f_ASAP7_75t_L g1200 ( 
.A(n_971),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_945),
.B(n_745),
.Y(n_1201)
);

HB1xp67_ASAP7_75t_L g1202 ( 
.A(n_962),
.Y(n_1202)
);

NOR2xp33_ASAP7_75t_L g1203 ( 
.A(n_991),
.B(n_760),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1109),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1111),
.Y(n_1205)
);

AOI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1023),
.A2(n_767),
.B1(n_782),
.B2(n_760),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1076),
.B(n_825),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1079),
.B(n_830),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1112),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_SL g1210 ( 
.A(n_945),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1093),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1093),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_L g1213 ( 
.A(n_1027),
.B(n_767),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_945),
.B(n_805),
.Y(n_1214)
);

INVx3_ASAP7_75t_L g1215 ( 
.A(n_952),
.Y(n_1215)
);

INVx2_ASAP7_75t_L g1216 ( 
.A(n_952),
.Y(n_1216)
);

INVx4_ASAP7_75t_L g1217 ( 
.A(n_1082),
.Y(n_1217)
);

INVx4_ASAP7_75t_SL g1218 ( 
.A(n_1052),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_SL g1219 ( 
.A(n_1108),
.B(n_384),
.Y(n_1219)
);

INVxp67_ASAP7_75t_SL g1220 ( 
.A(n_1020),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_996),
.B(n_881),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_952),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_1059),
.B(n_884),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1021),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_1024),
.B(n_782),
.Y(n_1225)
);

INVx3_ASAP7_75t_L g1226 ( 
.A(n_974),
.Y(n_1226)
);

INVx3_ASAP7_75t_L g1227 ( 
.A(n_974),
.Y(n_1227)
);

AND2x4_ASAP7_75t_L g1228 ( 
.A(n_963),
.B(n_884),
.Y(n_1228)
);

AND2x6_ASAP7_75t_L g1229 ( 
.A(n_1040),
.B(n_461),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1048),
.Y(n_1230)
);

AND2x2_ASAP7_75t_SL g1231 ( 
.A(n_969),
.B(n_538),
.Y(n_1231)
);

INVx4_ASAP7_75t_L g1232 ( 
.A(n_1084),
.Y(n_1232)
);

INVx1_ASAP7_75t_SL g1233 ( 
.A(n_1016),
.Y(n_1233)
);

INVx4_ASAP7_75t_SL g1234 ( 
.A(n_1020),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1055),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1088),
.B(n_834),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_974),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1056),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1018),
.Y(n_1239)
);

BUFx6f_ASAP7_75t_L g1240 ( 
.A(n_1020),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1066),
.Y(n_1241)
);

NAND2x1p5_ASAP7_75t_L g1242 ( 
.A(n_1068),
.B(n_471),
.Y(n_1242)
);

NAND2xp33_ASAP7_75t_SL g1243 ( 
.A(n_1041),
.B(n_799),
.Y(n_1243)
);

HB1xp67_ASAP7_75t_L g1244 ( 
.A(n_966),
.Y(n_1244)
);

BUFx10_ASAP7_75t_L g1245 ( 
.A(n_951),
.Y(n_1245)
);

BUFx6f_ASAP7_75t_L g1246 ( 
.A(n_1020),
.Y(n_1246)
);

AND2x2_ASAP7_75t_SL g1247 ( 
.A(n_970),
.B(n_573),
.Y(n_1247)
);

NOR2xp33_ASAP7_75t_L g1248 ( 
.A(n_1069),
.B(n_799),
.Y(n_1248)
);

AND2x6_ASAP7_75t_L g1249 ( 
.A(n_1072),
.B(n_471),
.Y(n_1249)
);

OR2x2_ASAP7_75t_L g1250 ( 
.A(n_979),
.B(n_805),
.Y(n_1250)
);

INVx1_ASAP7_75t_SL g1251 ( 
.A(n_1004),
.Y(n_1251)
);

AND2x2_ASAP7_75t_L g1252 ( 
.A(n_1008),
.B(n_807),
.Y(n_1252)
);

NAND2xp33_ASAP7_75t_L g1253 ( 
.A(n_1089),
.B(n_422),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1091),
.B(n_836),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1092),
.B(n_838),
.Y(n_1255)
);

BUFx6f_ASAP7_75t_L g1256 ( 
.A(n_1037),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1075),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1094),
.B(n_867),
.Y(n_1258)
);

INVx5_ASAP7_75t_L g1259 ( 
.A(n_1110),
.Y(n_1259)
);

INVx1_ASAP7_75t_SL g1260 ( 
.A(n_1010),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1078),
.Y(n_1261)
);

INVxp33_ASAP7_75t_L g1262 ( 
.A(n_947),
.Y(n_1262)
);

INVx3_ASAP7_75t_L g1263 ( 
.A(n_1018),
.Y(n_1263)
);

INVxp67_ASAP7_75t_SL g1264 ( 
.A(n_1037),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1081),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1085),
.Y(n_1266)
);

INVx3_ASAP7_75t_L g1267 ( 
.A(n_1018),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1099),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1103),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1025),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1061),
.B(n_807),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1025),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1030),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1061),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1061),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_SL g1276 ( 
.A(n_1095),
.B(n_384),
.Y(n_1276)
);

AO22x2_ASAP7_75t_L g1277 ( 
.A1(n_1003),
.A2(n_664),
.B1(n_576),
.B2(n_816),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1060),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_SL g1279 ( 
.A(n_1096),
.B(n_385),
.Y(n_1279)
);

NAND2xp33_ASAP7_75t_L g1280 ( 
.A(n_1100),
.B(n_423),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1054),
.Y(n_1281)
);

INVxp67_ASAP7_75t_SL g1282 ( 
.A(n_1037),
.Y(n_1282)
);

XOR2xp5_ASAP7_75t_L g1283 ( 
.A(n_944),
.B(n_704),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1058),
.Y(n_1284)
);

BUFx3_ASAP7_75t_L g1285 ( 
.A(n_1009),
.Y(n_1285)
);

INVx2_ASAP7_75t_L g1286 ( 
.A(n_1030),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1102),
.B(n_885),
.Y(n_1287)
);

AND2x4_ASAP7_75t_L g1288 ( 
.A(n_1046),
.B(n_885),
.Y(n_1288)
);

BUFx3_ASAP7_75t_L g1289 ( 
.A(n_943),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1105),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1107),
.Y(n_1291)
);

NAND2x1p5_ASAP7_75t_L g1292 ( 
.A(n_1030),
.B(n_471),
.Y(n_1292)
);

BUFx3_ASAP7_75t_L g1293 ( 
.A(n_992),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1074),
.B(n_896),
.Y(n_1294)
);

BUFx3_ASAP7_75t_L g1295 ( 
.A(n_994),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1086),
.Y(n_1296)
);

OR2x2_ASAP7_75t_L g1297 ( 
.A(n_1042),
.B(n_748),
.Y(n_1297)
);

OR2x2_ASAP7_75t_L g1298 ( 
.A(n_1042),
.B(n_1044),
.Y(n_1298)
);

AND2x4_ASAP7_75t_L g1299 ( 
.A(n_1041),
.B(n_896),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1086),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1086),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1069),
.Y(n_1302)
);

BUFx6f_ASAP7_75t_SL g1303 ( 
.A(n_967),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1070),
.Y(n_1304)
);

INVx4_ASAP7_75t_L g1305 ( 
.A(n_1037),
.Y(n_1305)
);

AO22x2_ASAP7_75t_L g1306 ( 
.A1(n_1036),
.A2(n_664),
.B1(n_816),
.B2(n_754),
.Y(n_1306)
);

CKINVDCx20_ASAP7_75t_R g1307 ( 
.A(n_944),
.Y(n_1307)
);

OA22x2_ASAP7_75t_L g1308 ( 
.A1(n_1034),
.A2(n_628),
.B1(n_629),
.B2(n_625),
.Y(n_1308)
);

NOR2xp67_ASAP7_75t_L g1309 ( 
.A(n_1119),
.B(n_1114),
.Y(n_1309)
);

INVxp67_ASAP7_75t_L g1310 ( 
.A(n_1250),
.Y(n_1310)
);

NAND2x1p5_ASAP7_75t_L g1311 ( 
.A(n_1133),
.B(n_1106),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_1133),
.B(n_982),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1172),
.B(n_1022),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1139),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1187),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1172),
.A2(n_1070),
.B1(n_1080),
.B2(n_1077),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1139),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1191),
.Y(n_1318)
);

NOR2xp33_ASAP7_75t_L g1319 ( 
.A(n_1118),
.B(n_956),
.Y(n_1319)
);

NAND2x1p5_ASAP7_75t_L g1320 ( 
.A(n_1133),
.B(n_1106),
.Y(n_1320)
);

INVxp67_ASAP7_75t_L g1321 ( 
.A(n_1202),
.Y(n_1321)
);

A2O1A1Ixp33_ASAP7_75t_L g1322 ( 
.A1(n_1129),
.A2(n_1077),
.B(n_1080),
.C(n_1019),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1194),
.Y(n_1323)
);

AOI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1144),
.A2(n_1014),
.B1(n_980),
.B2(n_389),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1179),
.Y(n_1325)
);

CKINVDCx5p33_ASAP7_75t_R g1326 ( 
.A(n_1289),
.Y(n_1326)
);

HB1xp67_ASAP7_75t_L g1327 ( 
.A(n_1202),
.Y(n_1327)
);

AND2x2_ASAP7_75t_SL g1328 ( 
.A(n_1156),
.B(n_953),
.Y(n_1328)
);

NAND2x1p5_ASAP7_75t_L g1329 ( 
.A(n_1169),
.B(n_1106),
.Y(n_1329)
);

AND2x4_ASAP7_75t_L g1330 ( 
.A(n_1169),
.B(n_984),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1179),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1148),
.A2(n_1144),
.B1(n_1114),
.B2(n_1298),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1127),
.B(n_1148),
.Y(n_1333)
);

AO22x2_ASAP7_75t_L g1334 ( 
.A1(n_1302),
.A2(n_980),
.B1(n_706),
.B2(n_705),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1198),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1175),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1178),
.Y(n_1337)
);

AO22x2_ASAP7_75t_L g1338 ( 
.A1(n_1304),
.A2(n_953),
.B1(n_755),
.B2(n_756),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1186),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_L g1340 ( 
.A(n_1127),
.B(n_1065),
.Y(n_1340)
);

NOR2xp33_ASAP7_75t_L g1341 ( 
.A(n_1193),
.B(n_1203),
.Y(n_1341)
);

BUFx4f_ASAP7_75t_L g1342 ( 
.A(n_1169),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_SL g1343 ( 
.A(n_1196),
.B(n_1026),
.Y(n_1343)
);

AO22x2_ASAP7_75t_L g1344 ( 
.A1(n_1283),
.A2(n_757),
.B1(n_759),
.B2(n_751),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1123),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1125),
.Y(n_1346)
);

AND2x4_ASAP7_75t_L g1347 ( 
.A(n_1196),
.B(n_987),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1201),
.B(n_1214),
.Y(n_1348)
);

BUFx6f_ASAP7_75t_L g1349 ( 
.A(n_1196),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1130),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1147),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_1154),
.Y(n_1352)
);

INVxp67_ASAP7_75t_L g1353 ( 
.A(n_1134),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1152),
.Y(n_1354)
);

A2O1A1Ixp33_ASAP7_75t_L g1355 ( 
.A1(n_1129),
.A2(n_908),
.B(n_909),
.C(n_901),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1155),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1158),
.Y(n_1357)
);

A2O1A1Ixp33_ASAP7_75t_L g1358 ( 
.A1(n_1270),
.A2(n_908),
.B(n_909),
.C(n_901),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1131),
.Y(n_1359)
);

INVxp67_ASAP7_75t_L g1360 ( 
.A(n_1244),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1128),
.B(n_1090),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1160),
.Y(n_1362)
);

BUFx3_ASAP7_75t_L g1363 ( 
.A(n_1180),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1164),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1193),
.B(n_997),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1165),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1166),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1161),
.Y(n_1368)
);

INVx3_ASAP7_75t_L g1369 ( 
.A(n_1215),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1132),
.Y(n_1370)
);

AND2x4_ASAP7_75t_L g1371 ( 
.A(n_1116),
.B(n_917),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1136),
.Y(n_1372)
);

AOI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1181),
.A2(n_389),
.B1(n_390),
.B2(n_385),
.Y(n_1373)
);

BUFx12f_ASAP7_75t_L g1374 ( 
.A(n_1154),
.Y(n_1374)
);

NAND2x1p5_ASAP7_75t_L g1375 ( 
.A(n_1120),
.B(n_1106),
.Y(n_1375)
);

AND2x4_ASAP7_75t_L g1376 ( 
.A(n_1116),
.B(n_917),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_L g1377 ( 
.A(n_1203),
.B(n_965),
.Y(n_1377)
);

OAI221xp5_ASAP7_75t_L g1378 ( 
.A1(n_1181),
.A2(n_641),
.B1(n_646),
.B2(n_629),
.C(n_628),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1137),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1161),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1145),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1204),
.B(n_968),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1149),
.Y(n_1383)
);

NAND3x1_ASAP7_75t_L g1384 ( 
.A(n_1206),
.B(n_955),
.C(n_764),
.Y(n_1384)
);

AND3x4_ASAP7_75t_L g1385 ( 
.A(n_1285),
.B(n_920),
.C(n_919),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1157),
.Y(n_1386)
);

AO22x2_ASAP7_75t_L g1387 ( 
.A1(n_1121),
.A2(n_1233),
.B1(n_1299),
.B2(n_1297),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1162),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1177),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1183),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1184),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1185),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1189),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1190),
.Y(n_1394)
);

OAI221xp5_ASAP7_75t_L g1395 ( 
.A1(n_1287),
.A2(n_653),
.B1(n_666),
.B2(n_646),
.C(n_641),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1192),
.Y(n_1396)
);

AO22x2_ASAP7_75t_L g1397 ( 
.A1(n_1233),
.A2(n_1299),
.B1(n_1306),
.B2(n_1277),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1170),
.Y(n_1398)
);

INVx2_ASAP7_75t_SL g1399 ( 
.A(n_1200),
.Y(n_1399)
);

AND2x4_ASAP7_75t_L g1400 ( 
.A(n_1116),
.B(n_919),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1128),
.B(n_920),
.Y(n_1401)
);

INVx2_ASAP7_75t_L g1402 ( 
.A(n_1215),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1223),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1223),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1224),
.Y(n_1405)
);

AOI22xp5_ASAP7_75t_L g1406 ( 
.A1(n_1272),
.A2(n_391),
.B1(n_392),
.B2(n_390),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1226),
.Y(n_1407)
);

AND2x4_ASAP7_75t_L g1408 ( 
.A(n_1124),
.B(n_928),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1230),
.Y(n_1409)
);

AND2x4_ASAP7_75t_L g1410 ( 
.A(n_1124),
.B(n_928),
.Y(n_1410)
);

OR2x2_ASAP7_75t_L g1411 ( 
.A(n_1251),
.B(n_972),
.Y(n_1411)
);

OAI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1126),
.A2(n_1231),
.B1(n_1119),
.B2(n_1211),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1235),
.Y(n_1413)
);

OAI221xp5_ASAP7_75t_L g1414 ( 
.A1(n_1287),
.A2(n_1126),
.B1(n_1208),
.B2(n_1236),
.C(n_1207),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1226),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1238),
.Y(n_1416)
);

INVxp67_ASAP7_75t_L g1417 ( 
.A(n_1244),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1205),
.B(n_975),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_1307),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1241),
.Y(n_1420)
);

OR2x2_ASAP7_75t_L g1421 ( 
.A(n_1251),
.B(n_933),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1199),
.B(n_933),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1227),
.Y(n_1423)
);

AO22x2_ASAP7_75t_L g1424 ( 
.A1(n_1306),
.A2(n_765),
.B1(n_763),
.B2(n_2),
.Y(n_1424)
);

AND2x4_ASAP7_75t_L g1425 ( 
.A(n_1124),
.B(n_934),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1257),
.Y(n_1426)
);

INVxp67_ASAP7_75t_L g1427 ( 
.A(n_1143),
.Y(n_1427)
);

INVxp67_ASAP7_75t_L g1428 ( 
.A(n_1209),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1261),
.Y(n_1429)
);

INVxp67_ASAP7_75t_L g1430 ( 
.A(n_1159),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1227),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1265),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1212),
.B(n_934),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1220),
.B(n_863),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1220),
.B(n_863),
.Y(n_1435)
);

INVxp67_ASAP7_75t_L g1436 ( 
.A(n_1159),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1266),
.Y(n_1437)
);

AND2x4_ASAP7_75t_L g1438 ( 
.A(n_1171),
.B(n_391),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1263),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1268),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1269),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1296),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_1153),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1300),
.Y(n_1444)
);

INVx4_ASAP7_75t_L g1445 ( 
.A(n_1173),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1263),
.Y(n_1446)
);

NOR2xp33_ASAP7_75t_L g1447 ( 
.A(n_1176),
.B(n_1262),
.Y(n_1447)
);

INVxp67_ASAP7_75t_L g1448 ( 
.A(n_1174),
.Y(n_1448)
);

INVxp67_ASAP7_75t_L g1449 ( 
.A(n_1174),
.Y(n_1449)
);

A2O1A1Ixp33_ASAP7_75t_L g1450 ( 
.A1(n_1294),
.A2(n_395),
.B(n_398),
.C(n_392),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1267),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1267),
.Y(n_1452)
);

INVx2_ASAP7_75t_L g1453 ( 
.A(n_1216),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1222),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1237),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1239),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1273),
.Y(n_1457)
);

BUFx2_ASAP7_75t_L g1458 ( 
.A(n_1200),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1286),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_1167),
.B(n_395),
.Y(n_1460)
);

A2O1A1Ixp33_ASAP7_75t_L g1461 ( 
.A1(n_1341),
.A2(n_1182),
.B(n_1167),
.C(n_1225),
.Y(n_1461)
);

AOI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1361),
.A2(n_1282),
.B(n_1264),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1348),
.B(n_1207),
.Y(n_1463)
);

AOI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1313),
.A2(n_1182),
.B1(n_1135),
.B2(n_1225),
.Y(n_1464)
);

BUFx3_ASAP7_75t_L g1465 ( 
.A(n_1363),
.Y(n_1465)
);

OAI21xp33_ASAP7_75t_SL g1466 ( 
.A1(n_1313),
.A2(n_1236),
.B(n_1208),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_SL g1467 ( 
.A(n_1319),
.B(n_1173),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1333),
.B(n_1254),
.Y(n_1468)
);

OAI21xp5_ASAP7_75t_L g1469 ( 
.A1(n_1309),
.A2(n_1115),
.B(n_1294),
.Y(n_1469)
);

OAI21xp5_ASAP7_75t_L g1470 ( 
.A1(n_1309),
.A2(n_1255),
.B(n_1254),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1365),
.B(n_1260),
.Y(n_1471)
);

AOI21xp5_ASAP7_75t_L g1472 ( 
.A1(n_1361),
.A2(n_1282),
.B(n_1264),
.Y(n_1472)
);

AOI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1340),
.A2(n_1259),
.B(n_1120),
.Y(n_1473)
);

OAI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1414),
.A2(n_1197),
.B1(n_1217),
.B2(n_1188),
.Y(n_1474)
);

AOI21xp5_ASAP7_75t_L g1475 ( 
.A1(n_1340),
.A2(n_1259),
.B(n_1120),
.Y(n_1475)
);

AOI21xp5_ASAP7_75t_L g1476 ( 
.A1(n_1333),
.A2(n_1259),
.B(n_1120),
.Y(n_1476)
);

NOR2xp33_ASAP7_75t_L g1477 ( 
.A(n_1447),
.B(n_1260),
.Y(n_1477)
);

NAND2xp33_ASAP7_75t_L g1478 ( 
.A(n_1349),
.B(n_1259),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1332),
.A2(n_1221),
.B1(n_1228),
.B2(n_1171),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1332),
.A2(n_1414),
.B1(n_1460),
.B2(n_1378),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_L g1481 ( 
.A(n_1345),
.B(n_1255),
.Y(n_1481)
);

OR2x6_ASAP7_75t_L g1482 ( 
.A(n_1374),
.B(n_1151),
.Y(n_1482)
);

INVx3_ASAP7_75t_L g1483 ( 
.A(n_1349),
.Y(n_1483)
);

AO21x1_ASAP7_75t_L g1484 ( 
.A1(n_1412),
.A2(n_1150),
.B(n_1258),
.Y(n_1484)
);

OAI321xp33_ASAP7_75t_L g1485 ( 
.A1(n_1378),
.A2(n_1206),
.A3(n_1248),
.B1(n_1213),
.B2(n_1113),
.C(n_1146),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1350),
.B(n_1258),
.Y(n_1486)
);

AOI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1353),
.A2(n_1142),
.B1(n_1228),
.B2(n_1290),
.Y(n_1487)
);

BUFx4f_ASAP7_75t_L g1488 ( 
.A(n_1349),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1351),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_SL g1490 ( 
.A(n_1428),
.B(n_1188),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_SL g1491 ( 
.A(n_1342),
.B(n_1197),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1403),
.Y(n_1492)
);

INVx2_ASAP7_75t_SL g1493 ( 
.A(n_1327),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1354),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1356),
.B(n_1217),
.Y(n_1495)
);

AOI21xp5_ASAP7_75t_L g1496 ( 
.A1(n_1401),
.A2(n_1305),
.B(n_1246),
.Y(n_1496)
);

AOI21xp5_ASAP7_75t_L g1497 ( 
.A1(n_1401),
.A2(n_1305),
.B(n_1246),
.Y(n_1497)
);

AO21x2_ASAP7_75t_L g1498 ( 
.A1(n_1412),
.A2(n_1301),
.B(n_1291),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1368),
.A2(n_1221),
.B1(n_1308),
.B2(n_1247),
.Y(n_1499)
);

O2A1O1Ixp33_ASAP7_75t_L g1500 ( 
.A1(n_1395),
.A2(n_1353),
.B(n_1450),
.C(n_1355),
.Y(n_1500)
);

AOI21xp5_ASAP7_75t_L g1501 ( 
.A1(n_1434),
.A2(n_1246),
.B(n_1240),
.Y(n_1501)
);

AOI21xp5_ASAP7_75t_L g1502 ( 
.A1(n_1434),
.A2(n_1435),
.B(n_1433),
.Y(n_1502)
);

NAND2x1p5_ASAP7_75t_L g1503 ( 
.A(n_1342),
.B(n_1232),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_SL g1504 ( 
.A(n_1324),
.B(n_1232),
.Y(n_1504)
);

BUFx8_ASAP7_75t_L g1505 ( 
.A(n_1458),
.Y(n_1505)
);

BUFx6f_ASAP7_75t_L g1506 ( 
.A(n_1311),
.Y(n_1506)
);

AOI21xp5_ASAP7_75t_L g1507 ( 
.A1(n_1435),
.A2(n_1256),
.B(n_1240),
.Y(n_1507)
);

NOR2xp67_ASAP7_75t_L g1508 ( 
.A(n_1445),
.B(n_1278),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_SL g1509 ( 
.A(n_1324),
.B(n_1288),
.Y(n_1509)
);

NAND3xp33_ASAP7_75t_L g1510 ( 
.A(n_1316),
.B(n_1213),
.C(n_1252),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1357),
.B(n_1362),
.Y(n_1511)
);

BUFx2_ASAP7_75t_L g1512 ( 
.A(n_1310),
.Y(n_1512)
);

O2A1O1Ixp5_ASAP7_75t_L g1513 ( 
.A1(n_1358),
.A2(n_1279),
.B(n_1276),
.C(n_1117),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_SL g1514 ( 
.A(n_1445),
.B(n_1288),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1364),
.B(n_1219),
.Y(n_1515)
);

AOI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1380),
.A2(n_1308),
.B1(n_1138),
.B2(n_1243),
.Y(n_1516)
);

OAI21xp5_ASAP7_75t_L g1517 ( 
.A1(n_1422),
.A2(n_1280),
.B(n_1253),
.Y(n_1517)
);

AO21x1_ASAP7_75t_L g1518 ( 
.A1(n_1422),
.A2(n_1150),
.B(n_1292),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1366),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_1427),
.B(n_1140),
.Y(n_1520)
);

AOI21xp5_ASAP7_75t_L g1521 ( 
.A1(n_1433),
.A2(n_1256),
.B(n_1240),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1421),
.B(n_1195),
.Y(n_1522)
);

CKINVDCx14_ASAP7_75t_R g1523 ( 
.A(n_1419),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1367),
.B(n_1274),
.Y(n_1524)
);

AOI21xp33_ASAP7_75t_L g1525 ( 
.A1(n_1321),
.A2(n_1284),
.B(n_1281),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1404),
.B(n_1275),
.Y(n_1526)
);

O2A1O1Ixp5_ASAP7_75t_L g1527 ( 
.A1(n_1315),
.A2(n_1271),
.B(n_1242),
.C(n_1292),
.Y(n_1527)
);

OAI22xp5_ASAP7_75t_L g1528 ( 
.A1(n_1398),
.A2(n_1210),
.B1(n_1256),
.B2(n_1168),
.Y(n_1528)
);

BUFx12f_ASAP7_75t_L g1529 ( 
.A(n_1326),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1373),
.B(n_1168),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1373),
.B(n_1168),
.Y(n_1531)
);

AOI21xp5_ASAP7_75t_L g1532 ( 
.A1(n_1375),
.A2(n_849),
.B(n_1234),
.Y(n_1532)
);

AOI21xp5_ASAP7_75t_L g1533 ( 
.A1(n_1375),
.A2(n_849),
.B(n_1234),
.Y(n_1533)
);

OAI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1369),
.A2(n_1210),
.B1(n_1295),
.B2(n_1293),
.Y(n_1534)
);

A2O1A1Ixp33_ASAP7_75t_L g1535 ( 
.A1(n_1325),
.A2(n_1163),
.B(n_409),
.C(n_410),
.Y(n_1535)
);

OAI321xp33_ASAP7_75t_L g1536 ( 
.A1(n_1395),
.A2(n_1146),
.A3(n_1138),
.B1(n_1277),
.B2(n_471),
.C(n_668),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1405),
.B(n_1234),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1409),
.B(n_1242),
.Y(n_1538)
);

AOI21xp5_ASAP7_75t_L g1539 ( 
.A1(n_1369),
.A2(n_849),
.B(n_862),
.Y(n_1539)
);

BUFx6f_ASAP7_75t_L g1540 ( 
.A(n_1311),
.Y(n_1540)
);

OAI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1413),
.A2(n_409),
.B1(n_410),
.B2(n_398),
.Y(n_1541)
);

AOI21xp5_ASAP7_75t_L g1542 ( 
.A1(n_1402),
.A2(n_849),
.B(n_862),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1416),
.B(n_1420),
.Y(n_1543)
);

OAI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1426),
.A2(n_636),
.B1(n_640),
.B2(n_623),
.Y(n_1544)
);

O2A1O1Ixp33_ASAP7_75t_L g1545 ( 
.A1(n_1322),
.A2(n_531),
.B(n_553),
.C(n_466),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1429),
.B(n_1432),
.Y(n_1546)
);

OAI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1437),
.A2(n_636),
.B1(n_640),
.B2(n_623),
.Y(n_1547)
);

OAI21xp5_ASAP7_75t_L g1548 ( 
.A1(n_1318),
.A2(n_1249),
.B(n_1229),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1468),
.B(n_1331),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1489),
.Y(n_1550)
);

INVx3_ASAP7_75t_L g1551 ( 
.A(n_1506),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1494),
.Y(n_1552)
);

AOI21xp5_ASAP7_75t_L g1553 ( 
.A1(n_1517),
.A2(n_1343),
.B(n_1329),
.Y(n_1553)
);

O2A1O1Ixp5_ASAP7_75t_L g1554 ( 
.A1(n_1484),
.A2(n_1336),
.B(n_1337),
.C(n_1323),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1463),
.B(n_1481),
.Y(n_1555)
);

BUFx6f_ASAP7_75t_L g1556 ( 
.A(n_1488),
.Y(n_1556)
);

O2A1O1Ixp33_ASAP7_75t_L g1557 ( 
.A1(n_1461),
.A2(n_1377),
.B(n_1436),
.C(n_1430),
.Y(n_1557)
);

INVxp67_ASAP7_75t_SL g1558 ( 
.A(n_1478),
.Y(n_1558)
);

BUFx2_ASAP7_75t_L g1559 ( 
.A(n_1512),
.Y(n_1559)
);

INVx1_ASAP7_75t_SL g1560 ( 
.A(n_1522),
.Y(n_1560)
);

OR2x6_ASAP7_75t_L g1561 ( 
.A(n_1482),
.B(n_1399),
.Y(n_1561)
);

NOR2xp33_ASAP7_75t_L g1562 ( 
.A(n_1477),
.B(n_1471),
.Y(n_1562)
);

HB1xp67_ASAP7_75t_L g1563 ( 
.A(n_1493),
.Y(n_1563)
);

BUFx6f_ASAP7_75t_L g1564 ( 
.A(n_1488),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1486),
.B(n_1387),
.Y(n_1565)
);

NOR2xp33_ASAP7_75t_L g1566 ( 
.A(n_1464),
.B(n_1360),
.Y(n_1566)
);

NOR3xp33_ASAP7_75t_L g1567 ( 
.A(n_1485),
.B(n_1418),
.C(n_1382),
.Y(n_1567)
);

O2A1O1Ixp33_ASAP7_75t_L g1568 ( 
.A1(n_1485),
.A2(n_1417),
.B(n_1449),
.C(n_1448),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1519),
.Y(n_1569)
);

BUFx3_ASAP7_75t_L g1570 ( 
.A(n_1465),
.Y(n_1570)
);

BUFx2_ASAP7_75t_SL g1571 ( 
.A(n_1508),
.Y(n_1571)
);

AOI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1510),
.A2(n_1328),
.B1(n_1334),
.B2(n_1352),
.Y(n_1572)
);

BUFx6f_ASAP7_75t_L g1573 ( 
.A(n_1506),
.Y(n_1573)
);

INVx2_ASAP7_75t_SL g1574 ( 
.A(n_1505),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_1529),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1483),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1470),
.B(n_1480),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1479),
.B(n_1387),
.Y(n_1578)
);

NOR2x1_ASAP7_75t_SL g1579 ( 
.A(n_1474),
.B(n_1446),
.Y(n_1579)
);

INVx1_ASAP7_75t_SL g1580 ( 
.A(n_1525),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1511),
.B(n_1371),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_SL g1582 ( 
.A(n_1520),
.B(n_1495),
.Y(n_1582)
);

AOI21xp5_ASAP7_75t_L g1583 ( 
.A1(n_1502),
.A2(n_1329),
.B(n_1320),
.Y(n_1583)
);

HB1xp67_ASAP7_75t_L g1584 ( 
.A(n_1483),
.Y(n_1584)
);

BUFx4f_ASAP7_75t_SL g1585 ( 
.A(n_1505),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1543),
.B(n_1371),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_SL g1587 ( 
.A(n_1530),
.B(n_1312),
.Y(n_1587)
);

O2A1O1Ixp5_ASAP7_75t_SL g1588 ( 
.A1(n_1504),
.A2(n_1339),
.B(n_1455),
.C(n_1454),
.Y(n_1588)
);

NOR2xp33_ASAP7_75t_R g1589 ( 
.A(n_1523),
.B(n_1443),
.Y(n_1589)
);

BUFx6f_ASAP7_75t_L g1590 ( 
.A(n_1506),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1509),
.B(n_1411),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1546),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1515),
.B(n_1467),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1492),
.Y(n_1594)
);

NOR2x1_ASAP7_75t_SL g1595 ( 
.A(n_1540),
.B(n_1452),
.Y(n_1595)
);

OAI22xp5_ASAP7_75t_L g1596 ( 
.A1(n_1487),
.A2(n_1440),
.B1(n_1441),
.B2(n_1406),
.Y(n_1596)
);

NOR3xp33_ASAP7_75t_SL g1597 ( 
.A(n_1536),
.B(n_1466),
.C(n_1535),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1526),
.Y(n_1598)
);

BUFx12f_ASAP7_75t_L g1599 ( 
.A(n_1482),
.Y(n_1599)
);

AND3x1_ASAP7_75t_SL g1600 ( 
.A(n_1536),
.B(n_1334),
.C(n_1384),
.Y(n_1600)
);

NOR2xp33_ASAP7_75t_L g1601 ( 
.A(n_1531),
.B(n_1438),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1554),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1554),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1555),
.B(n_1462),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1550),
.Y(n_1605)
);

INVx3_ASAP7_75t_L g1606 ( 
.A(n_1573),
.Y(n_1606)
);

INVx5_ASAP7_75t_L g1607 ( 
.A(n_1561),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_SL g1608 ( 
.A(n_1580),
.B(n_1503),
.Y(n_1608)
);

BUFx8_ASAP7_75t_L g1609 ( 
.A(n_1559),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1552),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1592),
.B(n_1472),
.Y(n_1611)
);

INVx6_ASAP7_75t_SL g1612 ( 
.A(n_1561),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1577),
.B(n_1498),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1569),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_1589),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_1585),
.Y(n_1616)
);

BUFx3_ASAP7_75t_L g1617 ( 
.A(n_1599),
.Y(n_1617)
);

BUFx2_ASAP7_75t_L g1618 ( 
.A(n_1576),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1597),
.B(n_1498),
.Y(n_1619)
);

INVx4_ASAP7_75t_L g1620 ( 
.A(n_1573),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1565),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1594),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1597),
.B(n_1469),
.Y(n_1623)
);

BUFx12f_ASAP7_75t_L g1624 ( 
.A(n_1575),
.Y(n_1624)
);

BUFx3_ASAP7_75t_L g1625 ( 
.A(n_1556),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1579),
.Y(n_1626)
);

BUFx6f_ASAP7_75t_L g1627 ( 
.A(n_1578),
.Y(n_1627)
);

BUFx3_ASAP7_75t_L g1628 ( 
.A(n_1556),
.Y(n_1628)
);

BUFx3_ASAP7_75t_L g1629 ( 
.A(n_1556),
.Y(n_1629)
);

INVx3_ASAP7_75t_L g1630 ( 
.A(n_1573),
.Y(n_1630)
);

BUFx3_ASAP7_75t_L g1631 ( 
.A(n_1556),
.Y(n_1631)
);

CKINVDCx8_ASAP7_75t_R g1632 ( 
.A(n_1571),
.Y(n_1632)
);

BUFx3_ASAP7_75t_L g1633 ( 
.A(n_1564),
.Y(n_1633)
);

INVx2_ASAP7_75t_SL g1634 ( 
.A(n_1573),
.Y(n_1634)
);

INVx5_ASAP7_75t_L g1635 ( 
.A(n_1561),
.Y(n_1635)
);

BUFx3_ASAP7_75t_L g1636 ( 
.A(n_1564),
.Y(n_1636)
);

BUFx3_ASAP7_75t_L g1637 ( 
.A(n_1564),
.Y(n_1637)
);

INVx5_ASAP7_75t_L g1638 ( 
.A(n_1590),
.Y(n_1638)
);

BUFx3_ASAP7_75t_L g1639 ( 
.A(n_1564),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1598),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1549),
.Y(n_1641)
);

BUFx3_ASAP7_75t_L g1642 ( 
.A(n_1590),
.Y(n_1642)
);

BUFx6f_ASAP7_75t_L g1643 ( 
.A(n_1590),
.Y(n_1643)
);

NOR2x1_ASAP7_75t_R g1644 ( 
.A(n_1570),
.B(n_1312),
.Y(n_1644)
);

INVx5_ASAP7_75t_L g1645 ( 
.A(n_1590),
.Y(n_1645)
);

BUFx3_ASAP7_75t_L g1646 ( 
.A(n_1551),
.Y(n_1646)
);

BUFx3_ASAP7_75t_L g1647 ( 
.A(n_1551),
.Y(n_1647)
);

INVx2_ASAP7_75t_SL g1648 ( 
.A(n_1576),
.Y(n_1648)
);

INVx1_ASAP7_75t_SL g1649 ( 
.A(n_1560),
.Y(n_1649)
);

BUFx6f_ASAP7_75t_L g1650 ( 
.A(n_1587),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1595),
.Y(n_1651)
);

OAI21x1_ASAP7_75t_SL g1652 ( 
.A1(n_1611),
.A2(n_1553),
.B(n_1500),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1605),
.Y(n_1653)
);

INVx3_ASAP7_75t_L g1654 ( 
.A(n_1620),
.Y(n_1654)
);

AO31x2_ASAP7_75t_L g1655 ( 
.A1(n_1602),
.A2(n_1518),
.A3(n_1583),
.B(n_1475),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_SL g1656 ( 
.A(n_1616),
.B(n_1122),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1605),
.Y(n_1657)
);

NOR2xp67_ASAP7_75t_L g1658 ( 
.A(n_1615),
.B(n_1534),
.Y(n_1658)
);

HB1xp67_ASAP7_75t_L g1659 ( 
.A(n_1627),
.Y(n_1659)
);

OA21x2_ASAP7_75t_L g1660 ( 
.A1(n_1602),
.A2(n_1469),
.B(n_1527),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1610),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1610),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1622),
.Y(n_1663)
);

INVx3_ASAP7_75t_SL g1664 ( 
.A(n_1649),
.Y(n_1664)
);

INVx3_ASAP7_75t_L g1665 ( 
.A(n_1620),
.Y(n_1665)
);

OAI211xp5_ASAP7_75t_L g1666 ( 
.A1(n_1623),
.A2(n_1567),
.B(n_1572),
.C(n_1557),
.Y(n_1666)
);

BUFx2_ASAP7_75t_L g1667 ( 
.A(n_1609),
.Y(n_1667)
);

OAI22xp5_ASAP7_75t_L g1668 ( 
.A1(n_1632),
.A2(n_1562),
.B1(n_1591),
.B2(n_1601),
.Y(n_1668)
);

AOI22xp33_ASAP7_75t_L g1669 ( 
.A1(n_1623),
.A2(n_1567),
.B1(n_1424),
.B2(n_1338),
.Y(n_1669)
);

BUFx2_ASAP7_75t_L g1670 ( 
.A(n_1609),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1614),
.Y(n_1671)
);

A2O1A1Ixp33_ASAP7_75t_L g1672 ( 
.A1(n_1623),
.A2(n_1566),
.B(n_1545),
.C(n_1568),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1614),
.Y(n_1673)
);

INVx2_ASAP7_75t_L g1674 ( 
.A(n_1622),
.Y(n_1674)
);

NOR2xp33_ASAP7_75t_L g1675 ( 
.A(n_1641),
.B(n_1627),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1641),
.B(n_1593),
.Y(n_1676)
);

OAI22xp33_ASAP7_75t_L g1677 ( 
.A1(n_1649),
.A2(n_1596),
.B1(n_1600),
.B2(n_1582),
.Y(n_1677)
);

OAI21x1_ASAP7_75t_L g1678 ( 
.A1(n_1626),
.A2(n_1588),
.B(n_1611),
.Y(n_1678)
);

BUFx2_ASAP7_75t_L g1679 ( 
.A(n_1609),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1640),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1640),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1618),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1618),
.Y(n_1683)
);

OAI21xp5_ASAP7_75t_L g1684 ( 
.A1(n_1604),
.A2(n_1513),
.B(n_1490),
.Y(n_1684)
);

NOR2xp67_ASAP7_75t_L g1685 ( 
.A(n_1624),
.B(n_1563),
.Y(n_1685)
);

OAI21x1_ASAP7_75t_L g1686 ( 
.A1(n_1626),
.A2(n_1497),
.B(n_1496),
.Y(n_1686)
);

INVx3_ASAP7_75t_L g1687 ( 
.A(n_1620),
.Y(n_1687)
);

BUFx12f_ASAP7_75t_L g1688 ( 
.A(n_1624),
.Y(n_1688)
);

CKINVDCx5p33_ASAP7_75t_R g1689 ( 
.A(n_1624),
.Y(n_1689)
);

INVx3_ASAP7_75t_L g1690 ( 
.A(n_1620),
.Y(n_1690)
);

HB1xp67_ASAP7_75t_L g1691 ( 
.A(n_1627),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1621),
.Y(n_1692)
);

O2A1O1Ixp33_ASAP7_75t_L g1693 ( 
.A1(n_1608),
.A2(n_1528),
.B(n_1491),
.C(n_1586),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1621),
.Y(n_1694)
);

OAI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1632),
.A2(n_1516),
.B1(n_1558),
.B2(n_1503),
.Y(n_1695)
);

BUFx12f_ASAP7_75t_L g1696 ( 
.A(n_1609),
.Y(n_1696)
);

AND2x4_ASAP7_75t_L g1697 ( 
.A(n_1607),
.B(n_1584),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1648),
.Y(n_1698)
);

OAI21x1_ASAP7_75t_L g1699 ( 
.A1(n_1603),
.A2(n_1507),
.B(n_1501),
.Y(n_1699)
);

OAI21x1_ASAP7_75t_L g1700 ( 
.A1(n_1603),
.A2(n_1473),
.B(n_1521),
.Y(n_1700)
);

A2O1A1Ixp33_ASAP7_75t_L g1701 ( 
.A1(n_1619),
.A2(n_1558),
.B(n_1581),
.C(n_1406),
.Y(n_1701)
);

OAI21x1_ASAP7_75t_L g1702 ( 
.A1(n_1604),
.A2(n_1476),
.B(n_1542),
.Y(n_1702)
);

AND2x4_ASAP7_75t_L g1703 ( 
.A(n_1607),
.B(n_1563),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1648),
.Y(n_1704)
);

OAI21x1_ASAP7_75t_L g1705 ( 
.A1(n_1651),
.A2(n_1539),
.B(n_1548),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1648),
.Y(n_1706)
);

A2O1A1Ixp33_ASAP7_75t_L g1707 ( 
.A1(n_1619),
.A2(n_1524),
.B(n_1499),
.C(n_1424),
.Y(n_1707)
);

O2A1O1Ixp33_ASAP7_75t_SL g1708 ( 
.A1(n_1651),
.A2(n_1514),
.B(n_1537),
.C(n_1538),
.Y(n_1708)
);

AO21x2_ASAP7_75t_L g1709 ( 
.A1(n_1619),
.A2(n_1548),
.B(n_1533),
.Y(n_1709)
);

OA21x2_ASAP7_75t_L g1710 ( 
.A1(n_1613),
.A2(n_1457),
.B(n_1456),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1627),
.B(n_1376),
.Y(n_1711)
);

OAI221xp5_ASAP7_75t_L g1712 ( 
.A1(n_1617),
.A2(n_1632),
.B1(n_1482),
.B2(n_1650),
.C(n_671),
.Y(n_1712)
);

AOI211xp5_ASAP7_75t_SL g1713 ( 
.A1(n_1613),
.A2(n_1544),
.B(n_1547),
.C(n_1541),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1627),
.B(n_1650),
.Y(n_1714)
);

AO21x1_ASAP7_75t_L g1715 ( 
.A1(n_1651),
.A2(n_1400),
.B(n_1376),
.Y(n_1715)
);

OAI22xp33_ASAP7_75t_L g1716 ( 
.A1(n_1627),
.A2(n_666),
.B1(n_671),
.B2(n_653),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1627),
.Y(n_1717)
);

AOI22xp33_ASAP7_75t_SL g1718 ( 
.A1(n_1650),
.A2(n_1338),
.B1(n_1397),
.B2(n_1344),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1650),
.Y(n_1719)
);

OR2x6_ASAP7_75t_L g1720 ( 
.A(n_1650),
.B(n_1574),
.Y(n_1720)
);

OAI21x1_ASAP7_75t_L g1721 ( 
.A1(n_1613),
.A2(n_1532),
.B(n_1444),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1650),
.Y(n_1722)
);

OAI21x1_ASAP7_75t_L g1723 ( 
.A1(n_1606),
.A2(n_1442),
.B(n_1320),
.Y(n_1723)
);

INVx1_ASAP7_75t_SL g1724 ( 
.A(n_1625),
.Y(n_1724)
);

AOI21x1_ASAP7_75t_L g1725 ( 
.A1(n_1634),
.A2(n_1397),
.B(n_1381),
.Y(n_1725)
);

OA21x2_ASAP7_75t_L g1726 ( 
.A1(n_1634),
.A2(n_1386),
.B(n_1335),
.Y(n_1726)
);

AOI22xp33_ASAP7_75t_SL g1727 ( 
.A1(n_1650),
.A2(n_1344),
.B1(n_531),
.B2(n_553),
.Y(n_1727)
);

OAI21x1_ASAP7_75t_L g1728 ( 
.A1(n_1606),
.A2(n_1415),
.B(n_1407),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1607),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1607),
.Y(n_1730)
);

NAND2x1p5_ASAP7_75t_L g1731 ( 
.A(n_1607),
.B(n_1540),
.Y(n_1731)
);

OAI21x1_ASAP7_75t_L g1732 ( 
.A1(n_1606),
.A2(n_1431),
.B(n_1423),
.Y(n_1732)
);

BUFx12f_ASAP7_75t_L g1733 ( 
.A(n_1617),
.Y(n_1733)
);

AND2x4_ASAP7_75t_L g1734 ( 
.A(n_1607),
.B(n_1540),
.Y(n_1734)
);

CKINVDCx14_ASAP7_75t_R g1735 ( 
.A(n_1617),
.Y(n_1735)
);

OAI21x1_ASAP7_75t_L g1736 ( 
.A1(n_1606),
.A2(n_1451),
.B(n_1439),
.Y(n_1736)
);

OAI21x1_ASAP7_75t_SL g1737 ( 
.A1(n_1634),
.A2(n_1459),
.B(n_1453),
.Y(n_1737)
);

OAI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1727),
.A2(n_1607),
.B1(n_1635),
.B2(n_1612),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1653),
.Y(n_1739)
);

BUFx4f_ASAP7_75t_SL g1740 ( 
.A(n_1688),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1657),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1675),
.B(n_1635),
.Y(n_1742)
);

INVx11_ASAP7_75t_L g1743 ( 
.A(n_1733),
.Y(n_1743)
);

AOI21xp5_ASAP7_75t_L g1744 ( 
.A1(n_1701),
.A2(n_1635),
.B(n_1638),
.Y(n_1744)
);

AOI22xp33_ASAP7_75t_L g1745 ( 
.A1(n_1669),
.A2(n_531),
.B1(n_553),
.B2(n_466),
.Y(n_1745)
);

OR2x6_ASAP7_75t_L g1746 ( 
.A(n_1720),
.B(n_1643),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1661),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1662),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1681),
.Y(n_1749)
);

BUFx8_ASAP7_75t_L g1750 ( 
.A(n_1696),
.Y(n_1750)
);

OAI222xp33_ASAP7_75t_L g1751 ( 
.A1(n_1669),
.A2(n_1635),
.B1(n_502),
.B2(n_495),
.C1(n_505),
.C2(n_499),
.Y(n_1751)
);

CKINVDCx6p67_ASAP7_75t_R g1752 ( 
.A(n_1664),
.Y(n_1752)
);

OR2x2_ASAP7_75t_L g1753 ( 
.A(n_1714),
.B(n_1635),
.Y(n_1753)
);

BUFx4f_ASAP7_75t_SL g1754 ( 
.A(n_1664),
.Y(n_1754)
);

INVx4_ASAP7_75t_L g1755 ( 
.A(n_1654),
.Y(n_1755)
);

BUFx2_ASAP7_75t_R g1756 ( 
.A(n_1689),
.Y(n_1756)
);

AOI22xp5_ASAP7_75t_L g1757 ( 
.A1(n_1666),
.A2(n_1385),
.B1(n_1635),
.B2(n_1330),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1663),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1719),
.B(n_1635),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1681),
.Y(n_1760)
);

CKINVDCx5p33_ASAP7_75t_R g1761 ( 
.A(n_1735),
.Y(n_1761)
);

AO21x2_ASAP7_75t_L g1762 ( 
.A1(n_1652),
.A2(n_1389),
.B(n_1388),
.Y(n_1762)
);

INVx2_ASAP7_75t_L g1763 ( 
.A(n_1674),
.Y(n_1763)
);

INVxp67_ASAP7_75t_L g1764 ( 
.A(n_1675),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1680),
.Y(n_1765)
);

AO21x2_ASAP7_75t_L g1766 ( 
.A1(n_1684),
.A2(n_1394),
.B(n_1393),
.Y(n_1766)
);

INVx1_ASAP7_75t_SL g1767 ( 
.A(n_1724),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1674),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1682),
.Y(n_1769)
);

INVx2_ASAP7_75t_SL g1770 ( 
.A(n_1667),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1683),
.Y(n_1771)
);

HB1xp67_ASAP7_75t_L g1772 ( 
.A(n_1710),
.Y(n_1772)
);

CKINVDCx5p33_ASAP7_75t_R g1773 ( 
.A(n_1735),
.Y(n_1773)
);

INVx3_ASAP7_75t_L g1774 ( 
.A(n_1703),
.Y(n_1774)
);

NAND2x1_ASAP7_75t_L g1775 ( 
.A(n_1726),
.B(n_1630),
.Y(n_1775)
);

BUFx2_ASAP7_75t_SL g1776 ( 
.A(n_1685),
.Y(n_1776)
);

BUFx8_ASAP7_75t_L g1777 ( 
.A(n_1670),
.Y(n_1777)
);

OAI21x1_ASAP7_75t_L g1778 ( 
.A1(n_1700),
.A2(n_1630),
.B(n_1317),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1671),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1671),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1673),
.Y(n_1781)
);

INVx1_ASAP7_75t_SL g1782 ( 
.A(n_1703),
.Y(n_1782)
);

AOI22xp33_ASAP7_75t_L g1783 ( 
.A1(n_1727),
.A2(n_466),
.B1(n_514),
.B2(n_492),
.Y(n_1783)
);

AOI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1666),
.A2(n_1347),
.B1(n_1330),
.B2(n_1400),
.Y(n_1784)
);

HB1xp67_ASAP7_75t_L g1785 ( 
.A(n_1710),
.Y(n_1785)
);

BUFx2_ASAP7_75t_L g1786 ( 
.A(n_1679),
.Y(n_1786)
);

AND2x4_ASAP7_75t_L g1787 ( 
.A(n_1722),
.B(n_1642),
.Y(n_1787)
);

OAI21x1_ASAP7_75t_SL g1788 ( 
.A1(n_1725),
.A2(n_1612),
.B(n_1314),
.Y(n_1788)
);

INVx2_ASAP7_75t_SL g1789 ( 
.A(n_1720),
.Y(n_1789)
);

INVx3_ASAP7_75t_L g1790 ( 
.A(n_1720),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1692),
.Y(n_1791)
);

HB1xp67_ASAP7_75t_L g1792 ( 
.A(n_1710),
.Y(n_1792)
);

AOI21x1_ASAP7_75t_L g1793 ( 
.A1(n_1668),
.A2(n_1347),
.B(n_1408),
.Y(n_1793)
);

OAI21x1_ASAP7_75t_L g1794 ( 
.A1(n_1678),
.A2(n_1630),
.B(n_1359),
.Y(n_1794)
);

AO21x1_ASAP7_75t_L g1795 ( 
.A1(n_1677),
.A2(n_1438),
.B(n_1410),
.Y(n_1795)
);

BUFx3_ASAP7_75t_L g1796 ( 
.A(n_1697),
.Y(n_1796)
);

OAI22xp33_ASAP7_75t_L g1797 ( 
.A1(n_1713),
.A2(n_1612),
.B1(n_1645),
.B2(n_1638),
.Y(n_1797)
);

AOI21xp33_ASAP7_75t_L g1798 ( 
.A1(n_1672),
.A2(n_1644),
.B(n_1643),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1673),
.Y(n_1799)
);

AOI22xp33_ASAP7_75t_L g1800 ( 
.A1(n_1718),
.A2(n_1677),
.B1(n_1716),
.B2(n_1712),
.Y(n_1800)
);

INVx4_ASAP7_75t_L g1801 ( 
.A(n_1654),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1694),
.Y(n_1802)
);

HB1xp67_ASAP7_75t_L g1803 ( 
.A(n_1659),
.Y(n_1803)
);

AOI22xp33_ASAP7_75t_L g1804 ( 
.A1(n_1718),
.A2(n_521),
.B1(n_524),
.B2(n_522),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1698),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1704),
.Y(n_1806)
);

AOI21xp5_ASAP7_75t_L g1807 ( 
.A1(n_1701),
.A2(n_1645),
.B(n_1638),
.Y(n_1807)
);

NAND2x1p5_ASAP7_75t_L g1808 ( 
.A(n_1726),
.B(n_1638),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1717),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_L g1810 ( 
.A1(n_1716),
.A2(n_525),
.B1(n_530),
.B2(n_526),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1717),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1706),
.Y(n_1812)
);

AOI21x1_ASAP7_75t_L g1813 ( 
.A1(n_1729),
.A2(n_1410),
.B(n_1408),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1659),
.Y(n_1814)
);

INVx1_ASAP7_75t_SL g1815 ( 
.A(n_1676),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1691),
.Y(n_1816)
);

AOI22xp5_ASAP7_75t_L g1817 ( 
.A1(n_1672),
.A2(n_1425),
.B1(n_1628),
.B2(n_1625),
.Y(n_1817)
);

INVx3_ASAP7_75t_L g1818 ( 
.A(n_1665),
.Y(n_1818)
);

OAI21x1_ASAP7_75t_L g1819 ( 
.A1(n_1702),
.A2(n_1630),
.B(n_1370),
.Y(n_1819)
);

AOI22xp33_ASAP7_75t_L g1820 ( 
.A1(n_1695),
.A2(n_532),
.B1(n_539),
.B2(n_534),
.Y(n_1820)
);

INVx2_ASAP7_75t_L g1821 ( 
.A(n_1691),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1726),
.Y(n_1822)
);

AOI21x1_ASAP7_75t_L g1823 ( 
.A1(n_1730),
.A2(n_1425),
.B(n_1372),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1697),
.B(n_1642),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1665),
.Y(n_1825)
);

AND2x6_ASAP7_75t_L g1826 ( 
.A(n_1734),
.B(n_1643),
.Y(n_1826)
);

HB1xp67_ASAP7_75t_L g1827 ( 
.A(n_1655),
.Y(n_1827)
);

INVx1_ASAP7_75t_SL g1828 ( 
.A(n_1687),
.Y(n_1828)
);

INVx3_ASAP7_75t_L g1829 ( 
.A(n_1687),
.Y(n_1829)
);

OAI21x1_ASAP7_75t_L g1830 ( 
.A1(n_1686),
.A2(n_1379),
.B(n_1346),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1660),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1721),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1660),
.Y(n_1833)
);

HB1xp67_ASAP7_75t_L g1834 ( 
.A(n_1655),
.Y(n_1834)
);

AOI22xp33_ASAP7_75t_SL g1835 ( 
.A1(n_1707),
.A2(n_542),
.B1(n_555),
.B2(n_547),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1655),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1655),
.Y(n_1837)
);

BUFx3_ASAP7_75t_L g1838 ( 
.A(n_1690),
.Y(n_1838)
);

OAI22xp33_ASAP7_75t_L g1839 ( 
.A1(n_1707),
.A2(n_1612),
.B1(n_1658),
.B2(n_1656),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1660),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1699),
.Y(n_1841)
);

AO21x2_ASAP7_75t_L g1842 ( 
.A1(n_1737),
.A2(n_1612),
.B(n_1390),
.Y(n_1842)
);

HB1xp67_ASAP7_75t_L g1843 ( 
.A(n_1709),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1711),
.B(n_1642),
.Y(n_1844)
);

AO21x2_ASAP7_75t_L g1845 ( 
.A1(n_1709),
.A2(n_1391),
.B(n_1383),
.Y(n_1845)
);

HB1xp67_ASAP7_75t_L g1846 ( 
.A(n_1711),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1715),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1690),
.Y(n_1848)
);

AOI22xp33_ASAP7_75t_SL g1849 ( 
.A1(n_1734),
.A2(n_558),
.B1(n_562),
.B2(n_561),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1723),
.Y(n_1850)
);

AOI22xp33_ASAP7_75t_SL g1851 ( 
.A1(n_1731),
.A2(n_569),
.B1(n_580),
.B2(n_579),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1708),
.Y(n_1852)
);

HB1xp67_ASAP7_75t_L g1853 ( 
.A(n_1705),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1728),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1732),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1708),
.Y(n_1856)
);

OAI22xp33_ASAP7_75t_L g1857 ( 
.A1(n_1731),
.A2(n_1645),
.B1(n_1638),
.B2(n_1628),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1736),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1693),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1693),
.Y(n_1860)
);

INVx2_ASAP7_75t_SL g1861 ( 
.A(n_1664),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1653),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1681),
.Y(n_1863)
);

CKINVDCx5p33_ASAP7_75t_R g1864 ( 
.A(n_1688),
.Y(n_1864)
);

INVx2_ASAP7_75t_L g1865 ( 
.A(n_1681),
.Y(n_1865)
);

BUFx6f_ASAP7_75t_L g1866 ( 
.A(n_1696),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1653),
.Y(n_1867)
);

AOI21x1_ASAP7_75t_L g1868 ( 
.A1(n_1668),
.A2(n_1396),
.B(n_1392),
.Y(n_1868)
);

AO21x2_ASAP7_75t_L g1869 ( 
.A1(n_1652),
.A2(n_1645),
.B(n_1638),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1675),
.B(n_1646),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1675),
.B(n_1646),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1681),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1653),
.Y(n_1873)
);

INVx3_ASAP7_75t_L g1874 ( 
.A(n_1703),
.Y(n_1874)
);

OR2x2_ASAP7_75t_L g1875 ( 
.A(n_1714),
.B(n_1647),
.Y(n_1875)
);

OAI21x1_ASAP7_75t_L g1876 ( 
.A1(n_1700),
.A2(n_1645),
.B(n_1638),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1653),
.Y(n_1877)
);

INVx3_ASAP7_75t_L g1878 ( 
.A(n_1703),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1653),
.Y(n_1879)
);

BUFx3_ASAP7_75t_L g1880 ( 
.A(n_1696),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1653),
.Y(n_1881)
);

BUFx6f_ASAP7_75t_L g1882 ( 
.A(n_1696),
.Y(n_1882)
);

BUFx3_ASAP7_75t_L g1883 ( 
.A(n_1696),
.Y(n_1883)
);

BUFx3_ASAP7_75t_L g1884 ( 
.A(n_1696),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1653),
.Y(n_1885)
);

INVx2_ASAP7_75t_SL g1886 ( 
.A(n_1664),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1653),
.Y(n_1887)
);

HB1xp67_ASAP7_75t_L g1888 ( 
.A(n_1803),
.Y(n_1888)
);

CKINVDCx5p33_ASAP7_75t_R g1889 ( 
.A(n_1752),
.Y(n_1889)
);

HB1xp67_ASAP7_75t_L g1890 ( 
.A(n_1803),
.Y(n_1890)
);

HB1xp67_ASAP7_75t_L g1891 ( 
.A(n_1814),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1809),
.Y(n_1892)
);

AND2x4_ASAP7_75t_L g1893 ( 
.A(n_1774),
.B(n_1643),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1764),
.B(n_1643),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1809),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1764),
.B(n_1643),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1739),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1741),
.Y(n_1898)
);

CKINVDCx5p33_ASAP7_75t_R g1899 ( 
.A(n_1864),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1747),
.Y(n_1900)
);

INVx2_ASAP7_75t_L g1901 ( 
.A(n_1811),
.Y(n_1901)
);

NOR2xp33_ASAP7_75t_R g1902 ( 
.A(n_1761),
.B(n_1245),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1782),
.B(n_1643),
.Y(n_1903)
);

NOR3xp33_ASAP7_75t_SL g1904 ( 
.A(n_1751),
.B(n_585),
.C(n_582),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1811),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1748),
.Y(n_1906)
);

NAND2xp33_ASAP7_75t_R g1907 ( 
.A(n_1773),
.B(n_0),
.Y(n_1907)
);

CKINVDCx16_ASAP7_75t_R g1908 ( 
.A(n_1880),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1758),
.Y(n_1909)
);

AOI22xp33_ASAP7_75t_L g1910 ( 
.A1(n_1835),
.A2(n_659),
.B1(n_668),
.B2(n_471),
.Y(n_1910)
);

NAND2xp33_ASAP7_75t_R g1911 ( 
.A(n_1786),
.B(n_1),
.Y(n_1911)
);

NAND2xp33_ASAP7_75t_SL g1912 ( 
.A(n_1783),
.B(n_1800),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1816),
.Y(n_1913)
);

BUFx3_ASAP7_75t_L g1914 ( 
.A(n_1754),
.Y(n_1914)
);

NOR2xp33_ASAP7_75t_L g1915 ( 
.A(n_1754),
.B(n_1644),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1815),
.B(n_1647),
.Y(n_1916)
);

BUFx4f_ASAP7_75t_SL g1917 ( 
.A(n_1750),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1846),
.B(n_1647),
.Y(n_1918)
);

BUFx6f_ASAP7_75t_L g1919 ( 
.A(n_1866),
.Y(n_1919)
);

NAND2xp33_ASAP7_75t_R g1920 ( 
.A(n_1787),
.B(n_2),
.Y(n_1920)
);

CKINVDCx5p33_ASAP7_75t_R g1921 ( 
.A(n_1750),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1774),
.B(n_1646),
.Y(n_1922)
);

CKINVDCx5p33_ASAP7_75t_R g1923 ( 
.A(n_1743),
.Y(n_1923)
);

INVx3_ASAP7_75t_L g1924 ( 
.A(n_1787),
.Y(n_1924)
);

HB1xp67_ASAP7_75t_L g1925 ( 
.A(n_1816),
.Y(n_1925)
);

BUFx3_ASAP7_75t_L g1926 ( 
.A(n_1777),
.Y(n_1926)
);

BUFx2_ASAP7_75t_L g1927 ( 
.A(n_1796),
.Y(n_1927)
);

NAND2xp33_ASAP7_75t_R g1928 ( 
.A(n_1874),
.B(n_3),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_L g1929 ( 
.A(n_1846),
.B(n_587),
.Y(n_1929)
);

NAND3xp33_ASAP7_75t_SL g1930 ( 
.A(n_1783),
.B(n_590),
.C(n_588),
.Y(n_1930)
);

OR2x6_ASAP7_75t_L g1931 ( 
.A(n_1744),
.B(n_1625),
.Y(n_1931)
);

BUFx2_ASAP7_75t_L g1932 ( 
.A(n_1796),
.Y(n_1932)
);

OR2x6_ASAP7_75t_L g1933 ( 
.A(n_1807),
.B(n_1628),
.Y(n_1933)
);

INVxp67_ASAP7_75t_L g1934 ( 
.A(n_1861),
.Y(n_1934)
);

NOR2xp33_ASAP7_75t_R g1935 ( 
.A(n_1740),
.B(n_1245),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1765),
.Y(n_1936)
);

NAND2xp33_ASAP7_75t_R g1937 ( 
.A(n_1874),
.B(n_3),
.Y(n_1937)
);

AND2x4_ASAP7_75t_L g1938 ( 
.A(n_1878),
.B(n_1629),
.Y(n_1938)
);

BUFx10_ASAP7_75t_L g1939 ( 
.A(n_1866),
.Y(n_1939)
);

BUFx3_ASAP7_75t_L g1940 ( 
.A(n_1777),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1862),
.Y(n_1941)
);

CKINVDCx16_ASAP7_75t_R g1942 ( 
.A(n_1880),
.Y(n_1942)
);

NAND2xp33_ASAP7_75t_R g1943 ( 
.A(n_1878),
.B(n_6),
.Y(n_1943)
);

AND2x6_ASAP7_75t_SL g1944 ( 
.A(n_1740),
.B(n_1303),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1867),
.Y(n_1945)
);

CKINVDCx5p33_ASAP7_75t_R g1946 ( 
.A(n_1756),
.Y(n_1946)
);

AND2x4_ASAP7_75t_L g1947 ( 
.A(n_1790),
.B(n_1629),
.Y(n_1947)
);

NAND2xp33_ASAP7_75t_R g1948 ( 
.A(n_1824),
.B(n_1875),
.Y(n_1948)
);

AND2x4_ASAP7_75t_SL g1949 ( 
.A(n_1886),
.B(n_1629),
.Y(n_1949)
);

AOI22xp33_ASAP7_75t_L g1950 ( 
.A1(n_1835),
.A2(n_668),
.B1(n_659),
.B2(n_1631),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1870),
.B(n_591),
.Y(n_1951)
);

OAI22xp5_ASAP7_75t_L g1952 ( 
.A1(n_1804),
.A2(n_1645),
.B1(n_1633),
.B2(n_1636),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1871),
.B(n_594),
.Y(n_1953)
);

AO21x2_ASAP7_75t_L g1954 ( 
.A1(n_1822),
.A2(n_1645),
.B(n_1633),
.Y(n_1954)
);

AND2x6_ASAP7_75t_L g1955 ( 
.A(n_1859),
.B(n_1631),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1770),
.B(n_1631),
.Y(n_1956)
);

NOR2xp33_ASAP7_75t_R g1957 ( 
.A(n_1866),
.B(n_1303),
.Y(n_1957)
);

BUFx4f_ASAP7_75t_SL g1958 ( 
.A(n_1883),
.Y(n_1958)
);

HB1xp67_ASAP7_75t_L g1959 ( 
.A(n_1821),
.Y(n_1959)
);

NAND2xp33_ASAP7_75t_R g1960 ( 
.A(n_1790),
.B(n_6),
.Y(n_1960)
);

NAND2xp33_ASAP7_75t_R g1961 ( 
.A(n_1759),
.B(n_7),
.Y(n_1961)
);

BUFx2_ASAP7_75t_L g1962 ( 
.A(n_1746),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1769),
.B(n_598),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1873),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1877),
.Y(n_1965)
);

AOI22xp33_ASAP7_75t_L g1966 ( 
.A1(n_1800),
.A2(n_668),
.B1(n_659),
.B2(n_1633),
.Y(n_1966)
);

CKINVDCx16_ASAP7_75t_R g1967 ( 
.A(n_1883),
.Y(n_1967)
);

AOI22xp33_ASAP7_75t_SL g1968 ( 
.A1(n_1738),
.A2(n_1860),
.B1(n_1751),
.B2(n_1795),
.Y(n_1968)
);

NOR2xp33_ASAP7_75t_R g1969 ( 
.A(n_1866),
.B(n_1636),
.Y(n_1969)
);

NAND2xp33_ASAP7_75t_R g1970 ( 
.A(n_1742),
.B(n_7),
.Y(n_1970)
);

INVx2_ASAP7_75t_L g1971 ( 
.A(n_1821),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1767),
.B(n_1636),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1771),
.B(n_604),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1806),
.B(n_605),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1879),
.Y(n_1975)
);

AOI22xp33_ASAP7_75t_L g1976 ( 
.A1(n_1745),
.A2(n_668),
.B1(n_659),
.B2(n_1637),
.Y(n_1976)
);

AO21x1_ASAP7_75t_L g1977 ( 
.A1(n_1839),
.A2(n_8),
.B(n_9),
.Y(n_1977)
);

NOR2xp33_ASAP7_75t_R g1978 ( 
.A(n_1882),
.B(n_1637),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1881),
.Y(n_1979)
);

CKINVDCx5p33_ASAP7_75t_R g1980 ( 
.A(n_1884),
.Y(n_1980)
);

NOR2xp33_ASAP7_75t_R g1981 ( 
.A(n_1882),
.B(n_1637),
.Y(n_1981)
);

CKINVDCx5p33_ASAP7_75t_R g1982 ( 
.A(n_1884),
.Y(n_1982)
);

BUFx3_ASAP7_75t_L g1983 ( 
.A(n_1882),
.Y(n_1983)
);

NOR2xp33_ASAP7_75t_R g1984 ( 
.A(n_1882),
.B(n_1639),
.Y(n_1984)
);

AND2x4_ASAP7_75t_SL g1985 ( 
.A(n_1844),
.B(n_1639),
.Y(n_1985)
);

OR2x4_ASAP7_75t_L g1986 ( 
.A(n_1753),
.B(n_659),
.Y(n_1986)
);

NOR2xp33_ASAP7_75t_R g1987 ( 
.A(n_1793),
.B(n_1639),
.Y(n_1987)
);

NAND2xp33_ASAP7_75t_R g1988 ( 
.A(n_1818),
.B(n_8),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1789),
.B(n_1805),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1885),
.Y(n_1990)
);

NAND2xp33_ASAP7_75t_R g1991 ( 
.A(n_1818),
.B(n_10),
.Y(n_1991)
);

OAI22xp5_ASAP7_75t_L g1992 ( 
.A1(n_1804),
.A2(n_609),
.B1(n_611),
.B2(n_606),
.Y(n_1992)
);

OAI21xp5_ASAP7_75t_L g1993 ( 
.A1(n_1745),
.A2(n_647),
.B(n_642),
.Y(n_1993)
);

AND2x2_ASAP7_75t_L g1994 ( 
.A(n_1749),
.B(n_10),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1749),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1760),
.B(n_12),
.Y(n_1996)
);

HB1xp67_ASAP7_75t_L g1997 ( 
.A(n_1812),
.Y(n_1997)
);

OAI22xp33_ASAP7_75t_L g1998 ( 
.A1(n_1839),
.A2(n_676),
.B1(n_614),
.B2(n_647),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1760),
.B(n_12),
.Y(n_1999)
);

OR2x2_ASAP7_75t_L g2000 ( 
.A(n_1812),
.B(n_13),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1791),
.B(n_13),
.Y(n_2001)
);

OR2x2_ASAP7_75t_L g2002 ( 
.A(n_1763),
.B(n_14),
.Y(n_2002)
);

CKINVDCx5p33_ASAP7_75t_R g2003 ( 
.A(n_1776),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1887),
.Y(n_2004)
);

NAND2xp33_ASAP7_75t_SL g2005 ( 
.A(n_1810),
.B(n_642),
.Y(n_2005)
);

CKINVDCx11_ASAP7_75t_R g2006 ( 
.A(n_1828),
.Y(n_2006)
);

AO31x2_ASAP7_75t_L g2007 ( 
.A1(n_1836),
.A2(n_19),
.A3(n_14),
.B(n_15),
.Y(n_2007)
);

NOR2xp33_ASAP7_75t_R g2008 ( 
.A(n_1829),
.B(n_15),
.Y(n_2008)
);

NAND4xp25_ASAP7_75t_L g2009 ( 
.A(n_1810),
.B(n_21),
.C(n_19),
.D(n_20),
.Y(n_2009)
);

CKINVDCx5p33_ASAP7_75t_R g2010 ( 
.A(n_1838),
.Y(n_2010)
);

NOR2xp33_ASAP7_75t_R g2011 ( 
.A(n_1829),
.B(n_21),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1802),
.B(n_22),
.Y(n_2012)
);

AND2x4_ASAP7_75t_L g2013 ( 
.A(n_1746),
.B(n_1141),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1763),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1768),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1860),
.B(n_22),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1768),
.Y(n_2017)
);

CKINVDCx8_ASAP7_75t_R g2018 ( 
.A(n_1826),
.Y(n_2018)
);

AOI22xp33_ASAP7_75t_L g2019 ( 
.A1(n_1820),
.A2(n_650),
.B1(n_655),
.B2(n_649),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1863),
.B(n_23),
.Y(n_2020)
);

OR2x2_ASAP7_75t_L g2021 ( 
.A(n_1863),
.B(n_23),
.Y(n_2021)
);

NOR2xp33_ASAP7_75t_R g2022 ( 
.A(n_1838),
.B(n_24),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_1865),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1779),
.B(n_25),
.Y(n_2024)
);

INVx3_ASAP7_75t_L g2025 ( 
.A(n_1755),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_1865),
.Y(n_2026)
);

AND2x2_ASAP7_75t_L g2027 ( 
.A(n_1872),
.B(n_26),
.Y(n_2027)
);

INVx3_ASAP7_75t_L g2028 ( 
.A(n_1755),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1872),
.Y(n_2029)
);

NOR3xp33_ASAP7_75t_SL g2030 ( 
.A(n_1797),
.B(n_650),
.C(n_649),
.Y(n_2030)
);

NOR2xp33_ASAP7_75t_L g2031 ( 
.A(n_1986),
.B(n_1798),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1924),
.B(n_1779),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1897),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_1924),
.B(n_1780),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1894),
.B(n_1780),
.Y(n_2035)
);

AND2x2_ASAP7_75t_L g2036 ( 
.A(n_1927),
.B(n_1781),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_1932),
.B(n_1781),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1898),
.Y(n_2038)
);

OR2x2_ASAP7_75t_L g2039 ( 
.A(n_1888),
.B(n_1843),
.Y(n_2039)
);

AOI22xp5_ASAP7_75t_L g2040 ( 
.A1(n_1912),
.A2(n_1797),
.B1(n_1820),
.B2(n_1817),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_1892),
.Y(n_2041)
);

AND2x4_ASAP7_75t_L g2042 ( 
.A(n_1962),
.B(n_1746),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1895),
.Y(n_2043)
);

INVx2_ASAP7_75t_L g2044 ( 
.A(n_1901),
.Y(n_2044)
);

AND2x2_ASAP7_75t_L g2045 ( 
.A(n_1989),
.B(n_1799),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1900),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1906),
.Y(n_2047)
);

INVx2_ASAP7_75t_L g2048 ( 
.A(n_1905),
.Y(n_2048)
);

INVx2_ASAP7_75t_SL g2049 ( 
.A(n_1890),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_1896),
.B(n_1799),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1909),
.Y(n_2051)
);

INVx2_ASAP7_75t_L g2052 ( 
.A(n_1913),
.Y(n_2052)
);

AND2x4_ASAP7_75t_L g2053 ( 
.A(n_1933),
.B(n_1850),
.Y(n_2053)
);

OR2x2_ASAP7_75t_L g2054 ( 
.A(n_1925),
.B(n_1843),
.Y(n_2054)
);

AND2x4_ASAP7_75t_L g2055 ( 
.A(n_1933),
.B(n_1825),
.Y(n_2055)
);

INVx2_ASAP7_75t_L g2056 ( 
.A(n_1971),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_1903),
.B(n_1908),
.Y(n_2057)
);

AND2x4_ASAP7_75t_L g2058 ( 
.A(n_1933),
.B(n_1848),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1936),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1941),
.Y(n_2060)
);

HB1xp67_ASAP7_75t_L g2061 ( 
.A(n_1959),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_1942),
.B(n_1853),
.Y(n_2062)
);

OA21x2_ASAP7_75t_L g2063 ( 
.A1(n_2001),
.A2(n_1833),
.B(n_1831),
.Y(n_2063)
);

INVxp67_ASAP7_75t_L g2064 ( 
.A(n_1961),
.Y(n_2064)
);

HB1xp67_ASAP7_75t_L g2065 ( 
.A(n_1997),
.Y(n_2065)
);

NAND3xp33_ASAP7_75t_L g2066 ( 
.A(n_1968),
.B(n_1847),
.C(n_1849),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_1894),
.B(n_1766),
.Y(n_2067)
);

OR2x2_ASAP7_75t_L g2068 ( 
.A(n_1891),
.B(n_1853),
.Y(n_2068)
);

AND2x2_ASAP7_75t_L g2069 ( 
.A(n_1967),
.B(n_1801),
.Y(n_2069)
);

AND2x2_ASAP7_75t_L g2070 ( 
.A(n_1934),
.B(n_1801),
.Y(n_2070)
);

NOR2x1_ASAP7_75t_SL g2071 ( 
.A(n_1931),
.B(n_1766),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_1985),
.B(n_1922),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1945),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_1995),
.B(n_1832),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1964),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_2014),
.Y(n_2076)
);

OR2x6_ASAP7_75t_L g2077 ( 
.A(n_1931),
.B(n_1808),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_1965),
.B(n_1852),
.Y(n_2078)
);

INVx3_ASAP7_75t_L g2079 ( 
.A(n_2025),
.Y(n_2079)
);

INVx2_ASAP7_75t_SL g2080 ( 
.A(n_2010),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1975),
.Y(n_2081)
);

OR2x2_ASAP7_75t_L g2082 ( 
.A(n_2015),
.B(n_1772),
.Y(n_2082)
);

OR2x2_ASAP7_75t_L g2083 ( 
.A(n_2029),
.B(n_1772),
.Y(n_2083)
);

INVxp67_ASAP7_75t_L g2084 ( 
.A(n_1970),
.Y(n_2084)
);

INVx2_ASAP7_75t_L g2085 ( 
.A(n_2017),
.Y(n_2085)
);

AND2x2_ASAP7_75t_L g2086 ( 
.A(n_2023),
.B(n_1845),
.Y(n_2086)
);

OR2x2_ASAP7_75t_L g2087 ( 
.A(n_2026),
.B(n_1785),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1979),
.Y(n_2088)
);

NOR2xp33_ASAP7_75t_L g2089 ( 
.A(n_1986),
.B(n_1757),
.Y(n_2089)
);

OR2x6_ASAP7_75t_L g2090 ( 
.A(n_1931),
.B(n_1808),
.Y(n_2090)
);

HB1xp67_ASAP7_75t_L g2091 ( 
.A(n_1990),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_2004),
.Y(n_2092)
);

HB1xp67_ASAP7_75t_L g2093 ( 
.A(n_1954),
.Y(n_2093)
);

INVx3_ASAP7_75t_SL g2094 ( 
.A(n_1921),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_1947),
.B(n_1845),
.Y(n_2095)
);

OR2x2_ASAP7_75t_L g2096 ( 
.A(n_1918),
.B(n_1785),
.Y(n_2096)
);

INVx2_ASAP7_75t_L g2097 ( 
.A(n_1954),
.Y(n_2097)
);

NOR2xp33_ASAP7_75t_L g2098 ( 
.A(n_1929),
.B(n_1856),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_2002),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_2021),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_2001),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2012),
.Y(n_2102)
);

AND2x2_ASAP7_75t_L g2103 ( 
.A(n_1947),
.B(n_1841),
.Y(n_2103)
);

AND2x2_ASAP7_75t_SL g2104 ( 
.A(n_1948),
.B(n_1792),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_2012),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_2000),
.Y(n_2106)
);

OAI22xp5_ASAP7_75t_L g2107 ( 
.A1(n_1966),
.A2(n_1851),
.B1(n_1849),
.B2(n_1784),
.Y(n_2107)
);

AND2x2_ASAP7_75t_L g2108 ( 
.A(n_2006),
.B(n_1792),
.Y(n_2108)
);

INVx2_ASAP7_75t_L g2109 ( 
.A(n_2025),
.Y(n_2109)
);

NAND2x1_ASAP7_75t_L g2110 ( 
.A(n_1955),
.B(n_1826),
.Y(n_2110)
);

OR2x2_ASAP7_75t_L g2111 ( 
.A(n_1916),
.B(n_1837),
.Y(n_2111)
);

NOR2xp33_ASAP7_75t_R g2112 ( 
.A(n_1920),
.B(n_1868),
.Y(n_2112)
);

AND2x2_ASAP7_75t_L g2113 ( 
.A(n_1893),
.B(n_1854),
.Y(n_2113)
);

INVx1_ASAP7_75t_L g2114 ( 
.A(n_2028),
.Y(n_2114)
);

AND2x2_ASAP7_75t_L g2115 ( 
.A(n_1893),
.B(n_1972),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_2028),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2024),
.Y(n_2117)
);

HB1xp67_ASAP7_75t_L g2118 ( 
.A(n_2007),
.Y(n_2118)
);

INVx3_ASAP7_75t_L g2119 ( 
.A(n_2018),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_1994),
.Y(n_2120)
);

INVx2_ASAP7_75t_L g2121 ( 
.A(n_2007),
.Y(n_2121)
);

INVx2_ASAP7_75t_L g2122 ( 
.A(n_2007),
.Y(n_2122)
);

AND2x2_ASAP7_75t_L g2123 ( 
.A(n_1938),
.B(n_1914),
.Y(n_2123)
);

INVx2_ASAP7_75t_L g2124 ( 
.A(n_1996),
.Y(n_2124)
);

AND2x2_ASAP7_75t_L g2125 ( 
.A(n_1938),
.B(n_1854),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_1999),
.Y(n_2126)
);

AOI21xp5_ASAP7_75t_L g2127 ( 
.A1(n_1910),
.A2(n_1857),
.B(n_1762),
.Y(n_2127)
);

INVx2_ASAP7_75t_SL g2128 ( 
.A(n_1949),
.Y(n_2128)
);

INVx8_ASAP7_75t_L g2129 ( 
.A(n_1944),
.Y(n_2129)
);

AO31x2_ASAP7_75t_L g2130 ( 
.A1(n_1977),
.A2(n_1831),
.A3(n_1840),
.B(n_1833),
.Y(n_2130)
);

AND2x2_ASAP7_75t_L g2131 ( 
.A(n_1956),
.B(n_1855),
.Y(n_2131)
);

BUFx3_ASAP7_75t_L g2132 ( 
.A(n_1926),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2020),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_2027),
.Y(n_2134)
);

INVx2_ASAP7_75t_L g2135 ( 
.A(n_1955),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_1955),
.Y(n_2136)
);

OAI31xp33_ASAP7_75t_L g2137 ( 
.A1(n_2009),
.A2(n_1857),
.A3(n_1834),
.B(n_1827),
.Y(n_2137)
);

BUFx2_ASAP7_75t_L g2138 ( 
.A(n_1955),
.Y(n_2138)
);

INVx3_ASAP7_75t_L g2139 ( 
.A(n_1939),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1974),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1963),
.Y(n_2141)
);

AND2x2_ASAP7_75t_L g2142 ( 
.A(n_1983),
.B(n_1855),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_1951),
.B(n_1762),
.Y(n_2143)
);

BUFx2_ASAP7_75t_L g2144 ( 
.A(n_1969),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_1973),
.Y(n_2145)
);

AND2x2_ASAP7_75t_L g2146 ( 
.A(n_2003),
.B(n_1858),
.Y(n_2146)
);

OAI22xp5_ASAP7_75t_L g2147 ( 
.A1(n_1950),
.A2(n_1851),
.B1(n_1813),
.B2(n_1775),
.Y(n_2147)
);

OR2x2_ASAP7_75t_L g2148 ( 
.A(n_1953),
.B(n_1827),
.Y(n_2148)
);

AOI22xp33_ASAP7_75t_L g2149 ( 
.A1(n_2009),
.A2(n_1993),
.B1(n_2005),
.B2(n_1930),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_2016),
.Y(n_2150)
);

HB1xp67_ASAP7_75t_L g2151 ( 
.A(n_1987),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_1919),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_1919),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_1919),
.Y(n_2154)
);

CKINVDCx5p33_ASAP7_75t_R g2155 ( 
.A(n_1946),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_1939),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2013),
.Y(n_2157)
);

AO31x2_ASAP7_75t_L g2158 ( 
.A1(n_1952),
.A2(n_1840),
.A3(n_1834),
.B(n_1794),
.Y(n_2158)
);

AND2x2_ASAP7_75t_L g2159 ( 
.A(n_1940),
.B(n_1869),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_1889),
.B(n_1869),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_2013),
.Y(n_2161)
);

HB1xp67_ASAP7_75t_L g2162 ( 
.A(n_1928),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2022),
.Y(n_2163)
);

AOI22xp33_ASAP7_75t_L g2164 ( 
.A1(n_1993),
.A2(n_658),
.B1(n_665),
.B2(n_655),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_1952),
.B(n_1826),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_1998),
.B(n_1826),
.Y(n_2166)
);

INVx2_ASAP7_75t_L g2167 ( 
.A(n_1958),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2008),
.Y(n_2168)
);

AND2x2_ASAP7_75t_L g2169 ( 
.A(n_1980),
.B(n_1876),
.Y(n_2169)
);

INVx3_ASAP7_75t_L g2170 ( 
.A(n_1917),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2091),
.Y(n_2171)
);

INVx2_ASAP7_75t_L g2172 ( 
.A(n_2109),
.Y(n_2172)
);

BUFx6f_ASAP7_75t_L g2173 ( 
.A(n_2094),
.Y(n_2173)
);

AOI21xp5_ASAP7_75t_L g2174 ( 
.A1(n_2107),
.A2(n_1976),
.B(n_1915),
.Y(n_2174)
);

NAND2x1p5_ASAP7_75t_SL g2175 ( 
.A(n_2159),
.B(n_1960),
.Y(n_2175)
);

OAI21xp5_ASAP7_75t_L g2176 ( 
.A1(n_2066),
.A2(n_2084),
.B(n_2162),
.Y(n_2176)
);

AO21x2_ASAP7_75t_L g2177 ( 
.A1(n_2093),
.A2(n_2011),
.B(n_1819),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2091),
.Y(n_2178)
);

INVx1_ASAP7_75t_L g2179 ( 
.A(n_2092),
.Y(n_2179)
);

INVxp67_ASAP7_75t_L g2180 ( 
.A(n_2162),
.Y(n_2180)
);

INVx2_ASAP7_75t_SL g2181 ( 
.A(n_2132),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2092),
.Y(n_2182)
);

OAI22xp33_ASAP7_75t_L g2183 ( 
.A1(n_2040),
.A2(n_1943),
.B1(n_1937),
.B2(n_1911),
.Y(n_2183)
);

INVxp67_ASAP7_75t_L g2184 ( 
.A(n_2098),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_2033),
.Y(n_2185)
);

INVx3_ASAP7_75t_L g2186 ( 
.A(n_2079),
.Y(n_2186)
);

AOI21xp5_ASAP7_75t_L g2187 ( 
.A1(n_2104),
.A2(n_1992),
.B(n_2019),
.Y(n_2187)
);

INVx2_ASAP7_75t_L g2188 ( 
.A(n_2109),
.Y(n_2188)
);

BUFx2_ASAP7_75t_L g2189 ( 
.A(n_2151),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_2038),
.Y(n_2190)
);

NAND4xp25_ASAP7_75t_L g2191 ( 
.A(n_2149),
.B(n_1907),
.C(n_1991),
.D(n_1988),
.Y(n_2191)
);

AOI21xp5_ASAP7_75t_L g2192 ( 
.A1(n_2104),
.A2(n_1992),
.B(n_1788),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2046),
.Y(n_2193)
);

INVx3_ASAP7_75t_L g2194 ( 
.A(n_2079),
.Y(n_2194)
);

OAI21x1_ASAP7_75t_L g2195 ( 
.A1(n_2110),
.A2(n_1778),
.B(n_1823),
.Y(n_2195)
);

OAI22xp5_ASAP7_75t_L g2196 ( 
.A1(n_2149),
.A2(n_1904),
.B1(n_2030),
.B2(n_1982),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2047),
.Y(n_2197)
);

OAI21x1_ASAP7_75t_L g2198 ( 
.A1(n_2097),
.A2(n_1830),
.B(n_1978),
.Y(n_2198)
);

O2A1O1Ixp33_ASAP7_75t_L g2199 ( 
.A1(n_2084),
.A2(n_1944),
.B(n_1842),
.C(n_1957),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2051),
.Y(n_2200)
);

OAI22xp5_ASAP7_75t_L g2201 ( 
.A1(n_2064),
.A2(n_1899),
.B1(n_1923),
.B2(n_1981),
.Y(n_2201)
);

AOI22xp33_ASAP7_75t_SL g2202 ( 
.A1(n_2112),
.A2(n_1984),
.B1(n_1902),
.B2(n_1935),
.Y(n_2202)
);

AND2x2_ASAP7_75t_L g2203 ( 
.A(n_2062),
.B(n_1842),
.Y(n_2203)
);

OA21x2_ASAP7_75t_L g2204 ( 
.A1(n_2097),
.A2(n_665),
.B(n_658),
.Y(n_2204)
);

OAI21xp33_ASAP7_75t_SL g2205 ( 
.A1(n_2064),
.A2(n_1826),
.B(n_27),
.Y(n_2205)
);

BUFx3_ASAP7_75t_L g2206 ( 
.A(n_2170),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_2059),
.Y(n_2207)
);

INVx2_ASAP7_75t_L g2208 ( 
.A(n_2076),
.Y(n_2208)
);

OAI222xp33_ASAP7_75t_L g2209 ( 
.A1(n_2147),
.A2(n_675),
.B1(n_674),
.B2(n_669),
.C1(n_433),
.C2(n_435),
.Y(n_2209)
);

INVx3_ASAP7_75t_L g2210 ( 
.A(n_2058),
.Y(n_2210)
);

INVxp67_ASAP7_75t_SL g2211 ( 
.A(n_2061),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2060),
.Y(n_2212)
);

NOR2x1_ASAP7_75t_SL g2213 ( 
.A(n_2077),
.B(n_1141),
.Y(n_2213)
);

AO31x2_ASAP7_75t_L g2214 ( 
.A1(n_2121),
.A2(n_29),
.A3(n_27),
.B(n_28),
.Y(n_2214)
);

AOI211xp5_ASAP7_75t_L g2215 ( 
.A1(n_2137),
.A2(n_674),
.B(n_675),
.C(n_669),
.Y(n_2215)
);

AND2x4_ASAP7_75t_L g2216 ( 
.A(n_2077),
.B(n_1141),
.Y(n_2216)
);

OAI21x1_ASAP7_75t_L g2217 ( 
.A1(n_2121),
.A2(n_1218),
.B(n_32),
.Y(n_2217)
);

AND2x2_ASAP7_75t_L g2218 ( 
.A(n_2108),
.B(n_32),
.Y(n_2218)
);

AOI21xp33_ASAP7_75t_L g2219 ( 
.A1(n_2143),
.A2(n_34),
.B(n_35),
.Y(n_2219)
);

INVx2_ASAP7_75t_L g2220 ( 
.A(n_2076),
.Y(n_2220)
);

BUFx3_ASAP7_75t_L g2221 ( 
.A(n_2170),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_2073),
.Y(n_2222)
);

AOI21xp5_ASAP7_75t_L g2223 ( 
.A1(n_2127),
.A2(n_427),
.B(n_426),
.Y(n_2223)
);

INVx2_ASAP7_75t_SL g2224 ( 
.A(n_2132),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2075),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2081),
.Y(n_2226)
);

AO31x2_ASAP7_75t_L g2227 ( 
.A1(n_2122),
.A2(n_39),
.A3(n_34),
.B(n_38),
.Y(n_2227)
);

INVx2_ASAP7_75t_L g2228 ( 
.A(n_2041),
.Y(n_2228)
);

OAI221xp5_ASAP7_75t_L g2229 ( 
.A1(n_2164),
.A2(n_428),
.B1(n_436),
.B2(n_438),
.C(n_440),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2088),
.Y(n_2230)
);

AO21x2_ASAP7_75t_L g2231 ( 
.A1(n_2093),
.A2(n_38),
.B(n_40),
.Y(n_2231)
);

AO31x2_ASAP7_75t_L g2232 ( 
.A1(n_2122),
.A2(n_43),
.A3(n_41),
.B(n_42),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_2150),
.B(n_41),
.Y(n_2233)
);

OAI211xp5_ASAP7_75t_L g2234 ( 
.A1(n_2112),
.A2(n_446),
.B(n_455),
.C(n_443),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2065),
.Y(n_2235)
);

INVx4_ASAP7_75t_L g2236 ( 
.A(n_2129),
.Y(n_2236)
);

INVx2_ASAP7_75t_L g2237 ( 
.A(n_2041),
.Y(n_2237)
);

INVx2_ASAP7_75t_L g2238 ( 
.A(n_2043),
.Y(n_2238)
);

OA21x2_ASAP7_75t_L g2239 ( 
.A1(n_2067),
.A2(n_464),
.B(n_463),
.Y(n_2239)
);

OA21x2_ASAP7_75t_L g2240 ( 
.A1(n_2053),
.A2(n_468),
.B(n_467),
.Y(n_2240)
);

AOI22xp33_ASAP7_75t_L g2241 ( 
.A1(n_2031),
.A2(n_473),
.B1(n_474),
.B2(n_470),
.Y(n_2241)
);

BUFx2_ASAP7_75t_L g2242 ( 
.A(n_2151),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2065),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2061),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2099),
.Y(n_2245)
);

OAI211xp5_ASAP7_75t_L g2246 ( 
.A1(n_2164),
.A2(n_483),
.B(n_484),
.C(n_475),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_2150),
.B(n_43),
.Y(n_2247)
);

OAI21xp33_ASAP7_75t_L g2248 ( 
.A1(n_2031),
.A2(n_490),
.B(n_486),
.Y(n_2248)
);

NAND4xp25_ASAP7_75t_L g2249 ( 
.A(n_2098),
.B(n_50),
.C(n_44),
.D(n_48),
.Y(n_2249)
);

INVx1_ASAP7_75t_L g2250 ( 
.A(n_2099),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_2101),
.B(n_48),
.Y(n_2251)
);

OAI22xp5_ASAP7_75t_SL g2252 ( 
.A1(n_2163),
.A2(n_1218),
.B1(n_52),
.B2(n_50),
.Y(n_2252)
);

OAI22xp33_ASAP7_75t_L g2253 ( 
.A1(n_2165),
.A2(n_496),
.B1(n_501),
.B2(n_493),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2100),
.Y(n_2254)
);

INVx1_ASAP7_75t_SL g2255 ( 
.A(n_2068),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_2100),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2078),
.Y(n_2257)
);

INVx2_ASAP7_75t_SL g2258 ( 
.A(n_2069),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2082),
.Y(n_2259)
);

NAND3xp33_ASAP7_75t_L g2260 ( 
.A(n_2118),
.B(n_509),
.C(n_508),
.Y(n_2260)
);

INVx1_ASAP7_75t_SL g2261 ( 
.A(n_2094),
.Y(n_2261)
);

AOI21xp33_ASAP7_75t_L g2262 ( 
.A1(n_2089),
.A2(n_51),
.B(n_52),
.Y(n_2262)
);

AOI22xp33_ASAP7_75t_L g2263 ( 
.A1(n_2089),
.A2(n_515),
.B1(n_516),
.B2(n_513),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_L g2264 ( 
.A(n_2102),
.B(n_2105),
.Y(n_2264)
);

HB1xp67_ASAP7_75t_L g2265 ( 
.A(n_2049),
.Y(n_2265)
);

OA21x2_ASAP7_75t_L g2266 ( 
.A1(n_2053),
.A2(n_518),
.B(n_517),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_2043),
.Y(n_2267)
);

INVx2_ASAP7_75t_L g2268 ( 
.A(n_2044),
.Y(n_2268)
);

OR2x2_ASAP7_75t_L g2269 ( 
.A(n_2148),
.B(n_53),
.Y(n_2269)
);

NAND3xp33_ASAP7_75t_L g2270 ( 
.A(n_2118),
.B(n_527),
.C(n_520),
.Y(n_2270)
);

A2O1A1Ixp33_ASAP7_75t_L g2271 ( 
.A1(n_2129),
.A2(n_2127),
.B(n_2166),
.C(n_2168),
.Y(n_2271)
);

OAI21x1_ASAP7_75t_L g2272 ( 
.A1(n_2086),
.A2(n_1218),
.B(n_53),
.Y(n_2272)
);

OR2x2_ASAP7_75t_L g2273 ( 
.A(n_2096),
.B(n_2106),
.Y(n_2273)
);

INVx2_ASAP7_75t_L g2274 ( 
.A(n_2044),
.Y(n_2274)
);

BUFx3_ASAP7_75t_L g2275 ( 
.A(n_2167),
.Y(n_2275)
);

NAND2xp5_ASAP7_75t_L g2276 ( 
.A(n_2117),
.B(n_56),
.Y(n_2276)
);

OAI221xp5_ASAP7_75t_L g2277 ( 
.A1(n_2140),
.A2(n_528),
.B1(n_533),
.B2(n_543),
.C(n_549),
.Y(n_2277)
);

INVxp67_ASAP7_75t_SL g2278 ( 
.A(n_2049),
.Y(n_2278)
);

OAI211xp5_ASAP7_75t_L g2279 ( 
.A1(n_2129),
.A2(n_550),
.B(n_557),
.C(n_559),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_L g2280 ( 
.A(n_2141),
.B(n_2145),
.Y(n_2280)
);

OA21x2_ASAP7_75t_L g2281 ( 
.A1(n_2053),
.A2(n_567),
.B(n_566),
.Y(n_2281)
);

AOI22xp5_ASAP7_75t_L g2282 ( 
.A1(n_2119),
.A2(n_575),
.B1(n_592),
.B2(n_593),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2083),
.Y(n_2283)
);

AND2x2_ASAP7_75t_L g2284 ( 
.A(n_2057),
.B(n_56),
.Y(n_2284)
);

AND2x2_ASAP7_75t_L g2285 ( 
.A(n_2160),
.B(n_57),
.Y(n_2285)
);

INVxp67_ASAP7_75t_L g2286 ( 
.A(n_2124),
.Y(n_2286)
);

OAI22xp33_ASAP7_75t_L g2287 ( 
.A1(n_2119),
.A2(n_595),
.B1(n_597),
.B2(n_603),
.Y(n_2287)
);

BUFx2_ASAP7_75t_L g2288 ( 
.A(n_2144),
.Y(n_2288)
);

NAND2xp5_ASAP7_75t_L g2289 ( 
.A(n_2124),
.B(n_57),
.Y(n_2289)
);

OAI21x1_ASAP7_75t_L g2290 ( 
.A1(n_2135),
.A2(n_58),
.B(n_59),
.Y(n_2290)
);

INVx1_ASAP7_75t_L g2291 ( 
.A(n_2048),
.Y(n_2291)
);

HB1xp67_ASAP7_75t_L g2292 ( 
.A(n_2180),
.Y(n_2292)
);

AOI211xp5_ASAP7_75t_SL g2293 ( 
.A1(n_2183),
.A2(n_2167),
.B(n_2156),
.C(n_2139),
.Y(n_2293)
);

AND2x2_ASAP7_75t_L g2294 ( 
.A(n_2288),
.B(n_2169),
.Y(n_2294)
);

HB1xp67_ASAP7_75t_L g2295 ( 
.A(n_2189),
.Y(n_2295)
);

OR2x2_ASAP7_75t_L g2296 ( 
.A(n_2273),
.B(n_2134),
.Y(n_2296)
);

AND2x2_ASAP7_75t_L g2297 ( 
.A(n_2242),
.B(n_2258),
.Y(n_2297)
);

HB1xp67_ASAP7_75t_L g2298 ( 
.A(n_2211),
.Y(n_2298)
);

AND2x2_ASAP7_75t_L g2299 ( 
.A(n_2210),
.B(n_2042),
.Y(n_2299)
);

OAI321xp33_ASAP7_75t_L g2300 ( 
.A1(n_2176),
.A2(n_2090),
.A3(n_2077),
.B1(n_2116),
.B2(n_2114),
.C(n_2153),
.Y(n_2300)
);

BUFx2_ASAP7_75t_L g2301 ( 
.A(n_2236),
.Y(n_2301)
);

BUFx3_ASAP7_75t_L g2302 ( 
.A(n_2173),
.Y(n_2302)
);

INVx2_ASAP7_75t_L g2303 ( 
.A(n_2210),
.Y(n_2303)
);

INVx2_ASAP7_75t_L g2304 ( 
.A(n_2186),
.Y(n_2304)
);

NAND2xp5_ASAP7_75t_L g2305 ( 
.A(n_2257),
.B(n_2063),
.Y(n_2305)
);

AOI221xp5_ASAP7_75t_L g2306 ( 
.A1(n_2191),
.A2(n_2120),
.B1(n_2126),
.B2(n_2133),
.C(n_2134),
.Y(n_2306)
);

HB1xp67_ASAP7_75t_L g2307 ( 
.A(n_2171),
.Y(n_2307)
);

CKINVDCx5p33_ASAP7_75t_R g2308 ( 
.A(n_2173),
.Y(n_2308)
);

INVx2_ASAP7_75t_L g2309 ( 
.A(n_2186),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_2185),
.Y(n_2310)
);

AND2x4_ASAP7_75t_L g2311 ( 
.A(n_2216),
.B(n_2090),
.Y(n_2311)
);

HB1xp67_ASAP7_75t_L g2312 ( 
.A(n_2178),
.Y(n_2312)
);

AND2x2_ASAP7_75t_L g2313 ( 
.A(n_2286),
.B(n_2042),
.Y(n_2313)
);

AND2x2_ASAP7_75t_L g2314 ( 
.A(n_2216),
.B(n_2042),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_2184),
.B(n_2063),
.Y(n_2315)
);

OR2x2_ASAP7_75t_L g2316 ( 
.A(n_2269),
.B(n_2255),
.Y(n_2316)
);

INVx2_ASAP7_75t_L g2317 ( 
.A(n_2194),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_2194),
.Y(n_2318)
);

OAI21x1_ASAP7_75t_L g2319 ( 
.A1(n_2198),
.A2(n_2087),
.B(n_2063),
.Y(n_2319)
);

AND2x2_ASAP7_75t_L g2320 ( 
.A(n_2236),
.B(n_2115),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2190),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2193),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2197),
.Y(n_2323)
);

HB1xp67_ASAP7_75t_L g2324 ( 
.A(n_2179),
.Y(n_2324)
);

AND2x4_ASAP7_75t_L g2325 ( 
.A(n_2213),
.B(n_2090),
.Y(n_2325)
);

AOI22xp33_ASAP7_75t_L g2326 ( 
.A1(n_2223),
.A2(n_2161),
.B1(n_2157),
.B2(n_2058),
.Y(n_2326)
);

AND2x2_ASAP7_75t_L g2327 ( 
.A(n_2181),
.B(n_2123),
.Y(n_2327)
);

AND2x2_ASAP7_75t_L g2328 ( 
.A(n_2224),
.B(n_2128),
.Y(n_2328)
);

AND2x2_ASAP7_75t_L g2329 ( 
.A(n_2255),
.B(n_2128),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_2235),
.B(n_2048),
.Y(n_2330)
);

AND2x4_ASAP7_75t_L g2331 ( 
.A(n_2275),
.B(n_2058),
.Y(n_2331)
);

AND2x4_ASAP7_75t_L g2332 ( 
.A(n_2206),
.B(n_2152),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_2243),
.B(n_2085),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_L g2334 ( 
.A(n_2244),
.B(n_2085),
.Y(n_2334)
);

AND2x2_ASAP7_75t_L g2335 ( 
.A(n_2221),
.B(n_2072),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_L g2336 ( 
.A(n_2200),
.B(n_2052),
.Y(n_2336)
);

NOR2xp33_ASAP7_75t_L g2337 ( 
.A(n_2173),
.B(n_2155),
.Y(n_2337)
);

INVx1_ASAP7_75t_L g2338 ( 
.A(n_2207),
.Y(n_2338)
);

BUFx2_ASAP7_75t_L g2339 ( 
.A(n_2175),
.Y(n_2339)
);

NAND3xp33_ASAP7_75t_L g2340 ( 
.A(n_2215),
.B(n_2095),
.C(n_2111),
.Y(n_2340)
);

AND2x4_ASAP7_75t_L g2341 ( 
.A(n_2278),
.B(n_2152),
.Y(n_2341)
);

AND2x2_ASAP7_75t_L g2342 ( 
.A(n_2203),
.B(n_2103),
.Y(n_2342)
);

HB1xp67_ASAP7_75t_L g2343 ( 
.A(n_2182),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_2212),
.B(n_2052),
.Y(n_2344)
);

INVx2_ASAP7_75t_L g2345 ( 
.A(n_2172),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2222),
.Y(n_2346)
);

OR2x2_ASAP7_75t_L g2347 ( 
.A(n_2259),
.B(n_2039),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_L g2348 ( 
.A(n_2225),
.B(n_2056),
.Y(n_2348)
);

NAND3xp33_ASAP7_75t_L g2349 ( 
.A(n_2215),
.B(n_2154),
.C(n_2146),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2226),
.Y(n_2350)
);

INVx2_ASAP7_75t_SL g2351 ( 
.A(n_2261),
.Y(n_2351)
);

AND2x2_ASAP7_75t_L g2352 ( 
.A(n_2245),
.B(n_2070),
.Y(n_2352)
);

INVx1_ASAP7_75t_L g2353 ( 
.A(n_2230),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2250),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2254),
.Y(n_2355)
);

INVx4_ASAP7_75t_L g2356 ( 
.A(n_2231),
.Y(n_2356)
);

BUFx2_ASAP7_75t_L g2357 ( 
.A(n_2205),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_L g2358 ( 
.A(n_2264),
.B(n_2056),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2256),
.Y(n_2359)
);

OR2x2_ASAP7_75t_L g2360 ( 
.A(n_2283),
.B(n_2130),
.Y(n_2360)
);

AND2x4_ASAP7_75t_L g2361 ( 
.A(n_2265),
.B(n_2154),
.Y(n_2361)
);

HB1xp67_ASAP7_75t_L g2362 ( 
.A(n_2231),
.Y(n_2362)
);

AND2x2_ASAP7_75t_L g2363 ( 
.A(n_2285),
.B(n_2055),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_2271),
.B(n_2130),
.Y(n_2364)
);

AND2x2_ASAP7_75t_L g2365 ( 
.A(n_2202),
.B(n_2055),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2208),
.Y(n_2366)
);

INVx1_ASAP7_75t_L g2367 ( 
.A(n_2220),
.Y(n_2367)
);

AND2x4_ASAP7_75t_L g2368 ( 
.A(n_2272),
.B(n_2138),
.Y(n_2368)
);

INVx1_ASAP7_75t_SL g2369 ( 
.A(n_2218),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_2291),
.Y(n_2370)
);

AND2x2_ASAP7_75t_L g2371 ( 
.A(n_2284),
.B(n_2055),
.Y(n_2371)
);

INVx2_ASAP7_75t_L g2372 ( 
.A(n_2188),
.Y(n_2372)
);

AOI33xp33_ASAP7_75t_L g2373 ( 
.A1(n_2199),
.A2(n_2080),
.A3(n_2074),
.B1(n_2036),
.B2(n_2037),
.B3(n_2032),
.Y(n_2373)
);

AND2x4_ASAP7_75t_L g2374 ( 
.A(n_2177),
.B(n_2135),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2280),
.Y(n_2375)
);

AO21x2_ASAP7_75t_L g2376 ( 
.A1(n_2233),
.A2(n_2071),
.B(n_2035),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_2247),
.B(n_2130),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2228),
.Y(n_2378)
);

INVx2_ASAP7_75t_L g2379 ( 
.A(n_2237),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_2238),
.B(n_2130),
.Y(n_2380)
);

AND2x2_ASAP7_75t_L g2381 ( 
.A(n_2177),
.B(n_2139),
.Y(n_2381)
);

HB1xp67_ASAP7_75t_L g2382 ( 
.A(n_2267),
.Y(n_2382)
);

HB1xp67_ASAP7_75t_L g2383 ( 
.A(n_2268),
.Y(n_2383)
);

INVx2_ASAP7_75t_L g2384 ( 
.A(n_2274),
.Y(n_2384)
);

OR2x2_ASAP7_75t_L g2385 ( 
.A(n_2289),
.B(n_2054),
.Y(n_2385)
);

BUFx2_ASAP7_75t_L g2386 ( 
.A(n_2205),
.Y(n_2386)
);

INVxp67_ASAP7_75t_L g2387 ( 
.A(n_2191),
.Y(n_2387)
);

INVx5_ASAP7_75t_SL g2388 ( 
.A(n_2252),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2214),
.Y(n_2389)
);

AND2x2_ASAP7_75t_SL g2390 ( 
.A(n_2239),
.B(n_2136),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2214),
.Y(n_2391)
);

NOR2xp33_ASAP7_75t_L g2392 ( 
.A(n_2276),
.B(n_2155),
.Y(n_2392)
);

INVx2_ASAP7_75t_L g2393 ( 
.A(n_2290),
.Y(n_2393)
);

INVx2_ASAP7_75t_L g2394 ( 
.A(n_2240),
.Y(n_2394)
);

INVx2_ASAP7_75t_L g2395 ( 
.A(n_2240),
.Y(n_2395)
);

NOR2xp33_ASAP7_75t_R g2396 ( 
.A(n_2251),
.B(n_2080),
.Y(n_2396)
);

HB1xp67_ASAP7_75t_L g2397 ( 
.A(n_2214),
.Y(n_2397)
);

AND2x4_ASAP7_75t_L g2398 ( 
.A(n_2192),
.B(n_2136),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_2239),
.B(n_2227),
.Y(n_2399)
);

OAI221xp5_ASAP7_75t_L g2400 ( 
.A1(n_2249),
.A2(n_608),
.B1(n_612),
.B2(n_616),
.C(n_618),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2227),
.Y(n_2401)
);

OR2x2_ASAP7_75t_L g2402 ( 
.A(n_2266),
.B(n_2045),
.Y(n_2402)
);

AOI22xp33_ASAP7_75t_L g2403 ( 
.A1(n_2187),
.A2(n_2125),
.B1(n_2142),
.B2(n_2113),
.Y(n_2403)
);

INVxp67_ASAP7_75t_SL g2404 ( 
.A(n_2204),
.Y(n_2404)
);

NAND2xp5_ASAP7_75t_L g2405 ( 
.A(n_2357),
.B(n_2174),
.Y(n_2405)
);

AND2x2_ASAP7_75t_L g2406 ( 
.A(n_2314),
.B(n_2266),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2292),
.Y(n_2407)
);

AND2x2_ASAP7_75t_L g2408 ( 
.A(n_2297),
.B(n_2281),
.Y(n_2408)
);

AND2x2_ASAP7_75t_L g2409 ( 
.A(n_2294),
.B(n_2281),
.Y(n_2409)
);

AND2x2_ASAP7_75t_L g2410 ( 
.A(n_2331),
.B(n_2301),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_L g2411 ( 
.A(n_2386),
.B(n_2249),
.Y(n_2411)
);

OR2x2_ASAP7_75t_L g2412 ( 
.A(n_2316),
.B(n_2204),
.Y(n_2412)
);

AOI22xp5_ASAP7_75t_L g2413 ( 
.A1(n_2388),
.A2(n_2260),
.B1(n_2270),
.B2(n_2248),
.Y(n_2413)
);

NOR2xp33_ASAP7_75t_R g2414 ( 
.A(n_2308),
.B(n_59),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2292),
.Y(n_2415)
);

AND2x2_ASAP7_75t_L g2416 ( 
.A(n_2339),
.B(n_2034),
.Y(n_2416)
);

AND2x2_ASAP7_75t_L g2417 ( 
.A(n_2299),
.B(n_2050),
.Y(n_2417)
);

OR2x2_ASAP7_75t_L g2418 ( 
.A(n_2385),
.B(n_2227),
.Y(n_2418)
);

HB1xp67_ASAP7_75t_L g2419 ( 
.A(n_2295),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_L g2420 ( 
.A(n_2351),
.B(n_2219),
.Y(n_2420)
);

AND2x2_ASAP7_75t_L g2421 ( 
.A(n_2295),
.B(n_2131),
.Y(n_2421)
);

AND2x2_ASAP7_75t_L g2422 ( 
.A(n_2398),
.B(n_2201),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2307),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_L g2424 ( 
.A(n_2306),
.B(n_2262),
.Y(n_2424)
);

OR2x2_ASAP7_75t_L g2425 ( 
.A(n_2296),
.B(n_2347),
.Y(n_2425)
);

AND2x4_ASAP7_75t_L g2426 ( 
.A(n_2356),
.B(n_2232),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_L g2427 ( 
.A(n_2306),
.B(n_2393),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2307),
.Y(n_2428)
);

AND2x2_ASAP7_75t_L g2429 ( 
.A(n_2398),
.B(n_2232),
.Y(n_2429)
);

AND2x2_ASAP7_75t_L g2430 ( 
.A(n_2303),
.B(n_2232),
.Y(n_2430)
);

AND2x2_ASAP7_75t_L g2431 ( 
.A(n_2325),
.B(n_2217),
.Y(n_2431)
);

AND2x2_ASAP7_75t_L g2432 ( 
.A(n_2331),
.B(n_2195),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2312),
.Y(n_2433)
);

NAND2x1_ASAP7_75t_L g2434 ( 
.A(n_2356),
.B(n_2260),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2312),
.Y(n_2435)
);

INVx2_ASAP7_75t_L g2436 ( 
.A(n_2374),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2310),
.Y(n_2437)
);

AND2x4_ASAP7_75t_L g2438 ( 
.A(n_2325),
.B(n_2270),
.Y(n_2438)
);

INVx2_ASAP7_75t_SL g2439 ( 
.A(n_2302),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2321),
.Y(n_2440)
);

INVx1_ASAP7_75t_L g2441 ( 
.A(n_2322),
.Y(n_2441)
);

NAND2xp5_ASAP7_75t_L g2442 ( 
.A(n_2293),
.B(n_2253),
.Y(n_2442)
);

AND2x2_ASAP7_75t_L g2443 ( 
.A(n_2320),
.B(n_2196),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_2293),
.B(n_2248),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2323),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2338),
.Y(n_2446)
);

AND2x2_ASAP7_75t_L g2447 ( 
.A(n_2365),
.B(n_2158),
.Y(n_2447)
);

AND2x2_ASAP7_75t_L g2448 ( 
.A(n_2329),
.B(n_2158),
.Y(n_2448)
);

OR2x2_ASAP7_75t_L g2449 ( 
.A(n_2375),
.B(n_2158),
.Y(n_2449)
);

OR2x2_ASAP7_75t_L g2450 ( 
.A(n_2402),
.B(n_2158),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2346),
.Y(n_2451)
);

AND2x2_ASAP7_75t_L g2452 ( 
.A(n_2313),
.B(n_2311),
.Y(n_2452)
);

AND2x2_ASAP7_75t_L g2453 ( 
.A(n_2311),
.B(n_2234),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_2350),
.Y(n_2454)
);

HB1xp67_ASAP7_75t_L g2455 ( 
.A(n_2298),
.Y(n_2455)
);

AND2x2_ASAP7_75t_L g2456 ( 
.A(n_2328),
.B(n_2241),
.Y(n_2456)
);

AND2x2_ASAP7_75t_L g2457 ( 
.A(n_2332),
.B(n_2282),
.Y(n_2457)
);

BUFx2_ASAP7_75t_L g2458 ( 
.A(n_2396),
.Y(n_2458)
);

INVx1_ASAP7_75t_L g2459 ( 
.A(n_2353),
.Y(n_2459)
);

OR2x2_ASAP7_75t_L g2460 ( 
.A(n_2298),
.B(n_2252),
.Y(n_2460)
);

AND2x2_ASAP7_75t_L g2461 ( 
.A(n_2332),
.B(n_2282),
.Y(n_2461)
);

OR2x2_ASAP7_75t_L g2462 ( 
.A(n_2377),
.B(n_2263),
.Y(n_2462)
);

INVx3_ASAP7_75t_L g2463 ( 
.A(n_2388),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2324),
.Y(n_2464)
);

NAND2x1p5_ASAP7_75t_L g2465 ( 
.A(n_2368),
.B(n_2209),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_2340),
.B(n_2287),
.Y(n_2466)
);

AND2x2_ASAP7_75t_L g2467 ( 
.A(n_2304),
.B(n_2309),
.Y(n_2467)
);

AND2x2_ASAP7_75t_L g2468 ( 
.A(n_2317),
.B(n_2279),
.Y(n_2468)
);

AND2x2_ASAP7_75t_L g2469 ( 
.A(n_2318),
.B(n_61),
.Y(n_2469)
);

AND2x2_ASAP7_75t_L g2470 ( 
.A(n_2341),
.B(n_62),
.Y(n_2470)
);

INVxp67_ASAP7_75t_SL g2471 ( 
.A(n_2362),
.Y(n_2471)
);

INVx2_ASAP7_75t_L g2472 ( 
.A(n_2374),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2324),
.Y(n_2473)
);

NAND4xp25_ASAP7_75t_L g2474 ( 
.A(n_2387),
.B(n_2277),
.C(n_2246),
.D(n_2229),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2343),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2343),
.Y(n_2476)
);

NAND4xp25_ASAP7_75t_L g2477 ( 
.A(n_2387),
.B(n_62),
.C(n_64),
.D(n_65),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_L g2478 ( 
.A(n_2369),
.B(n_65),
.Y(n_2478)
);

INVx2_ASAP7_75t_SL g2479 ( 
.A(n_2341),
.Y(n_2479)
);

AND2x2_ASAP7_75t_L g2480 ( 
.A(n_2342),
.B(n_71),
.Y(n_2480)
);

INVx2_ASAP7_75t_L g2481 ( 
.A(n_2319),
.Y(n_2481)
);

AND2x2_ASAP7_75t_L g2482 ( 
.A(n_2361),
.B(n_71),
.Y(n_2482)
);

BUFx2_ASAP7_75t_L g2483 ( 
.A(n_2368),
.Y(n_2483)
);

INVx2_ASAP7_75t_L g2484 ( 
.A(n_2361),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2362),
.Y(n_2485)
);

AND2x2_ASAP7_75t_L g2486 ( 
.A(n_2363),
.B(n_72),
.Y(n_2486)
);

NOR4xp25_ASAP7_75t_SL g2487 ( 
.A(n_2300),
.B(n_620),
.C(n_74),
.D(n_75),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_L g2488 ( 
.A(n_2394),
.B(n_73),
.Y(n_2488)
);

OR2x2_ASAP7_75t_L g2489 ( 
.A(n_2377),
.B(n_75),
.Y(n_2489)
);

INVx1_ASAP7_75t_SL g2490 ( 
.A(n_2335),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2370),
.Y(n_2491)
);

NAND2xp33_ASAP7_75t_SL g2492 ( 
.A(n_2388),
.B(n_77),
.Y(n_2492)
);

INVx2_ASAP7_75t_SL g2493 ( 
.A(n_2410),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_L g2494 ( 
.A(n_2419),
.B(n_2455),
.Y(n_2494)
);

AND2x2_ASAP7_75t_L g2495 ( 
.A(n_2422),
.B(n_2327),
.Y(n_2495)
);

NOR2xp33_ASAP7_75t_L g2496 ( 
.A(n_2463),
.B(n_2337),
.Y(n_2496)
);

AND2x2_ASAP7_75t_L g2497 ( 
.A(n_2422),
.B(n_2371),
.Y(n_2497)
);

OAI32xp33_ASAP7_75t_L g2498 ( 
.A1(n_2444),
.A2(n_2364),
.A3(n_2399),
.B1(n_2397),
.B2(n_2395),
.Y(n_2498)
);

OR2x2_ASAP7_75t_L g2499 ( 
.A(n_2460),
.B(n_2404),
.Y(n_2499)
);

INVx2_ASAP7_75t_L g2500 ( 
.A(n_2439),
.Y(n_2500)
);

OR2x2_ASAP7_75t_L g2501 ( 
.A(n_2411),
.B(n_2404),
.Y(n_2501)
);

INVx2_ASAP7_75t_SL g2502 ( 
.A(n_2479),
.Y(n_2502)
);

AND2x2_ASAP7_75t_L g2503 ( 
.A(n_2439),
.B(n_2352),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2419),
.Y(n_2504)
);

INVxp67_ASAP7_75t_L g2505 ( 
.A(n_2455),
.Y(n_2505)
);

OR2x2_ASAP7_75t_L g2506 ( 
.A(n_2425),
.B(n_2399),
.Y(n_2506)
);

AND2x4_ASAP7_75t_L g2507 ( 
.A(n_2483),
.B(n_2389),
.Y(n_2507)
);

OAI21xp33_ASAP7_75t_L g2508 ( 
.A1(n_2405),
.A2(n_2364),
.B(n_2400),
.Y(n_2508)
);

AND2x2_ASAP7_75t_L g2509 ( 
.A(n_2458),
.B(n_2390),
.Y(n_2509)
);

NOR2x1p5_ASAP7_75t_L g2510 ( 
.A(n_2463),
.B(n_2349),
.Y(n_2510)
);

INVx1_ASAP7_75t_L g2511 ( 
.A(n_2471),
.Y(n_2511)
);

OR2x2_ASAP7_75t_L g2512 ( 
.A(n_2489),
.B(n_2490),
.Y(n_2512)
);

CKINVDCx16_ASAP7_75t_R g2513 ( 
.A(n_2414),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2471),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2423),
.Y(n_2515)
);

INVx2_ASAP7_75t_L g2516 ( 
.A(n_2479),
.Y(n_2516)
);

INVx1_ASAP7_75t_L g2517 ( 
.A(n_2428),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_L g2518 ( 
.A(n_2407),
.B(n_2397),
.Y(n_2518)
);

INVx2_ASAP7_75t_SL g2519 ( 
.A(n_2414),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_2433),
.Y(n_2520)
);

AND2x2_ASAP7_75t_L g2521 ( 
.A(n_2452),
.B(n_2403),
.Y(n_2521)
);

INVxp67_ASAP7_75t_L g2522 ( 
.A(n_2492),
.Y(n_2522)
);

NAND2xp5_ASAP7_75t_L g2523 ( 
.A(n_2415),
.B(n_2391),
.Y(n_2523)
);

INVx1_ASAP7_75t_L g2524 ( 
.A(n_2435),
.Y(n_2524)
);

OAI21xp33_ASAP7_75t_L g2525 ( 
.A1(n_2424),
.A2(n_2400),
.B(n_2373),
.Y(n_2525)
);

AND2x2_ASAP7_75t_L g2526 ( 
.A(n_2457),
.B(n_2379),
.Y(n_2526)
);

INVx1_ASAP7_75t_L g2527 ( 
.A(n_2464),
.Y(n_2527)
);

INVx2_ASAP7_75t_L g2528 ( 
.A(n_2436),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2473),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2475),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2476),
.Y(n_2531)
);

AND2x2_ASAP7_75t_L g2532 ( 
.A(n_2461),
.B(n_2384),
.Y(n_2532)
);

OAI32xp33_ASAP7_75t_L g2533 ( 
.A1(n_2465),
.A2(n_2442),
.A3(n_2427),
.B1(n_2463),
.B2(n_2492),
.Y(n_2533)
);

OR2x2_ASAP7_75t_L g2534 ( 
.A(n_2412),
.B(n_2358),
.Y(n_2534)
);

OR2x2_ASAP7_75t_L g2535 ( 
.A(n_2420),
.B(n_2358),
.Y(n_2535)
);

OR2x2_ASAP7_75t_L g2536 ( 
.A(n_2418),
.B(n_2378),
.Y(n_2536)
);

AND2x2_ASAP7_75t_L g2537 ( 
.A(n_2453),
.B(n_2326),
.Y(n_2537)
);

INVx2_ASAP7_75t_L g2538 ( 
.A(n_2436),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_L g2539 ( 
.A(n_2437),
.B(n_2401),
.Y(n_2539)
);

INVx2_ASAP7_75t_L g2540 ( 
.A(n_2472),
.Y(n_2540)
);

NAND2x1_ASAP7_75t_L g2541 ( 
.A(n_2426),
.B(n_2381),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2485),
.Y(n_2542)
);

AND2x2_ASAP7_75t_L g2543 ( 
.A(n_2443),
.B(n_2345),
.Y(n_2543)
);

INVx2_ASAP7_75t_L g2544 ( 
.A(n_2472),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2491),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2440),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2441),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2445),
.Y(n_2548)
);

INVx2_ASAP7_75t_SL g2549 ( 
.A(n_2484),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2446),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2451),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2454),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2459),
.Y(n_2553)
);

INVx1_ASAP7_75t_SL g2554 ( 
.A(n_2470),
.Y(n_2554)
);

INVxp33_ASAP7_75t_L g2555 ( 
.A(n_2465),
.Y(n_2555)
);

INVx2_ASAP7_75t_L g2556 ( 
.A(n_2484),
.Y(n_2556)
);

INVx1_ASAP7_75t_L g2557 ( 
.A(n_2470),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2482),
.Y(n_2558)
);

INVx2_ASAP7_75t_L g2559 ( 
.A(n_2482),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2469),
.Y(n_2560)
);

NAND4xp75_ASAP7_75t_L g2561 ( 
.A(n_2413),
.B(n_2315),
.C(n_2392),
.D(n_2305),
.Y(n_2561)
);

INVx1_ASAP7_75t_SL g2562 ( 
.A(n_2434),
.Y(n_2562)
);

NOR2xp33_ASAP7_75t_L g2563 ( 
.A(n_2466),
.B(n_2354),
.Y(n_2563)
);

INVx2_ASAP7_75t_L g2564 ( 
.A(n_2417),
.Y(n_2564)
);

NAND2xp5_ASAP7_75t_L g2565 ( 
.A(n_2488),
.B(n_2355),
.Y(n_2565)
);

INVx1_ASAP7_75t_SL g2566 ( 
.A(n_2480),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2469),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2426),
.Y(n_2568)
);

AND2x4_ASAP7_75t_L g2569 ( 
.A(n_2468),
.B(n_2359),
.Y(n_2569)
);

INVx2_ASAP7_75t_L g2570 ( 
.A(n_2417),
.Y(n_2570)
);

OR2x2_ASAP7_75t_L g2571 ( 
.A(n_2462),
.B(n_2330),
.Y(n_2571)
);

NAND2xp5_ASAP7_75t_L g2572 ( 
.A(n_2426),
.B(n_2366),
.Y(n_2572)
);

INVx2_ASAP7_75t_L g2573 ( 
.A(n_2416),
.Y(n_2573)
);

INVx2_ASAP7_75t_L g2574 ( 
.A(n_2429),
.Y(n_2574)
);

AND2x2_ASAP7_75t_L g2575 ( 
.A(n_2497),
.B(n_2495),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2494),
.Y(n_2576)
);

INVx2_ASAP7_75t_L g2577 ( 
.A(n_2519),
.Y(n_2577)
);

OR2x2_ASAP7_75t_L g2578 ( 
.A(n_2566),
.B(n_2315),
.Y(n_2578)
);

AND2x2_ASAP7_75t_L g2579 ( 
.A(n_2509),
.B(n_2406),
.Y(n_2579)
);

HB1xp67_ASAP7_75t_L g2580 ( 
.A(n_2505),
.Y(n_2580)
);

INVx1_ASAP7_75t_SL g2581 ( 
.A(n_2513),
.Y(n_2581)
);

INVx2_ASAP7_75t_L g2582 ( 
.A(n_2541),
.Y(n_2582)
);

AND2x2_ASAP7_75t_L g2583 ( 
.A(n_2500),
.B(n_2408),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2494),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_L g2585 ( 
.A(n_2522),
.B(n_2468),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2505),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2504),
.Y(n_2587)
);

BUFx2_ASAP7_75t_L g2588 ( 
.A(n_2522),
.Y(n_2588)
);

INVx2_ASAP7_75t_SL g2589 ( 
.A(n_2507),
.Y(n_2589)
);

INVx2_ASAP7_75t_SL g2590 ( 
.A(n_2507),
.Y(n_2590)
);

AND2x2_ASAP7_75t_L g2591 ( 
.A(n_2503),
.B(n_2493),
.Y(n_2591)
);

INVx3_ASAP7_75t_L g2592 ( 
.A(n_2511),
.Y(n_2592)
);

AND2x2_ASAP7_75t_L g2593 ( 
.A(n_2566),
.B(n_2431),
.Y(n_2593)
);

AND2x2_ASAP7_75t_L g2594 ( 
.A(n_2496),
.B(n_2431),
.Y(n_2594)
);

AND2x4_ASAP7_75t_L g2595 ( 
.A(n_2502),
.B(n_2429),
.Y(n_2595)
);

HB1xp67_ASAP7_75t_L g2596 ( 
.A(n_2514),
.Y(n_2596)
);

AND2x2_ASAP7_75t_L g2597 ( 
.A(n_2496),
.B(n_2467),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2574),
.Y(n_2598)
);

AO21x1_ASAP7_75t_L g2599 ( 
.A1(n_2555),
.A2(n_2478),
.B(n_2438),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2574),
.Y(n_2600)
);

INVx2_ASAP7_75t_L g2601 ( 
.A(n_2549),
.Y(n_2601)
);

INVx2_ASAP7_75t_L g2602 ( 
.A(n_2516),
.Y(n_2602)
);

INVx2_ASAP7_75t_L g2603 ( 
.A(n_2573),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2518),
.Y(n_2604)
);

INVx1_ASAP7_75t_SL g2605 ( 
.A(n_2562),
.Y(n_2605)
);

INVx2_ASAP7_75t_L g2606 ( 
.A(n_2568),
.Y(n_2606)
);

INVx1_ASAP7_75t_SL g2607 ( 
.A(n_2562),
.Y(n_2607)
);

OAI21x1_ASAP7_75t_L g2608 ( 
.A1(n_2572),
.A2(n_2481),
.B(n_2430),
.Y(n_2608)
);

CKINVDCx16_ASAP7_75t_R g2609 ( 
.A(n_2499),
.Y(n_2609)
);

HB1xp67_ASAP7_75t_L g2610 ( 
.A(n_2554),
.Y(n_2610)
);

AOI22xp33_ASAP7_75t_L g2611 ( 
.A1(n_2525),
.A2(n_2474),
.B1(n_2438),
.B2(n_2409),
.Y(n_2611)
);

AND2x2_ASAP7_75t_L g2612 ( 
.A(n_2521),
.B(n_2467),
.Y(n_2612)
);

NOR2xp33_ASAP7_75t_L g2613 ( 
.A(n_2533),
.B(n_2456),
.Y(n_2613)
);

NAND2xp5_ASAP7_75t_L g2614 ( 
.A(n_2554),
.B(n_2486),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2518),
.Y(n_2615)
);

AND2x2_ASAP7_75t_L g2616 ( 
.A(n_2555),
.B(n_2543),
.Y(n_2616)
);

NOR2xp33_ASAP7_75t_L g2617 ( 
.A(n_2508),
.B(n_2560),
.Y(n_2617)
);

INVx2_ASAP7_75t_L g2618 ( 
.A(n_2512),
.Y(n_2618)
);

BUFx3_ASAP7_75t_L g2619 ( 
.A(n_2501),
.Y(n_2619)
);

OAI22xp5_ASAP7_75t_L g2620 ( 
.A1(n_2561),
.A2(n_2487),
.B1(n_2438),
.B2(n_2416),
.Y(n_2620)
);

AND2x2_ASAP7_75t_L g2621 ( 
.A(n_2526),
.B(n_2421),
.Y(n_2621)
);

INVx2_ASAP7_75t_L g2622 ( 
.A(n_2564),
.Y(n_2622)
);

AND2x2_ASAP7_75t_L g2623 ( 
.A(n_2532),
.B(n_2421),
.Y(n_2623)
);

BUFx2_ASAP7_75t_L g2624 ( 
.A(n_2569),
.Y(n_2624)
);

INVx2_ASAP7_75t_L g2625 ( 
.A(n_2570),
.Y(n_2625)
);

INVx2_ASAP7_75t_L g2626 ( 
.A(n_2569),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2539),
.Y(n_2627)
);

AND3x1_ASAP7_75t_L g2628 ( 
.A(n_2508),
.B(n_2480),
.C(n_2430),
.Y(n_2628)
);

INVx2_ASAP7_75t_L g2629 ( 
.A(n_2528),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_2539),
.Y(n_2630)
);

NOR2xp33_ASAP7_75t_L g2631 ( 
.A(n_2567),
.B(n_2477),
.Y(n_2631)
);

OR2x2_ASAP7_75t_L g2632 ( 
.A(n_2557),
.B(n_2382),
.Y(n_2632)
);

CKINVDCx16_ASAP7_75t_R g2633 ( 
.A(n_2537),
.Y(n_2633)
);

AND2x4_ASAP7_75t_L g2634 ( 
.A(n_2538),
.B(n_2481),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_L g2635 ( 
.A(n_2558),
.B(n_2447),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2523),
.Y(n_2636)
);

AND2x4_ASAP7_75t_L g2637 ( 
.A(n_2624),
.B(n_2559),
.Y(n_2637)
);

AOI31xp33_ASAP7_75t_L g2638 ( 
.A1(n_2599),
.A2(n_2525),
.A3(n_2563),
.B(n_2515),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2610),
.Y(n_2639)
);

INVx2_ASAP7_75t_L g2640 ( 
.A(n_2624),
.Y(n_2640)
);

INVx2_ASAP7_75t_L g2641 ( 
.A(n_2589),
.Y(n_2641)
);

NAND2xp5_ASAP7_75t_L g2642 ( 
.A(n_2581),
.B(n_2510),
.Y(n_2642)
);

AND2x2_ASAP7_75t_L g2643 ( 
.A(n_2581),
.B(n_2556),
.Y(n_2643)
);

AND2x4_ASAP7_75t_L g2644 ( 
.A(n_2589),
.B(n_2540),
.Y(n_2644)
);

AND2x4_ASAP7_75t_L g2645 ( 
.A(n_2590),
.B(n_2544),
.Y(n_2645)
);

AND2x4_ASAP7_75t_L g2646 ( 
.A(n_2590),
.B(n_2542),
.Y(n_2646)
);

INVx2_ASAP7_75t_L g2647 ( 
.A(n_2595),
.Y(n_2647)
);

AND2x2_ASAP7_75t_L g2648 ( 
.A(n_2575),
.B(n_2563),
.Y(n_2648)
);

INVxp67_ASAP7_75t_L g2649 ( 
.A(n_2588),
.Y(n_2649)
);

NAND2xp5_ASAP7_75t_L g2650 ( 
.A(n_2633),
.B(n_2517),
.Y(n_2650)
);

HB1xp67_ASAP7_75t_L g2651 ( 
.A(n_2588),
.Y(n_2651)
);

INVx1_ASAP7_75t_SL g2652 ( 
.A(n_2607),
.Y(n_2652)
);

OR2x2_ASAP7_75t_L g2653 ( 
.A(n_2609),
.B(n_2585),
.Y(n_2653)
);

BUFx2_ASAP7_75t_L g2654 ( 
.A(n_2619),
.Y(n_2654)
);

INVx2_ASAP7_75t_L g2655 ( 
.A(n_2595),
.Y(n_2655)
);

NAND2x1p5_ASAP7_75t_L g2656 ( 
.A(n_2619),
.B(n_2520),
.Y(n_2656)
);

NOR2xp33_ASAP7_75t_L g2657 ( 
.A(n_2633),
.B(n_2498),
.Y(n_2657)
);

INVx1_ASAP7_75t_SL g2658 ( 
.A(n_2607),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_SL g2659 ( 
.A(n_2599),
.B(n_2571),
.Y(n_2659)
);

NOR2xp33_ASAP7_75t_L g2660 ( 
.A(n_2609),
.B(n_2524),
.Y(n_2660)
);

AND2x2_ASAP7_75t_L g2661 ( 
.A(n_2575),
.B(n_2535),
.Y(n_2661)
);

AND2x2_ASAP7_75t_L g2662 ( 
.A(n_2597),
.B(n_2527),
.Y(n_2662)
);

NAND2xp5_ASAP7_75t_L g2663 ( 
.A(n_2605),
.B(n_2529),
.Y(n_2663)
);

NAND2xp5_ASAP7_75t_L g2664 ( 
.A(n_2597),
.B(n_2577),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2592),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2592),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2592),
.Y(n_2667)
);

INVx1_ASAP7_75t_SL g2668 ( 
.A(n_2616),
.Y(n_2668)
);

AND2x2_ASAP7_75t_L g2669 ( 
.A(n_2594),
.B(n_2530),
.Y(n_2669)
);

AND2x2_ASAP7_75t_L g2670 ( 
.A(n_2594),
.B(n_2531),
.Y(n_2670)
);

AND2x2_ASAP7_75t_L g2671 ( 
.A(n_2616),
.B(n_2506),
.Y(n_2671)
);

NAND2xp5_ASAP7_75t_L g2672 ( 
.A(n_2577),
.B(n_2565),
.Y(n_2672)
);

AND2x2_ASAP7_75t_L g2673 ( 
.A(n_2612),
.B(n_2565),
.Y(n_2673)
);

INVx1_ASAP7_75t_SL g2674 ( 
.A(n_2612),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2592),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2580),
.Y(n_2676)
);

AND2x2_ASAP7_75t_L g2677 ( 
.A(n_2621),
.B(n_2623),
.Y(n_2677)
);

INVx1_ASAP7_75t_SL g2678 ( 
.A(n_2591),
.Y(n_2678)
);

NAND2xp5_ASAP7_75t_L g2679 ( 
.A(n_2591),
.B(n_2545),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2596),
.Y(n_2680)
);

HB1xp67_ASAP7_75t_L g2681 ( 
.A(n_2619),
.Y(n_2681)
);

OR2x2_ASAP7_75t_L g2682 ( 
.A(n_2614),
.B(n_2534),
.Y(n_2682)
);

NOR2xp67_ASAP7_75t_L g2683 ( 
.A(n_2626),
.B(n_2536),
.Y(n_2683)
);

AOI222xp33_ASAP7_75t_L g2684 ( 
.A1(n_2659),
.A2(n_2617),
.B1(n_2613),
.B2(n_2611),
.C1(n_2620),
.C2(n_2631),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2681),
.Y(n_2685)
);

OAI22xp5_ASAP7_75t_L g2686 ( 
.A1(n_2638),
.A2(n_2628),
.B1(n_2618),
.B2(n_2601),
.Y(n_2686)
);

OR2x2_ASAP7_75t_L g2687 ( 
.A(n_2654),
.B(n_2618),
.Y(n_2687)
);

OAI221xp5_ASAP7_75t_L g2688 ( 
.A1(n_2657),
.A2(n_2628),
.B1(n_2635),
.B2(n_2586),
.C(n_2625),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_L g2689 ( 
.A(n_2677),
.B(n_2626),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_L g2690 ( 
.A(n_2677),
.B(n_2601),
.Y(n_2690)
);

INVx2_ASAP7_75t_L g2691 ( 
.A(n_2656),
.Y(n_2691)
);

NAND4xp75_ASAP7_75t_L g2692 ( 
.A(n_2659),
.B(n_2586),
.C(n_2584),
.D(n_2576),
.Y(n_2692)
);

INVx2_ASAP7_75t_L g2693 ( 
.A(n_2656),
.Y(n_2693)
);

OAI211xp5_ASAP7_75t_SL g2694 ( 
.A1(n_2642),
.A2(n_2576),
.B(n_2584),
.C(n_2604),
.Y(n_2694)
);

NAND2xp5_ASAP7_75t_L g2695 ( 
.A(n_2643),
.B(n_2602),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2651),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2640),
.Y(n_2697)
);

INVx2_ASAP7_75t_SL g2698 ( 
.A(n_2637),
.Y(n_2698)
);

NOR2xp33_ASAP7_75t_L g2699 ( 
.A(n_2668),
.B(n_2602),
.Y(n_2699)
);

NAND2xp5_ASAP7_75t_L g2700 ( 
.A(n_2643),
.B(n_2621),
.Y(n_2700)
);

NOR3xp33_ASAP7_75t_L g2701 ( 
.A(n_2650),
.B(n_2587),
.C(n_2604),
.Y(n_2701)
);

NOR2xp67_ASAP7_75t_SL g2702 ( 
.A(n_2653),
.B(n_2676),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2640),
.Y(n_2703)
);

OR2x2_ASAP7_75t_L g2704 ( 
.A(n_2652),
.B(n_2622),
.Y(n_2704)
);

NAND2xp33_ASAP7_75t_SL g2705 ( 
.A(n_2648),
.B(n_2593),
.Y(n_2705)
);

INVx3_ASAP7_75t_L g2706 ( 
.A(n_2644),
.Y(n_2706)
);

NAND2xp5_ASAP7_75t_L g2707 ( 
.A(n_2678),
.B(n_2623),
.Y(n_2707)
);

AND2x2_ASAP7_75t_L g2708 ( 
.A(n_2674),
.B(n_2593),
.Y(n_2708)
);

AND2x2_ASAP7_75t_L g2709 ( 
.A(n_2648),
.B(n_2583),
.Y(n_2709)
);

AOI21xp5_ASAP7_75t_L g2710 ( 
.A1(n_2657),
.A2(n_2579),
.B(n_2582),
.Y(n_2710)
);

NAND2x1_ASAP7_75t_L g2711 ( 
.A(n_2644),
.B(n_2595),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2665),
.Y(n_2712)
);

AOI21xp33_ASAP7_75t_SL g2713 ( 
.A1(n_2660),
.A2(n_2625),
.B(n_2622),
.Y(n_2713)
);

INVxp67_ASAP7_75t_L g2714 ( 
.A(n_2660),
.Y(n_2714)
);

AOI22xp33_ASAP7_75t_L g2715 ( 
.A1(n_2661),
.A2(n_2579),
.B1(n_2583),
.B2(n_2603),
.Y(n_2715)
);

INVxp67_ASAP7_75t_L g2716 ( 
.A(n_2644),
.Y(n_2716)
);

NAND4xp25_ASAP7_75t_L g2717 ( 
.A(n_2664),
.B(n_2587),
.C(n_2615),
.D(n_2603),
.Y(n_2717)
);

NAND3xp33_ASAP7_75t_SL g2718 ( 
.A(n_2658),
.B(n_2582),
.C(n_2578),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2666),
.Y(n_2719)
);

OAI21xp5_ASAP7_75t_SL g2720 ( 
.A1(n_2649),
.A2(n_2615),
.B(n_2636),
.Y(n_2720)
);

AOI22xp33_ASAP7_75t_L g2721 ( 
.A1(n_2671),
.A2(n_2636),
.B1(n_2595),
.B2(n_2629),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_L g2722 ( 
.A(n_2692),
.B(n_2637),
.Y(n_2722)
);

INVx2_ASAP7_75t_L g2723 ( 
.A(n_2706),
.Y(n_2723)
);

OAI21xp33_ASAP7_75t_L g2724 ( 
.A1(n_2684),
.A2(n_2671),
.B(n_2639),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2706),
.Y(n_2725)
);

NAND2xp5_ASAP7_75t_L g2726 ( 
.A(n_2698),
.B(n_2645),
.Y(n_2726)
);

OAI21xp33_ASAP7_75t_L g2727 ( 
.A1(n_2684),
.A2(n_2663),
.B(n_2673),
.Y(n_2727)
);

NAND2x1_ASAP7_75t_L g2728 ( 
.A(n_2691),
.B(n_2645),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2716),
.Y(n_2729)
);

NAND2xp5_ASAP7_75t_SL g2730 ( 
.A(n_2714),
.B(n_2637),
.Y(n_2730)
);

INVx3_ASAP7_75t_L g2731 ( 
.A(n_2711),
.Y(n_2731)
);

AND2x2_ASAP7_75t_L g2732 ( 
.A(n_2709),
.B(n_2673),
.Y(n_2732)
);

AND2x2_ASAP7_75t_L g2733 ( 
.A(n_2708),
.B(n_2662),
.Y(n_2733)
);

INVx1_ASAP7_75t_SL g2734 ( 
.A(n_2705),
.Y(n_2734)
);

AOI22xp5_ASAP7_75t_L g2735 ( 
.A1(n_2686),
.A2(n_2641),
.B1(n_2670),
.B2(n_2669),
.Y(n_2735)
);

NOR2xp33_ASAP7_75t_L g2736 ( 
.A(n_2700),
.B(n_2672),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2687),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2695),
.Y(n_2738)
);

OAI22xp33_ASAP7_75t_L g2739 ( 
.A1(n_2688),
.A2(n_2718),
.B1(n_2707),
.B2(n_2704),
.Y(n_2739)
);

AND2x2_ASAP7_75t_L g2740 ( 
.A(n_2715),
.B(n_2641),
.Y(n_2740)
);

NOR3xp33_ASAP7_75t_L g2741 ( 
.A(n_2694),
.B(n_2680),
.C(n_2679),
.Y(n_2741)
);

NAND2xp5_ASAP7_75t_L g2742 ( 
.A(n_2710),
.B(n_2645),
.Y(n_2742)
);

AOI21xp33_ASAP7_75t_SL g2743 ( 
.A1(n_2699),
.A2(n_2682),
.B(n_2646),
.Y(n_2743)
);

AOI22xp33_ASAP7_75t_L g2744 ( 
.A1(n_2702),
.A2(n_2701),
.B1(n_2685),
.B2(n_2696),
.Y(n_2744)
);

INVx1_ASAP7_75t_SL g2745 ( 
.A(n_2693),
.Y(n_2745)
);

NAND2x1_ASAP7_75t_SL g2746 ( 
.A(n_2697),
.B(n_2646),
.Y(n_2746)
);

INVxp67_ASAP7_75t_L g2747 ( 
.A(n_2690),
.Y(n_2747)
);

AND2x2_ASAP7_75t_L g2748 ( 
.A(n_2689),
.B(n_2669),
.Y(n_2748)
);

INVx2_ASAP7_75t_L g2749 ( 
.A(n_2703),
.Y(n_2749)
);

INVxp67_ASAP7_75t_L g2750 ( 
.A(n_2713),
.Y(n_2750)
);

NAND2xp5_ASAP7_75t_L g2751 ( 
.A(n_2721),
.B(n_2646),
.Y(n_2751)
);

OR2x2_ASAP7_75t_L g2752 ( 
.A(n_2717),
.B(n_2632),
.Y(n_2752)
);

NAND2xp5_ASAP7_75t_L g2753 ( 
.A(n_2712),
.B(n_2670),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_L g2754 ( 
.A(n_2732),
.B(n_2667),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2746),
.Y(n_2755)
);

OR2x2_ASAP7_75t_L g2756 ( 
.A(n_2726),
.B(n_2717),
.Y(n_2756)
);

NAND2xp5_ASAP7_75t_L g2757 ( 
.A(n_2734),
.B(n_2683),
.Y(n_2757)
);

AND2x2_ASAP7_75t_L g2758 ( 
.A(n_2733),
.B(n_2647),
.Y(n_2758)
);

NAND2xp5_ASAP7_75t_L g2759 ( 
.A(n_2734),
.B(n_2647),
.Y(n_2759)
);

AOI21xp5_ASAP7_75t_L g2760 ( 
.A1(n_2739),
.A2(n_2720),
.B(n_2675),
.Y(n_2760)
);

NAND2x1_ASAP7_75t_L g2761 ( 
.A(n_2731),
.B(n_2655),
.Y(n_2761)
);

INVxp67_ASAP7_75t_L g2762 ( 
.A(n_2742),
.Y(n_2762)
);

NAND2xp33_ASAP7_75t_SL g2763 ( 
.A(n_2728),
.B(n_2655),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_2723),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2725),
.Y(n_2765)
);

INVxp67_ASAP7_75t_L g2766 ( 
.A(n_2730),
.Y(n_2766)
);

OAI22xp33_ASAP7_75t_L g2767 ( 
.A1(n_2722),
.A2(n_2578),
.B1(n_2720),
.B2(n_2632),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2731),
.Y(n_2768)
);

NAND3xp33_ASAP7_75t_L g2769 ( 
.A(n_2741),
.B(n_2719),
.C(n_2629),
.Y(n_2769)
);

NOR2xp33_ASAP7_75t_L g2770 ( 
.A(n_2724),
.B(n_2606),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_SL g2771 ( 
.A(n_2743),
.B(n_2634),
.Y(n_2771)
);

INVx1_ASAP7_75t_L g2772 ( 
.A(n_2753),
.Y(n_2772)
);

AND2x2_ASAP7_75t_L g2773 ( 
.A(n_2748),
.B(n_2606),
.Y(n_2773)
);

AND2x2_ASAP7_75t_L g2774 ( 
.A(n_2740),
.B(n_2627),
.Y(n_2774)
);

NAND2xp5_ASAP7_75t_L g2775 ( 
.A(n_2745),
.B(n_2627),
.Y(n_2775)
);

NAND2xp5_ASAP7_75t_SL g2776 ( 
.A(n_2735),
.B(n_2634),
.Y(n_2776)
);

XNOR2xp5_ASAP7_75t_L g2777 ( 
.A(n_2744),
.B(n_2630),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2753),
.Y(n_2778)
);

NOR2xp33_ASAP7_75t_L g2779 ( 
.A(n_2766),
.B(n_2727),
.Y(n_2779)
);

NOR2xp33_ASAP7_75t_L g2780 ( 
.A(n_2762),
.B(n_2750),
.Y(n_2780)
);

CKINVDCx20_ASAP7_75t_L g2781 ( 
.A(n_2763),
.Y(n_2781)
);

NOR2x1_ASAP7_75t_L g2782 ( 
.A(n_2761),
.B(n_2722),
.Y(n_2782)
);

NAND2xp5_ASAP7_75t_L g2783 ( 
.A(n_2758),
.B(n_2745),
.Y(n_2783)
);

NAND2xp5_ASAP7_75t_L g2784 ( 
.A(n_2768),
.B(n_2737),
.Y(n_2784)
);

NOR2xp33_ASAP7_75t_L g2785 ( 
.A(n_2757),
.B(n_2747),
.Y(n_2785)
);

AND2x2_ASAP7_75t_L g2786 ( 
.A(n_2773),
.B(n_2729),
.Y(n_2786)
);

NAND2xp5_ASAP7_75t_L g2787 ( 
.A(n_2755),
.B(n_2751),
.Y(n_2787)
);

AO21x1_ASAP7_75t_L g2788 ( 
.A1(n_2760),
.A2(n_2767),
.B(n_2771),
.Y(n_2788)
);

NAND3xp33_ASAP7_75t_L g2789 ( 
.A(n_2770),
.B(n_2752),
.C(n_2736),
.Y(n_2789)
);

NAND3xp33_ASAP7_75t_L g2790 ( 
.A(n_2776),
.B(n_2769),
.C(n_2759),
.Y(n_2790)
);

AOI21xp5_ASAP7_75t_L g2791 ( 
.A1(n_2777),
.A2(n_2738),
.B(n_2749),
.Y(n_2791)
);

NAND2xp5_ASAP7_75t_L g2792 ( 
.A(n_2774),
.B(n_2630),
.Y(n_2792)
);

NAND3xp33_ASAP7_75t_L g2793 ( 
.A(n_2754),
.B(n_2600),
.C(n_2598),
.Y(n_2793)
);

INVx1_ASAP7_75t_L g2794 ( 
.A(n_2754),
.Y(n_2794)
);

AOI211x1_ASAP7_75t_SL g2795 ( 
.A1(n_2775),
.A2(n_2523),
.B(n_2572),
.C(n_2600),
.Y(n_2795)
);

OAI22xp5_ASAP7_75t_L g2796 ( 
.A1(n_2756),
.A2(n_2598),
.B1(n_2546),
.B2(n_2548),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2775),
.Y(n_2797)
);

O2A1O1Ixp33_ASAP7_75t_L g2798 ( 
.A1(n_2788),
.A2(n_2778),
.B(n_2772),
.C(n_2764),
.Y(n_2798)
);

AOI211xp5_ASAP7_75t_L g2799 ( 
.A1(n_2790),
.A2(n_2765),
.B(n_2547),
.C(n_2553),
.Y(n_2799)
);

AOI321xp33_ASAP7_75t_L g2800 ( 
.A1(n_2779),
.A2(n_2634),
.A3(n_2552),
.B1(n_2551),
.B2(n_2550),
.C(n_2608),
.Y(n_2800)
);

OAI21xp33_ASAP7_75t_L g2801 ( 
.A1(n_2780),
.A2(n_2634),
.B(n_2608),
.Y(n_2801)
);

AOI22xp33_ASAP7_75t_L g2802 ( 
.A1(n_2789),
.A2(n_2432),
.B1(n_2376),
.B2(n_2450),
.Y(n_2802)
);

OAI211xp5_ASAP7_75t_SL g2803 ( 
.A1(n_2787),
.A2(n_2449),
.B(n_2380),
.C(n_2305),
.Y(n_2803)
);

OAI22xp5_ASAP7_75t_L g2804 ( 
.A1(n_2783),
.A2(n_2360),
.B1(n_2380),
.B2(n_2382),
.Y(n_2804)
);

NOR2xp33_ASAP7_75t_L g2805 ( 
.A(n_2786),
.B(n_2376),
.Y(n_2805)
);

OAI321xp33_ASAP7_75t_L g2806 ( 
.A1(n_2784),
.A2(n_2448),
.A3(n_2330),
.B1(n_2334),
.B2(n_2333),
.C(n_2367),
.Y(n_2806)
);

NAND2xp5_ASAP7_75t_L g2807 ( 
.A(n_2782),
.B(n_2383),
.Y(n_2807)
);

OAI221xp5_ASAP7_75t_L g2808 ( 
.A1(n_2791),
.A2(n_2383),
.B1(n_2334),
.B2(n_2333),
.C(n_2372),
.Y(n_2808)
);

OAI211xp5_ASAP7_75t_L g2809 ( 
.A1(n_2785),
.A2(n_2348),
.B(n_2344),
.C(n_2336),
.Y(n_2809)
);

AOI222xp33_ASAP7_75t_L g2810 ( 
.A1(n_2797),
.A2(n_2348),
.B1(n_2344),
.B2(n_2336),
.C1(n_81),
.C2(n_82),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_L g2811 ( 
.A(n_2801),
.B(n_2794),
.Y(n_2811)
);

NAND2xp5_ASAP7_75t_L g2812 ( 
.A(n_2807),
.B(n_2795),
.Y(n_2812)
);

INVx1_ASAP7_75t_L g2813 ( 
.A(n_2800),
.Y(n_2813)
);

INVx1_ASAP7_75t_L g2814 ( 
.A(n_2798),
.Y(n_2814)
);

NAND2xp5_ASAP7_75t_L g2815 ( 
.A(n_2810),
.B(n_2792),
.Y(n_2815)
);

NOR3xp33_ASAP7_75t_L g2816 ( 
.A(n_2799),
.B(n_2793),
.C(n_2796),
.Y(n_2816)
);

OAI22x1_ASAP7_75t_L g2817 ( 
.A1(n_2805),
.A2(n_2781),
.B1(n_78),
.B2(n_79),
.Y(n_2817)
);

AOI322xp5_ASAP7_75t_L g2818 ( 
.A1(n_2802),
.A2(n_2806),
.A3(n_2803),
.B1(n_2809),
.B2(n_2808),
.C1(n_2804),
.C2(n_85),
.Y(n_2818)
);

OAI211xp5_ASAP7_75t_L g2819 ( 
.A1(n_2798),
.A2(n_77),
.B(n_78),
.C(n_81),
.Y(n_2819)
);

AOI22xp33_ASAP7_75t_SL g2820 ( 
.A1(n_2807),
.A2(n_82),
.B1(n_83),
.B2(n_87),
.Y(n_2820)
);

NAND4xp75_ASAP7_75t_L g2821 ( 
.A(n_2807),
.B(n_83),
.C(n_87),
.D(n_90),
.Y(n_2821)
);

INVx2_ASAP7_75t_SL g2822 ( 
.A(n_2807),
.Y(n_2822)
);

XNOR2xp5_ASAP7_75t_L g2823 ( 
.A(n_2799),
.B(n_91),
.Y(n_2823)
);

AOI21xp33_ASAP7_75t_L g2824 ( 
.A1(n_2813),
.A2(n_2814),
.B(n_2811),
.Y(n_2824)
);

OAI22xp33_ASAP7_75t_L g2825 ( 
.A1(n_2812),
.A2(n_92),
.B1(n_94),
.B2(n_95),
.Y(n_2825)
);

AOI221x1_ASAP7_75t_L g2826 ( 
.A1(n_2817),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.C(n_98),
.Y(n_2826)
);

OAI221xp5_ASAP7_75t_L g2827 ( 
.A1(n_2816),
.A2(n_96),
.B1(n_98),
.B2(n_99),
.C(n_100),
.Y(n_2827)
);

NAND2xp5_ASAP7_75t_L g2828 ( 
.A(n_2820),
.B(n_99),
.Y(n_2828)
);

OAI221xp5_ASAP7_75t_L g2829 ( 
.A1(n_2819),
.A2(n_101),
.B1(n_102),
.B2(n_103),
.C(n_104),
.Y(n_2829)
);

AOI21xp5_ASAP7_75t_L g2830 ( 
.A1(n_2815),
.A2(n_101),
.B(n_103),
.Y(n_2830)
);

AND2x2_ASAP7_75t_L g2831 ( 
.A(n_2822),
.B(n_104),
.Y(n_2831)
);

OAI211xp5_ASAP7_75t_SL g2832 ( 
.A1(n_2818),
.A2(n_105),
.B(n_106),
.C(n_108),
.Y(n_2832)
);

AOI22xp5_ASAP7_75t_L g2833 ( 
.A1(n_2821),
.A2(n_2823),
.B1(n_106),
.B2(n_110),
.Y(n_2833)
);

OAI21xp33_ASAP7_75t_L g2834 ( 
.A1(n_2813),
.A2(n_105),
.B(n_110),
.Y(n_2834)
);

AND2x4_ASAP7_75t_L g2835 ( 
.A(n_2822),
.B(n_111),
.Y(n_2835)
);

NOR3xp33_ASAP7_75t_SL g2836 ( 
.A(n_2819),
.B(n_112),
.C(n_113),
.Y(n_2836)
);

NAND3xp33_ASAP7_75t_L g2837 ( 
.A(n_2814),
.B(n_114),
.C(n_115),
.Y(n_2837)
);

AOI211xp5_ASAP7_75t_SL g2838 ( 
.A1(n_2819),
.A2(n_114),
.B(n_116),
.C(n_117),
.Y(n_2838)
);

OAI21xp33_ASAP7_75t_L g2839 ( 
.A1(n_2813),
.A2(n_116),
.B(n_119),
.Y(n_2839)
);

OAI22xp33_ASAP7_75t_L g2840 ( 
.A1(n_2814),
.A2(n_119),
.B1(n_121),
.B2(n_122),
.Y(n_2840)
);

AOI31xp33_ASAP7_75t_L g2841 ( 
.A1(n_2838),
.A2(n_122),
.A3(n_124),
.B(n_125),
.Y(n_2841)
);

NAND4xp25_ASAP7_75t_L g2842 ( 
.A(n_2824),
.B(n_124),
.C(n_126),
.D(n_127),
.Y(n_2842)
);

BUFx6f_ASAP7_75t_L g2843 ( 
.A(n_2835),
.Y(n_2843)
);

CKINVDCx5p33_ASAP7_75t_R g2844 ( 
.A(n_2831),
.Y(n_2844)
);

NOR2xp67_ASAP7_75t_L g2845 ( 
.A(n_2837),
.B(n_129),
.Y(n_2845)
);

NAND2xp5_ASAP7_75t_L g2846 ( 
.A(n_2835),
.B(n_129),
.Y(n_2846)
);

HB1xp67_ASAP7_75t_L g2847 ( 
.A(n_2826),
.Y(n_2847)
);

AOI22xp5_ASAP7_75t_L g2848 ( 
.A1(n_2832),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_2848)
);

NAND2xp5_ASAP7_75t_L g2849 ( 
.A(n_2840),
.B(n_130),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2828),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2829),
.Y(n_2851)
);

NOR2x1p5_ASAP7_75t_L g2852 ( 
.A(n_2836),
.B(n_131),
.Y(n_2852)
);

NAND3x2_ASAP7_75t_L g2853 ( 
.A(n_2834),
.B(n_132),
.C(n_133),
.Y(n_2853)
);

AOI211x1_ASAP7_75t_L g2854 ( 
.A1(n_2839),
.A2(n_134),
.B(n_135),
.C(n_137),
.Y(n_2854)
);

NAND3x1_ASAP7_75t_L g2855 ( 
.A(n_2833),
.B(n_134),
.C(n_138),
.Y(n_2855)
);

HB1xp67_ASAP7_75t_L g2856 ( 
.A(n_2843),
.Y(n_2856)
);

BUFx2_ASAP7_75t_L g2857 ( 
.A(n_2843),
.Y(n_2857)
);

HB1xp67_ASAP7_75t_L g2858 ( 
.A(n_2847),
.Y(n_2858)
);

CKINVDCx5p33_ASAP7_75t_R g2859 ( 
.A(n_2844),
.Y(n_2859)
);

XNOR2x2_ASAP7_75t_SL g2860 ( 
.A(n_2848),
.B(n_2827),
.Y(n_2860)
);

INVx1_ASAP7_75t_SL g2861 ( 
.A(n_2846),
.Y(n_2861)
);

CKINVDCx5p33_ASAP7_75t_R g2862 ( 
.A(n_2850),
.Y(n_2862)
);

NAND2xp5_ASAP7_75t_L g2863 ( 
.A(n_2841),
.B(n_2830),
.Y(n_2863)
);

NAND2xp33_ASAP7_75t_L g2864 ( 
.A(n_2855),
.B(n_2825),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2852),
.Y(n_2865)
);

HB1xp67_ASAP7_75t_L g2866 ( 
.A(n_2845),
.Y(n_2866)
);

CKINVDCx16_ASAP7_75t_R g2867 ( 
.A(n_2851),
.Y(n_2867)
);

AO22x2_ASAP7_75t_L g2868 ( 
.A1(n_2865),
.A2(n_2854),
.B1(n_2849),
.B2(n_2842),
.Y(n_2868)
);

CKINVDCx16_ASAP7_75t_R g2869 ( 
.A(n_2867),
.Y(n_2869)
);

AOI22xp33_ASAP7_75t_L g2870 ( 
.A1(n_2858),
.A2(n_2853),
.B1(n_143),
.B2(n_145),
.Y(n_2870)
);

AOI22xp5_ASAP7_75t_L g2871 ( 
.A1(n_2859),
.A2(n_139),
.B1(n_143),
.B2(n_147),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2856),
.Y(n_2872)
);

INVx2_ASAP7_75t_L g2873 ( 
.A(n_2857),
.Y(n_2873)
);

CKINVDCx11_ASAP7_75t_R g2874 ( 
.A(n_2861),
.Y(n_2874)
);

INVxp67_ASAP7_75t_L g2875 ( 
.A(n_2863),
.Y(n_2875)
);

XNOR2xp5_ASAP7_75t_L g2876 ( 
.A(n_2860),
.B(n_2862),
.Y(n_2876)
);

HB1xp67_ASAP7_75t_L g2877 ( 
.A(n_2866),
.Y(n_2877)
);

AOI22xp5_ASAP7_75t_L g2878 ( 
.A1(n_2864),
.A2(n_139),
.B1(n_1249),
.B2(n_1229),
.Y(n_2878)
);

HB1xp67_ASAP7_75t_L g2879 ( 
.A(n_2869),
.Y(n_2879)
);

OR3x1_ASAP7_75t_L g2880 ( 
.A(n_2872),
.B(n_149),
.C(n_153),
.Y(n_2880)
);

BUFx2_ASAP7_75t_L g2881 ( 
.A(n_2877),
.Y(n_2881)
);

OAI22xp5_ASAP7_75t_L g2882 ( 
.A1(n_2870),
.A2(n_863),
.B1(n_865),
.B2(n_165),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2868),
.Y(n_2883)
);

OAI22xp5_ASAP7_75t_SL g2884 ( 
.A1(n_2873),
.A2(n_156),
.B1(n_161),
.B2(n_167),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2868),
.Y(n_2885)
);

AND2x2_ASAP7_75t_L g2886 ( 
.A(n_2875),
.B(n_2874),
.Y(n_2886)
);

INVx2_ASAP7_75t_L g2887 ( 
.A(n_2876),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_2871),
.Y(n_2888)
);

BUFx3_ASAP7_75t_L g2889 ( 
.A(n_2878),
.Y(n_2889)
);

NOR2x1_ASAP7_75t_L g2890 ( 
.A(n_2872),
.B(n_176),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2879),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2881),
.Y(n_2892)
);

CKINVDCx20_ASAP7_75t_R g2893 ( 
.A(n_2886),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2883),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2885),
.Y(n_2895)
);

AOI22x1_ASAP7_75t_L g2896 ( 
.A1(n_2891),
.A2(n_2887),
.B1(n_2888),
.B2(n_2890),
.Y(n_2896)
);

CKINVDCx20_ASAP7_75t_R g2897 ( 
.A(n_2893),
.Y(n_2897)
);

INVx2_ASAP7_75t_L g2898 ( 
.A(n_2892),
.Y(n_2898)
);

AO22x1_ASAP7_75t_L g2899 ( 
.A1(n_2894),
.A2(n_2882),
.B1(n_2889),
.B2(n_2880),
.Y(n_2899)
);

CKINVDCx20_ASAP7_75t_R g2900 ( 
.A(n_2895),
.Y(n_2900)
);

OAI22xp5_ASAP7_75t_L g2901 ( 
.A1(n_2893),
.A2(n_2884),
.B1(n_863),
.B2(n_865),
.Y(n_2901)
);

AOI22x1_ASAP7_75t_SL g2902 ( 
.A1(n_2893),
.A2(n_177),
.B1(n_182),
.B2(n_184),
.Y(n_2902)
);

AO22x2_ASAP7_75t_L g2903 ( 
.A1(n_2892),
.A2(n_185),
.B1(n_190),
.B2(n_191),
.Y(n_2903)
);

NAND3xp33_ASAP7_75t_L g2904 ( 
.A(n_2896),
.B(n_865),
.C(n_194),
.Y(n_2904)
);

OAI21x1_ASAP7_75t_SL g2905 ( 
.A1(n_2901),
.A2(n_193),
.B(n_197),
.Y(n_2905)
);

NAND3xp33_ASAP7_75t_L g2906 ( 
.A(n_2898),
.B(n_865),
.C(n_203),
.Y(n_2906)
);

AOI22xp33_ASAP7_75t_L g2907 ( 
.A1(n_2897),
.A2(n_871),
.B1(n_1229),
.B2(n_1249),
.Y(n_2907)
);

AOI21xp5_ASAP7_75t_L g2908 ( 
.A1(n_2899),
.A2(n_202),
.B(n_207),
.Y(n_2908)
);

AND2x2_ASAP7_75t_L g2909 ( 
.A(n_2900),
.B(n_212),
.Y(n_2909)
);

AOI221xp5_ASAP7_75t_SL g2910 ( 
.A1(n_2908),
.A2(n_2902),
.B1(n_2903),
.B2(n_221),
.C(n_229),
.Y(n_2910)
);

OAI222xp33_ASAP7_75t_L g2911 ( 
.A1(n_2909),
.A2(n_2904),
.B1(n_2905),
.B2(n_2906),
.C1(n_2907),
.C2(n_235),
.Y(n_2911)
);

INVx1_ASAP7_75t_SL g2912 ( 
.A(n_2909),
.Y(n_2912)
);

OAI222xp33_ASAP7_75t_L g2913 ( 
.A1(n_2908),
.A2(n_214),
.B1(n_217),
.B2(n_231),
.C1(n_234),
.C2(n_240),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_2909),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2909),
.Y(n_2915)
);

AOI21x1_ASAP7_75t_L g2916 ( 
.A1(n_2914),
.A2(n_243),
.B(n_244),
.Y(n_2916)
);

NOR2xp67_ASAP7_75t_SL g2917 ( 
.A(n_2915),
.B(n_247),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2912),
.Y(n_2918)
);

AOI222xp33_ASAP7_75t_SL g2919 ( 
.A1(n_2910),
.A2(n_1249),
.B1(n_1229),
.B2(n_871),
.C1(n_251),
.C2(n_254),
.Y(n_2919)
);

OAI22xp5_ASAP7_75t_L g2920 ( 
.A1(n_2911),
.A2(n_248),
.B1(n_249),
.B2(n_250),
.Y(n_2920)
);

AOI22xp33_ASAP7_75t_L g2921 ( 
.A1(n_2918),
.A2(n_2913),
.B1(n_871),
.B2(n_1110),
.Y(n_2921)
);

AOI22xp5_ASAP7_75t_SL g2922 ( 
.A1(n_2920),
.A2(n_871),
.B1(n_262),
.B2(n_263),
.Y(n_2922)
);

AOI22xp5_ASAP7_75t_SL g2923 ( 
.A1(n_2917),
.A2(n_260),
.B1(n_264),
.B2(n_266),
.Y(n_2923)
);

OAI21xp5_ASAP7_75t_L g2924 ( 
.A1(n_2921),
.A2(n_2916),
.B(n_2919),
.Y(n_2924)
);

AO21x2_ASAP7_75t_L g2925 ( 
.A1(n_2923),
.A2(n_267),
.B(n_268),
.Y(n_2925)
);

OAI22x1_ASAP7_75t_L g2926 ( 
.A1(n_2925),
.A2(n_2922),
.B1(n_270),
.B2(n_273),
.Y(n_2926)
);

AOI211xp5_ASAP7_75t_L g2927 ( 
.A1(n_2926),
.A2(n_2924),
.B(n_274),
.C(n_278),
.Y(n_2927)
);


endmodule