module fake_jpeg_2226_n_579 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_579);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_579;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_18),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

INVxp33_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_6),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_17),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_15),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_9),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_62),
.B(n_78),
.Y(n_143)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_63),
.Y(n_148)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_64),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_19),
.B(n_9),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_65),
.B(n_69),
.Y(n_126)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_66),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_67),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_21),
.B(n_22),
.C(n_43),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_68),
.B(n_114),
.C(n_28),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_20),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_70),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_71),
.Y(n_164)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g198 ( 
.A(n_72),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_73),
.Y(n_168)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_74),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_75),
.Y(n_188)
);

BUFx8_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_76),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

INVx3_ASAP7_75t_SL g191 ( 
.A(n_77),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_29),
.B(n_10),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_30),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_79),
.B(n_1),
.Y(n_190)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_80),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_21),
.B(n_8),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_81),
.B(n_85),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_82),
.Y(n_154)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_83),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_25),
.Y(n_84)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_84),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_26),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_87),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_42),
.B(n_8),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_88),
.B(n_98),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_22),
.Y(n_89)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_89),
.Y(n_160)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_90),
.Y(n_145)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_91),
.Y(n_149)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_35),
.Y(n_92)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_92),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_23),
.Y(n_93)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_93),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_32),
.Y(n_94)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_94),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_32),
.Y(n_95)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_95),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_32),
.Y(n_96)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_96),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_26),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_97),
.B(n_101),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_43),
.B(n_18),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_47),
.B(n_1),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_99),
.B(n_110),
.Y(n_173)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_49),
.Y(n_100)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_26),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_102),
.Y(n_187)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_51),
.Y(n_104)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_104),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_50),
.B(n_8),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_105),
.B(n_111),
.Y(n_151)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_106),
.Y(n_200)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_107),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_40),
.Y(n_108)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_108),
.Y(n_178)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_46),
.Y(n_109)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_109),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_55),
.B(n_57),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_45),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_50),
.Y(n_112)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_112),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_27),
.B(n_18),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_113),
.B(n_117),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_54),
.B(n_18),
.C(n_8),
.Y(n_114)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_30),
.Y(n_115)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_115),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_52),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g159 ( 
.A(n_116),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_27),
.B(n_17),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_118),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_40),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_119),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_54),
.B(n_40),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_120),
.B(n_121),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_54),
.B(n_1),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_45),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_24),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_30),
.Y(n_123)
);

BUFx4f_ASAP7_75t_L g197 ( 
.A(n_123),
.Y(n_197)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_30),
.Y(n_124)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_124),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_76),
.B(n_58),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_125),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_127),
.B(n_128),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_68),
.B(n_28),
.C(n_58),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_121),
.A2(n_57),
.B1(n_39),
.B2(n_59),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_133),
.A2(n_176),
.B1(n_180),
.B2(n_144),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_99),
.A2(n_33),
.B1(n_59),
.B2(n_48),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_137),
.A2(n_189),
.B1(n_193),
.B2(n_124),
.Y(n_205)
);

OAI21xp33_ASAP7_75t_L g141 ( 
.A1(n_105),
.A2(n_39),
.B(n_37),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_141),
.B(n_3),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_76),
.A2(n_30),
.B1(n_37),
.B2(n_44),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_144),
.A2(n_147),
.B1(n_170),
.B2(n_180),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_81),
.A2(n_60),
.B1(n_19),
.B2(n_24),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_146),
.A2(n_157),
.B1(n_169),
.B2(n_201),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_79),
.A2(n_44),
.B1(n_48),
.B2(n_31),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_153),
.B(n_194),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_106),
.A2(n_33),
.B1(n_31),
.B2(n_56),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_72),
.B(n_13),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_166),
.B(n_172),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_112),
.A2(n_56),
.B1(n_46),
.B2(n_41),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_70),
.A2(n_56),
.B1(n_46),
.B2(n_34),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_70),
.B(n_12),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_82),
.B(n_12),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_174),
.B(n_175),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_82),
.B(n_7),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_120),
.A2(n_7),
.B1(n_16),
.B2(n_14),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_102),
.B(n_7),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_179),
.B(n_183),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_115),
.A2(n_34),
.B1(n_41),
.B2(n_7),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_66),
.B(n_13),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_77),
.A2(n_34),
.B1(n_41),
.B2(n_13),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_190),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_114),
.A2(n_41),
.B1(n_13),
.B2(n_4),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_123),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_84),
.A2(n_41),
.B1(n_5),
.B2(n_14),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_86),
.B(n_5),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_63),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_87),
.A2(n_16),
.B1(n_2),
.B2(n_3),
.Y(n_203)
);

OAI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_203),
.A2(n_94),
.B1(n_95),
.B2(n_71),
.Y(n_235)
);

INVx2_ASAP7_75t_SL g204 ( 
.A(n_198),
.Y(n_204)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_204),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_205),
.A2(n_269),
.B1(n_208),
.B2(n_242),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_92),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_206),
.B(n_219),
.Y(n_283)
);

AOI21xp33_ASAP7_75t_L g207 ( 
.A1(n_151),
.A2(n_109),
.B(n_89),
.Y(n_207)
);

OAI21xp33_ASAP7_75t_L g290 ( 
.A1(n_207),
.A2(n_213),
.B(n_238),
.Y(n_290)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_165),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_209),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_171),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g316 ( 
.A(n_210),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_139),
.A2(n_90),
.B1(n_74),
.B2(n_91),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_212),
.Y(n_287)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_156),
.Y(n_214)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_214),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_126),
.B(n_80),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_215),
.B(n_221),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_128),
.A2(n_195),
.B1(n_140),
.B2(n_61),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_216),
.A2(n_252),
.B1(n_258),
.B2(n_262),
.Y(n_284)
);

AO22x1_ASAP7_75t_L g217 ( 
.A1(n_190),
.A2(n_116),
.B1(n_93),
.B2(n_108),
.Y(n_217)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_217),
.Y(n_281)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_182),
.Y(n_218)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_218),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_127),
.B(n_96),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_132),
.Y(n_220)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_220),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_129),
.B(n_142),
.Y(n_221)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_155),
.Y(n_224)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_224),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_150),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_225),
.B(n_243),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_145),
.Y(n_227)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_227),
.Y(n_327)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_156),
.Y(n_228)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_228),
.Y(n_325)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_200),
.Y(n_230)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_230),
.Y(n_312)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_187),
.Y(n_231)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_231),
.Y(n_328)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_134),
.Y(n_232)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_232),
.Y(n_329)
);

AOI32xp33_ASAP7_75t_L g233 ( 
.A1(n_173),
.A2(n_75),
.A3(n_119),
.B1(n_73),
.B2(n_67),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_233),
.B(n_255),
.Y(n_285)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_145),
.Y(n_234)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_234),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_235),
.A2(n_265),
.B1(n_217),
.B2(n_241),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_163),
.B(n_2),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_236),
.B(n_240),
.Y(n_302)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_130),
.Y(n_237)
);

INVx4_ASAP7_75t_L g296 ( 
.A(n_237),
.Y(n_296)
);

A2O1A1Ixp33_ASAP7_75t_L g238 ( 
.A1(n_143),
.A2(n_3),
.B(n_16),
.C(n_181),
.Y(n_238)
);

BUFx12f_ASAP7_75t_L g239 ( 
.A(n_130),
.Y(n_239)
);

INVx11_ASAP7_75t_L g288 ( 
.A(n_239),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_141),
.B(n_3),
.Y(n_240)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_136),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_176),
.B(n_133),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_244),
.B(n_257),
.Y(n_304)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_149),
.Y(n_245)
);

INVx4_ASAP7_75t_L g332 ( 
.A(n_245),
.Y(n_332)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_158),
.Y(n_246)
);

BUFx12f_ASAP7_75t_L g313 ( 
.A(n_246),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_247),
.A2(n_160),
.B1(n_196),
.B2(n_167),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_177),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_248),
.B(n_254),
.Y(n_317)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_158),
.Y(n_249)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_249),
.Y(n_292)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_131),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_250),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_125),
.B(n_149),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_251),
.B(n_256),
.C(n_196),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_195),
.A2(n_140),
.B1(n_184),
.B2(n_138),
.Y(n_252)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_165),
.Y(n_253)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_253),
.Y(n_311)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_162),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_170),
.Y(n_255)
);

AND2x2_ASAP7_75t_SL g256 ( 
.A(n_199),
.B(n_140),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_146),
.B(n_147),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_161),
.A2(n_178),
.B1(n_198),
.B2(n_159),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_161),
.B(n_178),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_259),
.B(n_266),
.Y(n_305)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_135),
.Y(n_260)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_260),
.Y(n_323)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_191),
.Y(n_261)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_261),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_148),
.A2(n_152),
.B1(n_131),
.B2(n_188),
.Y(n_262)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_148),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_267),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_135),
.B(n_186),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_268),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_152),
.B(n_197),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_191),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_186),
.B(n_192),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_188),
.A2(n_197),
.B1(n_192),
.B2(n_154),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_167),
.B(n_164),
.Y(n_271)
);

OAI32xp33_ASAP7_75t_L g291 ( 
.A1(n_271),
.A2(n_168),
.A3(n_264),
.B1(n_268),
.B2(n_206),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_171),
.Y(n_272)
);

INVx8_ASAP7_75t_L g299 ( 
.A(n_272),
.Y(n_299)
);

INVx6_ASAP7_75t_L g273 ( 
.A(n_164),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_273),
.Y(n_275)
);

NAND2xp33_ASAP7_75t_SL g274 ( 
.A(n_154),
.B(n_160),
.Y(n_274)
);

BUFx8_ASAP7_75t_L g309 ( 
.A(n_274),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_276),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_277),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_255),
.A2(n_257),
.B1(n_265),
.B2(n_251),
.Y(n_278)
);

AO21x1_ASAP7_75t_L g373 ( 
.A1(n_278),
.A2(n_282),
.B(n_316),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_251),
.A2(n_168),
.B1(n_197),
.B2(n_217),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_291),
.B(n_239),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_300),
.A2(n_294),
.B1(n_324),
.B2(n_326),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_241),
.A2(n_219),
.B1(n_244),
.B2(n_205),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_303),
.A2(n_307),
.B1(n_315),
.B2(n_319),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_223),
.B(n_226),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_306),
.Y(n_354)
);

AO22x1_ASAP7_75t_SL g308 ( 
.A1(n_241),
.A2(n_247),
.B1(n_242),
.B2(n_229),
.Y(n_308)
);

OA21x2_ASAP7_75t_L g334 ( 
.A1(n_308),
.A2(n_204),
.B(n_261),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_270),
.B(n_211),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_310),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_232),
.B(n_243),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_314),
.B(n_331),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_240),
.A2(n_222),
.B1(n_247),
.B2(n_236),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_254),
.B(n_218),
.C(n_231),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_318),
.B(n_330),
.C(n_286),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_271),
.A2(n_273),
.B1(n_238),
.B2(n_260),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_256),
.A2(n_224),
.B1(n_220),
.B2(n_214),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_320),
.A2(n_322),
.B1(n_239),
.B2(n_280),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_256),
.A2(n_204),
.B(n_249),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g355 ( 
.A1(n_321),
.A2(n_309),
.B(n_287),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_210),
.A2(n_272),
.B1(n_230),
.B2(n_228),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_234),
.B(n_237),
.C(n_245),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_263),
.B(n_246),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_334),
.B(n_371),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_307),
.A2(n_267),
.B1(n_250),
.B2(n_253),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_335),
.A2(n_344),
.B1(n_348),
.B2(n_350),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_278),
.A2(n_239),
.B(n_209),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_336),
.A2(n_355),
.B(n_363),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_337),
.B(n_346),
.Y(n_389)
);

BUFx2_ASAP7_75t_L g394 ( 
.A(n_340),
.Y(n_394)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_280),
.Y(n_342)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_342),
.Y(n_381)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_292),
.Y(n_343)
);

INVx2_ASAP7_75t_SL g398 ( 
.A(n_343),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_304),
.A2(n_285),
.B1(n_283),
.B2(n_281),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_323),
.Y(n_345)
);

INVx1_ASAP7_75t_SL g411 ( 
.A(n_345),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_283),
.B(n_303),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_304),
.A2(n_281),
.B1(n_279),
.B2(n_291),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_329),
.Y(n_349)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_349),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_279),
.A2(n_282),
.B1(n_290),
.B2(n_308),
.Y(n_350)
);

O2A1O1Ixp33_ASAP7_75t_L g351 ( 
.A1(n_309),
.A2(n_287),
.B(n_277),
.C(n_308),
.Y(n_351)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_351),
.A2(n_373),
.B(n_350),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_302),
.B(n_319),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_352),
.B(n_356),
.Y(n_392)
);

BUFx24_ASAP7_75t_SL g353 ( 
.A(n_293),
.Y(n_353)
);

BUFx24_ASAP7_75t_SL g406 ( 
.A(n_353),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_302),
.B(n_305),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_321),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_357),
.B(n_359),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_318),
.B(n_317),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_358),
.B(n_364),
.Y(n_395)
);

INVx1_ASAP7_75t_SL g359 ( 
.A(n_309),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_326),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_360),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_295),
.B(n_327),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_361),
.B(n_373),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_329),
.B(n_320),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_362),
.B(n_313),
.C(n_288),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_L g363 ( 
.A1(n_284),
.A2(n_297),
.B(n_276),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_297),
.B(n_312),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_298),
.B(n_312),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_365),
.B(n_367),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_275),
.A2(n_328),
.B1(n_301),
.B2(n_298),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_366),
.A2(n_375),
.B1(n_342),
.B2(n_349),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_301),
.B(n_328),
.Y(n_367)
);

AOI32xp33_ASAP7_75t_L g368 ( 
.A1(n_289),
.A2(n_333),
.A3(n_332),
.B1(n_296),
.B2(n_286),
.Y(n_368)
);

A2O1A1O1Ixp25_ASAP7_75t_L g393 ( 
.A1(n_368),
.A2(n_313),
.B(n_351),
.C(n_337),
.D(n_369),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_333),
.A2(n_330),
.B(n_323),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_369),
.A2(n_357),
.B(n_355),
.Y(n_402)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_292),
.Y(n_370)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_370),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_316),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_374),
.B(n_376),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_299),
.A2(n_311),
.B1(n_324),
.B2(n_325),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_325),
.B(n_311),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_377),
.A2(n_378),
.B1(n_288),
.B2(n_313),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_299),
.A2(n_296),
.B1(n_332),
.B2(n_294),
.Y(n_378)
);

BUFx3_ASAP7_75t_L g423 ( 
.A(n_379),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_376),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_382),
.B(n_414),
.Y(n_442)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_383),
.Y(n_418)
);

CKINVDCx14_ASAP7_75t_R g385 ( 
.A(n_336),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_385),
.B(n_387),
.Y(n_422)
);

CKINVDCx14_ASAP7_75t_R g387 ( 
.A(n_338),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_388),
.B(n_390),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_SL g390 ( 
.A(n_346),
.B(n_313),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g434 ( 
.A1(n_393),
.A2(n_407),
.B(n_412),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_339),
.A2(n_352),
.B1(n_341),
.B2(n_348),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_396),
.A2(n_380),
.B1(n_395),
.B2(n_389),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_SL g399 ( 
.A(n_344),
.B(n_341),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_399),
.B(n_396),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_402),
.Y(n_419)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_366),
.Y(n_404)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_404),
.Y(n_421)
);

OA21x2_ASAP7_75t_L g417 ( 
.A1(n_405),
.A2(n_340),
.B(n_368),
.Y(n_417)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_351),
.A2(n_359),
.B(n_373),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_364),
.Y(n_408)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_408),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_334),
.A2(n_339),
.B(n_363),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_334),
.A2(n_335),
.B1(n_362),
.B2(n_377),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_413),
.A2(n_415),
.B1(n_391),
.B2(n_394),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_365),
.Y(n_414)
);

AOI22xp33_ASAP7_75t_L g415 ( 
.A1(n_347),
.A2(n_367),
.B1(n_372),
.B2(n_334),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_345),
.Y(n_416)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_416),
.Y(n_431)
);

OAI21xp5_ASAP7_75t_SL g465 ( 
.A1(n_417),
.A2(n_438),
.B(n_400),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_420),
.A2(n_385),
.B1(n_386),
.B2(n_393),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_403),
.B(n_374),
.C(n_358),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_424),
.B(n_430),
.C(n_446),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_387),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_426),
.B(n_435),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_410),
.B(n_356),
.Y(n_427)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_427),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_410),
.B(n_414),
.Y(n_428)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_428),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_408),
.B(n_343),
.Y(n_429)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_429),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_403),
.B(n_370),
.C(n_354),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_380),
.A2(n_378),
.B1(n_371),
.B2(n_360),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_432),
.A2(n_440),
.B1(n_413),
.B2(n_394),
.Y(n_449)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_381),
.Y(n_433)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_433),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_383),
.Y(n_435)
);

OA21x2_ASAP7_75t_L g437 ( 
.A1(n_405),
.A2(n_391),
.B(n_412),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_437),
.B(n_444),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_386),
.A2(n_375),
.B(n_360),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_SL g456 ( 
.A(n_439),
.B(n_390),
.Y(n_456)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_381),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_441),
.B(n_445),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_395),
.B(n_401),
.Y(n_443)
);

CKINVDCx14_ASAP7_75t_R g452 ( 
.A(n_443),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_382),
.B(n_404),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_398),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_399),
.B(n_389),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_397),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_447),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_392),
.B(n_397),
.Y(n_448)
);

CKINVDCx16_ASAP7_75t_R g451 ( 
.A(n_448),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_449),
.A2(n_450),
.B1(n_455),
.B2(n_462),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_418),
.A2(n_384),
.B1(n_407),
.B2(n_394),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_435),
.A2(n_392),
.B1(n_391),
.B2(n_402),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_SL g500 ( 
.A(n_456),
.B(n_438),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_424),
.B(n_388),
.C(n_384),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_457),
.B(n_467),
.C(n_468),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_461),
.A2(n_437),
.B1(n_438),
.B2(n_448),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_418),
.A2(n_393),
.B1(n_379),
.B2(n_400),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_444),
.A2(n_420),
.B1(n_440),
.B2(n_417),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_463),
.A2(n_476),
.B1(n_437),
.B2(n_425),
.Y(n_495)
);

A2O1A1Ixp33_ASAP7_75t_SL g481 ( 
.A1(n_465),
.A2(n_437),
.B(n_417),
.C(n_422),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_434),
.A2(n_401),
.B(n_398),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_466),
.A2(n_426),
.B(n_432),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_424),
.B(n_416),
.C(n_411),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_430),
.B(n_411),
.C(n_398),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_439),
.B(n_409),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_471),
.B(n_472),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_439),
.B(n_406),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_446),
.B(n_430),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_474),
.B(n_457),
.Y(n_496)
);

CKINVDCx16_ASAP7_75t_R g475 ( 
.A(n_422),
.Y(n_475)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_475),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_417),
.A2(n_425),
.B1(n_421),
.B2(n_442),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_464),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_478),
.B(n_481),
.Y(n_510)
);

FAx1_ASAP7_75t_SL g480 ( 
.A(n_456),
.B(n_434),
.CI(n_446),
.CON(n_480),
.SN(n_480)
);

XOR2x1_ASAP7_75t_L g522 ( 
.A(n_480),
.B(n_471),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_453),
.B(n_436),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g505 ( 
.A(n_482),
.B(n_487),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_452),
.B(n_442),
.Y(n_483)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_483),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_475),
.B(n_443),
.Y(n_484)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_484),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_458),
.B(n_427),
.Y(n_485)
);

NAND3xp33_ASAP7_75t_L g509 ( 
.A(n_485),
.B(n_492),
.C(n_458),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_453),
.B(n_436),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_467),
.B(n_436),
.C(n_419),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_488),
.B(n_490),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_464),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_470),
.Y(n_491)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_491),
.Y(n_507)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_454),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_470),
.Y(n_493)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_493),
.Y(n_508)
);

HAxp5_ASAP7_75t_SL g494 ( 
.A(n_454),
.B(n_428),
.CON(n_494),
.SN(n_494)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_494),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_495),
.A2(n_462),
.B1(n_463),
.B2(n_449),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_496),
.B(n_500),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g497 ( 
.A(n_466),
.Y(n_497)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_497),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g518 ( 
.A(n_498),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_474),
.B(n_429),
.C(n_421),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_499),
.B(n_468),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_SL g517 ( 
.A1(n_501),
.A2(n_465),
.B(n_473),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_483),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_504),
.B(n_506),
.Y(n_530)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_509),
.A2(n_511),
.B1(n_520),
.B2(n_459),
.Y(n_532)
);

AO221x1_ASAP7_75t_L g512 ( 
.A1(n_498),
.A2(n_450),
.B1(n_469),
.B2(n_476),
.C(n_451),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_512),
.B(n_486),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g515 ( 
.A(n_496),
.B(n_472),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_515),
.B(n_522),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_517),
.B(n_501),
.Y(n_527)
);

INVxp67_ASAP7_75t_SL g519 ( 
.A(n_484),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_519),
.B(n_459),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_477),
.A2(n_461),
.B1(n_473),
.B2(n_451),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_514),
.A2(n_479),
.B(n_488),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g546 ( 
.A1(n_523),
.A2(n_526),
.B1(n_528),
.B2(n_497),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_513),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_524),
.B(n_535),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g548 ( 
.A1(n_525),
.A2(n_532),
.B1(n_534),
.B2(n_460),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_502),
.A2(n_518),
.B1(n_503),
.B2(n_511),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g543 ( 
.A(n_527),
.B(n_529),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_518),
.A2(n_423),
.B1(n_469),
.B2(n_478),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_506),
.B(n_482),
.Y(n_529)
);

BUFx24_ASAP7_75t_SL g533 ( 
.A(n_515),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_533),
.B(n_505),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_505),
.B(n_479),
.C(n_487),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_516),
.B(n_489),
.Y(n_536)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_536),
.B(n_537),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_SL g537 ( 
.A(n_516),
.B(n_500),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_520),
.B(n_499),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_538),
.B(n_481),
.Y(n_539)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_539),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_540),
.B(n_544),
.Y(n_554)
);

XOR2xp5_ASAP7_75t_L g542 ( 
.A(n_536),
.B(n_522),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_542),
.B(n_547),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_538),
.A2(n_510),
.B1(n_521),
.B2(n_481),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_529),
.B(n_517),
.C(n_489),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_545),
.B(n_549),
.C(n_527),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_546),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_535),
.B(n_507),
.Y(n_547)
);

OAI22xp5_ASAP7_75t_L g560 ( 
.A1(n_548),
.A2(n_549),
.B1(n_551),
.B2(n_508),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_530),
.B(n_510),
.C(n_455),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_SL g550 ( 
.A1(n_524),
.A2(n_481),
.B1(n_423),
.B2(n_460),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_550),
.B(n_423),
.Y(n_556)
);

AO21x1_ASAP7_75t_L g552 ( 
.A1(n_539),
.A2(n_481),
.B(n_494),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_SL g564 ( 
.A1(n_552),
.A2(n_542),
.B(n_550),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_555),
.B(n_560),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_556),
.B(n_558),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_543),
.B(n_531),
.C(n_537),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_543),
.B(n_445),
.C(n_431),
.Y(n_561)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_561),
.A2(n_541),
.B(n_431),
.Y(n_567)
);

OAI21xp5_ASAP7_75t_L g562 ( 
.A1(n_559),
.A2(n_545),
.B(n_544),
.Y(n_562)
);

AOI21xp5_ASAP7_75t_L g572 ( 
.A1(n_562),
.A2(n_564),
.B(n_566),
.Y(n_572)
);

OAI21xp5_ASAP7_75t_SL g566 ( 
.A1(n_553),
.A2(n_541),
.B(n_493),
.Y(n_566)
);

INVxp67_ASAP7_75t_L g570 ( 
.A(n_567),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_SL g568 ( 
.A(n_554),
.B(n_558),
.Y(n_568)
);

NAND2xp33_ASAP7_75t_SL g571 ( 
.A(n_568),
.B(n_561),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g569 ( 
.A(n_565),
.B(n_555),
.C(n_557),
.Y(n_569)
);

AOI21xp5_ASAP7_75t_L g573 ( 
.A1(n_569),
.A2(n_563),
.B(n_552),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_571),
.Y(n_574)
);

INVxp33_ASAP7_75t_L g575 ( 
.A(n_573),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_574),
.B(n_572),
.C(n_563),
.Y(n_576)
);

OAI321xp33_ASAP7_75t_L g577 ( 
.A1(n_576),
.A2(n_570),
.A3(n_441),
.B1(n_447),
.B2(n_433),
.C(n_480),
.Y(n_577)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_577),
.B(n_575),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_578),
.B(n_480),
.Y(n_579)
);


endmodule