module fake_netlist_1_8318_n_13 (n_1, n_2, n_0, n_13);
input n_1;
input n_2;
input n_0;
output n_13;
wire n_11;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
BUFx6f_ASAP7_75t_L g3 ( .A(n_2), .Y(n_3) );
NOR2xp33_ASAP7_75t_L g4 ( .A(n_2), .B(n_0), .Y(n_4) );
AND2x2_ASAP7_75t_L g5 ( .A(n_3), .B(n_2), .Y(n_5) );
INVx2_ASAP7_75t_L g6 ( .A(n_3), .Y(n_6) );
OR2x2_ASAP7_75t_L g7 ( .A(n_5), .B(n_0), .Y(n_7) );
OR2x2_ASAP7_75t_L g8 ( .A(n_6), .B(n_0), .Y(n_8) );
OAI21xp5_ASAP7_75t_SL g9 ( .A1(n_7), .A2(n_4), .B(n_1), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_8), .Y(n_10) );
NAND3xp33_ASAP7_75t_L g11 ( .A(n_9), .B(n_1), .C(n_10), .Y(n_11) );
INVx2_ASAP7_75t_SL g12 ( .A(n_11), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_12), .Y(n_13) );
endmodule