module fake_jpeg_29144_n_367 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_367);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_367;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_21),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_8),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_25),
.B(n_0),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_50),
.Y(n_73)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_24),
.B(n_0),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_36),
.B(n_20),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_51),
.B(n_55),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_36),
.B(n_20),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g56 ( 
.A(n_29),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_56),
.Y(n_79)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_61),
.Y(n_108)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g64 ( 
.A(n_24),
.B(n_1),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_68),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_37),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_82),
.B(n_104),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_48),
.A2(n_44),
.B1(n_45),
.B2(n_22),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_83),
.A2(n_43),
.B1(n_42),
.B2(n_25),
.Y(n_121)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_84),
.Y(n_109)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_63),
.Y(n_87)
);

BUFx2_ASAP7_75t_SL g134 ( 
.A(n_87),
.Y(n_134)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_88),
.Y(n_129)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_94),
.Y(n_126)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_95),
.Y(n_124)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_54),
.Y(n_96)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

AO22x2_ASAP7_75t_L g97 ( 
.A1(n_49),
.A2(n_34),
.B1(n_23),
.B2(n_43),
.Y(n_97)
);

OA22x2_ASAP7_75t_L g118 ( 
.A1(n_97),
.A2(n_56),
.B1(n_23),
.B2(n_68),
.Y(n_118)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_58),
.Y(n_100)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_102),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_64),
.B(n_35),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_105),
.Y(n_110)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_107),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_97),
.A2(n_69),
.B1(n_65),
.B2(n_60),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_111),
.A2(n_121),
.B1(n_131),
.B2(n_139),
.Y(n_148)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_77),
.B(n_48),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_113),
.B(n_137),
.C(n_140),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_118),
.B(n_128),
.Y(n_157)
);

A2O1A1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_73),
.A2(n_41),
.B(n_40),
.C(n_32),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_L g160 ( 
.A1(n_123),
.A2(n_138),
.B(n_40),
.C(n_41),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_127),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_78),
.A2(n_27),
.B1(n_32),
.B2(n_31),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_101),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_130),
.B(n_135),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_73),
.A2(n_69),
.B1(n_65),
.B2(n_46),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_71),
.B(n_39),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_70),
.Y(n_136)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_42),
.Y(n_137)
);

HAxp5_ASAP7_75t_SL g138 ( 
.A(n_97),
.B(n_35),
.CON(n_138),
.SN(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_80),
.A2(n_38),
.B1(n_46),
.B2(n_45),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_93),
.B(n_39),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_101),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_141),
.B(n_79),
.Y(n_146)
);

O2A1O1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_138),
.A2(n_79),
.B(n_87),
.C(n_37),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_142),
.Y(n_176)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_143),
.B(n_144),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_134),
.Y(n_144)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_119),
.Y(n_145)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_145),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_146),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_93),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_147),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_137),
.A2(n_85),
.B(n_89),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_150),
.A2(n_160),
.B(n_137),
.Y(n_177)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_109),
.Y(n_151)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_151),
.Y(n_171)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_152),
.Y(n_173)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_122),
.Y(n_154)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_154),
.Y(n_185)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_156),
.B(n_159),
.Y(n_183)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_122),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_132),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_161),
.B(n_163),
.Y(n_172)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_119),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_166),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_135),
.Y(n_163)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_132),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_113),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_178),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_142),
.A2(n_128),
.B(n_110),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_170),
.A2(n_118),
.B(n_139),
.Y(n_195)
);

A2O1A1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_160),
.A2(n_113),
.B(n_118),
.C(n_123),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_174),
.A2(n_150),
.B(n_164),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_177),
.B(n_174),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_116),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_157),
.A2(n_148),
.B1(n_131),
.B2(n_118),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_181),
.A2(n_184),
.B1(n_80),
.B2(n_59),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_157),
.A2(n_148),
.B1(n_121),
.B2(n_164),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_186),
.B(n_179),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_166),
.C(n_154),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_187),
.B(n_191),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_188),
.A2(n_190),
.B(n_193),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_168),
.A2(n_162),
.B1(n_145),
.B2(n_149),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_184),
.B(n_112),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_185),
.Y(n_192)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_192),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_168),
.A2(n_149),
.B1(n_125),
.B2(n_165),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_185),
.Y(n_194)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_194),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_195),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_151),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_196),
.B(n_198),
.Y(n_209)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_197),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_174),
.B(n_153),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_178),
.B(n_117),
.C(n_156),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_199),
.B(n_167),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_201),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_176),
.A2(n_127),
.B1(n_133),
.B2(n_117),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_176),
.A2(n_125),
.B1(n_165),
.B2(n_158),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_202),
.A2(n_158),
.B1(n_167),
.B2(n_92),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_182),
.B(n_126),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_172),
.Y(n_221)
);

FAx1_ASAP7_75t_SL g204 ( 
.A(n_170),
.B(n_152),
.CI(n_75),
.CON(n_204),
.SN(n_204)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_204),
.B(n_172),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_207),
.A2(n_220),
.B1(n_167),
.B2(n_183),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_187),
.C(n_199),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_188),
.A2(n_177),
.B(n_181),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_212),
.A2(n_186),
.B(n_204),
.Y(n_234)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_197),
.Y(n_213)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_213),
.Y(n_226)
);

AO21x1_ASAP7_75t_L g240 ( 
.A1(n_214),
.A2(n_224),
.B(n_175),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_201),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_215),
.Y(n_245)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_192),
.Y(n_218)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_218),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_198),
.A2(n_200),
.B1(n_189),
.B2(n_202),
.Y(n_220)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_221),
.Y(n_236)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_194),
.Y(n_222)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_222),
.Y(n_238)
);

BUFx24_ASAP7_75t_SL g223 ( 
.A(n_203),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_223),
.Y(n_230)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_196),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_225),
.B(n_180),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g227 ( 
.A(n_225),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_227),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_228),
.B(n_237),
.C(n_211),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_215),
.A2(n_195),
.B1(n_189),
.B2(n_191),
.Y(n_229)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_229),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_231),
.A2(n_246),
.B1(n_208),
.B2(n_205),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_221),
.A2(n_209),
.B1(n_211),
.B2(n_224),
.Y(n_232)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_232),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_233),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_234),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_206),
.B(n_204),
.C(n_180),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_209),
.B(n_204),
.Y(n_239)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_239),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_240),
.B(n_244),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_206),
.B(n_175),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_247),
.Y(n_261)
);

AO22x1_ASAP7_75t_L g242 ( 
.A1(n_219),
.A2(n_167),
.B1(n_183),
.B2(n_171),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_242),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_210),
.B(n_183),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_243),
.B(n_234),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_173),
.Y(n_244)
);

OA22x2_ASAP7_75t_L g246 ( 
.A1(n_212),
.A2(n_173),
.B1(n_120),
.B2(n_115),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_120),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_244),
.A2(n_236),
.B1(n_207),
.B2(n_216),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_250),
.A2(n_246),
.B1(n_115),
.B2(n_92),
.Y(n_284)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_233),
.Y(n_254)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_254),
.Y(n_272)
);

INVxp33_ASAP7_75t_L g256 ( 
.A(n_239),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_256),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_257),
.B(n_264),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_230),
.B(n_218),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_258),
.Y(n_287)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_227),
.Y(n_259)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_259),
.Y(n_279)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_235),
.Y(n_263)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_263),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_228),
.B(n_241),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_264),
.B(n_271),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_222),
.C(n_217),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_266),
.C(n_247),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_237),
.B(n_217),
.C(n_208),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_238),
.Y(n_267)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_267),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_268),
.A2(n_269),
.B1(n_244),
.B2(n_245),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_231),
.A2(n_205),
.B1(n_136),
.B2(n_23),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_226),
.B(n_31),
.Y(n_270)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_270),
.Y(n_282)
);

NOR2xp67_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_240),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g295 ( 
.A(n_274),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_257),
.B(n_19),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_275),
.B(n_278),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_276),
.B(n_283),
.C(n_271),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_277),
.A2(n_255),
.B1(n_268),
.B2(n_269),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_246),
.C(n_242),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_284),
.B(n_256),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_261),
.B(n_265),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_285),
.B(n_261),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_248),
.A2(n_253),
.B1(n_250),
.B2(n_249),
.Y(n_286)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_286),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_262),
.A2(n_246),
.B(n_2),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_288),
.A2(n_290),
.B(n_291),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_262),
.A2(n_91),
.B(n_81),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_255),
.A2(n_91),
.B(n_81),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_252),
.Y(n_292)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_292),
.Y(n_297)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_280),
.Y(n_293)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_293),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_294),
.B(n_298),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_260),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_299),
.B(n_301),
.Y(n_321)
);

INVxp67_ASAP7_75t_SL g300 ( 
.A(n_272),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_300),
.B(n_305),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_307),
.Y(n_317)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_282),
.Y(n_304)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_304),
.Y(n_316)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_281),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_278),
.B(n_74),
.C(n_76),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_308),
.C(n_285),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_277),
.A2(n_28),
.B1(n_22),
.B2(n_45),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_276),
.B(n_76),
.C(n_28),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_302),
.Y(n_326)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_296),
.B(n_283),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_314),
.B(n_318),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_298),
.B(n_308),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_315),
.B(n_319),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_290),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_289),
.C(n_273),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_295),
.B(n_279),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_323),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_302),
.A2(n_288),
.B1(n_291),
.B2(n_289),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_322),
.A2(n_318),
.B1(n_310),
.B2(n_17),
.Y(n_335)
);

BUFx24_ASAP7_75t_SL g323 ( 
.A(n_297),
.Y(n_323)
);

FAx1_ASAP7_75t_SL g324 ( 
.A(n_314),
.B(n_303),
.CI(n_301),
.CON(n_324),
.SN(n_324)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_324),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_311),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_325),
.B(n_327),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_326),
.B(n_330),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_321),
.A2(n_305),
.B(n_293),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g329 ( 
.A1(n_316),
.A2(n_22),
.B1(n_28),
.B2(n_72),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_329),
.B(n_59),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_313),
.B(n_46),
.C(n_38),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_317),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_332),
.B(n_334),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_310),
.B(n_18),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_335),
.B(n_325),
.Y(n_339)
);

AOI21xp33_ASAP7_75t_L g336 ( 
.A1(n_331),
.A2(n_17),
.B(n_16),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_336),
.A2(n_4),
.B(n_5),
.Y(n_349)
);

OR2x2_ASAP7_75t_L g337 ( 
.A(n_333),
.B(n_1),
.Y(n_337)
);

AO21x1_ASAP7_75t_L g350 ( 
.A1(n_337),
.A2(n_342),
.B(n_346),
.Y(n_350)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_339),
.Y(n_348)
);

OR2x2_ASAP7_75t_L g342 ( 
.A(n_333),
.B(n_1),
.Y(n_342)
);

NOR2x1_ASAP7_75t_L g343 ( 
.A(n_324),
.B(n_2),
.Y(n_343)
);

NOR3xp33_ASAP7_75t_SL g351 ( 
.A(n_343),
.B(n_4),
.C(n_5),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_344),
.A2(n_59),
.B1(n_38),
.B2(n_10),
.Y(n_353)
);

INVxp33_ASAP7_75t_L g346 ( 
.A(n_328),
.Y(n_346)
);

INVxp33_ASAP7_75t_L g347 ( 
.A(n_338),
.Y(n_347)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_347),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_349),
.A2(n_340),
.B(n_9),
.Y(n_356)
);

NOR3xp33_ASAP7_75t_SL g357 ( 
.A(n_351),
.B(n_6),
.C(n_10),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_345),
.A2(n_6),
.B(n_7),
.Y(n_352)
);

AOI21x1_ASAP7_75t_L g359 ( 
.A1(n_352),
.A2(n_353),
.B(n_354),
.Y(n_359)
);

INVxp33_ASAP7_75t_L g354 ( 
.A(n_341),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_348),
.A2(n_342),
.B(n_337),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_355),
.B(n_356),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g360 ( 
.A(n_357),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g362 ( 
.A1(n_358),
.A2(n_350),
.B(n_11),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_362),
.B(n_10),
.C(n_11),
.Y(n_364)
);

AOI321xp33_ASAP7_75t_L g363 ( 
.A1(n_361),
.A2(n_350),
.A3(n_359),
.B1(n_12),
.B2(n_13),
.C(n_14),
.Y(n_363)
);

AO221x1_ASAP7_75t_L g365 ( 
.A1(n_363),
.A2(n_364),
.B1(n_360),
.B2(n_13),
.C(n_14),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_365),
.B(n_12),
.Y(n_366)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_366),
.B(n_14),
.Y(n_367)
);


endmodule