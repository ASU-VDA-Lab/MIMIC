module real_jpeg_5507_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_323;
wire n_215;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g62 ( 
.A(n_0),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_1),
.Y(n_75)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_1),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_1),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_2),
.A2(n_51),
.B1(n_129),
.B2(n_228),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_2),
.Y(n_228)
);

OAI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_2),
.A2(n_155),
.B1(n_228),
.B2(n_252),
.Y(n_251)
);

OAI22xp33_ASAP7_75t_SL g352 ( 
.A1(n_2),
.A2(n_228),
.B1(n_353),
.B2(n_354),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_L g376 ( 
.A1(n_2),
.A2(n_177),
.B1(n_228),
.B2(n_377),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_3),
.A2(n_27),
.B1(n_41),
.B2(n_44),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_3),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_3),
.A2(n_44),
.B1(n_120),
.B2(n_121),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_3),
.A2(n_44),
.B1(n_166),
.B2(n_168),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_3),
.A2(n_44),
.B1(n_218),
.B2(n_220),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_4),
.A2(n_27),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_4),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_4),
.A2(n_130),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_4),
.A2(n_130),
.B1(n_190),
.B2(n_192),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_4),
.A2(n_130),
.B1(n_271),
.B2(n_273),
.Y(n_270)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_5),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_6),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_6),
.Y(n_182)
);

INVx8_ASAP7_75t_L g213 ( 
.A(n_6),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_6),
.Y(n_286)
);

BUFx5_ASAP7_75t_L g392 ( 
.A(n_6),
.Y(n_392)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_7),
.Y(n_268)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_9),
.Y(n_443)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_10),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_10),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_11),
.A2(n_22),
.B1(n_83),
.B2(n_85),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_11),
.A2(n_22),
.B1(n_100),
.B2(n_102),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_11),
.A2(n_22),
.B1(n_184),
.B2(n_187),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_11),
.B(n_28),
.Y(n_281)
);

O2A1O1Ixp33_ASAP7_75t_L g337 ( 
.A1(n_11),
.A2(n_89),
.B(n_338),
.C(n_345),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_11),
.B(n_367),
.C(n_368),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_11),
.B(n_132),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_11),
.B(n_286),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_11),
.B(n_69),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_12),
.Y(n_446)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_13),
.Y(n_64)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_13),
.Y(n_67)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_13),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g367 ( 
.A(n_13),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_442),
.B(n_444),
.Y(n_14)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_138),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_137),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_52),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_19),
.B(n_53),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_39),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_20),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_28),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_21),
.B(n_45),
.Y(n_147)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_21),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B(n_25),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_22),
.B(n_26),
.Y(n_25)
);

OAI21xp33_ASAP7_75t_L g338 ( 
.A1(n_22),
.A2(n_339),
.B(n_342),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_23),
.A2(n_47),
.B1(n_49),
.B2(n_51),
.Y(n_46)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVxp33_ASAP7_75t_L g262 ( 
.A(n_25),
.Y(n_262)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2x1_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_28),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_28),
.B(n_40),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_28),
.B(n_227),
.Y(n_246)
);

AO22x2_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_31),
.B1(n_35),
.B2(n_37),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_34),
.Y(n_101)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_34),
.Y(n_105)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_34),
.Y(n_112)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_34),
.Y(n_124)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_36),
.Y(n_265)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_39),
.A2(n_127),
.B(n_128),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_39),
.B(n_246),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_45),
.Y(n_39)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_45),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_45),
.B(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_48),
.Y(n_258)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_131),
.C(n_134),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_54),
.B(n_438),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_86),
.C(n_125),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_55),
.A2(n_150),
.B1(n_151),
.B2(n_152),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_55),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_55),
.A2(n_86),
.B1(n_150),
.B2(n_236),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_55),
.A2(n_150),
.B1(n_248),
.B2(n_254),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_55),
.B(n_245),
.C(n_248),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_80),
.B(n_81),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_56),
.A2(n_189),
.B(n_196),
.Y(n_188)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_57),
.B(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_57),
.B(n_82),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_57),
.B(n_352),
.Y(n_351)
);

NOR2x1_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_69),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_63),
.B1(n_65),
.B2(n_68),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_61),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_61),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_61),
.Y(n_191)
);

INVx6_ASAP7_75t_L g344 ( 
.A(n_61),
.Y(n_344)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_62),
.Y(n_92)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_62),
.Y(n_170)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_62),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_62),
.Y(n_365)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AO22x2_ASAP7_75t_L g69 ( 
.A1(n_66),
.A2(n_70),
.B1(n_72),
.B2(n_76),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_69),
.B(n_165),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_69),
.B(n_352),
.Y(n_371)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g219 ( 
.A(n_75),
.Y(n_219)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx5_ASAP7_75t_L g221 ( 
.A(n_78),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_79),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_79),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_80),
.B(n_81),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_80),
.A2(n_164),
.B(n_189),
.Y(n_222)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_84),
.Y(n_85)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_86),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_106),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_87),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_98),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_91),
.B1(n_93),
.B2(n_94),
.Y(n_88)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_90),
.Y(n_97)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

INVx5_ASAP7_75t_L g353 ( 
.A(n_91),
.Y(n_353)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_96),
.Y(n_114)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVxp67_ASAP7_75t_SL g98 ( 
.A(n_99),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_99),
.A2(n_132),
.B(n_133),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_99),
.B(n_133),
.Y(n_224)
);

INVx6_ASAP7_75t_SL g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g156 ( 
.A(n_105),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_105),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_106),
.A2(n_132),
.B(n_153),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_106),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_118),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_107),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_111),
.B1(n_113),
.B2(n_115),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx4_ASAP7_75t_L g341 ( 
.A(n_110),
.Y(n_341)
);

AOI32xp33_ASAP7_75t_L g257 ( 
.A1(n_111),
.A2(n_258),
.A3(n_259),
.B1(n_262),
.B2(n_263),
.Y(n_257)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_116),
.Y(n_154)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_119),
.B(n_132),
.Y(n_158)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_120),
.Y(n_253)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_125),
.A2(n_126),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_127),
.A2(n_135),
.B(n_199),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_128),
.A2(n_135),
.B(n_136),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_131),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_131),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_131),
.A2(n_134),
.B1(n_310),
.B2(n_439),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_132),
.B(n_251),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_133),
.A2(n_153),
.B(n_157),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_133),
.B(n_251),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_134),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_136),
.B(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_136),
.B(n_226),
.Y(n_298)
);

A2O1A1O1Ixp25_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_239),
.B(n_433),
.C(n_436),
.D(n_441),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_229),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_141),
.B(n_200),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_141),
.B(n_200),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_172),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_159),
.B2(n_160),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_144),
.B(n_159),
.C(n_172),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_148),
.B2(n_149),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_145),
.A2(n_146),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_146),
.B(n_150),
.C(n_152),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_146),
.B(n_232),
.C(n_237),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_147),
.B(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_158),
.B(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_158),
.B(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_160),
.A2(n_161),
.B(n_171),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_161),
.B(n_171),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_163),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_162),
.Y(n_350)
);

INVxp67_ASAP7_75t_SL g163 ( 
.A(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_164),
.B(n_371),
.Y(n_413)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_170),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_197),
.B(n_198),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_173),
.A2(n_174),
.B1(n_202),
.B2(n_203),
.Y(n_201)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_188),
.Y(n_174)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_175),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_175),
.A2(n_197),
.B1(n_198),
.B2(n_204),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_175),
.A2(n_188),
.B1(n_197),
.B2(n_320),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_175),
.B(n_337),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_175),
.A2(n_197),
.B1(n_337),
.B2(n_416),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_181),
.B(n_183),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_176),
.B(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_176),
.B(n_183),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g292 ( 
.A(n_176),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_176),
.B(n_376),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_179),
.Y(n_176)
);

INVx8_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_178),
.Y(n_187)
);

INVx4_ASAP7_75t_L g378 ( 
.A(n_178),
.Y(n_378)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_183),
.Y(n_214)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_186),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_188),
.Y(n_320)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

AND2x2_ASAP7_75t_SL g293 ( 
.A(n_196),
.B(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_196),
.B(n_351),
.Y(n_380)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_198),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_205),
.C(n_207),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_201),
.A2(n_205),
.B1(n_206),
.B2(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_201),
.Y(n_324)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_207),
.B(n_323),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_223),
.C(n_225),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_208),
.A2(n_209),
.B1(n_317),
.B2(n_318),
.Y(n_316)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_222),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_210),
.B(n_222),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_215),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_211),
.B(n_374),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_214),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_213),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_215),
.B(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_216),
.A2(n_270),
.B(n_275),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_217),
.B(n_285),
.Y(n_284)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_219),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g274 ( 
.A(n_219),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_223),
.B(n_225),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_224),
.B(n_250),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_229),
.A2(n_434),
.B(n_435),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_238),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_230),
.B(n_238),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_237),
.Y(n_230)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_425),
.Y(n_239)
);

NAND3xp33_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_313),
.C(n_327),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_301),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_287),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_243),
.B(n_287),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_255),
.C(n_277),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_244),
.B(n_330),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_247),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_248),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_255),
.A2(n_256),
.B1(n_277),
.B2(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_269),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_257),
.B(n_269),
.Y(n_296)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx8_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

NAND2xp33_ASAP7_75t_SL g263 ( 
.A(n_264),
.B(n_266),
.Y(n_263)
);

INVx5_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_270),
.A2(n_284),
.B(n_292),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx8_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_277),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_280),
.C(n_282),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_278),
.B(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_300),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_280),
.A2(n_281),
.B1(n_282),
.B2(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_282),
.Y(n_335)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g401 ( 
.A(n_283),
.B(n_390),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_284),
.B(n_375),
.Y(n_403)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_295),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_289),
.B(n_290),
.C(n_295),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_293),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_293),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_294),
.B(n_371),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_298),
.C(n_299),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_301),
.A2(n_428),
.B(n_429),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_302),
.B(n_312),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_302),
.B(n_312),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_303),
.B(n_305),
.C(n_306),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_309),
.C(n_310),
.Y(n_321)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_309),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_325),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_314),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_322),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g325 ( 
.A(n_315),
.B(n_326),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_315),
.B(n_326),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_315),
.B(n_322),
.Y(n_432)
);

FAx1_ASAP7_75t_SL g315 ( 
.A(n_316),
.B(n_319),
.CI(n_321),
.CON(n_315),
.SN(n_315)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_325),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_328),
.A2(n_357),
.B(n_424),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g328 ( 
.A(n_329),
.B(n_332),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_329),
.B(n_332),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_336),
.C(n_348),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_333),
.B(n_420),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_336),
.A2(n_348),
.B1(n_349),
.B2(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_336),
.Y(n_421)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_337),
.Y(n_416)
);

INVx4_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx8_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx3_ASAP7_75t_SL g342 ( 
.A(n_343),
.Y(n_342)
);

INVx8_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

BUFx12f_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_351),
.Y(n_349)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_358),
.A2(n_418),
.B(n_423),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_359),
.A2(n_408),
.B(n_417),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_360),
.A2(n_384),
.B(n_407),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_372),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_361),
.B(n_372),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_370),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_362),
.A2(n_363),
.B1(n_370),
.B2(n_387),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_363),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_366),
.Y(n_363)
);

INVx5_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_370),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_379),
.Y(n_372)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_373),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_376),
.B(n_391),
.Y(n_390)
);

INVx3_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_380),
.A2(n_381),
.B1(n_382),
.B2(n_383),
.Y(n_379)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_380),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_381),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_381),
.B(n_382),
.C(n_410),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_385),
.A2(n_393),
.B(n_406),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_386),
.B(n_388),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_386),
.B(n_388),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_394),
.A2(n_402),
.B(n_405),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_401),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_400),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx6_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_403),
.B(n_404),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_403),
.B(n_404),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_411),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_409),
.B(n_411),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_415),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_413),
.B(n_414),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_413),
.B(n_414),
.C(n_415),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_419),
.B(n_422),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_419),
.B(n_422),
.Y(n_423)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g425 ( 
.A1(n_426),
.A2(n_427),
.B(n_430),
.C(n_431),
.D(n_432),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_440),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_437),
.B(n_440),
.Y(n_441)
);

INVx6_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx13_ASAP7_75t_L g445 ( 
.A(n_443),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_446),
.Y(n_444)
);


endmodule