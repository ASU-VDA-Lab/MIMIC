module fake_ariane_1186_n_106 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_17, n_4, n_2, n_18, n_9, n_11, n_26, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_25, n_106);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_26;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;
input n_25;

output n_106;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_90;
wire n_38;
wire n_47;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_34;
wire n_69;
wire n_95;
wire n_92;
wire n_98;
wire n_74;
wire n_33;
wire n_40;
wire n_53;
wire n_66;
wire n_71;
wire n_96;
wire n_49;
wire n_100;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_72;
wire n_105;
wire n_44;
wire n_30;
wire n_82;
wire n_42;
wire n_31;
wire n_57;
wire n_70;
wire n_85;
wire n_48;
wire n_94;
wire n_101;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_93;
wire n_61;
wire n_102;
wire n_43;
wire n_81;
wire n_87;
wire n_29;
wire n_41;
wire n_55;
wire n_28;
wire n_80;
wire n_97;
wire n_88;
wire n_68;
wire n_104;
wire n_78;
wire n_39;
wire n_63;
wire n_59;
wire n_99;
wire n_35;
wire n_54;

BUFx2_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_22),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_2),
.B(n_10),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_13),
.Y(n_44)
);

CKINVDCx5p33_ASAP7_75t_R g45 ( 
.A(n_0),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

CKINVDCx5p33_ASAP7_75t_R g47 ( 
.A(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_28),
.B(n_2),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_49),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_29),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_3),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_39),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_29),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

NAND3xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_3),
.C(n_8),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_32),
.Y(n_64)
);

AND2x4_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_35),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_52),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_50),
.A2(n_44),
.B1(n_37),
.B2(n_47),
.Y(n_67)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_55),
.A2(n_30),
.B(n_36),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_35),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_63),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_34),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_35),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_67),
.A2(n_54),
.B1(n_59),
.B2(n_61),
.Y(n_76)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

AOI21x1_ASAP7_75t_L g79 ( 
.A1(n_69),
.A2(n_58),
.B(n_62),
.Y(n_79)
);

INVx1_ASAP7_75t_SL g80 ( 
.A(n_66),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

AND2x4_ASAP7_75t_L g82 ( 
.A(n_74),
.B(n_56),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

BUFx10_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_73),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_80),
.B(n_65),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_76),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_80),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_82),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_90),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_87),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_92),
.A2(n_67),
.B1(n_87),
.B2(n_84),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_93),
.A2(n_84),
.B1(n_86),
.B2(n_85),
.Y(n_97)
);

AOI221xp5_ASAP7_75t_L g98 ( 
.A1(n_95),
.A2(n_71),
.B1(n_57),
.B2(n_70),
.C(n_94),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_96),
.B(n_97),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_75),
.Y(n_100)
);

AOI221xp5_ASAP7_75t_L g101 ( 
.A1(n_99),
.A2(n_57),
.B1(n_88),
.B2(n_41),
.C(n_34),
.Y(n_101)
);

NOR3xp33_ASAP7_75t_SL g102 ( 
.A(n_101),
.B(n_98),
.C(n_100),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_102),
.Y(n_103)
);

AO21x1_ASAP7_75t_SL g104 ( 
.A1(n_103),
.A2(n_11),
.B(n_12),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_38),
.Y(n_105)
);

AOI221xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_77),
.B1(n_18),
.B2(n_27),
.C(n_17),
.Y(n_106)
);


endmodule