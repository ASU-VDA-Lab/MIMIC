module fake_netlist_5_2558_n_801 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_801);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_801;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_785;
wire n_389;
wire n_549;
wire n_684;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_452;
wire n_397;
wire n_493;
wire n_525;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_173;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_373;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_779;
wire n_576;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_171;
wire n_756;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_752;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_782;
wire n_325;
wire n_449;
wire n_724;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_654;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_442;
wire n_192;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_771;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_183;
wire n_243;
wire n_185;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_670;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_521;
wire n_614;
wire n_663;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_432;
wire n_164;
wire n_395;
wire n_553;
wire n_727;
wire n_311;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_749;
wire n_772;
wire n_691;
wire n_717;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_796;
wire n_573;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_781;
wire n_474;
wire n_765;
wire n_542;
wire n_488;
wire n_463;
wire n_595;
wire n_736;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_745;
wire n_627;
wire n_767;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_176;
wire n_557;
wire n_182;
wire n_354;
wire n_575;
wire n_647;
wire n_480;
wire n_607;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_707;
wire n_710;
wire n_795;
wire n_695;
wire n_180;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_720;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_794;
wire n_768;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_791;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_566;
wire n_426;
wire n_520;
wire n_565;
wire n_409;
wire n_797;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_159;
wire n_334;
wire n_599;
wire n_766;
wire n_541;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_238;
wire n_639;
wire n_799;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_162;
wire n_759;
wire n_222;
wire n_438;
wire n_713;
wire n_324;
wire n_634;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;
wire n_784;

INVx1_ASAP7_75t_L g159 ( 
.A(n_100),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_151),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_155),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_137),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_123),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_35),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_70),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_74),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_60),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_7),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_54),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_12),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_23),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_112),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_107),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_27),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_113),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_32),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_157),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_62),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_84),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_52),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_14),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_64),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_79),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_109),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_135),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_122),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_106),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_99),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_68),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_152),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_101),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_50),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_44),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_8),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_117),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_104),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_120),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_61),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_108),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_37),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_6),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_63),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_66),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_111),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_41),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_69),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_145),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_42),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_49),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_72),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_26),
.Y(n_212)
);

NOR2xp67_ASAP7_75t_L g213 ( 
.A(n_148),
.B(n_127),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_83),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_168),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_174),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_174),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_0),
.Y(n_218)
);

BUFx12f_ASAP7_75t_L g219 ( 
.A(n_182),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_170),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_168),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_195),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_168),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_168),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_174),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_182),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_182),
.B(n_161),
.Y(n_227)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_174),
.Y(n_228)
);

AND2x4_ASAP7_75t_L g229 ( 
.A(n_192),
.B(n_0),
.Y(n_229)
);

AND2x4_ASAP7_75t_L g230 ( 
.A(n_191),
.B(n_1),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_175),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_166),
.B(n_1),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_171),
.B(n_2),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_202),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_159),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_162),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_207),
.B(n_2),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_3),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_175),
.Y(n_239)
);

NOR2xp67_ASAP7_75t_L g240 ( 
.A(n_163),
.B(n_3),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_175),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_165),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_167),
.Y(n_243)
);

INVxp67_ASAP7_75t_SL g244 ( 
.A(n_175),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_169),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_160),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_177),
.Y(n_247)
);

INVx5_ASAP7_75t_L g248 ( 
.A(n_172),
.Y(n_248)
);

AND2x4_ASAP7_75t_L g249 ( 
.A(n_180),
.B(n_181),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_186),
.B(n_4),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_213),
.B(n_4),
.Y(n_251)
);

OAI21x1_ASAP7_75t_L g252 ( 
.A1(n_187),
.A2(n_81),
.B(n_156),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_196),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_198),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_199),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_164),
.A2(n_188),
.B1(n_193),
.B2(n_206),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_200),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_204),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_246),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_215),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_221),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_222),
.Y(n_262)
);

NOR2xp67_ASAP7_75t_L g263 ( 
.A(n_248),
.B(n_214),
.Y(n_263)
);

AO21x2_ASAP7_75t_L g264 ( 
.A1(n_251),
.A2(n_237),
.B(n_233),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_256),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_256),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_248),
.Y(n_267)
);

CKINVDCx6p67_ASAP7_75t_R g268 ( 
.A(n_220),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_220),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_248),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_223),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_R g272 ( 
.A(n_219),
.B(n_205),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_216),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_226),
.Y(n_274)
);

INVx4_ASAP7_75t_L g275 ( 
.A(n_248),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_232),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_227),
.B(n_173),
.Y(n_277)
);

NAND2xp33_ASAP7_75t_R g278 ( 
.A(n_218),
.B(n_229),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_234),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_254),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_227),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_224),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_234),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_216),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_224),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_244),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_R g287 ( 
.A(n_235),
.B(n_176),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_254),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_249),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_216),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_R g291 ( 
.A(n_236),
.B(n_178),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_R g292 ( 
.A(n_242),
.B(n_179),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_249),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_243),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_R g295 ( 
.A(n_247),
.B(n_183),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_245),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_244),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_258),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_217),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_240),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_245),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_217),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_217),
.Y(n_303)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_225),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_245),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_257),
.Y(n_306)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_225),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_284),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_284),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_304),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_304),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_307),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_281),
.B(n_218),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_307),
.Y(n_314)
);

AND2x4_ASAP7_75t_L g315 ( 
.A(n_286),
.B(n_229),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_290),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_302),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_282),
.B(n_230),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_273),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_285),
.B(n_230),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_297),
.B(n_228),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_296),
.B(n_251),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_300),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_264),
.B(n_228),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_294),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_277),
.B(n_233),
.Y(n_326)
);

NAND3xp33_ASAP7_75t_L g327 ( 
.A(n_278),
.B(n_250),
.C(n_237),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_264),
.B(n_228),
.Y(n_328)
);

NOR2xp67_ASAP7_75t_L g329 ( 
.A(n_275),
.B(n_228),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_271),
.B(n_255),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_298),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_289),
.B(n_253),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_274),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_269),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_260),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_300),
.Y(n_336)
);

NOR2xp67_ASAP7_75t_L g337 ( 
.A(n_275),
.B(n_184),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_273),
.Y(n_338)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_273),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_261),
.B(n_255),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_273),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_299),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_301),
.B(n_305),
.Y(n_343)
);

NOR3xp33_ASAP7_75t_L g344 ( 
.A(n_265),
.B(n_250),
.C(n_238),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_293),
.B(n_257),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_299),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_259),
.B(n_257),
.Y(n_347)
);

AO221x1_ASAP7_75t_L g348 ( 
.A1(n_283),
.A2(n_255),
.B1(n_241),
.B2(n_239),
.C(n_231),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g349 ( 
.A1(n_279),
.A2(n_252),
.B(n_210),
.Y(n_349)
);

AOI221xp5_ASAP7_75t_L g350 ( 
.A1(n_266),
.A2(n_209),
.B1(n_189),
.B2(n_190),
.C(n_194),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_306),
.B(n_225),
.Y(n_351)
);

BUFx5_ASAP7_75t_L g352 ( 
.A(n_263),
.Y(n_352)
);

NAND2xp33_ASAP7_75t_L g353 ( 
.A(n_287),
.B(n_185),
.Y(n_353)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_299),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_299),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_267),
.B(n_231),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_270),
.B(n_231),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_303),
.B(n_239),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_279),
.B(n_262),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_276),
.B(n_255),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_280),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_303),
.B(n_239),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_303),
.B(n_241),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_303),
.B(n_197),
.Y(n_364)
);

BUFx6f_ASAP7_75t_SL g365 ( 
.A(n_268),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_288),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g367 ( 
.A(n_272),
.B(n_291),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_292),
.B(n_241),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_295),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_264),
.B(n_201),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_284),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_281),
.B(n_211),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_331),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_333),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_335),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_326),
.B(n_212),
.Y(n_376)
);

INVx2_ASAP7_75t_SL g377 ( 
.A(n_316),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_319),
.Y(n_378)
);

NAND3xp33_ASAP7_75t_SL g379 ( 
.A(n_350),
.B(n_5),
.C(n_6),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_318),
.B(n_5),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_319),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_317),
.Y(n_382)
);

INVx1_ASAP7_75t_SL g383 ( 
.A(n_361),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g384 ( 
.A(n_347),
.B(n_7),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_340),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_360),
.B(n_8),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_344),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_340),
.Y(n_388)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_323),
.B(n_9),
.Y(n_389)
);

NAND2x1p5_ASAP7_75t_L g390 ( 
.A(n_315),
.B(n_15),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_327),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_391)
);

BUFx4f_ASAP7_75t_L g392 ( 
.A(n_325),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_313),
.B(n_13),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_370),
.B(n_16),
.Y(n_394)
);

NAND3xp33_ASAP7_75t_SL g395 ( 
.A(n_361),
.B(n_13),
.C(n_14),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_309),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_372),
.B(n_17),
.Y(n_397)
);

INVx2_ASAP7_75t_SL g398 ( 
.A(n_311),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_312),
.Y(n_399)
);

NOR3xp33_ASAP7_75t_L g400 ( 
.A(n_359),
.B(n_18),
.C(n_19),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_334),
.Y(n_401)
);

OR2x2_ASAP7_75t_L g402 ( 
.A(n_320),
.B(n_20),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_330),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_330),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_315),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_370),
.B(n_324),
.Y(n_406)
);

AND2x4_ASAP7_75t_SL g407 ( 
.A(n_369),
.B(n_366),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_328),
.B(n_21),
.Y(n_408)
);

BUFx3_ASAP7_75t_L g409 ( 
.A(n_351),
.Y(n_409)
);

INVxp67_ASAP7_75t_SL g410 ( 
.A(n_362),
.Y(n_410)
);

AND2x4_ASAP7_75t_L g411 ( 
.A(n_314),
.B(n_22),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_371),
.Y(n_412)
);

INVx1_ASAP7_75t_SL g413 ( 
.A(n_322),
.Y(n_413)
);

AOI22xp33_ASAP7_75t_L g414 ( 
.A1(n_349),
.A2(n_24),
.B1(n_25),
.B2(n_28),
.Y(n_414)
);

HB1xp67_ASAP7_75t_L g415 ( 
.A(n_336),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_332),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_345),
.B(n_29),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_368),
.B(n_30),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_319),
.Y(n_419)
);

O2A1O1Ixp33_ASAP7_75t_L g420 ( 
.A1(n_349),
.A2(n_31),
.B(n_33),
.C(n_34),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_368),
.B(n_36),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_321),
.B(n_38),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_308),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_310),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_362),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_367),
.B(n_39),
.Y(n_426)
);

NOR2x1p5_ASAP7_75t_L g427 ( 
.A(n_356),
.B(n_40),
.Y(n_427)
);

INVx2_ASAP7_75t_SL g428 ( 
.A(n_357),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_363),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_363),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_358),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_338),
.Y(n_432)
);

AOI22xp33_ASAP7_75t_L g433 ( 
.A1(n_348),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_339),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_343),
.A2(n_158),
.B1(n_48),
.B2(n_51),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_364),
.B(n_47),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_365),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_353),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_355),
.B(n_57),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_341),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_342),
.B(n_58),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_346),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_378),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_401),
.Y(n_444)
);

INVx1_ASAP7_75t_SL g445 ( 
.A(n_383),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_406),
.A2(n_329),
.B(n_339),
.Y(n_446)
);

NOR3xp33_ASAP7_75t_L g447 ( 
.A(n_416),
.B(n_337),
.C(n_354),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_407),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_376),
.B(n_354),
.Y(n_449)
);

NOR2x1_ASAP7_75t_L g450 ( 
.A(n_379),
.B(n_365),
.Y(n_450)
);

A2O1A1Ixp33_ASAP7_75t_L g451 ( 
.A1(n_393),
.A2(n_59),
.B(n_65),
.C(n_67),
.Y(n_451)
);

OAI21x1_ASAP7_75t_L g452 ( 
.A1(n_408),
.A2(n_352),
.B(n_73),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_410),
.A2(n_352),
.B(n_75),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_383),
.B(n_415),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_375),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_429),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_401),
.Y(n_457)
);

BUFx4f_ASAP7_75t_L g458 ( 
.A(n_390),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_403),
.B(n_352),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_414),
.A2(n_71),
.B1(n_76),
.B2(n_77),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g461 ( 
.A1(n_394),
.A2(n_352),
.B(n_80),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_430),
.Y(n_462)
);

INVx3_ASAP7_75t_SL g463 ( 
.A(n_389),
.Y(n_463)
);

O2A1O1Ixp33_ASAP7_75t_L g464 ( 
.A1(n_386),
.A2(n_352),
.B(n_82),
.C(n_85),
.Y(n_464)
);

O2A1O1Ixp33_ASAP7_75t_L g465 ( 
.A1(n_391),
.A2(n_78),
.B(n_86),
.C(n_87),
.Y(n_465)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_385),
.A2(n_88),
.B(n_89),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_388),
.A2(n_90),
.B(n_91),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_404),
.A2(n_92),
.B(n_93),
.Y(n_468)
);

A2O1A1Ixp33_ASAP7_75t_SL g469 ( 
.A1(n_397),
.A2(n_94),
.B(n_95),
.C(n_96),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g470 ( 
.A(n_405),
.Y(n_470)
);

O2A1O1Ixp33_ASAP7_75t_L g471 ( 
.A1(n_391),
.A2(n_97),
.B(n_98),
.C(n_102),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_374),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_SL g473 ( 
.A(n_437),
.B(n_103),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_392),
.B(n_105),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_409),
.B(n_110),
.Y(n_475)
);

AO31x2_ASAP7_75t_L g476 ( 
.A1(n_425),
.A2(n_114),
.A3(n_115),
.B(n_116),
.Y(n_476)
);

A2O1A1Ixp33_ASAP7_75t_L g477 ( 
.A1(n_420),
.A2(n_118),
.B(n_119),
.C(n_121),
.Y(n_477)
);

O2A1O1Ixp33_ASAP7_75t_L g478 ( 
.A1(n_384),
.A2(n_124),
.B(n_125),
.C(n_126),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_392),
.B(n_128),
.Y(n_479)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_411),
.Y(n_480)
);

NAND3xp33_ASAP7_75t_SL g481 ( 
.A(n_387),
.B(n_413),
.C(n_380),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_413),
.B(n_129),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_428),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_411),
.Y(n_484)
);

A2O1A1Ixp33_ASAP7_75t_L g485 ( 
.A1(n_402),
.A2(n_130),
.B(n_131),
.C(n_132),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_431),
.A2(n_133),
.B(n_134),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g487 ( 
.A1(n_436),
.A2(n_136),
.B(n_138),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_373),
.Y(n_488)
);

NAND3xp33_ASAP7_75t_L g489 ( 
.A(n_387),
.B(n_140),
.C(n_141),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_390),
.A2(n_142),
.B1(n_143),
.B2(n_144),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_417),
.A2(n_146),
.B(n_147),
.Y(n_491)
);

O2A1O1Ixp5_ASAP7_75t_SL g492 ( 
.A1(n_435),
.A2(n_421),
.B(n_432),
.C(n_440),
.Y(n_492)
);

NOR3xp33_ASAP7_75t_SL g493 ( 
.A(n_395),
.B(n_149),
.C(n_150),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_396),
.Y(n_494)
);

CKINVDCx11_ASAP7_75t_R g495 ( 
.A(n_399),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_418),
.A2(n_153),
.B(n_154),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_378),
.A2(n_381),
.B(n_419),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_426),
.B(n_378),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_381),
.B(n_419),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_382),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_456),
.Y(n_501)
);

OAI21x1_ASAP7_75t_L g502 ( 
.A1(n_452),
.A2(n_441),
.B(n_439),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_448),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_455),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_445),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_492),
.A2(n_423),
.B(n_422),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g507 ( 
.A1(n_459),
.A2(n_381),
.B(n_419),
.Y(n_507)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_454),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_462),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_480),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_472),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_470),
.Y(n_512)
);

OAI21x1_ASAP7_75t_L g513 ( 
.A1(n_453),
.A2(n_434),
.B(n_442),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_480),
.Y(n_514)
);

AO21x2_ASAP7_75t_L g515 ( 
.A1(n_477),
.A2(n_449),
.B(n_446),
.Y(n_515)
);

BUFx2_ASAP7_75t_R g516 ( 
.A(n_444),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_484),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_484),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_488),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_494),
.Y(n_520)
);

BUFx3_ASAP7_75t_L g521 ( 
.A(n_457),
.Y(n_521)
);

BUFx2_ASAP7_75t_L g522 ( 
.A(n_483),
.Y(n_522)
);

BUFx12f_ASAP7_75t_L g523 ( 
.A(n_495),
.Y(n_523)
);

AO21x2_ASAP7_75t_L g524 ( 
.A1(n_469),
.A2(n_400),
.B(n_438),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_500),
.Y(n_525)
);

INVxp67_ASAP7_75t_SL g526 ( 
.A(n_443),
.Y(n_526)
);

AND2x2_ASAP7_75t_L g527 ( 
.A(n_482),
.B(n_427),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_498),
.B(n_377),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_463),
.Y(n_529)
);

AND2x4_ASAP7_75t_L g530 ( 
.A(n_450),
.B(n_424),
.Y(n_530)
);

INVx4_ASAP7_75t_L g531 ( 
.A(n_443),
.Y(n_531)
);

INVx5_ASAP7_75t_L g532 ( 
.A(n_443),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_476),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_499),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_475),
.Y(n_535)
);

BUFx12f_ASAP7_75t_L g536 ( 
.A(n_473),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_481),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_458),
.Y(n_538)
);

INVx3_ASAP7_75t_SL g539 ( 
.A(n_474),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_493),
.Y(n_540)
);

BUFx12f_ASAP7_75t_L g541 ( 
.A(n_458),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_489),
.Y(n_542)
);

BUFx2_ASAP7_75t_R g543 ( 
.A(n_479),
.Y(n_543)
);

INVx2_ASAP7_75t_SL g544 ( 
.A(n_476),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_490),
.Y(n_545)
);

CKINVDCx6p67_ASAP7_75t_R g546 ( 
.A(n_465),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_447),
.B(n_476),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_466),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_537),
.B(n_508),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_504),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_520),
.Y(n_551)
);

OAI21xp5_ASAP7_75t_L g552 ( 
.A1(n_542),
.A2(n_460),
.B(n_464),
.Y(n_552)
);

INVx2_ASAP7_75t_SL g553 ( 
.A(n_505),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_511),
.Y(n_554)
);

OAI22xp33_ASAP7_75t_L g555 ( 
.A1(n_536),
.A2(n_435),
.B1(n_438),
.B2(n_412),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_520),
.Y(n_556)
);

AO21x1_ASAP7_75t_L g557 ( 
.A1(n_547),
.A2(n_471),
.B(n_478),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_532),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_510),
.Y(n_559)
);

INVxp33_ASAP7_75t_L g560 ( 
.A(n_522),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_509),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_519),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_527),
.B(n_398),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_510),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_532),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_525),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_525),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_545),
.A2(n_468),
.B1(n_467),
.B2(n_486),
.Y(n_568)
);

BUFx2_ASAP7_75t_L g569 ( 
.A(n_521),
.Y(n_569)
);

AND2x4_ASAP7_75t_L g570 ( 
.A(n_538),
.B(n_485),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_518),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_501),
.Y(n_572)
);

BUFx2_ASAP7_75t_L g573 ( 
.A(n_521),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_534),
.Y(n_574)
);

AOI21x1_ASAP7_75t_L g575 ( 
.A1(n_533),
.A2(n_461),
.B(n_497),
.Y(n_575)
);

INVx4_ASAP7_75t_L g576 ( 
.A(n_532),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_538),
.B(n_451),
.Y(n_577)
);

CKINVDCx6p67_ASAP7_75t_R g578 ( 
.A(n_536),
.Y(n_578)
);

AOI21xp5_ASAP7_75t_L g579 ( 
.A1(n_548),
.A2(n_535),
.B(n_515),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_527),
.B(n_433),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_512),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_528),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_540),
.A2(n_530),
.B1(n_522),
.B2(n_539),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_518),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_531),
.Y(n_585)
);

HB1xp67_ASAP7_75t_L g586 ( 
.A(n_532),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_517),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_517),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_530),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_L g590 ( 
.A1(n_545),
.A2(n_487),
.B1(n_491),
.B2(n_496),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_530),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_514),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_582),
.B(n_546),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_R g594 ( 
.A(n_578),
.B(n_529),
.Y(n_594)
);

CKINVDCx16_ASAP7_75t_R g595 ( 
.A(n_569),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_550),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_573),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_580),
.B(n_546),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_563),
.B(n_540),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_578),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_574),
.B(n_545),
.Y(n_601)
);

OR2x6_ASAP7_75t_L g602 ( 
.A(n_570),
.B(n_545),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_560),
.B(n_516),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_560),
.B(n_529),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_566),
.B(n_545),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_R g606 ( 
.A(n_553),
.B(n_541),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_567),
.B(n_547),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_551),
.B(n_539),
.Y(n_608)
);

INVx8_ASAP7_75t_L g609 ( 
.A(n_558),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_583),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_549),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_554),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_551),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_589),
.B(n_503),
.Y(n_614)
);

HB1xp67_ASAP7_75t_L g615 ( 
.A(n_581),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_591),
.B(n_503),
.Y(n_616)
);

HB1xp67_ASAP7_75t_L g617 ( 
.A(n_561),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_556),
.Y(n_618)
);

AND2x4_ASAP7_75t_L g619 ( 
.A(n_570),
.B(n_531),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g620 ( 
.A(n_570),
.B(n_531),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_562),
.Y(n_621)
);

BUFx2_ASAP7_75t_L g622 ( 
.A(n_577),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_SL g623 ( 
.A1(n_552),
.A2(n_523),
.B1(n_541),
.B2(n_524),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_558),
.Y(n_624)
);

AO31x2_ASAP7_75t_L g625 ( 
.A1(n_557),
.A2(n_533),
.A3(n_507),
.B(n_544),
.Y(n_625)
);

NOR3xp33_ASAP7_75t_SL g626 ( 
.A(n_555),
.B(n_506),
.C(n_526),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_572),
.B(n_514),
.Y(n_627)
);

OR2x2_ASAP7_75t_L g628 ( 
.A(n_556),
.B(n_514),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_558),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_584),
.Y(n_630)
);

INVx3_ASAP7_75t_L g631 ( 
.A(n_558),
.Y(n_631)
);

INVx8_ASAP7_75t_L g632 ( 
.A(n_565),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_555),
.B(n_577),
.Y(n_633)
);

CKINVDCx11_ASAP7_75t_R g634 ( 
.A(n_565),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_565),
.Y(n_635)
);

HB1xp67_ASAP7_75t_L g636 ( 
.A(n_559),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_565),
.Y(n_637)
);

OA21x2_ASAP7_75t_L g638 ( 
.A1(n_579),
.A2(n_544),
.B(n_502),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_559),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_564),
.B(n_543),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_R g641 ( 
.A(n_585),
.B(n_523),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_564),
.Y(n_642)
);

NAND3xp33_ASAP7_75t_SL g643 ( 
.A(n_568),
.B(n_524),
.C(n_515),
.Y(n_643)
);

NOR3xp33_ASAP7_75t_SL g644 ( 
.A(n_587),
.B(n_524),
.C(n_532),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_588),
.Y(n_645)
);

AND3x2_ASAP7_75t_L g646 ( 
.A(n_577),
.B(n_515),
.C(n_513),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_571),
.B(n_513),
.Y(n_647)
);

OAI211xp5_ASAP7_75t_L g648 ( 
.A1(n_623),
.A2(n_568),
.B(n_590),
.C(n_548),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_617),
.Y(n_649)
);

AO21x2_ASAP7_75t_L g650 ( 
.A1(n_643),
.A2(n_575),
.B(n_502),
.Y(n_650)
);

NAND2xp33_ASAP7_75t_L g651 ( 
.A(n_611),
.B(n_590),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_640),
.B(n_571),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_639),
.Y(n_653)
);

AOI31xp33_ASAP7_75t_L g654 ( 
.A1(n_623),
.A2(n_592),
.A3(n_586),
.B(n_576),
.Y(n_654)
);

BUFx2_ASAP7_75t_SL g655 ( 
.A(n_597),
.Y(n_655)
);

INVx8_ASAP7_75t_L g656 ( 
.A(n_609),
.Y(n_656)
);

OAI221xp5_ASAP7_75t_L g657 ( 
.A1(n_593),
.A2(n_548),
.B1(n_592),
.B2(n_585),
.C(n_586),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_642),
.Y(n_658)
);

BUFx2_ASAP7_75t_L g659 ( 
.A(n_595),
.Y(n_659)
);

HB1xp67_ASAP7_75t_L g660 ( 
.A(n_647),
.Y(n_660)
);

BUFx5_ASAP7_75t_L g661 ( 
.A(n_630),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_613),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_645),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_598),
.A2(n_576),
.B1(n_602),
.B2(n_622),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_607),
.B(n_633),
.Y(n_665)
);

OR2x2_ASAP7_75t_L g666 ( 
.A(n_598),
.B(n_633),
.Y(n_666)
);

OAI221xp5_ASAP7_75t_L g667 ( 
.A1(n_593),
.A2(n_626),
.B1(n_610),
.B2(n_608),
.C(n_601),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_596),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_607),
.B(n_601),
.Y(n_669)
);

HB1xp67_ASAP7_75t_L g670 ( 
.A(n_615),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_612),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_621),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_614),
.B(n_616),
.Y(n_673)
);

HB1xp67_ASAP7_75t_L g674 ( 
.A(n_625),
.Y(n_674)
);

INVx4_ASAP7_75t_L g675 ( 
.A(n_609),
.Y(n_675)
);

AND2x4_ASAP7_75t_L g676 ( 
.A(n_619),
.B(n_620),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_636),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_609),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_618),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_599),
.B(n_627),
.Y(n_680)
);

HB1xp67_ASAP7_75t_L g681 ( 
.A(n_608),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_605),
.B(n_602),
.Y(n_682)
);

HB1xp67_ASAP7_75t_L g683 ( 
.A(n_605),
.Y(n_683)
);

OR2x2_ASAP7_75t_L g684 ( 
.A(n_602),
.B(n_604),
.Y(n_684)
);

AOI22xp5_ASAP7_75t_L g685 ( 
.A1(n_619),
.A2(n_620),
.B1(n_603),
.B2(n_600),
.Y(n_685)
);

INVx5_ASAP7_75t_L g686 ( 
.A(n_632),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_628),
.B(n_631),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_624),
.B(n_631),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_651),
.A2(n_643),
.B1(n_641),
.B2(n_606),
.Y(n_689)
);

AND2x4_ASAP7_75t_SL g690 ( 
.A(n_676),
.B(n_644),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_663),
.Y(n_691)
);

AOI22xp33_ASAP7_75t_SL g692 ( 
.A1(n_648),
.A2(n_594),
.B1(n_644),
.B2(n_637),
.Y(n_692)
);

INVxp67_ASAP7_75t_L g693 ( 
.A(n_670),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_661),
.Y(n_694)
);

INVx3_ASAP7_75t_SL g695 ( 
.A(n_656),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_673),
.B(n_624),
.Y(n_696)
);

AND2x4_ASAP7_75t_L g697 ( 
.A(n_660),
.B(n_646),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_649),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_681),
.B(n_629),
.Y(n_699)
);

OR2x2_ASAP7_75t_L g700 ( 
.A(n_666),
.B(n_625),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_680),
.B(n_625),
.Y(n_701)
);

OR2x2_ASAP7_75t_L g702 ( 
.A(n_660),
.B(n_638),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_665),
.B(n_635),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_665),
.B(n_682),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_668),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_661),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_671),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_683),
.B(n_634),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_684),
.B(n_638),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_672),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_669),
.B(n_677),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_682),
.Y(n_712)
);

NAND2x1p5_ASAP7_75t_L g713 ( 
.A(n_686),
.B(n_632),
.Y(n_713)
);

OR2x2_ASAP7_75t_L g714 ( 
.A(n_669),
.B(n_632),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_687),
.B(n_652),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_676),
.B(n_659),
.Y(n_716)
);

AND2x4_ASAP7_75t_L g717 ( 
.A(n_688),
.B(n_679),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_661),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_653),
.B(n_662),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_704),
.B(n_674),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_691),
.Y(n_721)
);

AND2x4_ASAP7_75t_L g722 ( 
.A(n_697),
.B(n_674),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_704),
.B(n_709),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_712),
.B(n_667),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_701),
.B(n_650),
.Y(n_725)
);

OR2x2_ASAP7_75t_L g726 ( 
.A(n_702),
.B(n_650),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_705),
.Y(n_727)
);

HB1xp67_ASAP7_75t_L g728 ( 
.A(n_693),
.Y(n_728)
);

INVx3_ASAP7_75t_L g729 ( 
.A(n_717),
.Y(n_729)
);

INVxp33_ASAP7_75t_SL g730 ( 
.A(n_715),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_707),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_710),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_700),
.B(n_664),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_698),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_697),
.B(n_648),
.Y(n_735)
);

BUFx2_ASAP7_75t_L g736 ( 
.A(n_697),
.Y(n_736)
);

INVx3_ASAP7_75t_L g737 ( 
.A(n_717),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_717),
.B(n_685),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_693),
.B(n_654),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_694),
.B(n_658),
.Y(n_740)
);

BUFx3_ASAP7_75t_L g741 ( 
.A(n_695),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_721),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_721),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_731),
.Y(n_744)
);

NOR2x1p5_ASAP7_75t_SL g745 ( 
.A(n_726),
.B(n_694),
.Y(n_745)
);

AND2x4_ASAP7_75t_L g746 ( 
.A(n_736),
.B(n_690),
.Y(n_746)
);

INVx1_ASAP7_75t_SL g747 ( 
.A(n_739),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_731),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_727),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_727),
.Y(n_750)
);

A2O1A1Ixp33_ASAP7_75t_L g751 ( 
.A1(n_724),
.A2(n_689),
.B(n_667),
.C(n_692),
.Y(n_751)
);

NAND4xp75_ASAP7_75t_L g752 ( 
.A(n_735),
.B(n_703),
.C(n_699),
.D(n_708),
.Y(n_752)
);

NOR3xp33_ASAP7_75t_L g753 ( 
.A(n_751),
.B(n_692),
.C(n_739),
.Y(n_753)
);

AOI211xp5_ASAP7_75t_L g754 ( 
.A1(n_747),
.A2(n_735),
.B(n_728),
.C(n_738),
.Y(n_754)
);

AOI21xp33_ASAP7_75t_L g755 ( 
.A1(n_747),
.A2(n_726),
.B(n_733),
.Y(n_755)
);

NOR3xp33_ASAP7_75t_L g756 ( 
.A(n_752),
.B(n_657),
.C(n_733),
.Y(n_756)
);

XNOR2xp5_ASAP7_75t_L g757 ( 
.A(n_746),
.B(n_716),
.Y(n_757)
);

AOI21xp33_ASAP7_75t_L g758 ( 
.A1(n_746),
.A2(n_689),
.B(n_711),
.Y(n_758)
);

INVxp67_ASAP7_75t_L g759 ( 
.A(n_742),
.Y(n_759)
);

OAI322xp33_ASAP7_75t_L g760 ( 
.A1(n_759),
.A2(n_743),
.A3(n_744),
.B1(n_748),
.B2(n_734),
.C1(n_749),
.C2(n_732),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_756),
.B(n_730),
.Y(n_761)
);

AOI22xp5_ASAP7_75t_L g762 ( 
.A1(n_753),
.A2(n_738),
.B1(n_736),
.B2(n_690),
.Y(n_762)
);

OR2x2_ASAP7_75t_L g763 ( 
.A(n_755),
.B(n_723),
.Y(n_763)
);

AOI221xp5_ASAP7_75t_L g764 ( 
.A1(n_754),
.A2(n_730),
.B1(n_725),
.B2(n_732),
.C(n_750),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_758),
.B(n_723),
.Y(n_765)
);

OR2x2_ASAP7_75t_L g766 ( 
.A(n_765),
.B(n_729),
.Y(n_766)
);

NAND3xp33_ASAP7_75t_SL g767 ( 
.A(n_764),
.B(n_714),
.C(n_725),
.Y(n_767)
);

OA22x2_ASAP7_75t_L g768 ( 
.A1(n_762),
.A2(n_757),
.B1(n_737),
.B2(n_729),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_761),
.B(n_741),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_769),
.B(n_763),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_766),
.Y(n_771)
);

OAI211xp5_ASAP7_75t_L g772 ( 
.A1(n_770),
.A2(n_767),
.B(n_768),
.C(n_741),
.Y(n_772)
);

OAI221xp5_ASAP7_75t_L g773 ( 
.A1(n_771),
.A2(n_655),
.B1(n_695),
.B2(n_729),
.C(n_737),
.Y(n_773)
);

NOR4xp25_ASAP7_75t_SL g774 ( 
.A(n_771),
.B(n_760),
.C(n_657),
.D(n_745),
.Y(n_774)
);

AOI22xp5_ASAP7_75t_L g775 ( 
.A1(n_772),
.A2(n_722),
.B1(n_737),
.B2(n_696),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_773),
.Y(n_776)
);

NOR2x1_ASAP7_75t_L g777 ( 
.A(n_774),
.B(n_675),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_773),
.Y(n_778)
);

NOR2x1_ASAP7_75t_L g779 ( 
.A(n_772),
.B(n_675),
.Y(n_779)
);

INVx2_ASAP7_75t_SL g780 ( 
.A(n_777),
.Y(n_780)
);

INVxp67_ASAP7_75t_L g781 ( 
.A(n_779),
.Y(n_781)
);

NOR4xp25_ASAP7_75t_L g782 ( 
.A(n_776),
.B(n_718),
.C(n_719),
.D(n_740),
.Y(n_782)
);

NAND4xp75_ASAP7_75t_L g783 ( 
.A(n_778),
.B(n_740),
.C(n_720),
.D(n_706),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_775),
.Y(n_784)
);

INVx2_ASAP7_75t_SL g785 ( 
.A(n_780),
.Y(n_785)
);

CKINVDCx16_ASAP7_75t_R g786 ( 
.A(n_784),
.Y(n_786)
);

INVx5_ASAP7_75t_L g787 ( 
.A(n_781),
.Y(n_787)
);

CKINVDCx20_ASAP7_75t_R g788 ( 
.A(n_783),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_785),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_787),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_786),
.Y(n_791)
);

OAI22xp5_ASAP7_75t_L g792 ( 
.A1(n_791),
.A2(n_788),
.B1(n_790),
.B2(n_789),
.Y(n_792)
);

BUFx2_ASAP7_75t_L g793 ( 
.A(n_791),
.Y(n_793)
);

BUFx2_ASAP7_75t_SL g794 ( 
.A(n_791),
.Y(n_794)
);

OAI22x1_ASAP7_75t_L g795 ( 
.A1(n_793),
.A2(n_782),
.B1(n_686),
.B2(n_713),
.Y(n_795)
);

CKINVDCx20_ASAP7_75t_R g796 ( 
.A(n_792),
.Y(n_796)
);

OAI22xp5_ASAP7_75t_SL g797 ( 
.A1(n_796),
.A2(n_794),
.B1(n_686),
.B2(n_713),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_797),
.B(n_795),
.Y(n_798)
);

AOI22xp5_ASAP7_75t_L g799 ( 
.A1(n_798),
.A2(n_656),
.B1(n_678),
.B2(n_722),
.Y(n_799)
);

OR2x6_ASAP7_75t_L g800 ( 
.A(n_799),
.B(n_656),
.Y(n_800)
);

AOI211xp5_ASAP7_75t_L g801 ( 
.A1(n_800),
.A2(n_678),
.B(n_722),
.C(n_720),
.Y(n_801)
);


endmodule