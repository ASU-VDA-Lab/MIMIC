module fake_aes_12424_n_742 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_742);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_742;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_199;
wire n_351;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_735;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_106;
wire n_553;
wire n_440;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_39), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_69), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_5), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_99), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_49), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_13), .Y(n_111) );
BUFx6f_ASAP7_75t_L g112 ( .A(n_3), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_96), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_86), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_25), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_32), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_12), .Y(n_117) );
INVxp67_ASAP7_75t_SL g118 ( .A(n_11), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_82), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_97), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_13), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_31), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_76), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_8), .Y(n_124) );
BUFx8_ASAP7_75t_SL g125 ( .A(n_98), .Y(n_125) );
BUFx3_ASAP7_75t_L g126 ( .A(n_0), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_41), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_65), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_89), .Y(n_129) );
BUFx2_ASAP7_75t_L g130 ( .A(n_79), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_58), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_37), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_102), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_38), .Y(n_134) );
INVxp67_ASAP7_75t_L g135 ( .A(n_10), .Y(n_135) );
INVx2_ASAP7_75t_SL g136 ( .A(n_83), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_77), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_62), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_19), .Y(n_139) );
BUFx2_ASAP7_75t_L g140 ( .A(n_57), .Y(n_140) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_66), .Y(n_141) );
BUFx8_ASAP7_75t_SL g142 ( .A(n_9), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_105), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g144 ( .A(n_71), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g145 ( .A(n_34), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_68), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_23), .Y(n_147) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_43), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_101), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g150 ( .A(n_29), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g151 ( .A(n_125), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_130), .B(n_0), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_126), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g154 ( .A(n_130), .B(n_1), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_140), .B(n_1), .Y(n_155) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_147), .Y(n_156) );
OAI22xp5_ASAP7_75t_SL g157 ( .A1(n_108), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_140), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_126), .Y(n_159) );
OAI22xp5_ASAP7_75t_SL g160 ( .A1(n_108), .A2(n_2), .B1(n_4), .B2(n_5), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_109), .Y(n_161) );
AND2x6_ASAP7_75t_L g162 ( .A(n_107), .B(n_24), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_110), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_107), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_147), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_111), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_115), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_115), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_128), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_121), .Y(n_170) );
AOI22xp33_ASAP7_75t_L g171 ( .A1(n_158), .A2(n_154), .B1(n_161), .B2(n_163), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_161), .B(n_136), .Y(n_172) );
BUFx2_ASAP7_75t_L g173 ( .A(n_152), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_163), .B(n_136), .Y(n_174) );
OR2x6_ASAP7_75t_L g175 ( .A(n_157), .B(n_139), .Y(n_175) );
AND2x2_ASAP7_75t_SL g176 ( .A(n_155), .B(n_128), .Y(n_176) );
AOI22xp33_ASAP7_75t_L g177 ( .A1(n_166), .A2(n_135), .B1(n_112), .B2(n_124), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_170), .B(n_106), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_164), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_156), .Y(n_180) );
INVx3_ASAP7_75t_L g181 ( .A(n_164), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_167), .Y(n_182) );
AND2x4_ASAP7_75t_L g183 ( .A(n_159), .B(n_112), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_156), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_167), .Y(n_185) );
AO22x2_ASAP7_75t_L g186 ( .A1(n_168), .A2(n_118), .B1(n_114), .B2(n_116), .Y(n_186) );
INVx3_ASAP7_75t_L g187 ( .A(n_168), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_169), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_153), .B(n_113), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_156), .Y(n_190) );
OAI22xp33_ASAP7_75t_L g191 ( .A1(n_151), .A2(n_117), .B1(n_124), .B2(n_112), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_153), .B(n_119), .Y(n_192) );
AND2x4_ASAP7_75t_L g193 ( .A(n_169), .B(n_112), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_156), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_156), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_162), .B(n_122), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_151), .B(n_117), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_165), .B(n_127), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_165), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_173), .B(n_106), .Y(n_200) );
HB1xp67_ASAP7_75t_L g201 ( .A(n_173), .Y(n_201) );
INVx8_ASAP7_75t_L g202 ( .A(n_183), .Y(n_202) );
HB1xp67_ASAP7_75t_L g203 ( .A(n_197), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_176), .B(n_120), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_179), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_176), .B(n_120), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_176), .B(n_123), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_179), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_174), .B(n_123), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_171), .B(n_134), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_174), .B(n_134), .Y(n_211) );
AOI22xp5_ASAP7_75t_L g212 ( .A1(n_186), .A2(n_160), .B1(n_144), .B2(n_145), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_172), .B(n_137), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_181), .Y(n_214) );
NOR2xp67_ASAP7_75t_L g215 ( .A(n_196), .B(n_26), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_178), .B(n_137), .Y(n_216) );
AOI22xp33_ASAP7_75t_L g217 ( .A1(n_186), .A2(n_162), .B1(n_112), .B2(n_131), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_182), .Y(n_218) );
AOI22xp33_ASAP7_75t_L g219 ( .A1(n_186), .A2(n_162), .B1(n_129), .B2(n_132), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_182), .Y(n_220) );
OAI21xp5_ASAP7_75t_L g221 ( .A1(n_196), .A2(n_162), .B(n_133), .Y(n_221) );
AND2x2_ASAP7_75t_L g222 ( .A(n_186), .B(n_141), .Y(n_222) );
OAI22xp5_ASAP7_75t_L g223 ( .A1(n_186), .A2(n_150), .B1(n_141), .B2(n_149), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_197), .B(n_143), .Y(n_224) );
AOI21x1_ASAP7_75t_L g225 ( .A1(n_194), .A2(n_138), .B(n_146), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_181), .Y(n_226) );
BUFx3_ASAP7_75t_L g227 ( .A(n_183), .Y(n_227) );
AOI22xp5_ASAP7_75t_L g228 ( .A1(n_175), .A2(n_149), .B1(n_143), .B2(n_162), .Y(n_228) );
AND2x2_ASAP7_75t_L g229 ( .A(n_185), .B(n_162), .Y(n_229) );
AND2x4_ASAP7_75t_L g230 ( .A(n_183), .B(n_6), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_191), .B(n_142), .Y(n_231) );
AOI22xp33_ASAP7_75t_SL g232 ( .A1(n_175), .A2(n_148), .B1(n_147), .B2(n_165), .Y(n_232) );
AOI22xp5_ASAP7_75t_L g233 ( .A1(n_177), .A2(n_148), .B1(n_147), .B2(n_165), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_192), .B(n_147), .Y(n_234) );
INVx3_ASAP7_75t_L g235 ( .A(n_183), .Y(n_235) );
AND2x2_ASAP7_75t_L g236 ( .A(n_185), .B(n_6), .Y(n_236) );
AOI22xp5_ASAP7_75t_L g237 ( .A1(n_175), .A2(n_148), .B1(n_165), .B2(n_9), .Y(n_237) );
AOI22xp5_ASAP7_75t_L g238 ( .A1(n_175), .A2(n_148), .B1(n_8), .B2(n_10), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_209), .B(n_189), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_221), .A2(n_192), .B(n_198), .Y(n_240) );
NOR2xp33_ASAP7_75t_SL g241 ( .A(n_223), .B(n_175), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_236), .Y(n_242) );
CKINVDCx14_ASAP7_75t_R g243 ( .A(n_222), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_219), .B(n_191), .Y(n_244) );
O2A1O1Ixp33_ASAP7_75t_L g245 ( .A1(n_203), .A2(n_188), .B(n_181), .C(n_187), .Y(n_245) );
AOI22x1_ASAP7_75t_L g246 ( .A1(n_229), .A2(n_188), .B1(n_187), .B2(n_181), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_205), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_211), .A2(n_193), .B(n_194), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_217), .B(n_187), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_201), .B(n_187), .Y(n_250) );
OAI21xp5_ASAP7_75t_L g251 ( .A1(n_229), .A2(n_193), .B(n_199), .Y(n_251) );
NAND2x1_ASAP7_75t_L g252 ( .A(n_205), .B(n_193), .Y(n_252) );
OAI22xp5_ASAP7_75t_L g253 ( .A1(n_238), .A2(n_193), .B1(n_148), .B2(n_199), .Y(n_253) );
A2O1A1Ixp33_ASAP7_75t_L g254 ( .A1(n_238), .A2(n_195), .B(n_190), .C(n_184), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_200), .B(n_224), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_222), .B(n_7), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_208), .A2(n_195), .B(n_190), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_236), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_230), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_204), .B(n_7), .Y(n_260) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_228), .B(n_180), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_206), .B(n_11), .Y(n_262) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_228), .B(n_180), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_207), .B(n_12), .Y(n_264) );
NAND3xp33_ASAP7_75t_L g265 ( .A(n_231), .B(n_190), .C(n_184), .Y(n_265) );
INVx3_ASAP7_75t_SL g266 ( .A(n_202), .Y(n_266) );
OAI21xp33_ASAP7_75t_SL g267 ( .A1(n_208), .A2(n_218), .B(n_220), .Y(n_267) );
BUFx6f_ASAP7_75t_L g268 ( .A(n_230), .Y(n_268) );
OAI22xp5_ASAP7_75t_L g269 ( .A1(n_237), .A2(n_195), .B1(n_184), .B2(n_180), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_218), .B(n_14), .Y(n_270) );
AOI21x1_ASAP7_75t_L g271 ( .A1(n_225), .A2(n_55), .B(n_103), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_230), .Y(n_272) );
AO31x2_ASAP7_75t_L g273 ( .A1(n_254), .A2(n_234), .A3(n_220), .B(n_214), .Y(n_273) );
AOI22xp5_ASAP7_75t_L g274 ( .A1(n_241), .A2(n_212), .B1(n_210), .B2(n_237), .Y(n_274) );
AND2x6_ASAP7_75t_L g275 ( .A(n_268), .B(n_235), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_247), .Y(n_276) );
AOI21xp5_ASAP7_75t_L g277 ( .A1(n_240), .A2(n_213), .B(n_216), .Y(n_277) );
A2O1A1Ixp33_ASAP7_75t_L g278 ( .A1(n_267), .A2(n_212), .B(n_232), .C(n_235), .Y(n_278) );
BUFx6f_ASAP7_75t_L g279 ( .A(n_266), .Y(n_279) );
OAI21x1_ASAP7_75t_L g280 ( .A1(n_246), .A2(n_225), .B(n_214), .Y(n_280) );
OAI22xp5_ASAP7_75t_L g281 ( .A1(n_268), .A2(n_227), .B1(n_235), .B2(n_202), .Y(n_281) );
NOR2xp33_ASAP7_75t_L g282 ( .A(n_255), .B(n_202), .Y(n_282) );
OAI21xp5_ASAP7_75t_L g283 ( .A1(n_261), .A2(n_226), .B(n_215), .Y(n_283) );
OAI21x1_ASAP7_75t_L g284 ( .A1(n_271), .A2(n_226), .B(n_215), .Y(n_284) );
OAI21xp5_ASAP7_75t_L g285 ( .A1(n_261), .A2(n_233), .B(n_227), .Y(n_285) );
A2O1A1Ixp33_ASAP7_75t_L g286 ( .A1(n_247), .A2(n_202), .B(n_15), .C(n_16), .Y(n_286) );
OAI21xp33_ASAP7_75t_L g287 ( .A1(n_239), .A2(n_14), .B(n_15), .Y(n_287) );
OA21x2_ASAP7_75t_L g288 ( .A1(n_254), .A2(n_56), .B(n_100), .Y(n_288) );
AOI21xp5_ASAP7_75t_L g289 ( .A1(n_263), .A2(n_54), .B(n_95), .Y(n_289) );
O2A1O1Ixp33_ASAP7_75t_SL g290 ( .A1(n_263), .A2(n_53), .B(n_94), .C(n_93), .Y(n_290) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_248), .A2(n_52), .B(n_92), .Y(n_291) );
NAND3xp33_ASAP7_75t_SL g292 ( .A(n_256), .B(n_264), .C(n_260), .Y(n_292) );
INVx2_ASAP7_75t_SL g293 ( .A(n_266), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_250), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_270), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_243), .B(n_16), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_242), .Y(n_297) );
OAI21x1_ASAP7_75t_L g298 ( .A1(n_284), .A2(n_249), .B(n_257), .Y(n_298) );
A2O1A1Ixp33_ASAP7_75t_L g299 ( .A1(n_278), .A2(n_258), .B(n_244), .C(n_245), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_276), .Y(n_300) );
NAND2x1_ASAP7_75t_L g301 ( .A(n_288), .B(n_268), .Y(n_301) );
AND2x4_ASAP7_75t_L g302 ( .A(n_279), .B(n_268), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_294), .B(n_272), .Y(n_303) );
AO21x2_ASAP7_75t_L g304 ( .A1(n_292), .A2(n_249), .B(n_244), .Y(n_304) );
AOI22xp33_ASAP7_75t_L g305 ( .A1(n_295), .A2(n_243), .B1(n_259), .B2(n_262), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_297), .B(n_251), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_273), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_286), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_286), .Y(n_309) );
AO21x2_ASAP7_75t_L g310 ( .A1(n_278), .A2(n_253), .B(n_265), .Y(n_310) );
OR2x2_ASAP7_75t_L g311 ( .A(n_274), .B(n_252), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_273), .Y(n_312) );
OAI21xp5_ASAP7_75t_L g313 ( .A1(n_277), .A2(n_269), .B(n_18), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g314 ( .A1(n_283), .A2(n_51), .B(n_91), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_273), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_282), .B(n_17), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_282), .B(n_17), .Y(n_317) );
OAI21x1_ASAP7_75t_L g318 ( .A1(n_280), .A2(n_59), .B(n_90), .Y(n_318) );
AND2x4_ASAP7_75t_L g319 ( .A(n_279), .B(n_50), .Y(n_319) );
INVx3_ASAP7_75t_L g320 ( .A(n_302), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_300), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_300), .Y(n_322) );
OA21x2_ASAP7_75t_L g323 ( .A1(n_313), .A2(n_287), .B(n_289), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_307), .Y(n_324) );
OA21x2_ASAP7_75t_L g325 ( .A1(n_313), .A2(n_285), .B(n_291), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_307), .Y(n_326) );
OAI21x1_ASAP7_75t_SL g327 ( .A1(n_314), .A2(n_288), .B(n_293), .Y(n_327) );
BUFx2_ASAP7_75t_L g328 ( .A(n_307), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_308), .B(n_273), .Y(n_329) );
BUFx2_ASAP7_75t_L g330 ( .A(n_307), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_312), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_312), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_312), .Y(n_333) );
INVx2_ASAP7_75t_SL g334 ( .A(n_302), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_312), .Y(n_335) );
INVx3_ASAP7_75t_L g336 ( .A(n_302), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_308), .B(n_288), .Y(n_337) );
AOI22xp33_ASAP7_75t_L g338 ( .A1(n_309), .A2(n_296), .B1(n_279), .B2(n_275), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_315), .Y(n_339) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_315), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_315), .Y(n_341) );
OR2x2_ASAP7_75t_L g342 ( .A(n_309), .B(n_279), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_315), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_303), .Y(n_344) );
INVx2_ASAP7_75t_SL g345 ( .A(n_302), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_317), .B(n_275), .Y(n_346) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_317), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_303), .Y(n_348) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_323), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_329), .B(n_304), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_326), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_324), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_324), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_329), .B(n_304), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_344), .B(n_304), .Y(n_355) );
AOI22xp5_ASAP7_75t_L g356 ( .A1(n_347), .A2(n_317), .B1(n_316), .B2(n_305), .Y(n_356) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_340), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_326), .Y(n_358) );
INVx2_ASAP7_75t_SL g359 ( .A(n_328), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_344), .B(n_304), .Y(n_360) );
INVx1_ASAP7_75t_SL g361 ( .A(n_328), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_348), .B(n_304), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_326), .Y(n_363) );
BUFx3_ASAP7_75t_L g364 ( .A(n_328), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_332), .Y(n_365) );
AND2x2_ASAP7_75t_SL g366 ( .A(n_347), .B(n_319), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_348), .B(n_329), .Y(n_367) );
OR2x2_ASAP7_75t_L g368 ( .A(n_340), .B(n_311), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_321), .B(n_299), .Y(n_369) );
INVx2_ASAP7_75t_SL g370 ( .A(n_330), .Y(n_370) );
AND2x4_ASAP7_75t_L g371 ( .A(n_332), .B(n_319), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_321), .B(n_299), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_326), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_322), .B(n_306), .Y(n_374) );
NOR2x1_ASAP7_75t_R g375 ( .A(n_346), .B(n_319), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_322), .B(n_306), .Y(n_376) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_330), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_341), .Y(n_378) );
AO21x2_ASAP7_75t_L g379 ( .A1(n_327), .A2(n_298), .B(n_318), .Y(n_379) );
BUFx2_ASAP7_75t_L g380 ( .A(n_330), .Y(n_380) );
AO21x2_ASAP7_75t_L g381 ( .A1(n_327), .A2(n_298), .B(n_318), .Y(n_381) );
INVx1_ASAP7_75t_SL g382 ( .A(n_342), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_335), .Y(n_383) );
AOI22xp5_ASAP7_75t_L g384 ( .A1(n_346), .A2(n_316), .B1(n_305), .B2(n_303), .Y(n_384) );
NOR2x1_ASAP7_75t_SL g385 ( .A(n_346), .B(n_311), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_341), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_335), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_335), .B(n_311), .Y(n_388) );
INVx3_ASAP7_75t_L g389 ( .A(n_335), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_331), .B(n_310), .Y(n_390) );
NOR2x1_ASAP7_75t_L g391 ( .A(n_342), .B(n_319), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_331), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_331), .B(n_333), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_333), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_333), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_351), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_350), .B(n_343), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_350), .B(n_343), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_352), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_367), .B(n_337), .Y(n_400) );
OR2x2_ASAP7_75t_L g401 ( .A(n_357), .B(n_343), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_352), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_367), .B(n_337), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_351), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_350), .B(n_339), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_354), .B(n_339), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_353), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_354), .B(n_339), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_354), .B(n_337), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_351), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_388), .B(n_320), .Y(n_411) );
AND2x4_ASAP7_75t_L g412 ( .A(n_371), .B(n_320), .Y(n_412) );
OR2x2_ASAP7_75t_L g413 ( .A(n_357), .B(n_368), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_388), .B(n_320), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_355), .B(n_320), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_353), .Y(n_416) );
INVxp67_ASAP7_75t_SL g417 ( .A(n_377), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_365), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_355), .B(n_320), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_365), .Y(n_420) );
INVx3_ASAP7_75t_L g421 ( .A(n_389), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_358), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_360), .B(n_336), .Y(n_423) );
NOR2xp33_ASAP7_75t_L g424 ( .A(n_384), .B(n_342), .Y(n_424) );
AND2x4_ASAP7_75t_SL g425 ( .A(n_377), .B(n_336), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_369), .B(n_336), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_378), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_358), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_378), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_386), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_358), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_363), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_384), .B(n_18), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_386), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_360), .B(n_336), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_368), .B(n_336), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_362), .B(n_345), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_369), .B(n_345), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_372), .B(n_345), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_363), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_363), .Y(n_441) );
INVx3_ASAP7_75t_L g442 ( .A(n_389), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_362), .B(n_334), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_393), .B(n_334), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_380), .B(n_334), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_393), .B(n_325), .Y(n_446) );
INVx3_ASAP7_75t_L g447 ( .A(n_389), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_387), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_393), .B(n_325), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_380), .B(n_338), .Y(n_450) );
OR2x2_ASAP7_75t_L g451 ( .A(n_359), .B(n_338), .Y(n_451) );
INVx3_ASAP7_75t_L g452 ( .A(n_389), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_387), .B(n_325), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_392), .Y(n_454) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_359), .Y(n_455) );
BUFx2_ASAP7_75t_L g456 ( .A(n_364), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_373), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_359), .B(n_325), .Y(n_458) );
AND3x2_ASAP7_75t_L g459 ( .A(n_371), .B(n_319), .C(n_302), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_373), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_356), .B(n_19), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_392), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_372), .B(n_325), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_394), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_390), .B(n_325), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_394), .Y(n_466) );
NOR2x1p5_ASAP7_75t_L g467 ( .A(n_417), .B(n_364), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_437), .B(n_364), .Y(n_468) );
OR2x2_ASAP7_75t_L g469 ( .A(n_413), .B(n_370), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_399), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_396), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_437), .B(n_385), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_399), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_413), .B(n_370), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_409), .B(n_356), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_409), .B(n_382), .Y(n_476) );
AND3x2_ASAP7_75t_L g477 ( .A(n_461), .B(n_371), .C(n_395), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_402), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_397), .B(n_390), .Y(n_479) );
NAND2x1p5_ASAP7_75t_L g480 ( .A(n_456), .B(n_366), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_402), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_396), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_397), .B(n_370), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_407), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_400), .B(n_361), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_443), .B(n_385), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_407), .Y(n_487) );
NOR2xp67_ASAP7_75t_L g488 ( .A(n_455), .B(n_421), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_398), .B(n_383), .Y(n_489) );
NAND2x1_ASAP7_75t_L g490 ( .A(n_456), .B(n_391), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_438), .B(n_382), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_400), .B(n_361), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_398), .B(n_373), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_403), .B(n_383), .Y(n_494) );
HB1xp67_ASAP7_75t_L g495 ( .A(n_455), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_443), .B(n_366), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_438), .B(n_376), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_444), .B(n_366), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_439), .B(n_374), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_444), .B(n_371), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_396), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_403), .B(n_383), .Y(n_502) );
AND2x4_ASAP7_75t_L g503 ( .A(n_412), .B(n_391), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_416), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_405), .B(n_395), .Y(n_505) );
INVx3_ASAP7_75t_L g506 ( .A(n_421), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_411), .B(n_376), .Y(n_507) );
BUFx2_ASAP7_75t_L g508 ( .A(n_417), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_416), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_405), .B(n_349), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_418), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_406), .B(n_374), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_418), .Y(n_513) );
NAND2xp67_ASAP7_75t_L g514 ( .A(n_425), .B(n_375), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_461), .B(n_375), .Y(n_515) );
HB1xp67_ASAP7_75t_L g516 ( .A(n_401), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_420), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_406), .B(n_349), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_439), .B(n_349), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_408), .B(n_349), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_408), .B(n_349), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_420), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_427), .Y(n_523) );
INVx2_ASAP7_75t_SL g524 ( .A(n_425), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_404), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_427), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_429), .B(n_349), .Y(n_527) );
INVxp67_ASAP7_75t_L g528 ( .A(n_401), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_415), .B(n_349), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_429), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_415), .B(n_381), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_430), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_430), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_404), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_433), .B(n_20), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_419), .B(n_381), .Y(n_536) );
AND2x4_ASAP7_75t_SL g537 ( .A(n_412), .B(n_411), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_404), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_419), .B(n_381), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_434), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_426), .B(n_379), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_414), .B(n_379), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_434), .B(n_310), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_414), .B(n_379), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_454), .Y(n_545) );
INVx2_ASAP7_75t_SL g546 ( .A(n_425), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_454), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_410), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_426), .B(n_379), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_410), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_436), .B(n_381), .Y(n_551) );
OR2x2_ASAP7_75t_L g552 ( .A(n_436), .B(n_20), .Y(n_552) );
INVxp67_ASAP7_75t_L g553 ( .A(n_516), .Y(n_553) );
INVx3_ASAP7_75t_L g554 ( .A(n_537), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_507), .B(n_475), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_516), .Y(n_556) );
INVxp67_ASAP7_75t_SL g557 ( .A(n_495), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_528), .B(n_479), .Y(n_558) );
OR2x6_ASAP7_75t_L g559 ( .A(n_480), .B(n_450), .Y(n_559) );
NAND3xp33_ASAP7_75t_L g560 ( .A(n_535), .B(n_463), .C(n_424), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_528), .B(n_424), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_470), .Y(n_562) );
AO22x1_ASAP7_75t_L g563 ( .A1(n_524), .A2(n_412), .B1(n_448), .B2(n_464), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_476), .B(n_423), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_508), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_473), .Y(n_566) );
INVxp67_ASAP7_75t_L g567 ( .A(n_495), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_478), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_497), .B(n_465), .Y(n_569) );
NAND2x1_ASAP7_75t_L g570 ( .A(n_524), .B(n_421), .Y(n_570) );
INVxp67_ASAP7_75t_SL g571 ( .A(n_467), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_481), .Y(n_572) );
BUFx2_ASAP7_75t_L g573 ( .A(n_546), .Y(n_573) );
NAND2xp33_ASAP7_75t_SL g574 ( .A(n_546), .B(n_445), .Y(n_574) );
NAND2x1_ASAP7_75t_L g575 ( .A(n_488), .B(n_421), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_515), .B(n_445), .Y(n_576) );
NAND2x1_ASAP7_75t_L g577 ( .A(n_506), .B(n_442), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_499), .B(n_465), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_484), .Y(n_579) );
OAI311xp33_ASAP7_75t_L g580 ( .A1(n_552), .A2(n_450), .A3(n_451), .B1(n_458), .C1(n_463), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_479), .B(n_446), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_487), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_504), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_512), .B(n_446), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_509), .Y(n_585) );
BUFx2_ASAP7_75t_L g586 ( .A(n_468), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_511), .Y(n_587) );
OR2x2_ASAP7_75t_L g588 ( .A(n_505), .B(n_423), .Y(n_588) );
OR2x2_ASAP7_75t_L g589 ( .A(n_494), .B(n_435), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_537), .B(n_435), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_542), .B(n_449), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_518), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_515), .A2(n_412), .B1(n_449), .B2(n_459), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_483), .B(n_453), .Y(n_594) );
INVx1_ASAP7_75t_SL g595 ( .A(n_469), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_483), .B(n_453), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_500), .B(n_442), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_513), .Y(n_598) );
OR2x2_ASAP7_75t_L g599 ( .A(n_502), .B(n_451), .Y(n_599) );
INVxp67_ASAP7_75t_L g600 ( .A(n_474), .Y(n_600) );
OR2x2_ASAP7_75t_L g601 ( .A(n_485), .B(n_458), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_535), .B(n_448), .Y(n_602) );
INVx1_ASAP7_75t_SL g603 ( .A(n_510), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_472), .B(n_442), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_517), .Y(n_605) );
OR2x2_ASAP7_75t_L g606 ( .A(n_492), .B(n_466), .Y(n_606) );
AND2x2_ASAP7_75t_SL g607 ( .A(n_486), .B(n_459), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g608 ( .A(n_491), .B(n_466), .Y(n_608) );
AOI32xp33_ASAP7_75t_L g609 ( .A1(n_498), .A2(n_442), .A3(n_447), .B1(n_452), .B2(n_462), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_522), .Y(n_610) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_489), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_544), .B(n_464), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_489), .B(n_493), .Y(n_613) );
OR2x6_ASAP7_75t_L g614 ( .A(n_480), .B(n_447), .Y(n_614) );
OR2x2_ASAP7_75t_L g615 ( .A(n_493), .B(n_462), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_529), .B(n_447), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_523), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_526), .Y(n_618) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_514), .B(n_21), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_530), .Y(n_620) );
AOI222xp33_ASAP7_75t_L g621 ( .A1(n_532), .A2(n_460), .B1(n_457), .B2(n_431), .C1(n_410), .C2(n_441), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_529), .B(n_447), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_510), .B(n_452), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_533), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_540), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_520), .B(n_452), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_545), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_547), .Y(n_628) );
OR2x2_ASAP7_75t_L g629 ( .A(n_521), .B(n_460), .Y(n_629) );
NAND2xp33_ASAP7_75t_SL g630 ( .A(n_490), .B(n_452), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_558), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_558), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_556), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_606), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g635 ( .A1(n_560), .A2(n_531), .B1(n_539), .B2(n_536), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_553), .B(n_531), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_562), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_566), .Y(n_638) );
INVxp33_ASAP7_75t_L g639 ( .A(n_602), .Y(n_639) );
INVx1_ASAP7_75t_SL g640 ( .A(n_586), .Y(n_640) );
AOI21xp5_ASAP7_75t_L g641 ( .A1(n_563), .A2(n_519), .B(n_527), .Y(n_641) );
NAND3xp33_ASAP7_75t_SL g642 ( .A(n_619), .B(n_496), .C(n_301), .Y(n_642) );
INVxp67_ASAP7_75t_L g643 ( .A(n_557), .Y(n_643) );
OAI21xp33_ASAP7_75t_L g644 ( .A1(n_609), .A2(n_549), .B(n_541), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_568), .Y(n_645) );
AOI221xp5_ASAP7_75t_L g646 ( .A1(n_580), .A2(n_539), .B1(n_536), .B2(n_520), .C(n_543), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_572), .Y(n_647) );
OAI22xp5_ASAP7_75t_L g648 ( .A1(n_571), .A2(n_503), .B1(n_551), .B2(n_506), .Y(n_648) );
NAND3xp33_ASAP7_75t_L g649 ( .A(n_567), .B(n_477), .C(n_506), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_608), .B(n_477), .Y(n_650) );
OAI221xp5_ASAP7_75t_L g651 ( .A1(n_560), .A2(n_550), .B1(n_548), .B2(n_538), .C(n_534), .Y(n_651) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_593), .A2(n_503), .B1(n_548), .B2(n_538), .Y(n_652) );
INVx1_ASAP7_75t_SL g653 ( .A(n_573), .Y(n_653) );
INVxp67_ASAP7_75t_L g654 ( .A(n_565), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_561), .B(n_569), .Y(n_655) );
AOI22xp5_ASAP7_75t_L g656 ( .A1(n_574), .A2(n_503), .B1(n_550), .B2(n_525), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_611), .B(n_525), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_590), .B(n_534), .Y(n_658) );
INVx2_ASAP7_75t_SL g659 ( .A(n_554), .Y(n_659) );
AOI21xp5_ASAP7_75t_L g660 ( .A1(n_630), .A2(n_501), .B(n_482), .Y(n_660) );
OR2x2_ASAP7_75t_L g661 ( .A(n_599), .B(n_482), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_579), .Y(n_662) );
A2O1A1Ixp33_ASAP7_75t_L g663 ( .A1(n_607), .A2(n_471), .B(n_314), .C(n_457), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_578), .B(n_471), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_582), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_595), .B(n_460), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_595), .B(n_457), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_629), .Y(n_668) );
INVx1_ASAP7_75t_SL g669 ( .A(n_615), .Y(n_669) );
AND2x2_ASAP7_75t_L g670 ( .A(n_594), .B(n_441), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_612), .B(n_441), .Y(n_671) );
NAND2xp5_ASAP7_75t_SL g672 ( .A(n_621), .B(n_440), .Y(n_672) );
OAI222xp33_ASAP7_75t_L g673 ( .A1(n_559), .A2(n_440), .B1(n_432), .B2(n_431), .C1(n_428), .C2(n_422), .Y(n_673) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_592), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g675 ( .A(n_555), .B(n_21), .Y(n_675) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_576), .A2(n_428), .B1(n_422), .B2(n_432), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_621), .B(n_422), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_583), .Y(n_678) );
AOI21xp5_ASAP7_75t_L g679 ( .A1(n_614), .A2(n_327), .B(n_301), .Y(n_679) );
NAND2xp33_ASAP7_75t_R g680 ( .A(n_675), .B(n_614), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_642), .A2(n_559), .B1(n_600), .B2(n_614), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g682 ( .A1(n_640), .A2(n_616), .B1(n_622), .B2(n_604), .Y(n_682) );
OAI21xp5_ASAP7_75t_L g683 ( .A1(n_643), .A2(n_642), .B(n_653), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_631), .Y(n_684) );
AOI22xp5_ASAP7_75t_L g685 ( .A1(n_652), .A2(n_626), .B1(n_623), .B2(n_603), .Y(n_685) );
OAI21xp33_ASAP7_75t_SL g686 ( .A1(n_656), .A2(n_581), .B(n_603), .Y(n_686) );
AOI221xp5_ASAP7_75t_L g687 ( .A1(n_644), .A2(n_580), .B1(n_627), .B2(n_625), .C(n_624), .Y(n_687) );
AOI321xp33_ASAP7_75t_L g688 ( .A1(n_635), .A2(n_591), .A3(n_584), .B1(n_601), .B2(n_617), .C(n_587), .Y(n_688) );
AOI22xp5_ASAP7_75t_L g689 ( .A1(n_659), .A2(n_597), .B1(n_620), .B2(n_618), .Y(n_689) );
OAI22xp5_ASAP7_75t_L g690 ( .A1(n_650), .A2(n_570), .B1(n_588), .B2(n_589), .Y(n_690) );
AOI21xp33_ASAP7_75t_L g691 ( .A1(n_639), .A2(n_577), .B(n_575), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_632), .A2(n_585), .B1(n_610), .B2(n_605), .Y(n_692) );
AOI31xp33_ASAP7_75t_SL g693 ( .A1(n_643), .A2(n_564), .A3(n_613), .B(n_22), .Y(n_693) );
OA21x2_ASAP7_75t_L g694 ( .A1(n_677), .A2(n_628), .B(n_598), .Y(n_694) );
AOI221x1_ASAP7_75t_L g695 ( .A1(n_648), .A2(n_596), .B1(n_281), .B2(n_301), .C(n_22), .Y(n_695) );
AOI221xp5_ASAP7_75t_L g696 ( .A1(n_672), .A2(n_290), .B1(n_310), .B2(n_323), .C(n_275), .Y(n_696) );
INVxp67_ASAP7_75t_L g697 ( .A(n_633), .Y(n_697) );
OAI221xp5_ASAP7_75t_SL g698 ( .A1(n_646), .A2(n_323), .B1(n_310), .B2(n_318), .C(n_275), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_669), .A2(n_323), .B1(n_28), .B2(n_30), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_655), .B(n_27), .Y(n_700) );
O2A1O1Ixp5_ASAP7_75t_L g701 ( .A1(n_673), .A2(n_663), .B(n_649), .C(n_660), .Y(n_701) );
AOI21xp5_ASAP7_75t_L g702 ( .A1(n_673), .A2(n_33), .B(n_35), .Y(n_702) );
AOI211xp5_ASAP7_75t_L g703 ( .A1(n_651), .A2(n_36), .B(n_40), .C(n_42), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_637), .Y(n_704) );
AOI211xp5_ASAP7_75t_SL g705 ( .A1(n_654), .A2(n_44), .B(n_45), .C(n_46), .Y(n_705) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_634), .A2(n_47), .B1(n_48), .B2(n_60), .Y(n_706) );
AOI322xp5_ASAP7_75t_L g707 ( .A1(n_636), .A2(n_61), .A3(n_63), .B1(n_64), .B2(n_67), .C1(n_70), .C2(n_72), .Y(n_707) );
AOI321xp33_ASAP7_75t_L g708 ( .A1(n_676), .A2(n_641), .A3(n_678), .B1(n_647), .B2(n_645), .C(n_665), .Y(n_708) );
NAND2xp5_ASAP7_75t_SL g709 ( .A(n_674), .B(n_73), .Y(n_709) );
AOI211xp5_ASAP7_75t_L g710 ( .A1(n_654), .A2(n_74), .B(n_75), .C(n_78), .Y(n_710) );
A2O1A1Ixp33_ASAP7_75t_L g711 ( .A1(n_679), .A2(n_80), .B(n_81), .C(n_84), .Y(n_711) );
NAND4xp25_ASAP7_75t_L g712 ( .A(n_638), .B(n_662), .C(n_664), .D(n_666), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_674), .B(n_85), .Y(n_713) );
OAI211xp5_ASAP7_75t_SL g714 ( .A1(n_667), .A2(n_87), .B(n_88), .C(n_104), .Y(n_714) );
OAI211xp5_ASAP7_75t_L g715 ( .A1(n_671), .A2(n_668), .B(n_661), .C(n_657), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_670), .B(n_658), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_631), .B(n_632), .Y(n_717) );
OA21x2_ASAP7_75t_L g718 ( .A1(n_643), .A2(n_677), .B(n_672), .Y(n_718) );
NAND2xp33_ASAP7_75t_L g719 ( .A(n_683), .B(n_681), .Y(n_719) );
NOR3xp33_ASAP7_75t_L g720 ( .A(n_701), .B(n_687), .C(n_686), .Y(n_720) );
NAND4xp25_ASAP7_75t_SL g721 ( .A(n_715), .B(n_691), .C(n_695), .D(n_685), .Y(n_721) );
NOR3xp33_ASAP7_75t_L g722 ( .A(n_714), .B(n_713), .C(n_700), .Y(n_722) );
OAI21xp5_ASAP7_75t_L g723 ( .A1(n_718), .A2(n_702), .B(n_690), .Y(n_723) );
NOR2x1_ASAP7_75t_L g724 ( .A(n_693), .B(n_711), .Y(n_724) );
NAND4xp25_ASAP7_75t_L g725 ( .A(n_680), .B(n_708), .C(n_688), .D(n_703), .Y(n_725) );
OR2x2_ASAP7_75t_L g726 ( .A(n_721), .B(n_712), .Y(n_726) );
NOR4xp25_ASAP7_75t_L g727 ( .A(n_725), .B(n_697), .C(n_698), .D(n_704), .Y(n_727) );
NAND3xp33_ASAP7_75t_L g728 ( .A(n_720), .B(n_718), .C(n_707), .Y(n_728) );
NOR3xp33_ASAP7_75t_L g729 ( .A(n_724), .B(n_710), .C(n_699), .Y(n_729) );
XOR2xp5_ASAP7_75t_L g730 ( .A(n_726), .B(n_723), .Y(n_730) );
NOR3xp33_ASAP7_75t_L g731 ( .A(n_728), .B(n_719), .C(n_722), .Y(n_731) );
AND3x4_ASAP7_75t_L g732 ( .A(n_727), .B(n_694), .C(n_705), .Y(n_732) );
NAND2xp33_ASAP7_75t_L g733 ( .A(n_731), .B(n_729), .Y(n_733) );
XOR2x1_ASAP7_75t_L g734 ( .A(n_730), .B(n_694), .Y(n_734) );
HB1xp67_ASAP7_75t_L g735 ( .A(n_734), .Y(n_735) );
NAND2xp33_ASAP7_75t_R g736 ( .A(n_733), .B(n_732), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_735), .Y(n_737) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_736), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g739 ( .A1(n_738), .A2(n_684), .B1(n_717), .B2(n_692), .Y(n_739) );
AO21x2_ASAP7_75t_L g740 ( .A1(n_739), .A2(n_737), .B(n_709), .Y(n_740) );
OA21x2_ASAP7_75t_L g741 ( .A1(n_740), .A2(n_706), .B(n_682), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_741), .A2(n_689), .B1(n_696), .B2(n_716), .Y(n_742) );
endmodule