module real_aes_15811_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_800;
wire n_618;
wire n_778;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_357;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_551;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_746;
wire n_656;
wire n_178;
wire n_409;
wire n_860;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_855;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
CKINVDCx5p33_ASAP7_75t_R g577 ( .A(n_0), .Y(n_577) );
AND2x4_ASAP7_75t_L g856 ( .A(n_1), .B(n_857), .Y(n_856) );
AOI22xp5_ASAP7_75t_L g257 ( .A1(n_2), .A2(n_4), .B1(n_258), .B2(n_259), .Y(n_257) );
AOI22xp33_ASAP7_75t_L g244 ( .A1(n_3), .A2(n_20), .B1(n_158), .B2(n_239), .Y(n_244) );
AOI22xp33_ASAP7_75t_L g194 ( .A1(n_5), .A2(n_52), .B1(n_166), .B2(n_195), .Y(n_194) );
BUFx3_ASAP7_75t_L g611 ( .A(n_6), .Y(n_611) );
AOI22xp5_ASAP7_75t_L g128 ( .A1(n_7), .A2(n_13), .B1(n_129), .B2(n_131), .Y(n_128) );
INVx1_ASAP7_75t_L g857 ( .A(n_8), .Y(n_857) );
CKINVDCx5p33_ASAP7_75t_R g238 ( .A(n_9), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_10), .B(n_164), .Y(n_625) );
OR2x2_ASAP7_75t_L g115 ( .A(n_11), .B(n_29), .Y(n_115) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_12), .Y(n_130) );
NAND2xp5_ASAP7_75t_SL g592 ( .A(n_14), .B(n_200), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_15), .B(n_173), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_16), .A2(n_84), .B1(n_200), .B2(n_239), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g116 ( .A1(n_17), .A2(n_117), .B1(n_503), .B2(n_504), .Y(n_116) );
INVx1_ASAP7_75t_L g503 ( .A(n_17), .Y(n_503) );
OAI21x1_ASAP7_75t_L g141 ( .A1(n_18), .A2(n_48), .B(n_142), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g248 ( .A(n_19), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_21), .B(n_158), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_22), .B(n_134), .Y(n_214) );
INVx4_ASAP7_75t_R g182 ( .A(n_23), .Y(n_182) );
AO32x2_ASAP7_75t_L g536 ( .A1(n_24), .A2(n_152), .A3(n_153), .B1(n_537), .B2(n_540), .Y(n_536) );
AO32x1_ASAP7_75t_L g641 ( .A1(n_24), .A2(n_152), .A3(n_153), .B1(n_537), .B2(n_540), .Y(n_641) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_25), .B(n_158), .Y(n_221) );
INVx1_ASAP7_75t_L g263 ( .A(n_26), .Y(n_263) );
A2O1A1Ixp33_ASAP7_75t_SL g236 ( .A1(n_27), .A2(n_129), .B(n_133), .C(n_237), .Y(n_236) );
AOI22xp33_ASAP7_75t_L g245 ( .A1(n_28), .A2(n_45), .B1(n_129), .B2(n_136), .Y(n_245) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_30), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_31), .A2(n_51), .B1(n_158), .B2(n_183), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g538 ( .A1(n_32), .A2(n_89), .B1(n_136), .B2(n_239), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_33), .B(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g553 ( .A(n_34), .B(n_549), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_35), .B(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g218 ( .A(n_36), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_37), .B(n_129), .Y(n_220) );
AOI22xp33_ASAP7_75t_L g561 ( .A1(n_38), .A2(n_67), .B1(n_136), .B2(n_562), .Y(n_561) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_39), .Y(n_156) );
INVx2_ASAP7_75t_L g105 ( .A(n_40), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g861 ( .A(n_41), .Y(n_861) );
INVx1_ASAP7_75t_L g111 ( .A(n_42), .Y(n_111) );
BUFx3_ASAP7_75t_L g517 ( .A(n_42), .Y(n_517) );
CKINVDCx5p33_ASAP7_75t_R g509 ( .A(n_43), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_44), .B(n_555), .Y(n_554) );
CKINVDCx5p33_ASAP7_75t_R g184 ( .A(n_46), .Y(n_184) );
AOI22xp33_ASAP7_75t_L g135 ( .A1(n_47), .A2(n_83), .B1(n_129), .B2(n_136), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g573 ( .A(n_49), .Y(n_573) );
CKINVDCx5p33_ASAP7_75t_R g602 ( .A(n_50), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g598 ( .A1(n_53), .A2(n_77), .B1(n_202), .B2(n_549), .Y(n_598) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_54), .Y(n_147) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_55), .A2(n_81), .B1(n_200), .B2(n_239), .Y(n_607) );
INVx1_ASAP7_75t_L g142 ( .A(n_56), .Y(n_142) );
AND2x4_ASAP7_75t_L g144 ( .A(n_57), .B(n_145), .Y(n_144) );
AOI22xp33_ASAP7_75t_L g255 ( .A1(n_58), .A2(n_88), .B1(n_136), .B2(n_256), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_59), .A2(n_525), .B1(n_851), .B2(n_852), .Y(n_524) );
INVx1_ASAP7_75t_L g851 ( .A(n_59), .Y(n_851) );
AO22x1_ASAP7_75t_L g198 ( .A1(n_60), .A2(n_72), .B1(n_199), .B2(n_201), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_61), .B(n_239), .Y(n_624) );
INVx1_ASAP7_75t_L g145 ( .A(n_62), .Y(n_145) );
AND2x2_ASAP7_75t_L g240 ( .A(n_63), .B(n_152), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_64), .B(n_152), .Y(n_630) );
A2O1A1Ixp33_ASAP7_75t_L g575 ( .A1(n_65), .A2(n_166), .B(n_193), .C(n_576), .Y(n_575) );
NAND3xp33_ASAP7_75t_L g629 ( .A(n_66), .B(n_239), .C(n_628), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_68), .B(n_166), .Y(n_165) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_69), .Y(n_231) );
AND2x2_ASAP7_75t_L g578 ( .A(n_70), .B(n_187), .Y(n_578) );
CKINVDCx5p33_ASAP7_75t_R g565 ( .A(n_71), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_73), .B(n_158), .Y(n_157) );
AOI22xp33_ASAP7_75t_L g600 ( .A1(n_74), .A2(n_94), .B1(n_200), .B2(n_202), .Y(n_600) );
INVx2_ASAP7_75t_L g134 ( .A(n_75), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_76), .B(n_159), .Y(n_590) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_78), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_79), .B(n_152), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g572 ( .A(n_80), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_82), .B(n_140), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_85), .B(n_628), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_86), .A2(n_98), .B1(n_136), .B2(n_183), .Y(n_608) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_87), .B(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_90), .B(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g113 ( .A(n_91), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_92), .B(n_173), .Y(n_556) );
A2O1A1Ixp33_ASAP7_75t_L g176 ( .A1(n_93), .A2(n_138), .B(n_166), .C(n_177), .Y(n_176) );
AND2x2_ASAP7_75t_L g186 ( .A(n_95), .B(n_187), .Y(n_186) );
NAND2xp33_ASAP7_75t_L g163 ( .A(n_96), .B(n_164), .Y(n_163) );
CKINVDCx5p33_ASAP7_75t_R g587 ( .A(n_97), .Y(n_587) );
AOI21xp5_ASAP7_75t_L g99 ( .A1(n_100), .A2(n_853), .B(n_860), .Y(n_99) );
OR2x6_ASAP7_75t_L g100 ( .A(n_101), .B(n_518), .Y(n_100) );
AO21x1_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_106), .B(n_508), .Y(n_101) );
CKINVDCx11_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
BUFx6f_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
INVx3_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_105), .B(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g521 ( .A(n_105), .Y(n_521) );
OAI21xp5_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_116), .B(n_505), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx4_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g507 ( .A(n_109), .Y(n_507) );
AND3x2_ASAP7_75t_L g109 ( .A(n_110), .B(n_112), .C(n_114), .Y(n_109) );
NOR3xp33_ASAP7_75t_L g854 ( .A(n_110), .B(n_112), .C(n_855), .Y(n_854) );
HB1xp67_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
BUFx2_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
INVx2_ASAP7_75t_L g515 ( .A(n_113), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_114), .B(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
NOR2x1_ASAP7_75t_L g516 ( .A(n_115), .B(n_517), .Y(n_516) );
BUFx2_ASAP7_75t_L g859 ( .A(n_115), .Y(n_859) );
HB1xp67_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx2_ASAP7_75t_L g504 ( .A(n_118), .Y(n_504) );
AND2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_412), .Y(n_118) );
NOR3xp33_ASAP7_75t_L g119 ( .A(n_120), .B(n_328), .C(n_359), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_294), .Y(n_120) );
AOI211x1_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_206), .B(n_249), .C(n_280), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_170), .Y(n_123) );
AND2x2_ASAP7_75t_L g435 ( .A(n_124), .B(n_310), .Y(n_435) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_149), .Y(n_124) );
INVx1_ASAP7_75t_L g320 ( .A(n_125), .Y(n_320) );
OR2x2_ASAP7_75t_L g441 ( .A(n_125), .B(n_292), .Y(n_441) );
INVx2_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_L g277 ( .A(n_126), .B(n_150), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_126), .B(n_292), .Y(n_291) );
INVx2_ASAP7_75t_L g309 ( .A(n_126), .Y(n_309) );
OR2x2_ASAP7_75t_L g340 ( .A(n_126), .B(n_171), .Y(n_340) );
AND2x2_ASAP7_75t_L g354 ( .A(n_126), .B(n_171), .Y(n_354) );
AND2x2_ASAP7_75t_L g391 ( .A(n_126), .B(n_347), .Y(n_391) );
AO31x2_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_139), .A3(n_143), .B(n_146), .Y(n_126) );
OAI22x1_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_132), .B1(n_135), .B2(n_137), .Y(n_127) );
INVx4_ASAP7_75t_L g131 ( .A(n_129), .Y(n_131) );
INVx3_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_130), .Y(n_136) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_130), .Y(n_158) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_130), .Y(n_164) );
INVx1_ASAP7_75t_L g166 ( .A(n_130), .Y(n_166) );
INVx1_ASAP7_75t_L g178 ( .A(n_130), .Y(n_178) );
INVx1_ASAP7_75t_L g183 ( .A(n_130), .Y(n_183) );
BUFx6f_ASAP7_75t_L g200 ( .A(n_130), .Y(n_200) );
INVx1_ASAP7_75t_L g202 ( .A(n_130), .Y(n_202) );
INVx1_ASAP7_75t_L g233 ( .A(n_130), .Y(n_233) );
INVx2_ASAP7_75t_L g239 ( .A(n_130), .Y(n_239) );
O2A1O1Ixp33_ASAP7_75t_L g155 ( .A1(n_131), .A2(n_156), .B(n_157), .C(n_159), .Y(n_155) );
OAI22xp5_ASAP7_75t_L g243 ( .A1(n_132), .A2(n_192), .B1(n_244), .B2(n_245), .Y(n_243) );
OAI22xp5_ASAP7_75t_L g254 ( .A1(n_132), .A2(n_137), .B1(n_255), .B2(n_257), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_132), .A2(n_553), .B(n_554), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g560 ( .A1(n_132), .A2(n_192), .B1(n_561), .B2(n_563), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g597 ( .A1(n_132), .A2(n_598), .B1(n_599), .B2(n_600), .Y(n_597) );
OAI22xp5_ASAP7_75t_L g606 ( .A1(n_132), .A2(n_133), .B1(n_607), .B2(n_608), .Y(n_606) );
INVx6_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_133), .A2(n_163), .B(n_165), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_133), .B(n_198), .Y(n_197) );
A2O1A1Ixp33_ASAP7_75t_L g293 ( .A1(n_133), .A2(n_191), .B(n_198), .C(n_204), .Y(n_293) );
OAI22xp5_ASAP7_75t_L g537 ( .A1(n_133), .A2(n_235), .B1(n_538), .B2(n_539), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g623 ( .A1(n_133), .A2(n_624), .B(n_625), .Y(n_623) );
BUFx8_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g138 ( .A(n_134), .Y(n_138) );
INVx2_ASAP7_75t_L g161 ( .A(n_134), .Y(n_161) );
INVx1_ASAP7_75t_L g217 ( .A(n_134), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_136), .B(n_216), .Y(n_215) );
INVx2_ASAP7_75t_L g258 ( .A(n_136), .Y(n_258) );
INVx2_ASAP7_75t_L g551 ( .A(n_136), .Y(n_551) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_137), .B(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g574 ( .A(n_138), .Y(n_574) );
INVx1_ASAP7_75t_SL g599 ( .A(n_138), .Y(n_599) );
INVx2_ASAP7_75t_L g621 ( .A(n_139), .Y(n_621) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g148 ( .A(n_140), .Y(n_148) );
INVx2_ASAP7_75t_L g174 ( .A(n_140), .Y(n_174) );
OAI21xp33_ASAP7_75t_L g204 ( .A1(n_140), .A2(n_196), .B(n_205), .Y(n_204) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_141), .Y(n_153) );
INVx2_ASAP7_75t_L g185 ( .A(n_143), .Y(n_185) );
BUFx10_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx10_ASAP7_75t_L g169 ( .A(n_144), .Y(n_169) );
INVx1_ASAP7_75t_L g205 ( .A(n_144), .Y(n_205) );
INVx1_ASAP7_75t_L g261 ( .A(n_144), .Y(n_261) );
AO31x2_ASAP7_75t_L g558 ( .A1(n_144), .A2(n_559), .A3(n_560), .B(n_564), .Y(n_558) );
NOR2xp33_ASAP7_75t_L g146 ( .A(n_147), .B(n_148), .Y(n_146) );
INVx2_ASAP7_75t_L g187 ( .A(n_148), .Y(n_187) );
BUFx2_ASAP7_75t_L g227 ( .A(n_148), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_148), .B(n_248), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_148), .B(n_263), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_148), .B(n_602), .Y(n_601) );
BUFx2_ASAP7_75t_L g271 ( .A(n_149), .Y(n_271) );
AND2x2_ASAP7_75t_L g322 ( .A(n_149), .B(n_188), .Y(n_322) );
AND2x2_ASAP7_75t_L g465 ( .A(n_149), .B(n_171), .Y(n_465) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx3_ASAP7_75t_L g289 ( .A(n_150), .Y(n_289) );
AND2x2_ASAP7_75t_L g308 ( .A(n_150), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g345 ( .A(n_150), .Y(n_345) );
AND2x2_ASAP7_75t_L g369 ( .A(n_150), .B(n_171), .Y(n_369) );
NAND2x1p5_ASAP7_75t_L g150 ( .A(n_151), .B(n_154), .Y(n_150) );
NOR2x1_ASAP7_75t_L g167 ( .A(n_152), .B(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g246 ( .A(n_152), .Y(n_246) );
INVx4_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
AND2x2_ASAP7_75t_L g222 ( .A(n_153), .B(n_169), .Y(n_222) );
INVx2_ASAP7_75t_SL g545 ( .A(n_153), .Y(n_545) );
BUFx3_ASAP7_75t_L g559 ( .A(n_153), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_153), .B(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g584 ( .A(n_153), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_153), .B(n_610), .Y(n_609) );
OAI21x1_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_162), .B(n_167), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_158), .B(n_231), .Y(n_230) );
INVx2_ASAP7_75t_L g562 ( .A(n_158), .Y(n_562) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_158), .A2(n_183), .B1(n_572), .B2(n_573), .Y(n_571) );
INVx2_ASAP7_75t_SL g159 ( .A(n_160), .Y(n_159) );
OAI22xp5_ASAP7_75t_L g589 ( .A1(n_160), .A2(n_590), .B1(n_591), .B2(n_592), .Y(n_589) );
INVx2_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
BUFx3_ASAP7_75t_L g193 ( .A(n_161), .Y(n_193) );
OAI22xp33_ASAP7_75t_L g181 ( .A1(n_164), .A2(n_182), .B1(n_183), .B2(n_184), .Y(n_181) );
INVx2_ASAP7_75t_L g256 ( .A(n_164), .Y(n_256) );
INVx1_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
AO31x2_ASAP7_75t_L g242 ( .A1(n_169), .A2(n_243), .A3(n_246), .B(n_247), .Y(n_242) );
OAI21x1_ASAP7_75t_L g585 ( .A1(n_169), .A2(n_586), .B(n_589), .Y(n_585) );
AOI31xp67_ASAP7_75t_L g605 ( .A1(n_169), .A2(n_246), .A3(n_606), .B(n_609), .Y(n_605) );
OAI21x1_ASAP7_75t_L g622 ( .A1(n_169), .A2(n_623), .B(n_626), .Y(n_622) );
HB1xp67_ASAP7_75t_L g269 ( .A(n_170), .Y(n_269) );
AND2x2_ASAP7_75t_L g330 ( .A(n_170), .B(n_319), .Y(n_330) );
INVx2_ASAP7_75t_L g462 ( .A(n_170), .Y(n_462) );
AND2x2_ASAP7_75t_L g170 ( .A(n_171), .B(n_188), .Y(n_170) );
INVx1_ASAP7_75t_L g267 ( .A(n_171), .Y(n_267) );
AND2x4_ASAP7_75t_L g279 ( .A(n_171), .B(n_189), .Y(n_279) );
INVx2_ASAP7_75t_L g347 ( .A(n_171), .Y(n_347) );
AO21x2_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_175), .B(n_186), .Y(n_171) );
AOI21x1_ASAP7_75t_L g568 ( .A1(n_172), .A2(n_569), .B(n_578), .Y(n_568) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_180), .B(n_185), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_178), .B(n_179), .Y(n_177) );
INVx2_ASAP7_75t_L g195 ( .A(n_178), .Y(n_195) );
INVx1_ASAP7_75t_L g591 ( .A(n_183), .Y(n_591) );
AND2x2_ASAP7_75t_L g346 ( .A(n_188), .B(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g353 ( .A(n_188), .Y(n_353) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AND2x2_ASAP7_75t_L g431 ( .A(n_189), .B(n_347), .Y(n_431) );
AOI21x1_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_197), .B(n_203), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
OAI21x1_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_194), .B(n_196), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g219 ( .A1(n_192), .A2(n_220), .B(n_221), .Y(n_219) );
AOI21x1_ASAP7_75t_L g547 ( .A1(n_192), .A2(n_548), .B(n_550), .Y(n_547) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVxp67_ASAP7_75t_SL g199 ( .A(n_200), .Y(n_199) );
INVx3_ASAP7_75t_L g555 ( .A(n_200), .Y(n_555) );
OAI21xp33_ASAP7_75t_SL g213 ( .A1(n_201), .A2(n_214), .B(n_215), .Y(n_213) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g576 ( .A(n_202), .B(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_205), .A2(n_229), .B(n_236), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g569 ( .A1(n_205), .A2(n_570), .B(n_575), .Y(n_569) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_208), .B(n_223), .Y(n_207) );
OR2x2_ASAP7_75t_L g336 ( .A(n_208), .B(n_224), .Y(n_336) );
AND2x2_ASAP7_75t_L g474 ( .A(n_208), .B(n_418), .Y(n_474) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
AND2x4_ASAP7_75t_L g251 ( .A(n_209), .B(n_252), .Y(n_251) );
OR2x2_ASAP7_75t_L g356 ( .A(n_209), .B(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_209), .B(n_298), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_209), .B(n_274), .Y(n_411) );
INVx3_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx1_ASAP7_75t_L g268 ( .A(n_210), .Y(n_268) );
AND2x2_ASAP7_75t_L g284 ( .A(n_210), .B(n_285), .Y(n_284) );
NAND2x1p5_ASAP7_75t_SL g297 ( .A(n_210), .B(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g305 ( .A(n_210), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_210), .B(n_274), .Y(n_376) );
AND2x2_ASAP7_75t_L g424 ( .A(n_210), .B(n_253), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_210), .B(n_252), .Y(n_467) );
BUFx2_ASAP7_75t_L g486 ( .A(n_210), .Y(n_486) );
AND2x4_ASAP7_75t_L g210 ( .A(n_211), .B(n_212), .Y(n_210) );
OAI21xp5_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_219), .B(n_222), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_217), .B(n_218), .Y(n_216) );
BUFx4f_ASAP7_75t_L g235 ( .A(n_217), .Y(n_235) );
INVx1_ASAP7_75t_L g628 ( .A(n_217), .Y(n_628) );
INVx1_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
OR2x2_ASAP7_75t_L g270 ( .A(n_224), .B(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g383 ( .A(n_224), .Y(n_383) );
OR2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_241), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g286 ( .A(n_225), .B(n_253), .Y(n_286) );
INVx2_ASAP7_75t_L g298 ( .A(n_225), .Y(n_298) );
AND2x2_ASAP7_75t_L g334 ( .A(n_225), .B(n_242), .Y(n_334) );
INVx2_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx1_ASAP7_75t_L g274 ( .A(n_226), .Y(n_274) );
AOI21x1_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_228), .B(n_240), .Y(n_226) );
AO31x2_ASAP7_75t_L g253 ( .A1(n_227), .A2(n_254), .A3(n_260), .B(n_262), .Y(n_253) );
OAI21xp5_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_232), .B(n_235), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_233), .B(n_234), .Y(n_232) );
INVx2_ASAP7_75t_L g259 ( .A(n_233), .Y(n_259) );
O2A1O1Ixp5_ASAP7_75t_L g586 ( .A1(n_235), .A2(n_259), .B(n_587), .C(n_588), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_238), .B(n_239), .Y(n_237) );
INVx2_ASAP7_75t_SL g549 ( .A(n_239), .Y(n_549) );
INVx1_ASAP7_75t_L g358 ( .A(n_241), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_241), .B(n_253), .Y(n_375) );
INVx2_ASAP7_75t_SL g241 ( .A(n_242), .Y(n_241) );
BUFx2_ASAP7_75t_L g285 ( .A(n_242), .Y(n_285) );
OR2x2_ASAP7_75t_L g317 ( .A(n_242), .B(n_253), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_242), .B(n_253), .Y(n_395) );
OAI22xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_270), .B1(n_272), .B2(n_276), .Y(n_249) );
AOI22xp5_ASAP7_75t_L g250 ( .A1(n_251), .A2(n_264), .B1(n_268), .B2(n_269), .Y(n_250) );
INVx2_ASAP7_75t_L g275 ( .A(n_251), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_251), .B(n_334), .Y(n_348) );
AND2x2_ASAP7_75t_L g382 ( .A(n_251), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g300 ( .A(n_253), .Y(n_300) );
INVx1_ASAP7_75t_L g306 ( .A(n_253), .Y(n_306) );
AO31x2_ASAP7_75t_L g596 ( .A1(n_260), .A2(n_559), .A3(n_597), .B(n_601), .Y(n_596) );
INVx2_ASAP7_75t_SL g260 ( .A(n_261), .Y(n_260) );
INVx2_ASAP7_75t_SL g540 ( .A(n_261), .Y(n_540) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
OR2x2_ASAP7_75t_L g440 ( .A(n_266), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g321 ( .A(n_267), .Y(n_321) );
AND3x1_ASAP7_75t_L g425 ( .A(n_267), .B(n_288), .C(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g381 ( .A(n_268), .Y(n_381) );
AND2x4_ASAP7_75t_L g417 ( .A(n_268), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g455 ( .A(n_271), .Y(n_455) );
INVx1_ASAP7_75t_L g459 ( .A(n_272), .Y(n_459) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
OR2x2_ASAP7_75t_L g432 ( .A(n_273), .B(n_433), .Y(n_432) );
INVxp67_ASAP7_75t_SL g480 ( .A(n_273), .Y(n_480) );
INVxp67_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g380 ( .A(n_274), .B(n_358), .Y(n_380) );
AND2x2_ASAP7_75t_L g422 ( .A(n_274), .B(n_289), .Y(n_422) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_274), .Y(n_426) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_277), .B(n_278), .Y(n_276) );
O2A1O1Ixp33_ASAP7_75t_L g341 ( .A1(n_277), .A2(n_278), .B(n_342), .C(n_348), .Y(n_341) );
NAND2x1_ASAP7_75t_L g385 ( .A(n_277), .B(n_386), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_277), .B(n_435), .Y(n_481) );
INVx3_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_279), .B(n_308), .Y(n_327) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
NAND2xp5_ASAP7_75t_SL g281 ( .A(n_282), .B(n_287), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
INVx2_ASAP7_75t_L g303 ( .A(n_285), .Y(n_303) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_286), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g428 ( .A(n_287), .B(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g287 ( .A(n_288), .B(n_290), .Y(n_287) );
AND2x2_ASAP7_75t_L g337 ( .A(n_288), .B(n_338), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_288), .B(n_354), .Y(n_401) );
NAND2x1p5_ASAP7_75t_L g407 ( .A(n_288), .B(n_408), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_288), .B(n_346), .Y(n_502) );
INVx3_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
BUFx2_ASAP7_75t_L g485 ( .A(n_289), .Y(n_485) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g311 ( .A(n_292), .Y(n_311) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AOI21xp5_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_307), .B(n_312), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_301), .Y(n_295) );
OR2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_299), .Y(n_296) );
OAI33xp33_ASAP7_75t_L g361 ( .A1(n_297), .A2(n_302), .A3(n_362), .B1(n_363), .B2(n_365), .B3(n_366), .Y(n_361) );
OR2x2_ASAP7_75t_L g493 ( .A(n_297), .B(n_317), .Y(n_493) );
INVx2_ASAP7_75t_L g495 ( .A(n_297), .Y(n_495) );
INVx1_ASAP7_75t_L g316 ( .A(n_298), .Y(n_316) );
OR2x2_ASAP7_75t_L g357 ( .A(n_298), .B(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_302), .B(n_304), .Y(n_301) );
INVx1_ASAP7_75t_L g365 ( .A(n_302), .Y(n_365) );
NOR3xp33_ASAP7_75t_L g483 ( .A(n_302), .B(n_484), .C(n_486), .Y(n_483) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_303), .B(n_443), .Y(n_442) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_303), .B(n_467), .Y(n_471) );
AND2x4_ASAP7_75t_L g500 ( .A(n_303), .B(n_501), .Y(n_500) );
INVxp67_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g326 ( .A(n_305), .Y(n_326) );
OR2x2_ASAP7_75t_L g332 ( .A(n_305), .B(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g445 ( .A(n_305), .B(n_380), .Y(n_445) );
INVx1_ASAP7_75t_L g501 ( .A(n_305), .Y(n_501) );
AND2x4_ASAP7_75t_SL g307 ( .A(n_308), .B(n_310), .Y(n_307) );
INVx1_ASAP7_75t_L g324 ( .A(n_308), .Y(n_324) );
INVx1_ASAP7_75t_L g367 ( .A(n_309), .Y(n_367) );
AND2x2_ASAP7_75t_L g408 ( .A(n_309), .B(n_311), .Y(n_408) );
INVx1_ASAP7_75t_L g448 ( .A(n_310), .Y(n_448) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g339 ( .A(n_311), .B(n_340), .Y(n_339) );
OAI22xp33_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_318), .B1(n_325), .B2(n_327), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
OR2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_317), .Y(n_315) );
INVx2_ASAP7_75t_L g404 ( .A(n_317), .Y(n_404) );
INVx2_ASAP7_75t_L g418 ( .A(n_317), .Y(n_418) );
AOI211xp5_ASAP7_75t_L g318 ( .A1(n_319), .A2(n_321), .B(n_322), .C(n_323), .Y(n_318) );
INVx1_ASAP7_75t_L g362 ( .A(n_319), .Y(n_362) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_320), .B(n_345), .Y(n_447) );
OR2x2_ASAP7_75t_L g463 ( .A(n_320), .B(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g476 ( .A(n_320), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_322), .B(n_390), .Y(n_451) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_SL g328 ( .A(n_329), .B(n_349), .Y(n_328) );
AOI221xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_331), .B1(n_335), .B2(n_337), .C(n_341), .Y(n_329) );
INVx2_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OAI32xp33_ASAP7_75t_L g498 ( .A1(n_332), .A2(n_429), .A3(n_447), .B1(n_499), .B2(n_502), .Y(n_498) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g468 ( .A(n_334), .Y(n_468) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
OAI21xp5_ASAP7_75t_L g349 ( .A1(n_337), .A2(n_350), .B(n_355), .Y(n_349) );
NAND2x1_ASAP7_75t_L g497 ( .A(n_338), .B(n_485), .Y(n_497) );
INVx2_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
INVx2_ASAP7_75t_L g372 ( .A(n_340), .Y(n_372) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_346), .Y(n_343) );
AND2x2_ASAP7_75t_L g491 ( .A(n_344), .B(n_372), .Y(n_491) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g439 ( .A(n_345), .Y(n_439) );
INVx2_ASAP7_75t_L g392 ( .A(n_346), .Y(n_392) );
INVx2_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_352), .B(n_354), .Y(n_351) );
AND2x2_ASAP7_75t_L g368 ( .A(n_352), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g387 ( .A(n_353), .Y(n_387) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NAND4xp25_ASAP7_75t_L g359 ( .A(n_360), .B(n_377), .C(n_388), .D(n_399), .Y(n_359) );
AOI22xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_368), .B1(n_370), .B2(n_373), .Y(n_360) );
OAI22xp5_ASAP7_75t_L g489 ( .A1(n_362), .A2(n_490), .B1(n_492), .B2(n_493), .Y(n_489) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AND2x2_ASAP7_75t_L g472 ( .A(n_367), .B(n_431), .Y(n_472) );
AND2x2_ASAP7_75t_L g475 ( .A(n_369), .B(n_476), .Y(n_475) );
AOI22xp5_ASAP7_75t_L g388 ( .A1(n_370), .A2(n_389), .B1(n_393), .B2(n_396), .Y(n_388) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OR2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
OR2x2_ASAP7_75t_L g410 ( .A(n_375), .B(n_411), .Y(n_410) );
OR2x2_ASAP7_75t_L g394 ( .A(n_376), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g405 ( .A(n_376), .Y(n_405) );
OAI21xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_382), .B(n_384), .Y(n_377) );
O2A1O1Ixp33_ASAP7_75t_L g482 ( .A1(n_378), .A2(n_483), .B(n_487), .C(n_489), .Y(n_482) );
AND2x2_ASAP7_75t_L g378 ( .A(n_379), .B(n_381), .Y(n_378) );
INVxp67_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g457 ( .A(n_380), .Y(n_457) );
AND2x4_ASAP7_75t_L g450 ( .A(n_383), .B(n_424), .Y(n_450) );
INVx2_ASAP7_75t_SL g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_390), .B(n_392), .Y(n_389) );
OAI21xp33_ASAP7_75t_L g415 ( .A1(n_390), .A2(n_416), .B(n_419), .Y(n_415) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g421 ( .A(n_391), .B(n_422), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_391), .B(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
OR2x2_ASAP7_75t_L g397 ( .A(n_395), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g427 ( .A1(n_397), .A2(n_428), .B1(n_432), .B2(n_434), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_402), .B1(n_406), .B2(n_409), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_404), .Y(n_420) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_413), .B(n_477), .Y(n_412) );
NAND4xp25_ASAP7_75t_L g413 ( .A(n_414), .B(n_436), .C(n_452), .D(n_469), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_415), .B(n_427), .Y(n_414) );
INVx2_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
AND2x2_ASAP7_75t_L g479 ( .A(n_417), .B(n_480), .Y(n_479) );
AOI22xp5_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_421), .B1(n_423), .B2(n_425), .Y(n_419) );
INVxp67_ASAP7_75t_L g443 ( .A(n_423), .Y(n_443) );
BUFx2_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g433 ( .A(n_424), .Y(n_433) );
AND2x2_ASAP7_75t_L g456 ( .A(n_424), .B(n_457), .Y(n_456) );
INVx3_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
AOI21xp5_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_442), .B(n_444), .Y(n_436) );
NOR2x1_ASAP7_75t_L g437 ( .A(n_438), .B(n_440), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
OR2x6_ASAP7_75t_L g461 ( .A(n_439), .B(n_462), .Y(n_461) );
INVx3_ASAP7_75t_L g458 ( .A(n_440), .Y(n_458) );
OAI32xp33_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_446), .A3(n_448), .B1(n_449), .B2(n_451), .Y(n_444) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AOI221xp5_ASAP7_75t_L g452 ( .A1(n_453), .A2(n_456), .B1(n_458), .B2(n_459), .C(n_460), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_463), .B(n_466), .Y(n_460) );
INVx2_ASAP7_75t_SL g464 ( .A(n_465), .Y(n_464) );
OR2x2_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
NOR2x1_ASAP7_75t_L g469 ( .A(n_470), .B(n_473), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_472), .Y(n_470) );
INVx1_ASAP7_75t_L g492 ( .A(n_471), .Y(n_492) );
INVx1_ASAP7_75t_L g488 ( .A(n_472), .Y(n_488) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
OAI211xp5_ASAP7_75t_SL g477 ( .A1(n_478), .A2(n_481), .B(n_482), .C(n_494), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVxp67_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_SL g490 ( .A(n_491), .Y(n_490) );
AOI21xp33_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_496), .B(n_498), .Y(n_494) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
AOI22x1_ASAP7_75t_L g525 ( .A1(n_504), .A2(n_526), .B1(n_528), .B2(n_848), .Y(n_525) );
OAI21xp33_ASAP7_75t_L g518 ( .A1(n_505), .A2(n_519), .B(n_524), .Y(n_518) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_509), .B(n_510), .Y(n_508) );
INVx5_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
BUFx10_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_516), .Y(n_514) );
BUFx8_ASAP7_75t_SL g527 ( .A(n_515), .Y(n_527) );
CKINVDCx5p33_ASAP7_75t_R g850 ( .A(n_515), .Y(n_850) );
INVx1_ASAP7_75t_L g523 ( .A(n_517), .Y(n_523) );
INVx6_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
AND2x6_ASAP7_75t_SL g520 ( .A(n_521), .B(n_522), .Y(n_520) );
INVx1_ASAP7_75t_L g852 ( .A(n_525), .Y(n_852) );
CKINVDCx5p33_ASAP7_75t_R g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
NOR2x1p5_ASAP7_75t_L g529 ( .A(n_530), .B(n_756), .Y(n_529) );
NAND4xp75_ASAP7_75t_L g530 ( .A(n_531), .B(n_653), .C(n_687), .D(n_736), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_532), .A2(n_579), .B(n_612), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_541), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx2_ASAP7_75t_L g732 ( .A(n_535), .Y(n_732) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g617 ( .A(n_536), .B(n_543), .Y(n_617) );
AND2x4_ASAP7_75t_L g648 ( .A(n_536), .B(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g669 ( .A(n_536), .Y(n_669) );
OAI21x1_ASAP7_75t_L g546 ( .A1(n_540), .A2(n_547), .B(n_552), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g769 ( .A(n_541), .B(n_770), .Y(n_769) );
AND2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_557), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_542), .B(n_683), .Y(n_760) );
HB1xp67_ASAP7_75t_L g787 ( .A(n_542), .Y(n_787) );
OR2x2_ASAP7_75t_L g836 ( .A(n_542), .B(n_640), .Y(n_836) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g652 ( .A(n_543), .Y(n_652) );
INVx3_ASAP7_75t_L g660 ( .A(n_543), .Y(n_660) );
OR2x2_ASAP7_75t_L g668 ( .A(n_543), .B(n_669), .Y(n_668) );
OR2x2_ASAP7_75t_L g696 ( .A(n_543), .B(n_666), .Y(n_696) );
INVx1_ASAP7_75t_L g707 ( .A(n_543), .Y(n_707) );
AND2x2_ASAP7_75t_L g728 ( .A(n_543), .B(n_669), .Y(n_728) );
INVxp67_ASAP7_75t_L g752 ( .A(n_543), .Y(n_752) );
BUFx2_ASAP7_75t_L g796 ( .A(n_543), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_543), .B(n_558), .Y(n_805) );
AND2x2_ASAP7_75t_L g812 ( .A(n_543), .B(n_813), .Y(n_812) );
BUFx6f_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
OAI21x1_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_546), .B(n_556), .Y(n_544) );
OAI21xp5_ASAP7_75t_L g626 ( .A1(n_551), .A2(n_627), .B(n_629), .Y(n_626) );
AND2x2_ASAP7_75t_L g670 ( .A(n_557), .B(n_671), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g824 ( .A1(n_557), .A2(n_582), .B1(n_786), .B2(n_825), .Y(n_824) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_566), .Y(n_557) );
OR2x2_ASAP7_75t_L g640 ( .A(n_558), .B(n_641), .Y(n_640) );
INVx3_ASAP7_75t_L g649 ( .A(n_558), .Y(n_649) );
AND2x2_ASAP7_75t_L g661 ( .A(n_558), .B(n_641), .Y(n_661) );
AND2x2_ASAP7_75t_L g719 ( .A(n_558), .B(n_567), .Y(n_719) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g616 ( .A(n_567), .Y(n_616) );
INVx1_ASAP7_75t_L g710 ( .A(n_567), .Y(n_710) );
HB1xp67_ASAP7_75t_L g813 ( .A(n_567), .Y(n_813) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g666 ( .A(n_568), .Y(n_666) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_571), .B(n_574), .Y(n_570) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_594), .Y(n_580) );
AND2x2_ASAP7_75t_L g767 ( .A(n_581), .B(n_713), .Y(n_767) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
AOI32xp33_ASAP7_75t_L g797 ( .A1(n_582), .A2(n_690), .A3(n_764), .B1(n_798), .B2(n_800), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_582), .B(n_827), .Y(n_826) );
INVx2_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
OR2x2_ASAP7_75t_L g619 ( .A(n_583), .B(n_620), .Y(n_619) );
OR2x2_ASAP7_75t_L g636 ( .A(n_583), .B(n_596), .Y(n_636) );
BUFx2_ASAP7_75t_L g655 ( .A(n_583), .Y(n_655) );
INVx1_ASAP7_75t_L g702 ( .A(n_583), .Y(n_702) );
AND2x2_ASAP7_75t_L g735 ( .A(n_583), .B(n_714), .Y(n_735) );
OA21x2_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_585), .B(n_593), .Y(n_583) );
OA21x2_ASAP7_75t_L g681 ( .A1(n_584), .A2(n_585), .B(n_593), .Y(n_681) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
OR2x2_ASAP7_75t_L g618 ( .A(n_595), .B(n_619), .Y(n_618) );
OR2x2_ASAP7_75t_L g823 ( .A(n_595), .B(n_707), .Y(n_823) );
INVx1_ASAP7_75t_L g827 ( .A(n_595), .Y(n_827) );
OR2x2_ASAP7_75t_L g595 ( .A(n_596), .B(n_603), .Y(n_595) );
INVx2_ASAP7_75t_L g651 ( .A(n_596), .Y(n_651) );
AND2x2_ASAP7_75t_L g675 ( .A(n_596), .B(n_634), .Y(n_675) );
AND2x2_ASAP7_75t_L g686 ( .A(n_596), .B(n_681), .Y(n_686) );
INVx1_ASAP7_75t_L g693 ( .A(n_596), .Y(n_693) );
AND2x2_ASAP7_75t_L g701 ( .A(n_596), .B(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g714 ( .A(n_596), .Y(n_714) );
AND2x2_ASAP7_75t_L g780 ( .A(n_596), .B(n_603), .Y(n_780) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
OR2x2_ASAP7_75t_L g644 ( .A(n_604), .B(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g634 ( .A(n_605), .Y(n_634) );
CKINVDCx5p33_ASAP7_75t_R g610 ( .A(n_611), .Y(n_610) );
OAI221xp5_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_618), .B1(n_631), .B2(n_637), .C(n_642), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
OAI21xp5_ASAP7_75t_L g763 ( .A1(n_614), .A2(n_764), .B(n_767), .Y(n_763) );
AND2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_617), .Y(n_614) );
AND2x4_ASAP7_75t_L g839 ( .A(n_615), .B(n_639), .Y(n_839) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
AND2x4_ASAP7_75t_L g683 ( .A(n_616), .B(n_649), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_617), .B(n_718), .Y(n_717) );
BUFx2_ASAP7_75t_L g748 ( .A(n_617), .Y(n_748) );
OR2x2_ASAP7_75t_L g692 ( .A(n_619), .B(n_693), .Y(n_692) );
OR2x2_ASAP7_75t_L g754 ( .A(n_619), .B(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g825 ( .A(n_619), .Y(n_825) );
AND2x2_ASAP7_75t_L g633 ( .A(n_620), .B(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g782 ( .A(n_620), .B(n_681), .Y(n_782) );
OAI21xp5_ASAP7_75t_L g620 ( .A1(n_621), .A2(n_622), .B(n_630), .Y(n_620) );
OAI21x1_ASAP7_75t_L g645 ( .A1(n_621), .A2(n_622), .B(n_630), .Y(n_645) );
OAI221xp5_ASAP7_75t_L g662 ( .A1(n_631), .A2(n_663), .B1(n_664), .B2(n_673), .C(n_682), .Y(n_662) );
OAI221xp5_ASAP7_75t_L g758 ( .A1(n_631), .A2(n_746), .B1(n_759), .B2(n_761), .C(n_763), .Y(n_758) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_633), .B(n_635), .Y(n_632) );
AND2x2_ASAP7_75t_L g685 ( .A(n_633), .B(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g698 ( .A(n_634), .B(n_681), .Y(n_698) );
INVx2_ASAP7_75t_L g704 ( .A(n_634), .Y(n_704) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OAI221xp5_ASAP7_75t_L g768 ( .A1(n_637), .A2(n_769), .B1(n_774), .B2(n_778), .C(n_783), .Y(n_768) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OR2x2_ASAP7_75t_L g820 ( .A(n_640), .B(n_790), .Y(n_820) );
INVx1_ASAP7_75t_L g672 ( .A(n_641), .Y(n_672) );
INVx1_ASAP7_75t_L g709 ( .A(n_641), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_643), .B(n_646), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g658 ( .A(n_644), .Y(n_658) );
OR2x2_ASAP7_75t_L g721 ( .A(n_644), .B(n_657), .Y(n_721) );
INVx2_ASAP7_75t_L g734 ( .A(n_644), .Y(n_734) );
INVx2_ASAP7_75t_L g679 ( .A(n_645), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_647), .B(n_650), .Y(n_646) );
INVx3_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
BUFx2_ASAP7_75t_L g684 ( .A(n_648), .Y(n_684) );
AND2x4_ASAP7_75t_L g690 ( .A(n_648), .B(n_691), .Y(n_690) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_648), .B(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g764 ( .A(n_648), .B(n_765), .Y(n_764) );
AND2x2_ASAP7_75t_L g841 ( .A(n_648), .B(n_796), .Y(n_841) );
AND2x2_ASAP7_75t_L g665 ( .A(n_649), .B(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g727 ( .A(n_649), .Y(n_727) );
INVx1_ASAP7_75t_L g786 ( .A(n_649), .Y(n_786) );
OR2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_652), .Y(n_650) );
INVx2_ASAP7_75t_SL g657 ( .A(n_651), .Y(n_657) );
AND2x2_ASAP7_75t_L g699 ( .A(n_651), .B(n_678), .Y(n_699) );
AND2x2_ASAP7_75t_L g773 ( .A(n_652), .B(n_727), .Y(n_773) );
AOI21xp5_ASAP7_75t_L g653 ( .A1(n_654), .A2(n_659), .B(n_662), .Y(n_653) );
AND2x2_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .Y(n_654) );
INVx1_ASAP7_75t_L g739 ( .A(n_655), .Y(n_739) );
AND2x2_ASAP7_75t_L g806 ( .A(n_655), .B(n_734), .Y(n_806) );
AND2x2_ASAP7_75t_L g821 ( .A(n_655), .B(n_780), .Y(n_821) );
AND2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
INVx2_ASAP7_75t_L g775 ( .A(n_657), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_657), .B(n_782), .Y(n_792) );
OAI33xp33_ASAP7_75t_L g829 ( .A1(n_657), .A2(n_731), .A3(n_799), .B1(n_830), .B2(n_831), .B3(n_832), .Y(n_829) );
AND2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_660), .B(n_666), .Y(n_790) );
AND2x2_ASAP7_75t_L g818 ( .A(n_661), .B(n_766), .Y(n_818) );
AOI21xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_667), .B(n_670), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g691 ( .A(n_666), .Y(n_691) );
INVx1_ASAP7_75t_L g766 ( .A(n_666), .Y(n_766) );
OAI32xp33_ASAP7_75t_L g711 ( .A1(n_667), .A2(n_692), .A3(n_712), .B1(n_715), .B2(n_717), .Y(n_711) );
INVx2_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
OR2x2_ASAP7_75t_L g746 ( .A(n_668), .B(n_691), .Y(n_746) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g724 ( .A(n_672), .Y(n_724) );
INVx2_ASAP7_75t_L g772 ( .A(n_672), .Y(n_772) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
AND2x4_ASAP7_75t_L g674 ( .A(n_675), .B(n_676), .Y(n_674) );
INVx2_ASAP7_75t_L g755 ( .A(n_675), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_676), .B(n_713), .Y(n_712) );
AND2x2_ASAP7_75t_L g815 ( .A(n_676), .B(n_762), .Y(n_815) );
INVx2_ASAP7_75t_L g846 ( .A(n_676), .Y(n_846) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
OR2x2_ASAP7_75t_L g761 ( .A(n_677), .B(n_762), .Y(n_761) );
NAND2x1p5_ASAP7_75t_L g677 ( .A(n_678), .B(n_680), .Y(n_677) );
AND2x2_ASAP7_75t_L g703 ( .A(n_678), .B(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g745 ( .A(n_679), .Y(n_745) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
OAI21xp5_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_684), .B(n_685), .Y(n_682) );
INVx2_ASAP7_75t_L g753 ( .A(n_683), .Y(n_753) );
AND2x2_ASAP7_75t_L g737 ( .A(n_684), .B(n_738), .Y(n_737) );
NOR3x1_ASAP7_75t_L g687 ( .A(n_688), .B(n_711), .C(n_720), .Y(n_687) );
OAI21xp5_ASAP7_75t_SL g688 ( .A1(n_689), .A2(n_692), .B(n_694), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
NAND2xp5_ASAP7_75t_SL g832 ( .A(n_691), .B(n_833), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_693), .B(n_744), .Y(n_743) );
AOI22xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_697), .B1(n_700), .B2(n_705), .Y(n_694) );
INVx3_ASAP7_75t_L g729 ( .A(n_696), .Y(n_729) );
AND2x2_ASAP7_75t_L g697 ( .A(n_698), .B(n_699), .Y(n_697) );
INVxp67_ASAP7_75t_L g742 ( .A(n_698), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_698), .B(n_777), .Y(n_776) );
AND2x4_ASAP7_75t_L g700 ( .A(n_701), .B(n_703), .Y(n_700) );
AND2x2_ASAP7_75t_L g843 ( .A(n_701), .B(n_734), .Y(n_843) );
AND2x2_ASAP7_75t_L g713 ( .A(n_704), .B(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g762 ( .A(n_704), .Y(n_762) );
INVx1_ASAP7_75t_L g799 ( .A(n_704), .Y(n_799) );
NOR2xp33_ASAP7_75t_L g833 ( .A(n_704), .B(n_745), .Y(n_833) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
NAND2x1p5_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
INVx1_ASAP7_75t_L g830 ( .A(n_708), .Y(n_830) );
AND2x2_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
INVx1_ASAP7_75t_L g716 ( .A(n_710), .Y(n_716) );
AND2x2_ASAP7_75t_L g842 ( .A(n_713), .B(n_782), .Y(n_842) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
BUFx2_ASAP7_75t_L g750 ( .A(n_719), .Y(n_750) );
AND2x2_ASAP7_75t_L g847 ( .A(n_719), .B(n_728), .Y(n_847) );
OAI22xp33_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_722), .B1(n_730), .B2(n_733), .Y(n_720) );
AOI211xp5_ASAP7_75t_SL g722 ( .A1(n_723), .A2(n_725), .B(n_728), .C(n_729), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
OR2x2_ASAP7_75t_L g804 ( .A(n_724), .B(n_805), .Y(n_804) );
INVxp67_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVxp33_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_734), .B(n_735), .Y(n_733) );
AND2x2_ASAP7_75t_L g738 ( .A(n_734), .B(n_739), .Y(n_738) );
AND2x2_ASAP7_75t_L g816 ( .A(n_735), .B(n_777), .Y(n_816) );
INVx1_ASAP7_75t_L g831 ( .A(n_735), .Y(n_831) );
NOR3xp33_ASAP7_75t_L g736 ( .A(n_737), .B(n_740), .C(n_747), .Y(n_736) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_741), .B(n_746), .Y(n_740) );
OR2x2_ASAP7_75t_L g741 ( .A(n_742), .B(n_743), .Y(n_741) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx2_ASAP7_75t_L g777 ( .A(n_745), .Y(n_777) );
O2A1O1Ixp33_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_749), .B(n_751), .C(n_754), .Y(n_747) );
AOI22xp5_ASAP7_75t_L g840 ( .A1(n_748), .A2(n_841), .B1(n_842), .B2(n_843), .Y(n_840) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
OR2x2_ASAP7_75t_L g751 ( .A(n_752), .B(n_753), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_757), .B(n_808), .Y(n_756) );
NOR3xp33_ASAP7_75t_SL g757 ( .A(n_758), .B(n_768), .C(n_793), .Y(n_757) );
HB1xp67_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
AOI22xp5_ASAP7_75t_L g802 ( .A1(n_764), .A2(n_803), .B1(n_806), .B2(n_807), .Y(n_802) );
INVx1_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
AND2x2_ASAP7_75t_L g770 ( .A(n_771), .B(n_773), .Y(n_770) );
AND2x2_ASAP7_75t_L g788 ( .A(n_771), .B(n_789), .Y(n_788) );
AND2x4_ASAP7_75t_L g811 ( .A(n_771), .B(n_812), .Y(n_811) );
INVx2_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
OR2x2_ASAP7_75t_L g774 ( .A(n_775), .B(n_776), .Y(n_774) );
INVx1_ASAP7_75t_L g807 ( .A(n_776), .Y(n_807) );
OR2x2_ASAP7_75t_L g778 ( .A(n_779), .B(n_781), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_782), .B(n_799), .Y(n_801) );
OAI21xp5_ASAP7_75t_L g783 ( .A1(n_784), .A2(n_788), .B(n_791), .Y(n_783) );
AND2x2_ASAP7_75t_L g784 ( .A(n_785), .B(n_787), .Y(n_784) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
AOI22xp5_ASAP7_75t_L g844 ( .A1(n_788), .A2(n_843), .B1(n_845), .B2(n_847), .Y(n_844) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
OAI21xp33_ASAP7_75t_SL g793 ( .A1(n_794), .A2(n_797), .B(n_802), .Y(n_793) );
INVx1_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_795), .B(n_839), .Y(n_838) );
BUFx2_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g800 ( .A(n_801), .Y(n_800) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g834 ( .A(n_805), .Y(n_834) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_807), .A2(n_829), .B1(n_834), .B2(n_835), .Y(n_828) );
NOR2xp33_ASAP7_75t_L g808 ( .A(n_809), .B(n_837), .Y(n_808) );
OAI211xp5_ASAP7_75t_SL g809 ( .A1(n_810), .A2(n_814), .B(n_817), .C(n_828), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
NOR2x1_ASAP7_75t_L g814 ( .A(n_815), .B(n_816), .Y(n_814) );
O2A1O1Ixp5_ASAP7_75t_L g817 ( .A1(n_818), .A2(n_819), .B(n_821), .C(n_822), .Y(n_817) );
INVx1_ASAP7_75t_L g819 ( .A(n_820), .Y(n_819) );
OAI22xp5_ASAP7_75t_L g822 ( .A1(n_820), .A2(n_823), .B1(n_824), .B2(n_826), .Y(n_822) );
OAI211xp5_ASAP7_75t_L g837 ( .A1(n_831), .A2(n_838), .B(n_840), .C(n_844), .Y(n_837) );
INVx2_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx8_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
BUFx12f_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
BUFx6f_ASAP7_75t_L g862 ( .A(n_853), .Y(n_862) );
AND2x2_ASAP7_75t_SL g853 ( .A(n_854), .B(n_858), .Y(n_853) );
INVx2_ASAP7_75t_SL g855 ( .A(n_856), .Y(n_855) );
CKINVDCx5p33_ASAP7_75t_R g858 ( .A(n_859), .Y(n_858) );
NOR2xp33_ASAP7_75t_L g860 ( .A(n_861), .B(n_862), .Y(n_860) );
endmodule