module fake_jpeg_19705_n_328 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_328);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx4f_ASAP7_75t_SL g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_9),
.B(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_5),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_42),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_17),
.B(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_27),
.B(n_0),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_43),
.Y(n_46)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_41),
.A2(n_31),
.B1(n_33),
.B2(n_18),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_53),
.A2(n_24),
.B1(n_29),
.B2(n_32),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_31),
.B1(n_33),
.B2(n_18),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_55),
.A2(n_43),
.B1(n_24),
.B2(n_29),
.Y(n_85)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_60),
.B(n_36),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_62),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_64),
.B(n_66),
.Y(n_124)
);

BUFx2_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_48),
.B(n_42),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_35),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_68),
.B(n_70),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_27),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_60),
.B(n_26),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_71),
.B(n_73),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_26),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_63),
.A2(n_33),
.B1(n_44),
.B2(n_38),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_74),
.A2(n_85),
.B1(n_46),
.B2(n_20),
.Y(n_119)
);

BUFx6f_ASAP7_75t_SL g75 ( 
.A(n_47),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_75),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_39),
.Y(n_77)
);

FAx1_ASAP7_75t_SL g108 ( 
.A(n_77),
.B(n_19),
.CI(n_34),
.CON(n_108),
.SN(n_108)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_50),
.A2(n_44),
.B1(n_38),
.B2(n_43),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_78),
.A2(n_91),
.B1(n_57),
.B2(n_32),
.Y(n_107)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_79),
.B(n_83),
.Y(n_121)
);

BUFx6f_ASAP7_75t_SL g82 ( 
.A(n_47),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_82),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_51),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_88),
.Y(n_100)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_92),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_90),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_45),
.B(n_17),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_45),
.Y(n_93)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_49),
.B(n_20),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_59),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_34),
.Y(n_98)
);

XNOR2x1_ASAP7_75t_L g150 ( 
.A(n_98),
.B(n_108),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_101),
.Y(n_131)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_69),
.B(n_39),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_103),
.A2(n_110),
.B(n_120),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_91),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_106),
.B(n_109),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_107),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_77),
.B(n_40),
.C(n_30),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_89),
.A2(n_39),
.B(n_2),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_65),
.Y(n_114)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_114),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_40),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_116),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_67),
.B(n_21),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_67),
.B(n_21),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_118),
.B(n_82),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_119),
.A2(n_123),
.B1(n_86),
.B2(n_95),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_25),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_86),
.A2(n_21),
.B1(n_28),
.B2(n_20),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_125),
.A2(n_148),
.B1(n_103),
.B2(n_120),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_100),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_126),
.B(n_127),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_117),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_129),
.B(n_136),
.Y(n_171)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_96),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_132),
.B(n_143),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_104),
.Y(n_133)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

O2A1O1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_106),
.A2(n_87),
.B(n_80),
.C(n_75),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_134),
.A2(n_142),
.B(n_152),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_121),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_137),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_110),
.A2(n_19),
.B(n_25),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_138),
.A2(n_147),
.B(n_131),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_113),
.B(n_88),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_139),
.Y(n_170)
);

AND2x2_ASAP7_75t_SL g142 ( 
.A(n_116),
.B(n_90),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_144),
.Y(n_159)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_146),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_120),
.A2(n_25),
.B(n_20),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_119),
.A2(n_107),
.B1(n_101),
.B2(n_105),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_109),
.A2(n_84),
.B1(n_23),
.B2(n_22),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_149),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_113),
.B(n_30),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_112),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_101),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_97),
.Y(n_153)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_96),
.Y(n_154)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_154),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_98),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_157),
.B(n_163),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_160),
.A2(n_172),
.B1(n_141),
.B2(n_132),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_161),
.B(n_169),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_140),
.B(n_105),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_176),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_128),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_165),
.A2(n_166),
.B(n_23),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_135),
.A2(n_131),
.B(n_152),
.Y(n_166)
);

OAI21xp33_ASAP7_75t_L g167 ( 
.A1(n_128),
.A2(n_124),
.B(n_108),
.Y(n_167)
);

OAI21xp33_ASAP7_75t_L g206 ( 
.A1(n_167),
.A2(n_12),
.B(n_14),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_130),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_129),
.A2(n_104),
.B1(n_111),
.B2(n_112),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_108),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_173),
.B(n_149),
.C(n_147),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_126),
.B(n_124),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_174),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_144),
.B(n_102),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_175),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_140),
.B(n_103),
.Y(n_176)
);

AO21x1_ASAP7_75t_L g178 ( 
.A1(n_138),
.A2(n_123),
.B(n_102),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_178),
.A2(n_142),
.B(n_134),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_145),
.A2(n_114),
.B1(n_97),
.B2(n_99),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_179),
.A2(n_185),
.B1(n_187),
.B2(n_143),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_137),
.B(n_30),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_180),
.B(n_182),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_146),
.B(n_30),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_130),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_122),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_145),
.A2(n_99),
.B1(n_28),
.B2(n_22),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_136),
.B(n_148),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_133),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_125),
.A2(n_28),
.B1(n_22),
.B2(n_30),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_190),
.B(n_206),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_186),
.A2(n_160),
.B1(n_181),
.B2(n_156),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_191),
.A2(n_194),
.B1(n_198),
.B2(n_207),
.Y(n_226)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_192),
.Y(n_240)
);

XOR2x2_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_142),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_193),
.B(n_209),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_156),
.A2(n_142),
.B1(n_153),
.B2(n_141),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_171),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_203),
.Y(n_219)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_158),
.Y(n_196)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_196),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_197),
.A2(n_216),
.B1(n_218),
.B2(n_180),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_157),
.B(n_81),
.C(n_76),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_210),
.C(n_215),
.Y(n_228)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_188),
.Y(n_204)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_204),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_164),
.A2(n_133),
.B1(n_154),
.B2(n_122),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_173),
.B(n_81),
.C(n_76),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_166),
.A2(n_23),
.B(n_8),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_211),
.B(n_214),
.Y(n_223)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_212),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_181),
.A2(n_7),
.B1(n_13),
.B2(n_12),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_213),
.A2(n_155),
.B1(n_182),
.B2(n_188),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_162),
.B(n_159),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_165),
.B(n_28),
.C(n_7),
.Y(n_215)
);

OAI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_170),
.A2(n_13),
.B1(n_11),
.B2(n_10),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_184),
.Y(n_217)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_217),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_170),
.A2(n_13),
.B1(n_10),
.B2(n_8),
.Y(n_218)
);

NOR3xp33_ASAP7_75t_L g224 ( 
.A(n_195),
.B(n_159),
.C(n_183),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_224),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_214),
.B(n_164),
.Y(n_225)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_225),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_177),
.C(n_176),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_238),
.C(n_190),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_208),
.B(n_201),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_242),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_189),
.B(n_169),
.Y(n_231)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_231),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_189),
.B(n_168),
.Y(n_233)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_233),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_234),
.A2(n_237),
.B1(n_241),
.B2(n_243),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_205),
.Y(n_235)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_235),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_177),
.C(n_184),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_217),
.Y(n_239)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_239),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_199),
.A2(n_178),
.B1(n_179),
.B2(n_155),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_193),
.B(n_178),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_203),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_223),
.A2(n_226),
.B1(n_197),
.B2(n_233),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_245),
.A2(n_246),
.B1(n_10),
.B2(n_7),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_223),
.A2(n_213),
.B1(n_200),
.B2(n_192),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_219),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_247),
.B(n_255),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_253),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_230),
.B(n_209),
.C(n_191),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_221),
.C(n_220),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_202),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_242),
.B(n_202),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_260),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_228),
.B(n_196),
.C(n_215),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_219),
.Y(n_259)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_259),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_238),
.B(n_211),
.Y(n_260)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_231),
.Y(n_262)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_262),
.Y(n_266)
);

A2O1A1Ixp33_ASAP7_75t_SL g263 ( 
.A1(n_240),
.A2(n_194),
.B(n_207),
.C(n_204),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_263),
.A2(n_226),
.B1(n_236),
.B2(n_225),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_228),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_265),
.B(n_268),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_221),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_257),
.A2(n_222),
.B(n_232),
.Y(n_269)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_269),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_244),
.B(n_232),
.Y(n_270)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_270),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_256),
.B(n_220),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_271),
.Y(n_282)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_272),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_273),
.B(n_275),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_237),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_253),
.B(n_248),
.C(n_260),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_276),
.B(n_280),
.C(n_263),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_261),
.A2(n_236),
.B1(n_227),
.B2(n_243),
.Y(n_278)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_278),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_279),
.A2(n_252),
.B1(n_249),
.B2(n_247),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_1),
.C(n_2),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_258),
.Y(n_281)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_281),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_284),
.A2(n_285),
.B1(n_4),
.B2(n_5),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_266),
.A2(n_263),
.B1(n_3),
.B2(n_4),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_275),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_280),
.Y(n_289)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_289),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_274),
.B(n_263),
.C(n_4),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_291),
.B(n_294),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_264),
.B(n_2),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_286),
.A2(n_265),
.B(n_273),
.Y(n_295)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_295),
.Y(n_315)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_288),
.A2(n_276),
.B(n_274),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_299),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_283),
.C(n_292),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_268),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_301),
.B(n_302),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_277),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_283),
.B(n_277),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_304),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_4),
.Y(n_304)
);

OAI21xp33_ASAP7_75t_L g306 ( 
.A1(n_282),
.A2(n_6),
.B(n_290),
.Y(n_306)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_306),
.B(n_294),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_287),
.Y(n_307)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_307),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_301),
.C(n_302),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_312),
.Y(n_318)
);

INVx6_ASAP7_75t_L g312 ( 
.A(n_305),
.Y(n_312)
);

NOR2xp67_ASAP7_75t_L g313 ( 
.A(n_306),
.B(n_284),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_313),
.B(n_304),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_316),
.B(n_317),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_297),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_319),
.A2(n_314),
.B(n_315),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_321),
.B(n_316),
.C(n_320),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_322),
.C(n_318),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_324),
.A2(n_312),
.B(n_309),
.Y(n_325)
);

MAJx2_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_310),
.C(n_308),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_6),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_6),
.B(n_318),
.Y(n_328)
);


endmodule