module fake_jpeg_2611_n_134 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_134);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_134;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_22),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_31),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_5),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_19),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_52),
.Y(n_69)
);

OAI21xp33_ASAP7_75t_L g53 ( 
.A1(n_46),
.A2(n_39),
.B(n_43),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_53),
.B(n_54),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_42),
.B(n_0),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

OAI21xp33_ASAP7_75t_L g56 ( 
.A1(n_46),
.A2(n_0),
.B(n_1),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_57),
.Y(n_67)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_43),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g68 ( 
.A1(n_58),
.A2(n_47),
.B1(n_49),
.B2(n_41),
.Y(n_68)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_62),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_57),
.A2(n_45),
.B1(n_39),
.B2(n_49),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_63),
.A2(n_60),
.B1(n_67),
.B2(n_38),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_54),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_64),
.B(n_44),
.Y(n_70)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_68),
.A2(n_51),
.B1(n_50),
.B2(n_44),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_72),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_61),
.B(n_40),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_74),
.B(n_78),
.Y(n_84)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_68),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_61),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_69),
.A2(n_50),
.B(n_42),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_SL g94 ( 
.A(n_79),
.B(n_68),
.Y(n_94)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_79),
.B(n_41),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_83),
.B(n_85),
.Y(n_105)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_82),
.B(n_40),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_89),
.Y(n_108)
);

OAI32xp33_ASAP7_75t_L g88 ( 
.A1(n_77),
.A2(n_68),
.A3(n_75),
.B1(n_76),
.B2(n_65),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_90),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_71),
.B(n_48),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_73),
.B(n_66),
.Y(n_91)
);

NAND3xp33_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_7),
.C(n_8),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_94),
.B(n_73),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_99),
.Y(n_110)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_97),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_90),
.A2(n_47),
.B1(n_51),
.B2(n_5),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_98),
.B(n_100),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_14),
.C(n_29),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_88),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_93),
.A2(n_4),
.B(n_7),
.C(n_8),
.Y(n_101)
);

A2O1A1Ixp33_ASAP7_75t_SL g112 ( 
.A1(n_101),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_112)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_9),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_103),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g104 ( 
.A(n_95),
.B(n_21),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_109),
.C(n_99),
.Y(n_119)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_106),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_9),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_116),
.Y(n_120)
);

NOR2xp67_ASAP7_75t_L g116 ( 
.A(n_105),
.B(n_23),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_108),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_117),
.A2(n_107),
.B(n_102),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_119),
.B(n_104),
.C(n_101),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g121 ( 
.A(n_110),
.B(n_107),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_121),
.B(n_122),
.Y(n_127)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_123),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_114),
.A2(n_24),
.B(n_28),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_124),
.A2(n_115),
.B1(n_112),
.B2(n_32),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_26),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_126),
.A2(n_120),
.B(n_111),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_128),
.A2(n_129),
.B1(n_112),
.B2(n_113),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_118),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_131),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_132),
.A2(n_127),
.B(n_110),
.Y(n_133)
);

AOI221xp5_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_118),
.B1(n_13),
.B2(n_16),
.C(n_27),
.Y(n_134)
);


endmodule