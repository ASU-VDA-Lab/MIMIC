module fake_jpeg_6041_n_58 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_58);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_58;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx2_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_5),
.B(n_4),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_13),
.B(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_17),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_18),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_15),
.B(n_2),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_20),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_14),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_7),
.C(n_9),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_8),
.B(n_3),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g31 ( 
.A1(n_22),
.A2(n_25),
.B(n_6),
.Y(n_31)
);

NOR2x1_ASAP7_75t_L g23 ( 
.A(n_10),
.B(n_3),
.Y(n_23)
);

NOR2x1_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_10),
.Y(n_29)
);

AND2x6_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_5),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_24),
.A2(n_16),
.B(n_8),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_11),
.B(n_6),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_27),
.A2(n_35),
.B1(n_25),
.B2(n_20),
.Y(n_38)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_19),
.Y(n_36)
);

AO21x1_ASAP7_75t_L g40 ( 
.A1(n_29),
.A2(n_31),
.B(n_10),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_SL g30 ( 
.A1(n_24),
.A2(n_16),
.B(n_9),
.C(n_10),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_30),
.A2(n_22),
.B(n_21),
.Y(n_37)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_12),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_38),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_39),
.Y(n_44)
);

AO21x1_ASAP7_75t_L g42 ( 
.A1(n_28),
.A2(n_12),
.B(n_31),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_27),
.B(n_35),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_43),
.B(n_34),
.C(n_32),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_48),
.Y(n_52)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_39),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_34),
.C(n_30),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g54 ( 
.A1(n_50),
.A2(n_51),
.B(n_53),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_47),
.A2(n_30),
.B1(n_33),
.B2(n_42),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_26),
.Y(n_53)
);

NOR2xp67_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_48),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g57 ( 
.A1(n_55),
.A2(n_56),
.B(n_30),
.Y(n_57)
);

A2O1A1O1Ixp25_ASAP7_75t_L g56 ( 
.A1(n_50),
.A2(n_45),
.B(n_46),
.C(n_40),
.D(n_44),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_54),
.Y(n_58)
);


endmodule