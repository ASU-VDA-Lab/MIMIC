module fake_jpeg_12684_n_69 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_69);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_69;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_67;
wire n_66;

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_4),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_7),
.B(n_5),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_12),
.B(n_23),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_28),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_33),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_0),
.Y(n_33)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_25),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_34),
.B(n_35),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_1),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_36),
.A2(n_26),
.B(n_25),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_1),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_2),
.Y(n_46)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_31),
.C(n_24),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_44),
.C(n_43),
.Y(n_52)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_42),
.B(n_46),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_14),
.C(n_20),
.Y(n_44)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_13),
.B1(n_19),
.B2(n_18),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_50),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_47),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_52),
.A2(n_3),
.B(n_6),
.Y(n_58)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_53),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_44),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_52),
.Y(n_63)
);

O2A1O1Ixp33_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_56),
.B(n_48),
.C(n_54),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_63),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_64),
.B(n_57),
.C(n_59),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_61),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

A2O1A1O1Ixp25_ASAP7_75t_L g68 ( 
.A1(n_67),
.A2(n_55),
.B(n_11),
.C(n_15),
.D(n_16),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_68),
.A2(n_9),
.B(n_17),
.Y(n_69)
);


endmodule