module fake_netlist_6_4050_n_1843 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1843);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1843;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_236;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g186 ( 
.A(n_128),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_126),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_96),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_115),
.Y(n_189)
);

BUFx8_ASAP7_75t_SL g190 ( 
.A(n_166),
.Y(n_190)
);

BUFx10_ASAP7_75t_L g191 ( 
.A(n_6),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_170),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_23),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_12),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_179),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_64),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_155),
.Y(n_197)
);

BUFx10_ASAP7_75t_L g198 ( 
.A(n_124),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_52),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_130),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_32),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_56),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_72),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_26),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_178),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_135),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_121),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_80),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_88),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_149),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_46),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_136),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_117),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_10),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_41),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_181),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_140),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_12),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_54),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_46),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_78),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_169),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_11),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_141),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_24),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_61),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_35),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_22),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_185),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_68),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_120),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_113),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_70),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_142),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_83),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_8),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_26),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_160),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_37),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_125),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_165),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_77),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_73),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_98),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_29),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_97),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_60),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_184),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_17),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_74),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_139),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_145),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_47),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_32),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_15),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_13),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_87),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_131),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_19),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_23),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_38),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_175),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_48),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_101),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_109),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_65),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_52),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_7),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_0),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_0),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_150),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_156),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_8),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_114),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_34),
.Y(n_275)
);

BUFx10_ASAP7_75t_L g276 ( 
.A(n_81),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_91),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_40),
.Y(n_278)
);

BUFx2_ASAP7_75t_L g279 ( 
.A(n_174),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_9),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_90),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_63),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_108),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_29),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_92),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_66),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_38),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_75),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_148),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_99),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_106),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_40),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_45),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_5),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_89),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_47),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_62),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_162),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_11),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_173),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_82),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_25),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_102),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_84),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_27),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_144),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_50),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_55),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_79),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_48),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_104),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_20),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_58),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_133),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_105),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_107),
.Y(n_316)
);

BUFx10_ASAP7_75t_L g317 ( 
.A(n_182),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_183),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_111),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_119),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_159),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_2),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_44),
.Y(n_323)
);

BUFx10_ASAP7_75t_L g324 ( 
.A(n_122),
.Y(n_324)
);

BUFx5_ASAP7_75t_L g325 ( 
.A(n_36),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_176),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_51),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_158),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_137),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_134),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_147),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_24),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_100),
.Y(n_333)
);

INVx2_ASAP7_75t_SL g334 ( 
.A(n_21),
.Y(n_334)
);

BUFx10_ASAP7_75t_L g335 ( 
.A(n_34),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_95),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_118),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_6),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_127),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_54),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_4),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_2),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_27),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_16),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_154),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_9),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_44),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_56),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_19),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_85),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_152),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_171),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_13),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_22),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_172),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_20),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_36),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_61),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_58),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_163),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_31),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_123),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_93),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_57),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_116),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g366 ( 
.A(n_10),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_7),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_325),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_197),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_325),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_190),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_325),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_325),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_325),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_325),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_229),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_191),
.Y(n_377)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_291),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_325),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_325),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_239),
.Y(n_381)
);

CKINVDCx14_ASAP7_75t_R g382 ( 
.A(n_260),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_208),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_239),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_239),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_230),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_231),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_233),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_239),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_239),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_209),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_268),
.Y(n_392)
);

INVxp67_ASAP7_75t_SL g393 ( 
.A(n_189),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_312),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_235),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_312),
.Y(n_396)
);

INVxp33_ASAP7_75t_L g397 ( 
.A(n_194),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_312),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_238),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_312),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_242),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_244),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_248),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_312),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_367),
.Y(n_405)
);

INVxp67_ASAP7_75t_SL g406 ( 
.A(n_283),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_247),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_191),
.Y(n_408)
);

INVxp67_ASAP7_75t_SL g409 ( 
.A(n_210),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_247),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_251),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_366),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_258),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_367),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_366),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_240),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_191),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_262),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_266),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_199),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_220),
.Y(n_421)
);

INVxp67_ASAP7_75t_SL g422 ( 
.A(n_224),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_249),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_253),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_271),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_272),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_254),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_255),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_256),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_273),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_275),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_292),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_294),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_299),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_305),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_340),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_282),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_349),
.Y(n_438)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_335),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_285),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_264),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_354),
.Y(n_442)
);

INVxp33_ASAP7_75t_SL g443 ( 
.A(n_201),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_357),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_359),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_193),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_193),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_334),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_334),
.Y(n_449)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_335),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_257),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_257),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_274),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_316),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_316),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_337),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_243),
.Y(n_457)
);

INVx2_ASAP7_75t_SL g458 ( 
.A(n_335),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_286),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_289),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_243),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_374),
.Y(n_462)
);

INVx2_ASAP7_75t_SL g463 ( 
.A(n_394),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_381),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_457),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_457),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_409),
.B(n_279),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_381),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_461),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_376),
.Y(n_470)
);

NAND3xp33_ASAP7_75t_L g471 ( 
.A(n_407),
.B(n_364),
.C(n_227),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_414),
.B(n_200),
.Y(n_472)
);

INVx6_ASAP7_75t_L g473 ( 
.A(n_392),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_414),
.B(n_200),
.Y(n_474)
);

BUFx2_ASAP7_75t_L g475 ( 
.A(n_382),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_384),
.B(n_187),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_384),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_385),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_461),
.Y(n_479)
);

NOR3xp33_ASAP7_75t_L g480 ( 
.A(n_393),
.B(n_284),
.C(n_226),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_385),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_386),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_383),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_374),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_369),
.B(n_201),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_389),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_389),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_390),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_394),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_410),
.B(n_328),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_390),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_396),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_396),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_368),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_398),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_398),
.B(n_187),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_400),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_400),
.B(n_188),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_404),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_368),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_404),
.B(n_188),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_370),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_370),
.B(n_192),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_372),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_372),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g506 ( 
.A(n_378),
.B(n_198),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_373),
.Y(n_507)
);

OAI21x1_ASAP7_75t_L g508 ( 
.A1(n_373),
.A2(n_379),
.B(n_375),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_375),
.B(n_379),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_380),
.B(n_192),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_380),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_451),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_451),
.B(n_195),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g514 ( 
.A(n_391),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_420),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_452),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_420),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_452),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_424),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_454),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_424),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_454),
.B(n_195),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_412),
.B(n_328),
.Y(n_523)
);

INVx3_ASAP7_75t_L g524 ( 
.A(n_455),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_455),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_405),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_405),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_428),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_428),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_458),
.B(n_198),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_429),
.Y(n_531)
);

BUFx2_ASAP7_75t_L g532 ( 
.A(n_377),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_429),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_415),
.B(n_203),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_430),
.Y(n_535)
);

AND3x2_ASAP7_75t_L g536 ( 
.A(n_408),
.B(n_365),
.C(n_306),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_430),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_387),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_421),
.B(n_203),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_416),
.A2(n_327),
.B1(n_263),
.B2(n_313),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_490),
.B(n_406),
.Y(n_541)
);

NAND3xp33_ASAP7_75t_L g542 ( 
.A(n_503),
.B(n_427),
.C(n_423),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_507),
.Y(n_543)
);

INVx2_ASAP7_75t_SL g544 ( 
.A(n_473),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_489),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_470),
.Y(n_546)
);

INVx5_ASAP7_75t_L g547 ( 
.A(n_484),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_484),
.Y(n_548)
);

INVx4_ASAP7_75t_L g549 ( 
.A(n_484),
.Y(n_549)
);

NAND2xp33_ASAP7_75t_SL g550 ( 
.A(n_530),
.B(n_458),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_503),
.B(n_388),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_507),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_494),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_489),
.Y(n_554)
);

INVx2_ASAP7_75t_SL g555 ( 
.A(n_473),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_472),
.Y(n_556)
);

INVxp67_ASAP7_75t_SL g557 ( 
.A(n_508),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_494),
.Y(n_558)
);

BUFx3_ASAP7_75t_L g559 ( 
.A(n_472),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_489),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_530),
.B(n_395),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_494),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_500),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_465),
.Y(n_564)
);

BUFx3_ASAP7_75t_L g565 ( 
.A(n_474),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_484),
.Y(n_566)
);

INVx2_ASAP7_75t_SL g567 ( 
.A(n_473),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_465),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_465),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_484),
.Y(n_570)
);

BUFx2_ASAP7_75t_L g571 ( 
.A(n_532),
.Y(n_571)
);

NAND2xp33_ASAP7_75t_L g572 ( 
.A(n_510),
.B(n_399),
.Y(n_572)
);

INVx1_ASAP7_75t_SL g573 ( 
.A(n_483),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_467),
.B(n_401),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_467),
.B(n_402),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_484),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_L g577 ( 
.A1(n_510),
.A2(n_422),
.B1(n_443),
.B2(n_365),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_502),
.B(n_403),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_470),
.B(n_411),
.Y(n_579)
);

OR2x6_ASAP7_75t_L g580 ( 
.A(n_473),
.B(n_221),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_466),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_466),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_466),
.Y(n_583)
);

OR2x2_ASAP7_75t_L g584 ( 
.A(n_476),
.B(n_496),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_500),
.Y(n_585)
);

NAND2xp33_ASAP7_75t_L g586 ( 
.A(n_534),
.B(n_413),
.Y(n_586)
);

AO21x2_ASAP7_75t_L g587 ( 
.A1(n_508),
.A2(n_196),
.B(n_186),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_L g588 ( 
.A1(n_508),
.A2(n_397),
.B1(n_243),
.B2(n_431),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_502),
.B(n_418),
.Y(n_589)
);

INVx2_ASAP7_75t_SL g590 ( 
.A(n_473),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_469),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_502),
.B(n_419),
.Y(n_592)
);

INVx4_ASAP7_75t_SL g593 ( 
.A(n_484),
.Y(n_593)
);

OAI21xp33_ASAP7_75t_SL g594 ( 
.A1(n_506),
.A2(n_447),
.B(n_446),
.Y(n_594)
);

AOI22xp33_ASAP7_75t_L g595 ( 
.A1(n_490),
.A2(n_243),
.B1(n_431),
.B2(n_432),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_500),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_504),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_502),
.B(n_425),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_469),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_504),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_469),
.Y(n_601)
);

NAND3xp33_ASAP7_75t_L g602 ( 
.A(n_509),
.B(n_433),
.C(n_432),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_473),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_504),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_479),
.Y(n_605)
);

INVx4_ASAP7_75t_L g606 ( 
.A(n_535),
.Y(n_606)
);

BUFx2_ASAP7_75t_L g607 ( 
.A(n_532),
.Y(n_607)
);

NAND2xp33_ASAP7_75t_SL g608 ( 
.A(n_532),
.B(n_506),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_R g609 ( 
.A(n_482),
.B(n_371),
.Y(n_609)
);

AND2x4_ASAP7_75t_L g610 ( 
.A(n_474),
.B(n_490),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_479),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_482),
.B(n_426),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_505),
.Y(n_613)
);

NAND3xp33_ASAP7_75t_L g614 ( 
.A(n_509),
.B(n_434),
.C(n_433),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_479),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_505),
.Y(n_616)
);

INVx1_ASAP7_75t_SL g617 ( 
.A(n_483),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_463),
.Y(n_618)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_535),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_463),
.Y(n_620)
);

AND2x4_ASAP7_75t_L g621 ( 
.A(n_474),
.B(n_206),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_505),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_502),
.Y(n_623)
);

OR2x2_ASAP7_75t_L g624 ( 
.A(n_476),
.B(n_417),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_511),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_463),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_462),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_538),
.B(n_437),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_538),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_511),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_511),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_462),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_485),
.B(n_440),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_462),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_534),
.B(n_459),
.Y(n_635)
);

NAND2xp33_ASAP7_75t_SL g636 ( 
.A(n_475),
.B(n_308),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_464),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_523),
.B(n_446),
.Y(n_638)
);

BUFx4f_ASAP7_75t_L g639 ( 
.A(n_535),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_485),
.B(n_460),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_464),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_514),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_468),
.Y(n_643)
);

BUFx10_ASAP7_75t_L g644 ( 
.A(n_536),
.Y(n_644)
);

AOI22xp5_ASAP7_75t_L g645 ( 
.A1(n_480),
.A2(n_353),
.B1(n_218),
.B2(n_215),
.Y(n_645)
);

AO22x2_ASAP7_75t_L g646 ( 
.A1(n_480),
.A2(n_265),
.B1(n_216),
.B2(n_232),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_462),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_468),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_462),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_477),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_516),
.Y(n_651)
);

BUFx4f_ASAP7_75t_L g652 ( 
.A(n_535),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_477),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_478),
.Y(n_654)
);

INVx4_ASAP7_75t_L g655 ( 
.A(n_535),
.Y(n_655)
);

BUFx6f_ASAP7_75t_SL g656 ( 
.A(n_528),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_475),
.B(n_439),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_516),
.Y(n_658)
);

INVx4_ASAP7_75t_L g659 ( 
.A(n_535),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_523),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_539),
.B(n_450),
.Y(n_661)
);

BUFx3_ASAP7_75t_L g662 ( 
.A(n_523),
.Y(n_662)
);

BUFx6f_ASAP7_75t_SL g663 ( 
.A(n_528),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_496),
.B(n_205),
.Y(n_664)
);

INVx4_ASAP7_75t_L g665 ( 
.A(n_535),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_478),
.Y(n_666)
);

OR2x6_ASAP7_75t_L g667 ( 
.A(n_471),
.B(n_241),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_475),
.B(n_198),
.Y(n_668)
);

BUFx10_ASAP7_75t_L g669 ( 
.A(n_536),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_498),
.B(n_303),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_498),
.B(n_329),
.Y(n_671)
);

INVxp33_ASAP7_75t_L g672 ( 
.A(n_540),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_525),
.B(n_447),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_481),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_481),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_486),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_486),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_501),
.B(n_350),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_487),
.Y(n_679)
);

AOI22xp33_ASAP7_75t_L g680 ( 
.A1(n_513),
.A2(n_522),
.B1(n_501),
.B2(n_529),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_487),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_488),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_513),
.A2(n_243),
.B1(n_434),
.B2(n_435),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_488),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_516),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_491),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_491),
.Y(n_687)
);

OR2x2_ASAP7_75t_L g688 ( 
.A(n_522),
.B(n_448),
.Y(n_688)
);

INVx4_ASAP7_75t_L g689 ( 
.A(n_516),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_492),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_492),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_584),
.B(n_471),
.Y(n_692)
);

INVxp67_ASAP7_75t_L g693 ( 
.A(n_661),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_545),
.Y(n_694)
);

INVx2_ASAP7_75t_SL g695 ( 
.A(n_638),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_556),
.Y(n_696)
);

AND2x4_ASAP7_75t_L g697 ( 
.A(n_559),
.B(n_533),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_584),
.B(n_520),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_680),
.B(n_520),
.Y(n_699)
);

NAND2x1p5_ASAP7_75t_L g700 ( 
.A(n_610),
.B(n_246),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_635),
.B(n_520),
.Y(n_701)
);

AOI22xp5_ASAP7_75t_SL g702 ( 
.A1(n_672),
.A2(n_441),
.B1(n_456),
.B2(n_453),
.Y(n_702)
);

A2O1A1Ixp33_ASAP7_75t_L g703 ( 
.A1(n_660),
.A2(n_288),
.B(n_331),
.C(n_250),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_545),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_565),
.Y(n_705)
);

BUFx3_ASAP7_75t_L g706 ( 
.A(n_638),
.Y(n_706)
);

O2A1O1Ixp33_ASAP7_75t_L g707 ( 
.A1(n_688),
.A2(n_537),
.B(n_533),
.C(n_525),
.Y(n_707)
);

NOR2xp33_ASAP7_75t_L g708 ( 
.A(n_624),
.B(n_551),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_610),
.B(n_252),
.Y(n_709)
);

INVxp67_ASAP7_75t_L g710 ( 
.A(n_571),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_610),
.B(n_277),
.Y(n_711)
);

OAI22xp33_ASAP7_75t_L g712 ( 
.A1(n_667),
.A2(n_223),
.B1(n_361),
.B2(n_219),
.Y(n_712)
);

INVx2_ASAP7_75t_SL g713 ( 
.A(n_541),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_554),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_664),
.B(n_520),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_670),
.B(n_520),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_554),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_671),
.B(n_524),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_624),
.B(n_207),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_673),
.Y(n_720)
);

NOR3xp33_ASAP7_75t_L g721 ( 
.A(n_608),
.B(n_540),
.C(n_537),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_678),
.B(n_524),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_543),
.B(n_524),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_560),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_660),
.B(n_281),
.Y(n_725)
);

OAI22xp33_ASAP7_75t_L g726 ( 
.A1(n_667),
.A2(n_202),
.B1(n_361),
.B2(n_358),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_588),
.B(n_295),
.Y(n_727)
);

AND2x4_ASAP7_75t_L g728 ( 
.A(n_662),
.B(n_435),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_574),
.B(n_207),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_578),
.B(n_298),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_673),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_609),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_637),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_552),
.B(n_524),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_552),
.B(n_493),
.Y(n_735)
);

INVx2_ASAP7_75t_SL g736 ( 
.A(n_541),
.Y(n_736)
);

OAI22xp5_ASAP7_75t_L g737 ( 
.A1(n_662),
.A2(n_352),
.B1(n_309),
.B2(n_311),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_575),
.B(n_493),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_560),
.Y(n_739)
);

BUFx2_ASAP7_75t_L g740 ( 
.A(n_571),
.Y(n_740)
);

OAI22xp5_ASAP7_75t_L g741 ( 
.A1(n_557),
.A2(n_355),
.B1(n_314),
.B2(n_315),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_688),
.B(n_212),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_589),
.B(n_495),
.Y(n_743)
);

NOR2x1p5_ASAP7_75t_L g744 ( 
.A(n_546),
.B(n_202),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_564),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_592),
.B(n_321),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_564),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_568),
.Y(n_748)
);

OAI22xp5_ASAP7_75t_L g749 ( 
.A1(n_577),
.A2(n_544),
.B1(n_567),
.B2(n_555),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_637),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_598),
.B(n_495),
.Y(n_751)
);

BUFx5_ASAP7_75t_L g752 ( 
.A(n_623),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_568),
.Y(n_753)
);

OAI22xp33_ASAP7_75t_L g754 ( 
.A1(n_667),
.A2(n_204),
.B1(n_358),
.B2(n_356),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_569),
.Y(n_755)
);

NAND2xp33_ASAP7_75t_L g756 ( 
.A(n_544),
.B(n_290),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_641),
.B(n_497),
.Y(n_757)
);

HB1xp67_ASAP7_75t_L g758 ( 
.A(n_607),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_641),
.B(n_497),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_561),
.B(n_212),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_569),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_643),
.Y(n_762)
);

NAND2x1p5_ASAP7_75t_L g763 ( 
.A(n_555),
.B(n_326),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_643),
.B(n_499),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_623),
.B(n_339),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_581),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_572),
.A2(n_300),
.B1(n_301),
.B2(n_304),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_648),
.B(n_499),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_648),
.B(n_526),
.Y(n_769)
);

BUFx5_ASAP7_75t_L g770 ( 
.A(n_553),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_548),
.Y(n_771)
);

NOR3xp33_ASAP7_75t_L g772 ( 
.A(n_633),
.B(n_449),
.C(n_448),
.Y(n_772)
);

NOR3xp33_ASAP7_75t_L g773 ( 
.A(n_640),
.B(n_449),
.C(n_438),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_654),
.B(n_679),
.Y(n_774)
);

NOR2x1p5_ASAP7_75t_L g775 ( 
.A(n_546),
.B(n_629),
.Y(n_775)
);

NAND3xp33_ASAP7_75t_L g776 ( 
.A(n_586),
.B(n_228),
.C(n_225),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_654),
.B(n_526),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_679),
.B(n_526),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_639),
.A2(n_512),
.B(n_529),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_581),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_681),
.B(n_526),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_582),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_582),
.Y(n_783)
);

INVxp67_ASAP7_75t_L g784 ( 
.A(n_607),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_548),
.Y(n_785)
);

NAND2x1p5_ASAP7_75t_L g786 ( 
.A(n_567),
.B(n_526),
.Y(n_786)
);

OR2x2_ASAP7_75t_L g787 ( 
.A(n_573),
.B(n_436),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_681),
.B(n_512),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_583),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_583),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_550),
.A2(n_318),
.B1(n_319),
.B2(n_320),
.Y(n_791)
);

INVxp67_ASAP7_75t_L g792 ( 
.A(n_579),
.Y(n_792)
);

HB1xp67_ASAP7_75t_L g793 ( 
.A(n_667),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_591),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_682),
.Y(n_795)
);

INVx5_ASAP7_75t_L g796 ( 
.A(n_548),
.Y(n_796)
);

AOI22xp33_ASAP7_75t_L g797 ( 
.A1(n_667),
.A2(n_223),
.B1(n_356),
.B2(n_348),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_594),
.B(n_627),
.Y(n_798)
);

BUFx6f_ASAP7_75t_L g799 ( 
.A(n_548),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_682),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_594),
.B(n_213),
.Y(n_801)
);

NAND2xp33_ASAP7_75t_L g802 ( 
.A(n_590),
.B(n_603),
.Y(n_802)
);

HB1xp67_ASAP7_75t_L g803 ( 
.A(n_621),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_591),
.Y(n_804)
);

OAI22xp5_ASAP7_75t_L g805 ( 
.A1(n_590),
.A2(n_603),
.B1(n_580),
.B2(n_595),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_686),
.B(n_512),
.Y(n_806)
);

NAND2xp33_ASAP7_75t_L g807 ( 
.A(n_686),
.B(n_330),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_627),
.B(n_333),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_621),
.B(n_516),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_SL g810 ( 
.A(n_629),
.B(n_514),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_599),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_621),
.B(n_650),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_621),
.B(n_516),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_599),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_612),
.B(n_213),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_650),
.B(n_516),
.Y(n_816)
);

BUFx3_ASAP7_75t_L g817 ( 
.A(n_642),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_628),
.B(n_217),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_653),
.B(n_518),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_653),
.B(n_666),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_666),
.B(n_674),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_642),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_674),
.B(n_518),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_675),
.B(n_518),
.Y(n_824)
);

INVx2_ASAP7_75t_SL g825 ( 
.A(n_669),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_675),
.B(n_518),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_601),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_668),
.B(n_217),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_676),
.B(n_518),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_587),
.A2(n_218),
.B1(n_348),
.B2(n_347),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_676),
.B(n_518),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_677),
.B(n_518),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_684),
.B(n_529),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_684),
.B(n_531),
.Y(n_834)
);

INVx2_ASAP7_75t_SL g835 ( 
.A(n_669),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_687),
.B(n_531),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_657),
.B(n_542),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_601),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_617),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_687),
.B(n_531),
.Y(n_840)
);

BUFx3_ASAP7_75t_L g841 ( 
.A(n_644),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_690),
.B(n_222),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_690),
.B(n_527),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_691),
.B(n_222),
.Y(n_844)
);

OAI22xp33_ASAP7_75t_L g845 ( 
.A1(n_645),
.A2(n_211),
.B1(n_214),
.B2(n_215),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_548),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_691),
.B(n_234),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_587),
.A2(n_211),
.B1(n_214),
.B2(n_219),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_639),
.A2(n_527),
.B(n_521),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_566),
.B(n_570),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_618),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_566),
.B(n_234),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_542),
.B(n_336),
.Y(n_853)
);

OR2x2_ASAP7_75t_SL g854 ( 
.A(n_793),
.B(n_645),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_708),
.B(n_576),
.Y(n_855)
);

INVx5_ASAP7_75t_L g856 ( 
.A(n_771),
.Y(n_856)
);

OR2x2_ASAP7_75t_L g857 ( 
.A(n_693),
.B(n_636),
.Y(n_857)
);

AND2x6_ASAP7_75t_L g858 ( 
.A(n_699),
.B(n_576),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_708),
.B(n_656),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_L g860 ( 
.A1(n_692),
.A2(n_646),
.B1(n_587),
.B2(n_614),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_697),
.Y(n_861)
);

INVx3_ASAP7_75t_L g862 ( 
.A(n_697),
.Y(n_862)
);

INVx3_ASAP7_75t_L g863 ( 
.A(n_771),
.Y(n_863)
);

AO22x1_ASAP7_75t_L g864 ( 
.A1(n_729),
.A2(n_342),
.B1(n_341),
.B2(n_338),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_713),
.B(n_644),
.Y(n_865)
);

INVx3_ASAP7_75t_L g866 ( 
.A(n_771),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_R g867 ( 
.A(n_732),
.B(n_656),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_696),
.Y(n_868)
);

BUFx6f_ASAP7_75t_SL g869 ( 
.A(n_817),
.Y(n_869)
);

OR2x2_ASAP7_75t_L g870 ( 
.A(n_758),
.B(n_580),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_SL g871 ( 
.A1(n_729),
.A2(n_663),
.B1(n_656),
.B2(n_646),
.Y(n_871)
);

HB1xp67_ASAP7_75t_L g872 ( 
.A(n_758),
.Y(n_872)
);

HB1xp67_ASAP7_75t_L g873 ( 
.A(n_740),
.Y(n_873)
);

AOI22xp33_ASAP7_75t_L g874 ( 
.A1(n_692),
.A2(n_646),
.B1(n_602),
.B2(n_614),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_736),
.B(n_576),
.Y(n_875)
);

HB1xp67_ASAP7_75t_L g876 ( 
.A(n_706),
.Y(n_876)
);

BUFx2_ASAP7_75t_L g877 ( 
.A(n_839),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_SL g878 ( 
.A(n_810),
.B(n_663),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_738),
.B(n_618),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_701),
.B(n_566),
.Y(n_880)
);

AOI22xp5_ASAP7_75t_L g881 ( 
.A1(n_837),
.A2(n_663),
.B1(n_580),
.B2(n_646),
.Y(n_881)
);

BUFx2_ASAP7_75t_L g882 ( 
.A(n_710),
.Y(n_882)
);

AOI21xp33_ASAP7_75t_L g883 ( 
.A1(n_815),
.A2(n_580),
.B(n_683),
.Y(n_883)
);

INVx1_ASAP7_75t_SL g884 ( 
.A(n_787),
.Y(n_884)
);

INVxp33_ASAP7_75t_SL g885 ( 
.A(n_822),
.Y(n_885)
);

INVx4_ASAP7_75t_L g886 ( 
.A(n_771),
.Y(n_886)
);

OAI22xp33_ASAP7_75t_L g887 ( 
.A1(n_720),
.A2(n_602),
.B1(n_580),
.B2(n_338),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_705),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_698),
.B(n_620),
.Y(n_889)
);

AND2x4_ASAP7_75t_L g890 ( 
.A(n_695),
.B(n_436),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_815),
.B(n_620),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_742),
.B(n_644),
.Y(n_892)
);

BUFx6f_ASAP7_75t_L g893 ( 
.A(n_785),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_792),
.B(n_644),
.Y(n_894)
);

HB1xp67_ASAP7_75t_L g895 ( 
.A(n_784),
.Y(n_895)
);

BUFx3_ASAP7_75t_L g896 ( 
.A(n_841),
.Y(n_896)
);

A2O1A1Ixp33_ASAP7_75t_L g897 ( 
.A1(n_837),
.A2(n_553),
.B(n_596),
.C(n_597),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_742),
.B(n_626),
.Y(n_898)
);

OAI22xp5_ASAP7_75t_L g899 ( 
.A1(n_803),
.A2(n_639),
.B1(n_652),
.B2(n_626),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_702),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_733),
.B(n_558),
.Y(n_901)
);

INVx2_ASAP7_75t_SL g902 ( 
.A(n_728),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_803),
.Y(n_903)
);

INVx3_ASAP7_75t_L g904 ( 
.A(n_785),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_750),
.B(n_558),
.Y(n_905)
);

AOI22xp33_ASAP7_75t_L g906 ( 
.A1(n_830),
.A2(n_597),
.B1(n_562),
.B2(n_563),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_694),
.Y(n_907)
);

AND2x4_ASAP7_75t_L g908 ( 
.A(n_731),
.B(n_442),
.Y(n_908)
);

AND2x2_ASAP7_75t_SL g909 ( 
.A(n_830),
.B(n_652),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_775),
.Y(n_910)
);

AND2x2_ASAP7_75t_L g911 ( 
.A(n_719),
.B(n_669),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_719),
.B(n_562),
.Y(n_912)
);

AOI22xp5_ASAP7_75t_L g913 ( 
.A1(n_793),
.A2(n_596),
.B1(n_600),
.B2(n_604),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_762),
.Y(n_914)
);

BUFx3_ASAP7_75t_L g915 ( 
.A(n_825),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_795),
.B(n_563),
.Y(n_916)
);

INVx3_ASAP7_75t_L g917 ( 
.A(n_785),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_845),
.B(n_853),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_704),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_800),
.B(n_585),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_820),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_851),
.Y(n_922)
);

NOR2xp33_ASAP7_75t_L g923 ( 
.A(n_853),
.B(n_585),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_821),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_714),
.Y(n_925)
);

INVx3_ASAP7_75t_L g926 ( 
.A(n_785),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_743),
.B(n_600),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_770),
.B(n_566),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_751),
.B(n_604),
.Y(n_929)
);

AOI22xp5_ASAP7_75t_L g930 ( 
.A1(n_721),
.A2(n_613),
.B1(n_630),
.B2(n_616),
.Y(n_930)
);

OAI22xp5_ASAP7_75t_L g931 ( 
.A1(n_749),
.A2(n_652),
.B1(n_616),
.B2(n_622),
.Y(n_931)
);

NAND2x1p5_ASAP7_75t_L g932 ( 
.A(n_812),
.B(n_606),
.Y(n_932)
);

AND2x2_ASAP7_75t_L g933 ( 
.A(n_828),
.B(n_442),
.Y(n_933)
);

AOI22xp5_ASAP7_75t_L g934 ( 
.A1(n_812),
.A2(n_631),
.B1(n_613),
.B2(n_622),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_821),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_774),
.B(n_625),
.Y(n_936)
);

AOI22xp33_ASAP7_75t_L g937 ( 
.A1(n_848),
.A2(n_625),
.B1(n_630),
.B2(n_631),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_770),
.B(n_566),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_788),
.Y(n_939)
);

BUFx3_ASAP7_75t_L g940 ( 
.A(n_835),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_802),
.A2(n_549),
.B(n_665),
.Y(n_941)
);

INVx3_ASAP7_75t_L g942 ( 
.A(n_799),
.Y(n_942)
);

INVx3_ASAP7_75t_L g943 ( 
.A(n_799),
.Y(n_943)
);

INVx5_ASAP7_75t_L g944 ( 
.A(n_799),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_806),
.Y(n_945)
);

AOI22xp33_ASAP7_75t_L g946 ( 
.A1(n_848),
.A2(n_343),
.B1(n_280),
.B2(n_347),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_770),
.B(n_570),
.Y(n_947)
);

INVx5_ASAP7_75t_L g948 ( 
.A(n_799),
.Y(n_948)
);

INVx2_ASAP7_75t_L g949 ( 
.A(n_717),
.Y(n_949)
);

BUFx2_ASAP7_75t_L g950 ( 
.A(n_700),
.Y(n_950)
);

AOI22xp33_ASAP7_75t_L g951 ( 
.A1(n_727),
.A2(n_343),
.B1(n_346),
.B2(n_344),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_715),
.B(n_570),
.Y(n_952)
);

AO22x1_ASAP7_75t_L g953 ( 
.A1(n_828),
.A2(n_341),
.B1(n_342),
.B2(n_344),
.Y(n_953)
);

AOI22xp5_ASAP7_75t_L g954 ( 
.A1(n_709),
.A2(n_549),
.B1(n_651),
.B2(n_658),
.Y(n_954)
);

INVxp67_ASAP7_75t_L g955 ( 
.A(n_760),
.Y(n_955)
);

INVx2_ASAP7_75t_SL g956 ( 
.A(n_744),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_716),
.B(n_570),
.Y(n_957)
);

NOR2x1p5_ASAP7_75t_L g958 ( 
.A(n_776),
.B(n_346),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_770),
.B(n_570),
.Y(n_959)
);

BUFx3_ASAP7_75t_L g960 ( 
.A(n_700),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_718),
.B(n_549),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_770),
.B(n_606),
.Y(n_962)
);

AND2x4_ASAP7_75t_L g963 ( 
.A(n_773),
.B(n_444),
.Y(n_963)
);

BUFx3_ASAP7_75t_L g964 ( 
.A(n_763),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_724),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_735),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_722),
.B(n_632),
.Y(n_967)
);

INVx2_ASAP7_75t_SL g968 ( 
.A(n_842),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_846),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_770),
.B(n_606),
.Y(n_970)
);

NAND2x1p5_ASAP7_75t_L g971 ( 
.A(n_809),
.B(n_619),
.Y(n_971)
);

INVx3_ASAP7_75t_L g972 ( 
.A(n_846),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_757),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_759),
.Y(n_974)
);

OAI21xp5_ASAP7_75t_L g975 ( 
.A1(n_798),
.A2(n_647),
.B(n_634),
.Y(n_975)
);

INVx3_ASAP7_75t_L g976 ( 
.A(n_846),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_764),
.Y(n_977)
);

AND2x4_ASAP7_75t_L g978 ( 
.A(n_725),
.B(n_444),
.Y(n_978)
);

AOI22xp5_ASAP7_75t_L g979 ( 
.A1(n_709),
.A2(n_658),
.B1(n_651),
.B2(n_647),
.Y(n_979)
);

AOI22xp33_ASAP7_75t_L g980 ( 
.A1(n_727),
.A2(n_276),
.B1(n_317),
.B2(n_324),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_707),
.B(n_632),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_739),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_712),
.B(n_619),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_745),
.Y(n_984)
);

AOI22xp5_ASAP7_75t_L g985 ( 
.A1(n_711),
.A2(n_658),
.B1(n_651),
.B2(n_634),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_752),
.B(n_619),
.Y(n_986)
);

BUFx3_ASAP7_75t_L g987 ( 
.A(n_763),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_752),
.B(n_655),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_768),
.Y(n_989)
);

INVx2_ASAP7_75t_SL g990 ( 
.A(n_842),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_747),
.Y(n_991)
);

AND2x4_ASAP7_75t_L g992 ( 
.A(n_725),
.B(n_445),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_796),
.A2(n_655),
.B(n_665),
.Y(n_993)
);

INVxp67_ASAP7_75t_L g994 ( 
.A(n_760),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_752),
.B(n_655),
.Y(n_995)
);

AOI22xp33_ASAP7_75t_L g996 ( 
.A1(n_797),
.A2(n_324),
.B1(n_276),
.B2(n_317),
.Y(n_996)
);

INVx3_ASAP7_75t_SL g997 ( 
.A(n_844),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_833),
.Y(n_998)
);

AOI22xp33_ASAP7_75t_L g999 ( 
.A1(n_797),
.A2(n_324),
.B1(n_276),
.B2(n_317),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_818),
.B(n_445),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_711),
.B(n_649),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_752),
.B(n_659),
.Y(n_1002)
);

INVx2_ASAP7_75t_SL g1003 ( 
.A(n_844),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_752),
.B(n_659),
.Y(n_1004)
);

HB1xp67_ASAP7_75t_L g1005 ( 
.A(n_798),
.Y(n_1005)
);

AOI22xp5_ASAP7_75t_L g1006 ( 
.A1(n_730),
.A2(n_659),
.B1(n_665),
.B2(n_689),
.Y(n_1006)
);

AOI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_730),
.A2(n_746),
.B1(n_808),
.B2(n_805),
.Y(n_1007)
);

AOI22xp33_ASAP7_75t_L g1008 ( 
.A1(n_726),
.A2(n_605),
.B1(n_611),
.B2(n_615),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_748),
.Y(n_1009)
);

AOI22xp33_ASAP7_75t_SL g1010 ( 
.A1(n_801),
.A2(n_336),
.B1(n_345),
.B2(n_351),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_801),
.B(n_605),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_746),
.B(n_723),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_834),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_836),
.Y(n_1014)
);

INVx2_ASAP7_75t_SL g1015 ( 
.A(n_847),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_726),
.B(n_236),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_753),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_767),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_840),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_786),
.A2(n_351),
.B1(n_362),
.B2(n_360),
.Y(n_1020)
);

AOI22xp33_ASAP7_75t_L g1021 ( 
.A1(n_754),
.A2(n_615),
.B1(n_237),
.B2(n_322),
.Y(n_1021)
);

HB1xp67_ASAP7_75t_L g1022 ( 
.A(n_741),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_734),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_754),
.B(n_245),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_769),
.Y(n_1025)
);

INVx4_ASAP7_75t_L g1026 ( 
.A(n_846),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_786),
.A2(n_345),
.B1(n_360),
.B2(n_362),
.Y(n_1027)
);

CKINVDCx20_ASAP7_75t_R g1028 ( 
.A(n_791),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_755),
.Y(n_1029)
);

INVx3_ASAP7_75t_L g1030 ( 
.A(n_752),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_777),
.B(n_593),
.Y(n_1031)
);

HB1xp67_ASAP7_75t_L g1032 ( 
.A(n_778),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_781),
.B(n_593),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_847),
.B(n_593),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_955),
.B(n_852),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_949),
.Y(n_1036)
);

AND2x2_ASAP7_75t_SL g1037 ( 
.A(n_918),
.B(n_772),
.Y(n_1037)
);

O2A1O1Ixp5_ASAP7_75t_L g1038 ( 
.A1(n_918),
.A2(n_852),
.B(n_808),
.C(n_765),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_1030),
.A2(n_796),
.B(n_850),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_1030),
.A2(n_796),
.B(n_850),
.Y(n_1040)
);

BUFx12f_ASAP7_75t_L g1041 ( 
.A(n_877),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_884),
.B(n_765),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_966),
.B(n_843),
.Y(n_1043)
);

INVx3_ASAP7_75t_L g1044 ( 
.A(n_893),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_856),
.A2(n_796),
.B(n_809),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_973),
.B(n_737),
.Y(n_1046)
);

BUFx6f_ASAP7_75t_L g1047 ( 
.A(n_893),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_974),
.B(n_761),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_893),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_994),
.B(n_807),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_914),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_859),
.B(n_813),
.Y(n_1052)
);

A2O1A1Ixp33_ASAP7_75t_SL g1053 ( 
.A1(n_859),
.A2(n_756),
.B(n_849),
.C(n_779),
.Y(n_1053)
);

HB1xp67_ASAP7_75t_L g1054 ( 
.A(n_873),
.Y(n_1054)
);

HB1xp67_ASAP7_75t_L g1055 ( 
.A(n_873),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_977),
.B(n_766),
.Y(n_1056)
);

BUFx2_ASAP7_75t_L g1057 ( 
.A(n_872),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_885),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_933),
.B(n_515),
.Y(n_1059)
);

CKINVDCx12_ASAP7_75t_R g1060 ( 
.A(n_857),
.Y(n_1060)
);

BUFx12f_ASAP7_75t_L g1061 ( 
.A(n_910),
.Y(n_1061)
);

O2A1O1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_1022),
.A2(n_1016),
.B(n_1024),
.C(n_892),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_989),
.B(n_780),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_912),
.B(n_782),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_949),
.Y(n_1065)
);

INVx2_ASAP7_75t_SL g1066 ( 
.A(n_872),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_912),
.B(n_783),
.Y(n_1067)
);

CKINVDCx14_ASAP7_75t_R g1068 ( 
.A(n_867),
.Y(n_1068)
);

NOR3xp33_ASAP7_75t_SL g1069 ( 
.A(n_900),
.B(n_287),
.C(n_278),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_965),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_856),
.A2(n_813),
.B(n_689),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_965),
.Y(n_1072)
);

A2O1A1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_1007),
.A2(n_703),
.B(n_838),
.C(n_789),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_894),
.B(n_790),
.Y(n_1074)
);

AO22x1_ASAP7_75t_L g1075 ( 
.A1(n_1016),
.A2(n_259),
.B1(n_261),
.B2(n_267),
.Y(n_1075)
);

OAI21xp33_ASAP7_75t_L g1076 ( 
.A1(n_996),
.A2(n_269),
.B(n_270),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_911),
.B(n_816),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1005),
.B(n_794),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_903),
.Y(n_1079)
);

AOI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_1018),
.A2(n_811),
.B1(n_804),
.B2(n_814),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_874),
.A2(n_827),
.B1(n_831),
.B2(n_829),
.Y(n_1081)
);

CKINVDCx20_ASAP7_75t_R g1082 ( 
.A(n_867),
.Y(n_1082)
);

BUFx3_ASAP7_75t_L g1083 ( 
.A(n_882),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_874),
.A2(n_826),
.B1(n_824),
.B2(n_823),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_879),
.B(n_819),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_894),
.B(n_832),
.Y(n_1086)
);

INVx3_ASAP7_75t_L g1087 ( 
.A(n_893),
.Y(n_1087)
);

HB1xp67_ASAP7_75t_L g1088 ( 
.A(n_876),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_876),
.B(n_515),
.Y(n_1089)
);

AO32x1_ASAP7_75t_L g1090 ( 
.A1(n_931),
.A2(n_521),
.A3(n_519),
.B1(n_517),
.B2(n_527),
.Y(n_1090)
);

OAI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_1005),
.A2(n_909),
.B1(n_860),
.B2(n_996),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_923),
.B(n_517),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_883),
.A2(n_363),
.B(n_296),
.C(n_297),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_856),
.A2(n_689),
.B(n_547),
.Y(n_1094)
);

O2A1O1Ixp33_ASAP7_75t_L g1095 ( 
.A1(n_1022),
.A2(n_519),
.B(n_302),
.C(n_307),
.Y(n_1095)
);

O2A1O1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_1024),
.A2(n_293),
.B(n_310),
.C(n_323),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_L g1097 ( 
.A(n_923),
.B(n_363),
.Y(n_1097)
);

BUFx12f_ASAP7_75t_L g1098 ( 
.A(n_956),
.Y(n_1098)
);

BUFx2_ASAP7_75t_L g1099 ( 
.A(n_895),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_921),
.B(n_593),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_969),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_862),
.B(n_685),
.Y(n_1102)
);

AOI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_902),
.A2(n_685),
.B1(n_332),
.B2(n_547),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_939),
.B(n_685),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_945),
.B(n_1032),
.Y(n_1105)
);

OAI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_909),
.A2(n_685),
.B1(n_547),
.B2(n_4),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_856),
.A2(n_547),
.B(n_685),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_944),
.A2(n_547),
.B(n_180),
.Y(n_1108)
);

BUFx6f_ASAP7_75t_L g1109 ( 
.A(n_969),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_897),
.A2(n_547),
.B(n_177),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_968),
.A2(n_1003),
.B(n_990),
.C(n_1015),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_944),
.A2(n_168),
.B(n_167),
.Y(n_1112)
);

O2A1O1Ixp5_ASAP7_75t_SL g1113 ( 
.A1(n_855),
.A2(n_1),
.B(n_3),
.C(n_5),
.Y(n_1113)
);

AO32x1_ASAP7_75t_L g1114 ( 
.A1(n_899),
.A2(n_1),
.A3(n_3),
.B1(n_14),
.B2(n_15),
.Y(n_1114)
);

AO21x1_ASAP7_75t_L g1115 ( 
.A1(n_1011),
.A2(n_14),
.B(n_16),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1032),
.B(n_17),
.Y(n_1116)
);

BUFx2_ASAP7_75t_L g1117 ( 
.A(n_854),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_R g1118 ( 
.A(n_878),
.B(n_164),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_898),
.B(n_18),
.Y(n_1119)
);

O2A1O1Ixp33_ASAP7_75t_L g1120 ( 
.A1(n_887),
.A2(n_18),
.B(n_21),
.C(n_25),
.Y(n_1120)
);

OAI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_860),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_999),
.A2(n_28),
.B1(n_30),
.B2(n_33),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_862),
.B(n_71),
.Y(n_1123)
);

OAI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_897),
.A2(n_161),
.B(n_69),
.Y(n_1124)
);

BUFx4f_ASAP7_75t_L g1125 ( 
.A(n_997),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_997),
.B(n_33),
.Y(n_1126)
);

O2A1O1Ixp33_ASAP7_75t_L g1127 ( 
.A1(n_887),
.A2(n_35),
.B(n_39),
.C(n_41),
.Y(n_1127)
);

OAI22xp33_ASAP7_75t_L g1128 ( 
.A1(n_870),
.A2(n_39),
.B1(n_42),
.B2(n_43),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_999),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_1129)
);

NOR3xp33_ASAP7_75t_SL g1130 ( 
.A(n_1020),
.B(n_1027),
.C(n_888),
.Y(n_1130)
);

BUFx4f_ASAP7_75t_L g1131 ( 
.A(n_950),
.Y(n_1131)
);

XOR2x2_ASAP7_75t_L g1132 ( 
.A(n_946),
.B(n_49),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_983),
.A2(n_51),
.B1(n_53),
.B2(n_55),
.Y(n_1133)
);

INVx4_ASAP7_75t_L g1134 ( 
.A(n_944),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_865),
.B(n_112),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_891),
.B(n_57),
.Y(n_1136)
);

BUFx6f_ASAP7_75t_L g1137 ( 
.A(n_969),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_998),
.B(n_59),
.Y(n_1138)
);

BUFx2_ASAP7_75t_L g1139 ( 
.A(n_896),
.Y(n_1139)
);

OR2x6_ASAP7_75t_L g1140 ( 
.A(n_960),
.B(n_129),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_896),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_969),
.Y(n_1142)
);

OAI22xp5_ASAP7_75t_L g1143 ( 
.A1(n_983),
.A2(n_67),
.B1(n_76),
.B2(n_86),
.Y(n_1143)
);

BUFx12f_ASAP7_75t_L g1144 ( 
.A(n_958),
.Y(n_1144)
);

AO22x1_ASAP7_75t_L g1145 ( 
.A1(n_960),
.A2(n_94),
.B1(n_103),
.B2(n_110),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_944),
.A2(n_132),
.B(n_138),
.Y(n_1146)
);

BUFx4f_ASAP7_75t_L g1147 ( 
.A(n_861),
.Y(n_1147)
);

INVx4_ASAP7_75t_L g1148 ( 
.A(n_948),
.Y(n_1148)
);

OR2x6_ASAP7_75t_SL g1149 ( 
.A(n_868),
.B(n_143),
.Y(n_1149)
);

A2O1A1Ixp33_ASAP7_75t_L g1150 ( 
.A1(n_881),
.A2(n_146),
.B(n_151),
.C(n_153),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_948),
.A2(n_157),
.B(n_961),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_1028),
.B(n_1000),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1013),
.B(n_1014),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_948),
.A2(n_962),
.B(n_970),
.Y(n_1154)
);

OA21x2_ASAP7_75t_L g1155 ( 
.A1(n_880),
.A2(n_975),
.B(n_952),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_901),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_984),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_948),
.A2(n_962),
.B(n_970),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_1009),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_871),
.B(n_964),
.Y(n_1160)
);

INVx5_ASAP7_75t_L g1161 ( 
.A(n_886),
.Y(n_1161)
);

AND2x2_ASAP7_75t_L g1162 ( 
.A(n_890),
.B(n_978),
.Y(n_1162)
);

INVx1_ASAP7_75t_SL g1163 ( 
.A(n_890),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_957),
.A2(n_988),
.B(n_1002),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1019),
.B(n_1023),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_905),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1009),
.Y(n_1167)
);

OR2x6_ASAP7_75t_L g1168 ( 
.A(n_964),
.B(n_987),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1025),
.B(n_927),
.Y(n_1169)
);

BUFx6f_ASAP7_75t_L g1170 ( 
.A(n_915),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_916),
.Y(n_1171)
);

INVx3_ASAP7_75t_L g1172 ( 
.A(n_886),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_987),
.B(n_908),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_929),
.B(n_978),
.Y(n_1174)
);

O2A1O1Ixp33_ASAP7_75t_L g1175 ( 
.A1(n_855),
.A2(n_980),
.B(n_875),
.C(n_922),
.Y(n_1175)
);

HB1xp67_ASAP7_75t_L g1176 ( 
.A(n_869),
.Y(n_1176)
);

AO21x1_ASAP7_75t_L g1177 ( 
.A1(n_880),
.A2(n_1012),
.B(n_981),
.Y(n_1177)
);

BUFx6f_ASAP7_75t_L g1178 ( 
.A(n_940),
.Y(n_1178)
);

BUFx2_ASAP7_75t_L g1179 ( 
.A(n_908),
.Y(n_1179)
);

NAND2x1_ASAP7_75t_L g1180 ( 
.A(n_1026),
.B(n_863),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1029),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_R g1182 ( 
.A(n_869),
.B(n_940),
.Y(n_1182)
);

INVx1_ASAP7_75t_L g1183 ( 
.A(n_920),
.Y(n_1183)
);

NOR2xp33_ASAP7_75t_L g1184 ( 
.A(n_864),
.B(n_1010),
.Y(n_1184)
);

BUFx3_ASAP7_75t_L g1185 ( 
.A(n_963),
.Y(n_1185)
);

O2A1O1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_980),
.A2(n_875),
.B(n_889),
.C(n_963),
.Y(n_1186)
);

NAND3xp33_ASAP7_75t_L g1187 ( 
.A(n_1062),
.B(n_946),
.C(n_953),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1156),
.B(n_992),
.Y(n_1188)
);

OA21x2_ASAP7_75t_L g1189 ( 
.A1(n_1110),
.A2(n_967),
.B(n_936),
.Y(n_1189)
);

INVx3_ASAP7_75t_L g1190 ( 
.A(n_1134),
.Y(n_1190)
);

AO31x2_ASAP7_75t_L g1191 ( 
.A1(n_1177),
.A2(n_941),
.A3(n_1033),
.B(n_1034),
.Y(n_1191)
);

NAND3xp33_ASAP7_75t_L g1192 ( 
.A(n_1184),
.B(n_951),
.C(n_1021),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1051),
.Y(n_1193)
);

AOI221xp5_ASAP7_75t_SL g1194 ( 
.A1(n_1076),
.A2(n_951),
.B1(n_1021),
.B2(n_937),
.C(n_906),
.Y(n_1194)
);

INVxp67_ASAP7_75t_SL g1195 ( 
.A(n_1054),
.Y(n_1195)
);

AO22x2_ASAP7_75t_L g1196 ( 
.A1(n_1091),
.A2(n_935),
.B1(n_924),
.B2(n_992),
.Y(n_1196)
);

BUFx2_ASAP7_75t_L g1197 ( 
.A(n_1083),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1053),
.A2(n_995),
.B(n_986),
.Y(n_1198)
);

INVxp67_ASAP7_75t_L g1199 ( 
.A(n_1055),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1052),
.A2(n_913),
.B1(n_971),
.B2(n_932),
.Y(n_1200)
);

OAI21xp5_ASAP7_75t_SL g1201 ( 
.A1(n_1122),
.A2(n_930),
.B(n_937),
.Y(n_1201)
);

OAI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1038),
.A2(n_1001),
.B(n_985),
.Y(n_1202)
);

OAI22xp5_ASAP7_75t_L g1203 ( 
.A1(n_1169),
.A2(n_971),
.B1(n_932),
.B2(n_1006),
.Y(n_1203)
);

BUFx2_ASAP7_75t_L g1204 ( 
.A(n_1099),
.Y(n_1204)
);

OAI22xp5_ASAP7_75t_L g1205 ( 
.A1(n_1169),
.A2(n_954),
.B1(n_1026),
.B2(n_959),
.Y(n_1205)
);

OAI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_1163),
.A2(n_991),
.B1(n_925),
.B2(n_1017),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1162),
.B(n_982),
.Y(n_1207)
);

AO21x1_ASAP7_75t_L g1208 ( 
.A1(n_1091),
.A2(n_1031),
.B(n_959),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1164),
.A2(n_986),
.B(n_988),
.Y(n_1209)
);

NOR2xp67_ASAP7_75t_L g1210 ( 
.A(n_1161),
.B(n_943),
.Y(n_1210)
);

OAI21xp5_ASAP7_75t_SL g1211 ( 
.A1(n_1122),
.A2(n_906),
.B(n_1008),
.Y(n_1211)
);

A2O1A1Ixp33_ASAP7_75t_L g1212 ( 
.A1(n_1096),
.A2(n_919),
.B(n_907),
.C(n_934),
.Y(n_1212)
);

AND2x4_ASAP7_75t_L g1213 ( 
.A(n_1185),
.B(n_1168),
.Y(n_1213)
);

AO21x1_ASAP7_75t_L g1214 ( 
.A1(n_1106),
.A2(n_1031),
.B(n_928),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1166),
.B(n_1171),
.Y(n_1215)
);

AOI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1077),
.A2(n_947),
.B(n_938),
.Y(n_1216)
);

OAI21xp33_ASAP7_75t_SL g1217 ( 
.A1(n_1110),
.A2(n_947),
.B(n_938),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_1058),
.Y(n_1218)
);

OAI22x1_ASAP7_75t_L g1219 ( 
.A1(n_1117),
.A2(n_928),
.B1(n_1029),
.B2(n_979),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1036),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_1168),
.B(n_972),
.Y(n_1221)
);

INVxp67_ASAP7_75t_L g1222 ( 
.A(n_1057),
.Y(n_1222)
);

CKINVDCx20_ASAP7_75t_R g1223 ( 
.A(n_1082),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1085),
.A2(n_1004),
.B(n_1002),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_SL g1225 ( 
.A(n_1041),
.B(n_942),
.Y(n_1225)
);

AOI21xp33_ASAP7_75t_L g1226 ( 
.A1(n_1037),
.A2(n_1004),
.B(n_995),
.Y(n_1226)
);

INVx3_ASAP7_75t_SL g1227 ( 
.A(n_1170),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1154),
.A2(n_993),
.B(n_863),
.Y(n_1228)
);

BUFx3_ASAP7_75t_L g1229 ( 
.A(n_1139),
.Y(n_1229)
);

AND2x4_ASAP7_75t_L g1230 ( 
.A(n_1168),
.B(n_926),
.Y(n_1230)
);

OR2x2_ASAP7_75t_L g1231 ( 
.A(n_1163),
.B(n_1105),
.Y(n_1231)
);

AOI221x1_ASAP7_75t_L g1232 ( 
.A1(n_1106),
.A2(n_926),
.B1(n_866),
.B2(n_904),
.C(n_917),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1158),
.A2(n_942),
.B(n_866),
.Y(n_1233)
);

INVx3_ASAP7_75t_L g1234 ( 
.A(n_1134),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_SL g1235 ( 
.A(n_1125),
.B(n_904),
.Y(n_1235)
);

AO31x2_ASAP7_75t_L g1236 ( 
.A1(n_1073),
.A2(n_858),
.A3(n_917),
.B(n_943),
.Y(n_1236)
);

OAI21x1_ASAP7_75t_L g1237 ( 
.A1(n_1039),
.A2(n_976),
.B(n_972),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1040),
.A2(n_976),
.B(n_858),
.Y(n_1238)
);

OAI21xp33_ASAP7_75t_L g1239 ( 
.A1(n_1132),
.A2(n_858),
.B(n_1126),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1065),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1042),
.B(n_858),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1070),
.Y(n_1242)
);

CKINVDCx5p33_ASAP7_75t_R g1243 ( 
.A(n_1061),
.Y(n_1243)
);

AO31x2_ASAP7_75t_L g1244 ( 
.A1(n_1084),
.A2(n_858),
.A3(n_1115),
.B(n_1081),
.Y(n_1244)
);

INVx8_ASAP7_75t_L g1245 ( 
.A(n_1161),
.Y(n_1245)
);

NAND2x1p5_ASAP7_75t_L g1246 ( 
.A(n_1161),
.B(n_1131),
.Y(n_1246)
);

AO31x2_ASAP7_75t_L g1247 ( 
.A1(n_1084),
.A2(n_1081),
.A3(n_1086),
.B(n_1093),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1183),
.B(n_1153),
.Y(n_1248)
);

NAND3xp33_ASAP7_75t_L g1249 ( 
.A(n_1097),
.B(n_1129),
.C(n_1035),
.Y(n_1249)
);

AOI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1129),
.A2(n_1121),
.B1(n_1174),
.B2(n_1160),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1072),
.Y(n_1251)
);

NAND2xp33_ASAP7_75t_L g1252 ( 
.A(n_1046),
.B(n_1153),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1151),
.A2(n_1071),
.B(n_1094),
.Y(n_1253)
);

AOI21x1_ASAP7_75t_L g1254 ( 
.A1(n_1064),
.A2(n_1067),
.B(n_1092),
.Y(n_1254)
);

AO31x2_ASAP7_75t_L g1255 ( 
.A1(n_1150),
.A2(n_1121),
.A3(n_1111),
.B(n_1074),
.Y(n_1255)
);

HB1xp67_ASAP7_75t_L g1256 ( 
.A(n_1088),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1165),
.B(n_1059),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1043),
.B(n_1050),
.Y(n_1258)
);

AO22x2_ASAP7_75t_L g1259 ( 
.A1(n_1133),
.A2(n_1124),
.B1(n_1143),
.B2(n_1136),
.Y(n_1259)
);

NAND3xp33_ASAP7_75t_L g1260 ( 
.A(n_1130),
.B(n_1075),
.C(n_1095),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1089),
.B(n_1048),
.Y(n_1261)
);

OAI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1175),
.A2(n_1119),
.B(n_1124),
.Y(n_1262)
);

AND2x4_ASAP7_75t_L g1263 ( 
.A(n_1173),
.B(n_1179),
.Y(n_1263)
);

HB1xp67_ASAP7_75t_SL g1264 ( 
.A(n_1176),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1107),
.A2(n_1045),
.B(n_1078),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1157),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1048),
.B(n_1116),
.Y(n_1267)
);

INVx3_ASAP7_75t_L g1268 ( 
.A(n_1148),
.Y(n_1268)
);

NAND2xp33_ASAP7_75t_R g1269 ( 
.A(n_1182),
.B(n_1118),
.Y(n_1269)
);

INVxp67_ASAP7_75t_L g1270 ( 
.A(n_1066),
.Y(n_1270)
);

NOR2xp33_ASAP7_75t_L g1271 ( 
.A(n_1060),
.B(n_1079),
.Y(n_1271)
);

AOI211x1_ASAP7_75t_L g1272 ( 
.A1(n_1133),
.A2(n_1128),
.B(n_1138),
.C(n_1056),
.Y(n_1272)
);

BUFx2_ASAP7_75t_L g1273 ( 
.A(n_1141),
.Y(n_1273)
);

AOI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1155),
.A2(n_1078),
.B(n_1102),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1148),
.A2(n_1155),
.B(n_1104),
.Y(n_1275)
);

OAI21xp33_ASAP7_75t_SL g1276 ( 
.A1(n_1063),
.A2(n_1113),
.B(n_1140),
.Y(n_1276)
);

HB1xp67_ASAP7_75t_L g1277 ( 
.A(n_1170),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1159),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1108),
.A2(n_1100),
.B(n_1167),
.Y(n_1279)
);

OA21x2_ASAP7_75t_L g1280 ( 
.A1(n_1181),
.A2(n_1123),
.B(n_1112),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1180),
.A2(n_1146),
.B(n_1044),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1147),
.A2(n_1080),
.B1(n_1172),
.B2(n_1140),
.Y(n_1282)
);

O2A1O1Ixp5_ASAP7_75t_SL g1283 ( 
.A1(n_1135),
.A2(n_1114),
.B(n_1044),
.C(n_1087),
.Y(n_1283)
);

O2A1O1Ixp33_ASAP7_75t_SL g1284 ( 
.A1(n_1120),
.A2(n_1127),
.B(n_1103),
.C(n_1087),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1147),
.B(n_1178),
.Y(n_1285)
);

AOI21xp33_ASAP7_75t_L g1286 ( 
.A1(n_1178),
.A2(n_1140),
.B(n_1068),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1178),
.B(n_1149),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1172),
.A2(n_1090),
.B(n_1145),
.Y(n_1288)
);

BUFx2_ASAP7_75t_L g1289 ( 
.A(n_1098),
.Y(n_1289)
);

OAI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1069),
.A2(n_1090),
.B(n_1114),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1047),
.A2(n_1049),
.B(n_1101),
.Y(n_1291)
);

INVx3_ASAP7_75t_L g1292 ( 
.A(n_1047),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_L g1293 ( 
.A(n_1144),
.B(n_1047),
.Y(n_1293)
);

NOR2x1_ASAP7_75t_SL g1294 ( 
.A(n_1049),
.B(n_1101),
.Y(n_1294)
);

OAI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1114),
.A2(n_1049),
.B(n_1101),
.Y(n_1295)
);

INVx4_ASAP7_75t_L g1296 ( 
.A(n_1109),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1109),
.B(n_1137),
.Y(n_1297)
);

INVx2_ASAP7_75t_SL g1298 ( 
.A(n_1142),
.Y(n_1298)
);

A2O1A1Ixp33_ASAP7_75t_L g1299 ( 
.A1(n_1109),
.A2(n_918),
.B(n_1062),
.C(n_729),
.Y(n_1299)
);

AOI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1137),
.A2(n_1053),
.B(n_944),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1137),
.B(n_1142),
.Y(n_1301)
);

OAI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1038),
.A2(n_918),
.B(n_1186),
.Y(n_1302)
);

AOI21xp5_ASAP7_75t_L g1303 ( 
.A1(n_1053),
.A2(n_944),
.B(n_856),
.Y(n_1303)
);

AOI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1164),
.A2(n_880),
.B(n_1077),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1053),
.A2(n_944),
.B(n_856),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1053),
.A2(n_944),
.B(n_856),
.Y(n_1306)
);

A2O1A1Ixp33_ASAP7_75t_L g1307 ( 
.A1(n_1062),
.A2(n_918),
.B(n_729),
.C(n_692),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1053),
.A2(n_944),
.B(n_856),
.Y(n_1308)
);

AO31x2_ASAP7_75t_L g1309 ( 
.A1(n_1177),
.A2(n_1091),
.A3(n_897),
.B(n_1106),
.Y(n_1309)
);

INVx5_ASAP7_75t_L g1310 ( 
.A(n_1134),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1053),
.A2(n_944),
.B(n_856),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1053),
.A2(n_944),
.B(n_856),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1053),
.A2(n_944),
.B(n_856),
.Y(n_1313)
);

CKINVDCx20_ASAP7_75t_R g1314 ( 
.A(n_1082),
.Y(n_1314)
);

AO32x2_ASAP7_75t_L g1315 ( 
.A1(n_1091),
.A2(n_1106),
.A3(n_1121),
.B1(n_1133),
.B2(n_1129),
.Y(n_1315)
);

INVx1_ASAP7_75t_SL g1316 ( 
.A(n_1083),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1053),
.A2(n_944),
.B(n_856),
.Y(n_1317)
);

OAI21x1_ASAP7_75t_L g1318 ( 
.A1(n_1164),
.A2(n_1158),
.B(n_1154),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1053),
.A2(n_944),
.B(n_856),
.Y(n_1319)
);

AO31x2_ASAP7_75t_L g1320 ( 
.A1(n_1177),
.A2(n_1091),
.A3(n_897),
.B(n_1106),
.Y(n_1320)
);

OAI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1038),
.A2(n_918),
.B(n_1186),
.Y(n_1321)
);

OAI21xp5_ASAP7_75t_SL g1322 ( 
.A1(n_1152),
.A2(n_918),
.B(n_672),
.Y(n_1322)
);

AO21x1_ASAP7_75t_L g1323 ( 
.A1(n_1091),
.A2(n_1106),
.B(n_1110),
.Y(n_1323)
);

AND2x4_ASAP7_75t_L g1324 ( 
.A(n_1185),
.B(n_1162),
.Y(n_1324)
);

NOR2xp67_ASAP7_75t_SL g1325 ( 
.A(n_1058),
.B(n_732),
.Y(n_1325)
);

NOR2xp67_ASAP7_75t_SL g1326 ( 
.A(n_1058),
.B(n_732),
.Y(n_1326)
);

INVx4_ASAP7_75t_L g1327 ( 
.A(n_1161),
.Y(n_1327)
);

INVx3_ASAP7_75t_L g1328 ( 
.A(n_1134),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_1058),
.Y(n_1329)
);

NOR2xp33_ASAP7_75t_L g1330 ( 
.A(n_1152),
.B(n_693),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1053),
.A2(n_944),
.B(n_856),
.Y(n_1331)
);

AND2x4_ASAP7_75t_L g1332 ( 
.A(n_1185),
.B(n_1162),
.Y(n_1332)
);

AND2x4_ASAP7_75t_L g1333 ( 
.A(n_1185),
.B(n_1162),
.Y(n_1333)
);

O2A1O1Ixp5_ASAP7_75t_L g1334 ( 
.A1(n_1110),
.A2(n_729),
.B(n_918),
.C(n_859),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1053),
.A2(n_944),
.B(n_856),
.Y(n_1335)
);

AO32x2_ASAP7_75t_L g1336 ( 
.A1(n_1091),
.A2(n_1106),
.A3(n_1121),
.B1(n_1133),
.B2(n_1129),
.Y(n_1336)
);

OAI21x1_ASAP7_75t_L g1337 ( 
.A1(n_1164),
.A2(n_1158),
.B(n_1154),
.Y(n_1337)
);

BUFx3_ASAP7_75t_L g1338 ( 
.A(n_1083),
.Y(n_1338)
);

NOR3xp33_ASAP7_75t_L g1339 ( 
.A(n_1062),
.B(n_918),
.C(n_729),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_1228),
.A2(n_1279),
.B(n_1238),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_1218),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_SL g1342 ( 
.A1(n_1192),
.A2(n_1187),
.B1(n_1260),
.B2(n_1330),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1207),
.B(n_1324),
.Y(n_1343)
);

CKINVDCx6p67_ASAP7_75t_R g1344 ( 
.A(n_1227),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1257),
.B(n_1248),
.Y(n_1345)
);

AO21x2_ASAP7_75t_L g1346 ( 
.A1(n_1262),
.A2(n_1339),
.B(n_1321),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_SL g1347 ( 
.A1(n_1192),
.A2(n_1187),
.B1(n_1260),
.B2(n_1249),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1304),
.A2(n_1209),
.B(n_1265),
.Y(n_1348)
);

INVx2_ASAP7_75t_SL g1349 ( 
.A(n_1338),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1198),
.A2(n_1275),
.B(n_1237),
.Y(n_1350)
);

OR2x2_ASAP7_75t_L g1351 ( 
.A(n_1231),
.B(n_1215),
.Y(n_1351)
);

OR2x2_ASAP7_75t_L g1352 ( 
.A(n_1256),
.B(n_1261),
.Y(n_1352)
);

OR2x6_ASAP7_75t_L g1353 ( 
.A(n_1245),
.B(n_1272),
.Y(n_1353)
);

A2O1A1Ixp33_ASAP7_75t_L g1354 ( 
.A1(n_1334),
.A2(n_1307),
.B(n_1211),
.C(n_1217),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1252),
.A2(n_1302),
.B(n_1217),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1300),
.A2(n_1308),
.B(n_1312),
.Y(n_1356)
);

BUFx6f_ASAP7_75t_L g1357 ( 
.A(n_1245),
.Y(n_1357)
);

OA21x2_ASAP7_75t_L g1358 ( 
.A1(n_1232),
.A2(n_1323),
.B(n_1288),
.Y(n_1358)
);

OAI21x1_ASAP7_75t_L g1359 ( 
.A1(n_1303),
.A2(n_1313),
.B(n_1317),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1305),
.A2(n_1306),
.B(n_1311),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1239),
.A2(n_1250),
.B1(n_1259),
.B2(n_1267),
.Y(n_1361)
);

OAI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1212),
.A2(n_1203),
.B(n_1200),
.Y(n_1362)
);

INVx2_ASAP7_75t_SL g1363 ( 
.A(n_1229),
.Y(n_1363)
);

NOR2xp67_ASAP7_75t_L g1364 ( 
.A(n_1329),
.B(n_1270),
.Y(n_1364)
);

OR2x6_ASAP7_75t_L g1365 ( 
.A(n_1245),
.B(n_1272),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1319),
.A2(n_1335),
.B(n_1331),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1281),
.A2(n_1233),
.B(n_1224),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_SL g1368 ( 
.A1(n_1259),
.A2(n_1282),
.B1(n_1196),
.B2(n_1271),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1274),
.A2(n_1216),
.B(n_1202),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1254),
.A2(n_1205),
.B(n_1280),
.Y(n_1370)
);

AOI221xp5_ASAP7_75t_L g1371 ( 
.A1(n_1201),
.A2(n_1194),
.B1(n_1250),
.B2(n_1284),
.C(n_1196),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1324),
.B(n_1332),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1332),
.B(n_1333),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1295),
.A2(n_1283),
.B(n_1280),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1188),
.B(n_1263),
.Y(n_1375)
);

OA21x2_ASAP7_75t_L g1376 ( 
.A1(n_1290),
.A2(n_1208),
.B(n_1214),
.Y(n_1376)
);

NAND2x1p5_ASAP7_75t_L g1377 ( 
.A(n_1310),
.B(n_1327),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1189),
.A2(n_1291),
.B(n_1201),
.Y(n_1378)
);

AOI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1219),
.A2(n_1189),
.B(n_1241),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1240),
.A2(n_1266),
.B(n_1278),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1242),
.A2(n_1251),
.B(n_1268),
.Y(n_1381)
);

AO31x2_ASAP7_75t_L g1382 ( 
.A1(n_1244),
.A2(n_1236),
.A3(n_1320),
.B(n_1309),
.Y(n_1382)
);

OAI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1190),
.A2(n_1268),
.B(n_1234),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1297),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1301),
.Y(n_1385)
);

BUFx5_ASAP7_75t_L g1386 ( 
.A(n_1221),
.Y(n_1386)
);

NOR2xp67_ASAP7_75t_L g1387 ( 
.A(n_1199),
.B(n_1285),
.Y(n_1387)
);

AOI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1269),
.A2(n_1263),
.B1(n_1287),
.B2(n_1326),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1206),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1190),
.A2(n_1234),
.B(n_1328),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1195),
.Y(n_1391)
);

OA21x2_ASAP7_75t_L g1392 ( 
.A1(n_1226),
.A2(n_1244),
.B(n_1320),
.Y(n_1392)
);

AND2x4_ASAP7_75t_L g1393 ( 
.A(n_1221),
.B(n_1230),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_SL g1394 ( 
.A(n_1325),
.B(n_1243),
.Y(n_1394)
);

OR2x2_ASAP7_75t_L g1395 ( 
.A(n_1222),
.B(n_1273),
.Y(n_1395)
);

OAI21xp5_ASAP7_75t_L g1396 ( 
.A1(n_1276),
.A2(n_1235),
.B(n_1210),
.Y(n_1396)
);

AO32x2_ASAP7_75t_L g1397 ( 
.A1(n_1315),
.A2(n_1336),
.A3(n_1320),
.B1(n_1309),
.B2(n_1276),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1247),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1328),
.A2(n_1292),
.B(n_1246),
.Y(n_1399)
);

OAI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1225),
.A2(n_1336),
.B1(n_1315),
.B2(n_1286),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1310),
.A2(n_1230),
.B(n_1294),
.Y(n_1401)
);

AO21x2_ASAP7_75t_L g1402 ( 
.A1(n_1247),
.A2(n_1191),
.B(n_1309),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1191),
.A2(n_1293),
.B(n_1277),
.Y(n_1403)
);

INVx2_ASAP7_75t_SL g1404 ( 
.A(n_1197),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1247),
.Y(n_1405)
);

CKINVDCx20_ASAP7_75t_R g1406 ( 
.A(n_1223),
.Y(n_1406)
);

O2A1O1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1316),
.A2(n_1213),
.B(n_1289),
.C(n_1298),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1255),
.Y(n_1408)
);

BUFx3_ASAP7_75t_L g1409 ( 
.A(n_1314),
.Y(n_1409)
);

AOI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1264),
.A2(n_1327),
.B1(n_1296),
.B2(n_1315),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1255),
.Y(n_1411)
);

AO32x2_ASAP7_75t_L g1412 ( 
.A1(n_1203),
.A2(n_1121),
.A3(n_1091),
.B1(n_1133),
.B2(n_1129),
.Y(n_1412)
);

OAI211xp5_ASAP7_75t_L g1413 ( 
.A1(n_1322),
.A2(n_918),
.B(n_999),
.C(n_996),
.Y(n_1413)
);

NOR2xp33_ASAP7_75t_L g1414 ( 
.A(n_1330),
.B(n_918),
.Y(n_1414)
);

OR2x2_ASAP7_75t_L g1415 ( 
.A(n_1231),
.B(n_1258),
.Y(n_1415)
);

OR2x2_ASAP7_75t_L g1416 ( 
.A(n_1231),
.B(n_1258),
.Y(n_1416)
);

AO21x2_ASAP7_75t_L g1417 ( 
.A1(n_1262),
.A2(n_1339),
.B(n_1321),
.Y(n_1417)
);

NOR2x1_ASAP7_75t_R g1418 ( 
.A(n_1218),
.B(n_642),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1192),
.A2(n_918),
.B1(n_1132),
.B2(n_1339),
.Y(n_1419)
);

AO21x2_ASAP7_75t_L g1420 ( 
.A1(n_1262),
.A2(n_1339),
.B(n_1321),
.Y(n_1420)
);

AO32x2_ASAP7_75t_L g1421 ( 
.A1(n_1203),
.A2(n_1121),
.A3(n_1091),
.B1(n_1133),
.B2(n_1129),
.Y(n_1421)
);

OAI21x1_ASAP7_75t_L g1422 ( 
.A1(n_1253),
.A2(n_1337),
.B(n_1318),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1192),
.A2(n_918),
.B1(n_1132),
.B2(n_1339),
.Y(n_1423)
);

NAND3xp33_ASAP7_75t_L g1424 ( 
.A(n_1339),
.B(n_729),
.C(n_1307),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1330),
.B(n_918),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1207),
.B(n_1152),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1220),
.Y(n_1427)
);

AOI221xp5_ASAP7_75t_L g1428 ( 
.A1(n_1192),
.A2(n_918),
.B1(n_845),
.B2(n_693),
.C(n_1307),
.Y(n_1428)
);

AND2x4_ASAP7_75t_L g1429 ( 
.A(n_1221),
.B(n_1230),
.Y(n_1429)
);

BUFx12f_ASAP7_75t_L g1430 ( 
.A(n_1243),
.Y(n_1430)
);

O2A1O1Ixp33_ASAP7_75t_SL g1431 ( 
.A1(n_1307),
.A2(n_1299),
.B(n_1124),
.C(n_1150),
.Y(n_1431)
);

BUFx2_ASAP7_75t_SL g1432 ( 
.A(n_1338),
.Y(n_1432)
);

AOI22xp33_ASAP7_75t_L g1433 ( 
.A1(n_1192),
.A2(n_918),
.B1(n_1132),
.B2(n_1339),
.Y(n_1433)
);

A2O1A1Ixp33_ASAP7_75t_L g1434 ( 
.A1(n_1334),
.A2(n_918),
.B(n_1307),
.C(n_1062),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1220),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1193),
.Y(n_1436)
);

OAI21xp5_ASAP7_75t_L g1437 ( 
.A1(n_1334),
.A2(n_729),
.B(n_1307),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1330),
.A2(n_918),
.B1(n_729),
.B2(n_1192),
.Y(n_1438)
);

OA21x2_ASAP7_75t_L g1439 ( 
.A1(n_1262),
.A2(n_1321),
.B(n_1302),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1192),
.A2(n_918),
.B1(n_1132),
.B2(n_1339),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1220),
.Y(n_1441)
);

OR2x2_ASAP7_75t_L g1442 ( 
.A(n_1231),
.B(n_1258),
.Y(n_1442)
);

NAND2x1p5_ASAP7_75t_L g1443 ( 
.A(n_1310),
.B(n_1327),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1262),
.A2(n_1252),
.B(n_1302),
.Y(n_1444)
);

NAND2x1p5_ASAP7_75t_L g1445 ( 
.A(n_1310),
.B(n_1327),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1220),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1192),
.A2(n_918),
.B1(n_1132),
.B2(n_1339),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1192),
.A2(n_918),
.B1(n_1132),
.B2(n_1339),
.Y(n_1448)
);

INVx4_ASAP7_75t_L g1449 ( 
.A(n_1245),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1220),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1192),
.A2(n_918),
.B1(n_1132),
.B2(n_1339),
.Y(n_1451)
);

BUFx3_ASAP7_75t_L g1452 ( 
.A(n_1227),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1192),
.A2(n_918),
.B1(n_1132),
.B2(n_1339),
.Y(n_1453)
);

INVx1_ASAP7_75t_SL g1454 ( 
.A(n_1204),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1192),
.A2(n_918),
.B1(n_1132),
.B2(n_1339),
.Y(n_1455)
);

OAI21x1_ASAP7_75t_SL g1456 ( 
.A1(n_1214),
.A2(n_1115),
.B(n_1124),
.Y(n_1456)
);

BUFx2_ASAP7_75t_L g1457 ( 
.A(n_1197),
.Y(n_1457)
);

OA21x2_ASAP7_75t_L g1458 ( 
.A1(n_1262),
.A2(n_1321),
.B(n_1302),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_1341),
.Y(n_1459)
);

OA21x2_ASAP7_75t_L g1460 ( 
.A1(n_1362),
.A2(n_1355),
.B(n_1374),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1426),
.B(n_1343),
.Y(n_1461)
);

INVxp67_ASAP7_75t_L g1462 ( 
.A(n_1395),
.Y(n_1462)
);

BUFx2_ASAP7_75t_SL g1463 ( 
.A(n_1364),
.Y(n_1463)
);

HB1xp67_ASAP7_75t_L g1464 ( 
.A(n_1352),
.Y(n_1464)
);

AOI21xp5_ASAP7_75t_L g1465 ( 
.A1(n_1431),
.A2(n_1424),
.B(n_1438),
.Y(n_1465)
);

AND2x4_ASAP7_75t_L g1466 ( 
.A(n_1393),
.B(n_1429),
.Y(n_1466)
);

AOI21xp5_ASAP7_75t_SL g1467 ( 
.A1(n_1345),
.A2(n_1425),
.B(n_1414),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1347),
.B(n_1361),
.Y(n_1468)
);

BUFx6f_ASAP7_75t_L g1469 ( 
.A(n_1452),
.Y(n_1469)
);

OAI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1419),
.A2(n_1451),
.B1(n_1423),
.B2(n_1448),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1419),
.A2(n_1451),
.B1(n_1423),
.B2(n_1448),
.Y(n_1471)
);

O2A1O1Ixp33_ASAP7_75t_L g1472 ( 
.A1(n_1413),
.A2(n_1425),
.B(n_1414),
.C(n_1434),
.Y(n_1472)
);

OR2x2_ASAP7_75t_L g1473 ( 
.A(n_1415),
.B(n_1416),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1442),
.B(n_1351),
.Y(n_1474)
);

O2A1O1Ixp33_ASAP7_75t_L g1475 ( 
.A1(n_1433),
.A2(n_1447),
.B(n_1453),
.C(n_1455),
.Y(n_1475)
);

AOI21xp5_ASAP7_75t_SL g1476 ( 
.A1(n_1428),
.A2(n_1407),
.B(n_1439),
.Y(n_1476)
);

OA21x2_ASAP7_75t_L g1477 ( 
.A1(n_1374),
.A2(n_1370),
.B(n_1360),
.Y(n_1477)
);

AOI21xp5_ASAP7_75t_SL g1478 ( 
.A1(n_1458),
.A2(n_1418),
.B(n_1377),
.Y(n_1478)
);

NAND4xp25_ASAP7_75t_L g1479 ( 
.A(n_1433),
.B(n_1440),
.C(n_1453),
.D(n_1455),
.Y(n_1479)
);

OR2x2_ASAP7_75t_L g1480 ( 
.A(n_1361),
.B(n_1391),
.Y(n_1480)
);

BUFx2_ASAP7_75t_L g1481 ( 
.A(n_1457),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1342),
.B(n_1440),
.Y(n_1482)
);

OR2x2_ASAP7_75t_L g1483 ( 
.A(n_1375),
.B(n_1454),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1384),
.Y(n_1484)
);

O2A1O1Ixp33_ASAP7_75t_L g1485 ( 
.A1(n_1447),
.A2(n_1354),
.B(n_1456),
.C(n_1400),
.Y(n_1485)
);

A2O1A1Ixp33_ASAP7_75t_L g1486 ( 
.A1(n_1354),
.A2(n_1371),
.B(n_1368),
.C(n_1396),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1372),
.B(n_1373),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1400),
.A2(n_1410),
.B1(n_1388),
.B2(n_1436),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1385),
.B(n_1346),
.Y(n_1489)
);

AND2x4_ASAP7_75t_SL g1490 ( 
.A(n_1344),
.B(n_1406),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1346),
.B(n_1417),
.Y(n_1491)
);

INVx1_ASAP7_75t_SL g1492 ( 
.A(n_1406),
.Y(n_1492)
);

CKINVDCx20_ASAP7_75t_R g1493 ( 
.A(n_1341),
.Y(n_1493)
);

CKINVDCx20_ASAP7_75t_R g1494 ( 
.A(n_1409),
.Y(n_1494)
);

OAI31xp33_ASAP7_75t_L g1495 ( 
.A1(n_1394),
.A2(n_1389),
.A3(n_1404),
.B(n_1409),
.Y(n_1495)
);

INVxp67_ASAP7_75t_L g1496 ( 
.A(n_1363),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1417),
.B(n_1420),
.Y(n_1497)
);

O2A1O1Ixp5_ASAP7_75t_L g1498 ( 
.A1(n_1379),
.A2(n_1405),
.B(n_1398),
.C(n_1411),
.Y(n_1498)
);

A2O1A1Ixp33_ASAP7_75t_SL g1499 ( 
.A1(n_1398),
.A2(n_1405),
.B(n_1408),
.C(n_1411),
.Y(n_1499)
);

AOI21xp5_ASAP7_75t_SL g1500 ( 
.A1(n_1377),
.A2(n_1443),
.B(n_1445),
.Y(n_1500)
);

A2O1A1Ixp33_ASAP7_75t_L g1501 ( 
.A1(n_1387),
.A2(n_1378),
.B(n_1401),
.C(n_1403),
.Y(n_1501)
);

INVx1_ASAP7_75t_SL g1502 ( 
.A(n_1432),
.Y(n_1502)
);

OA21x2_ASAP7_75t_L g1503 ( 
.A1(n_1359),
.A2(n_1366),
.B(n_1369),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1450),
.B(n_1427),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1380),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1402),
.B(n_1382),
.Y(n_1506)
);

OAI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1353),
.A2(n_1365),
.B1(n_1421),
.B2(n_1412),
.Y(n_1507)
);

OAI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1353),
.A2(n_1365),
.B1(n_1421),
.B2(n_1412),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1380),
.Y(n_1509)
);

OAI22xp5_ASAP7_75t_SL g1510 ( 
.A1(n_1430),
.A2(n_1365),
.B1(n_1353),
.B2(n_1349),
.Y(n_1510)
);

AOI21xp5_ASAP7_75t_SL g1511 ( 
.A1(n_1443),
.A2(n_1445),
.B(n_1449),
.Y(n_1511)
);

AOI21xp5_ASAP7_75t_SL g1512 ( 
.A1(n_1449),
.A2(n_1357),
.B(n_1446),
.Y(n_1512)
);

OAI22xp5_ASAP7_75t_L g1513 ( 
.A1(n_1412),
.A2(n_1421),
.B1(n_1441),
.B2(n_1435),
.Y(n_1513)
);

OAI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1412),
.A2(n_1421),
.B1(n_1446),
.B2(n_1441),
.Y(n_1514)
);

OAI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1376),
.A2(n_1392),
.B1(n_1358),
.B2(n_1357),
.Y(n_1515)
);

HB1xp67_ASAP7_75t_L g1516 ( 
.A(n_1381),
.Y(n_1516)
);

OR2x2_ASAP7_75t_L g1517 ( 
.A(n_1392),
.B(n_1376),
.Y(n_1517)
);

OA22x2_ASAP7_75t_L g1518 ( 
.A1(n_1399),
.A2(n_1381),
.B1(n_1390),
.B2(n_1383),
.Y(n_1518)
);

AOI221x1_ASAP7_75t_SL g1519 ( 
.A1(n_1397),
.A2(n_1358),
.B1(n_1386),
.B2(n_1369),
.C(n_1357),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1386),
.B(n_1383),
.Y(n_1520)
);

O2A1O1Ixp33_ASAP7_75t_L g1521 ( 
.A1(n_1356),
.A2(n_1397),
.B(n_1348),
.C(n_1350),
.Y(n_1521)
);

OAI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1397),
.A2(n_1367),
.B1(n_1422),
.B2(n_1340),
.Y(n_1522)
);

O2A1O1Ixp5_ASAP7_75t_L g1523 ( 
.A1(n_1397),
.A2(n_1334),
.B(n_1444),
.C(n_1437),
.Y(n_1523)
);

OAI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1422),
.A2(n_918),
.B1(n_1423),
.B2(n_1419),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1345),
.B(n_1415),
.Y(n_1525)
);

AOI21xp5_ASAP7_75t_SL g1526 ( 
.A1(n_1438),
.A2(n_1307),
.B(n_1299),
.Y(n_1526)
);

OA21x2_ASAP7_75t_L g1527 ( 
.A1(n_1362),
.A2(n_1355),
.B(n_1374),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1345),
.B(n_1415),
.Y(n_1528)
);

AOI21xp5_ASAP7_75t_SL g1529 ( 
.A1(n_1438),
.A2(n_1307),
.B(n_1299),
.Y(n_1529)
);

OR2x2_ASAP7_75t_L g1530 ( 
.A(n_1352),
.B(n_1415),
.Y(n_1530)
);

OAI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1419),
.A2(n_918),
.B1(n_1433),
.B2(n_1423),
.Y(n_1531)
);

AOI221xp5_ASAP7_75t_L g1532 ( 
.A1(n_1438),
.A2(n_918),
.B1(n_1419),
.B2(n_1433),
.C(n_1423),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1352),
.B(n_1415),
.Y(n_1533)
);

OAI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1419),
.A2(n_918),
.B1(n_1433),
.B2(n_1423),
.Y(n_1534)
);

AOI21xp5_ASAP7_75t_SL g1535 ( 
.A1(n_1438),
.A2(n_1307),
.B(n_1299),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1426),
.B(n_1343),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1345),
.B(n_1415),
.Y(n_1537)
);

OAI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1419),
.A2(n_918),
.B1(n_1433),
.B2(n_1423),
.Y(n_1538)
);

OAI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1419),
.A2(n_918),
.B1(n_1433),
.B2(n_1423),
.Y(n_1539)
);

AOI221x1_ASAP7_75t_SL g1540 ( 
.A1(n_1414),
.A2(n_845),
.B1(n_1425),
.B2(n_754),
.C(n_726),
.Y(n_1540)
);

O2A1O1Ixp5_ASAP7_75t_L g1541 ( 
.A1(n_1444),
.A2(n_1334),
.B(n_1437),
.C(n_1323),
.Y(n_1541)
);

OAI22xp5_ASAP7_75t_L g1542 ( 
.A1(n_1419),
.A2(n_918),
.B1(n_1433),
.B2(n_1423),
.Y(n_1542)
);

O2A1O1Ixp5_ASAP7_75t_L g1543 ( 
.A1(n_1444),
.A2(n_1334),
.B(n_1437),
.C(n_1323),
.Y(n_1543)
);

O2A1O1Ixp5_ASAP7_75t_L g1544 ( 
.A1(n_1444),
.A2(n_1334),
.B(n_1437),
.C(n_1323),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_L g1545 ( 
.A(n_1467),
.B(n_1473),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1505),
.Y(n_1546)
);

BUFx2_ASAP7_75t_L g1547 ( 
.A(n_1520),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1489),
.B(n_1513),
.Y(n_1548)
);

OR2x2_ASAP7_75t_L g1549 ( 
.A(n_1497),
.B(n_1491),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1509),
.Y(n_1550)
);

OAI21x1_ASAP7_75t_L g1551 ( 
.A1(n_1521),
.A2(n_1522),
.B(n_1498),
.Y(n_1551)
);

INVx2_ASAP7_75t_L g1552 ( 
.A(n_1517),
.Y(n_1552)
);

HB1xp67_ASAP7_75t_L g1553 ( 
.A(n_1516),
.Y(n_1553)
);

OR2x6_ASAP7_75t_L g1554 ( 
.A(n_1526),
.B(n_1529),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1477),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1460),
.B(n_1527),
.Y(n_1556)
);

BUFx4f_ASAP7_75t_SL g1557 ( 
.A(n_1493),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1460),
.B(n_1527),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1506),
.B(n_1515),
.Y(n_1559)
);

AOI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1535),
.A2(n_1465),
.B(n_1476),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1477),
.Y(n_1561)
);

OA21x2_ASAP7_75t_L g1562 ( 
.A1(n_1523),
.A2(n_1544),
.B(n_1543),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1507),
.B(n_1508),
.Y(n_1563)
);

INVx3_ASAP7_75t_L g1564 ( 
.A(n_1518),
.Y(n_1564)
);

AO21x2_ASAP7_75t_L g1565 ( 
.A1(n_1499),
.A2(n_1501),
.B(n_1524),
.Y(n_1565)
);

NOR2xp33_ASAP7_75t_L g1566 ( 
.A(n_1492),
.B(n_1474),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1503),
.Y(n_1567)
);

INVxp33_ASAP7_75t_L g1568 ( 
.A(n_1461),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1480),
.B(n_1507),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1519),
.Y(n_1570)
);

INVxp67_ASAP7_75t_L g1571 ( 
.A(n_1484),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1513),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1508),
.B(n_1514),
.Y(n_1573)
);

OR2x6_ASAP7_75t_L g1574 ( 
.A(n_1478),
.B(n_1510),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1541),
.B(n_1488),
.Y(n_1575)
);

BUFx2_ASAP7_75t_L g1576 ( 
.A(n_1464),
.Y(n_1576)
);

HB1xp67_ASAP7_75t_L g1577 ( 
.A(n_1488),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1530),
.B(n_1533),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1504),
.B(n_1486),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1485),
.Y(n_1580)
);

OR2x6_ASAP7_75t_L g1581 ( 
.A(n_1500),
.B(n_1512),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1483),
.B(n_1462),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1468),
.B(n_1528),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1468),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1472),
.B(n_1536),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1525),
.Y(n_1586)
);

BUFx2_ASAP7_75t_L g1587 ( 
.A(n_1481),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1537),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1482),
.Y(n_1589)
);

BUFx4f_ASAP7_75t_L g1590 ( 
.A(n_1554),
.Y(n_1590)
);

NOR2x1_ASAP7_75t_L g1591 ( 
.A(n_1581),
.B(n_1511),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1546),
.Y(n_1592)
);

NOR2x1_ASAP7_75t_L g1593 ( 
.A(n_1581),
.B(n_1463),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1552),
.B(n_1487),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1550),
.Y(n_1595)
);

NOR2xp33_ASAP7_75t_L g1596 ( 
.A(n_1580),
.B(n_1471),
.Y(n_1596)
);

OR2x2_ASAP7_75t_L g1597 ( 
.A(n_1549),
.B(n_1479),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1588),
.B(n_1532),
.Y(n_1598)
);

BUFx6f_ASAP7_75t_L g1599 ( 
.A(n_1554),
.Y(n_1599)
);

BUFx2_ASAP7_75t_L g1600 ( 
.A(n_1564),
.Y(n_1600)
);

CKINVDCx5p33_ASAP7_75t_R g1601 ( 
.A(n_1557),
.Y(n_1601)
);

AOI22xp33_ASAP7_75t_L g1602 ( 
.A1(n_1554),
.A2(n_1471),
.B1(n_1470),
.B2(n_1531),
.Y(n_1602)
);

OAI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1554),
.A2(n_1470),
.B1(n_1534),
.B2(n_1539),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1588),
.B(n_1542),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1573),
.B(n_1556),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1548),
.B(n_1542),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1548),
.B(n_1539),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_L g1608 ( 
.A(n_1580),
.B(n_1531),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1556),
.B(n_1466),
.Y(n_1609)
);

INVx1_ASAP7_75t_SL g1610 ( 
.A(n_1547),
.Y(n_1610)
);

AO21x2_ASAP7_75t_L g1611 ( 
.A1(n_1565),
.A2(n_1538),
.B(n_1534),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1555),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1556),
.B(n_1466),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1561),
.Y(n_1614)
);

HB1xp67_ASAP7_75t_L g1615 ( 
.A(n_1553),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1597),
.B(n_1576),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1605),
.B(n_1547),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1610),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1605),
.B(n_1563),
.Y(n_1619)
);

AOI221xp5_ASAP7_75t_L g1620 ( 
.A1(n_1596),
.A2(n_1475),
.B1(n_1538),
.B2(n_1560),
.C(n_1540),
.Y(n_1620)
);

AOI22xp33_ASAP7_75t_L g1621 ( 
.A1(n_1603),
.A2(n_1554),
.B1(n_1560),
.B2(n_1577),
.Y(n_1621)
);

AOI21xp5_ASAP7_75t_L g1622 ( 
.A1(n_1603),
.A2(n_1554),
.B(n_1575),
.Y(n_1622)
);

AOI31xp33_ASAP7_75t_L g1623 ( 
.A1(n_1602),
.A2(n_1577),
.A3(n_1575),
.B(n_1545),
.Y(n_1623)
);

CKINVDCx20_ASAP7_75t_R g1624 ( 
.A(n_1601),
.Y(n_1624)
);

AOI221xp5_ASAP7_75t_L g1625 ( 
.A1(n_1596),
.A2(n_1575),
.B1(n_1570),
.B2(n_1589),
.C(n_1585),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_L g1626 ( 
.A(n_1601),
.B(n_1578),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1595),
.Y(n_1627)
);

NAND2xp33_ASAP7_75t_R g1628 ( 
.A(n_1597),
.B(n_1459),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1605),
.B(n_1563),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_1610),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1597),
.B(n_1576),
.Y(n_1631)
);

OAI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1602),
.A2(n_1589),
.B1(n_1570),
.B2(n_1563),
.Y(n_1632)
);

NAND4xp25_ASAP7_75t_L g1633 ( 
.A(n_1608),
.B(n_1495),
.C(n_1566),
.D(n_1585),
.Y(n_1633)
);

OR2x6_ASAP7_75t_L g1634 ( 
.A(n_1599),
.B(n_1574),
.Y(n_1634)
);

A2O1A1Ixp33_ASAP7_75t_L g1635 ( 
.A1(n_1608),
.A2(n_1569),
.B(n_1585),
.C(n_1579),
.Y(n_1635)
);

AOI221xp5_ASAP7_75t_L g1636 ( 
.A1(n_1606),
.A2(n_1586),
.B1(n_1571),
.B2(n_1568),
.C(n_1584),
.Y(n_1636)
);

NAND4xp25_ASAP7_75t_SL g1637 ( 
.A(n_1607),
.B(n_1502),
.C(n_1569),
.D(n_1579),
.Y(n_1637)
);

AOI22xp33_ASAP7_75t_L g1638 ( 
.A1(n_1611),
.A2(n_1607),
.B1(n_1590),
.B2(n_1599),
.Y(n_1638)
);

OAI31xp33_ASAP7_75t_L g1639 ( 
.A1(n_1598),
.A2(n_1579),
.A3(n_1583),
.B(n_1490),
.Y(n_1639)
);

OAI221xp5_ASAP7_75t_SL g1640 ( 
.A1(n_1598),
.A2(n_1583),
.B1(n_1574),
.B2(n_1559),
.C(n_1582),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1609),
.B(n_1572),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1595),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1595),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1604),
.B(n_1578),
.Y(n_1644)
);

OAI211xp5_ASAP7_75t_SL g1645 ( 
.A1(n_1604),
.A2(n_1582),
.B(n_1496),
.C(n_1584),
.Y(n_1645)
);

OR2x6_ASAP7_75t_L g1646 ( 
.A(n_1599),
.B(n_1574),
.Y(n_1646)
);

NAND4xp25_ASAP7_75t_L g1647 ( 
.A(n_1593),
.B(n_1584),
.C(n_1582),
.D(n_1587),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1592),
.Y(n_1648)
);

OAI211xp5_ASAP7_75t_L g1649 ( 
.A1(n_1593),
.A2(n_1562),
.B(n_1559),
.C(n_1587),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1613),
.B(n_1572),
.Y(n_1650)
);

AOI211xp5_ASAP7_75t_L g1651 ( 
.A1(n_1599),
.A2(n_1559),
.B(n_1558),
.C(n_1551),
.Y(n_1651)
);

BUFx3_ASAP7_75t_L g1652 ( 
.A(n_1624),
.Y(n_1652)
);

INVxp67_ASAP7_75t_SL g1653 ( 
.A(n_1618),
.Y(n_1653)
);

INVx4_ASAP7_75t_SL g1654 ( 
.A(n_1634),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1619),
.B(n_1629),
.Y(n_1655)
);

HB1xp67_ASAP7_75t_L g1656 ( 
.A(n_1630),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1627),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1616),
.Y(n_1658)
);

INVxp67_ASAP7_75t_L g1659 ( 
.A(n_1644),
.Y(n_1659)
);

AND2x6_ASAP7_75t_L g1660 ( 
.A(n_1619),
.B(n_1591),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1642),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1631),
.B(n_1594),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1642),
.Y(n_1663)
);

NAND2x1p5_ASAP7_75t_SL g1664 ( 
.A(n_1620),
.B(n_1591),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1636),
.B(n_1635),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1643),
.Y(n_1666)
);

AOI21x1_ASAP7_75t_L g1667 ( 
.A1(n_1648),
.A2(n_1612),
.B(n_1614),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1643),
.Y(n_1668)
);

OR2x6_ASAP7_75t_L g1669 ( 
.A(n_1634),
.B(n_1574),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1625),
.B(n_1594),
.Y(n_1670)
);

OR2x6_ASAP7_75t_L g1671 ( 
.A(n_1634),
.B(n_1574),
.Y(n_1671)
);

OA21x2_ASAP7_75t_L g1672 ( 
.A1(n_1649),
.A2(n_1614),
.B(n_1612),
.Y(n_1672)
);

OA21x2_ASAP7_75t_L g1673 ( 
.A1(n_1638),
.A2(n_1614),
.B(n_1567),
.Y(n_1673)
);

INVx1_ASAP7_75t_SL g1674 ( 
.A(n_1626),
.Y(n_1674)
);

NAND3xp33_ASAP7_75t_SL g1675 ( 
.A(n_1639),
.B(n_1600),
.C(n_1494),
.Y(n_1675)
);

INVx5_ASAP7_75t_L g1676 ( 
.A(n_1634),
.Y(n_1676)
);

NAND2xp33_ASAP7_75t_L g1677 ( 
.A(n_1665),
.B(n_1599),
.Y(n_1677)
);

HB1xp67_ASAP7_75t_L g1678 ( 
.A(n_1656),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1655),
.B(n_1617),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1658),
.B(n_1647),
.Y(n_1680)
);

AND2x4_ASAP7_75t_L g1681 ( 
.A(n_1654),
.B(n_1634),
.Y(n_1681)
);

BUFx2_ASAP7_75t_L g1682 ( 
.A(n_1654),
.Y(n_1682)
);

NAND3xp33_ASAP7_75t_SL g1683 ( 
.A(n_1674),
.B(n_1639),
.C(n_1651),
.Y(n_1683)
);

BUFx2_ASAP7_75t_L g1684 ( 
.A(n_1654),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1657),
.Y(n_1685)
);

AND2x4_ASAP7_75t_L g1686 ( 
.A(n_1676),
.B(n_1646),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_L g1687 ( 
.A(n_1652),
.B(n_1557),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_SL g1688 ( 
.A(n_1676),
.B(n_1623),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1676),
.B(n_1641),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1676),
.B(n_1641),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1657),
.Y(n_1691)
);

HB1xp67_ASAP7_75t_L g1692 ( 
.A(n_1653),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1670),
.B(n_1647),
.Y(n_1693)
);

NOR2x1_ASAP7_75t_L g1694 ( 
.A(n_1675),
.B(n_1637),
.Y(n_1694)
);

OR2x2_ASAP7_75t_L g1695 ( 
.A(n_1662),
.B(n_1650),
.Y(n_1695)
);

INVx1_ASAP7_75t_SL g1696 ( 
.A(n_1652),
.Y(n_1696)
);

OR2x2_ASAP7_75t_L g1697 ( 
.A(n_1659),
.B(n_1615),
.Y(n_1697)
);

AOI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1664),
.A2(n_1611),
.B1(n_1633),
.B2(n_1632),
.Y(n_1698)
);

NOR3xp33_ASAP7_75t_L g1699 ( 
.A(n_1652),
.B(n_1633),
.C(n_1623),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1667),
.Y(n_1700)
);

NAND4xp25_ASAP7_75t_L g1701 ( 
.A(n_1664),
.B(n_1640),
.C(n_1622),
.D(n_1651),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1669),
.B(n_1646),
.Y(n_1702)
);

HB1xp67_ASAP7_75t_L g1703 ( 
.A(n_1661),
.Y(n_1703)
);

AOI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1664),
.A2(n_1611),
.B1(n_1632),
.B2(n_1621),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1669),
.B(n_1646),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1663),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1667),
.Y(n_1707)
);

OAI21xp33_ASAP7_75t_L g1708 ( 
.A1(n_1698),
.A2(n_1671),
.B(n_1645),
.Y(n_1708)
);

NOR2xp33_ASAP7_75t_L g1709 ( 
.A(n_1696),
.B(n_1469),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1703),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1685),
.Y(n_1711)
);

HB1xp67_ASAP7_75t_L g1712 ( 
.A(n_1692),
.Y(n_1712)
);

INVx1_ASAP7_75t_SL g1713 ( 
.A(n_1682),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1689),
.Y(n_1714)
);

OR2x2_ASAP7_75t_L g1715 ( 
.A(n_1678),
.B(n_1673),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1682),
.B(n_1671),
.Y(n_1716)
);

NOR2x1p5_ASAP7_75t_SL g1717 ( 
.A(n_1700),
.B(n_1707),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1680),
.B(n_1693),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1689),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1691),
.Y(n_1720)
);

INVx1_ASAP7_75t_SL g1721 ( 
.A(n_1684),
.Y(n_1721)
);

OAI21xp5_ASAP7_75t_L g1722 ( 
.A1(n_1694),
.A2(n_1672),
.B(n_1673),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1684),
.B(n_1671),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1690),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1681),
.B(n_1671),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1699),
.B(n_1660),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1681),
.B(n_1660),
.Y(n_1727)
);

O2A1O1Ixp33_ASAP7_75t_SL g1728 ( 
.A1(n_1688),
.A2(n_1628),
.B(n_1668),
.C(n_1666),
.Y(n_1728)
);

OR2x2_ASAP7_75t_L g1729 ( 
.A(n_1680),
.B(n_1673),
.Y(n_1729)
);

INVx2_ASAP7_75t_SL g1730 ( 
.A(n_1681),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1681),
.B(n_1660),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1693),
.B(n_1673),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1695),
.B(n_1697),
.Y(n_1733)
);

NOR2xp67_ASAP7_75t_L g1734 ( 
.A(n_1683),
.B(n_1666),
.Y(n_1734)
);

HB1xp67_ASAP7_75t_L g1735 ( 
.A(n_1697),
.Y(n_1735)
);

OAI211xp5_ASAP7_75t_L g1736 ( 
.A1(n_1698),
.A2(n_1672),
.B(n_1562),
.C(n_1600),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1722),
.B(n_1686),
.Y(n_1737)
);

INVx2_ASAP7_75t_L g1738 ( 
.A(n_1715),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1727),
.B(n_1731),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1712),
.B(n_1704),
.Y(n_1740)
);

INVxp67_ASAP7_75t_L g1741 ( 
.A(n_1713),
.Y(n_1741)
);

AND3x2_ASAP7_75t_L g1742 ( 
.A(n_1710),
.B(n_1687),
.C(n_1686),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1727),
.B(n_1686),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1735),
.B(n_1734),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1731),
.B(n_1686),
.Y(n_1745)
);

INVx1_ASAP7_75t_SL g1746 ( 
.A(n_1721),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1730),
.B(n_1702),
.Y(n_1747)
);

INVx2_ASAP7_75t_SL g1748 ( 
.A(n_1716),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1730),
.B(n_1716),
.Y(n_1749)
);

BUFx3_ASAP7_75t_L g1750 ( 
.A(n_1710),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1720),
.Y(n_1751)
);

AOI22xp33_ASAP7_75t_L g1752 ( 
.A1(n_1708),
.A2(n_1694),
.B1(n_1701),
.B2(n_1704),
.Y(n_1752)
);

INVx2_ASAP7_75t_SL g1753 ( 
.A(n_1723),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1723),
.B(n_1702),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1715),
.Y(n_1755)
);

INVx1_ASAP7_75t_SL g1756 ( 
.A(n_1718),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1720),
.Y(n_1757)
);

NOR2xp33_ASAP7_75t_L g1758 ( 
.A(n_1718),
.B(n_1677),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1714),
.B(n_1705),
.Y(n_1759)
);

CKINVDCx16_ASAP7_75t_R g1760 ( 
.A(n_1732),
.Y(n_1760)
);

BUFx3_ASAP7_75t_L g1761 ( 
.A(n_1714),
.Y(n_1761)
);

OR2x2_ASAP7_75t_L g1762 ( 
.A(n_1733),
.B(n_1706),
.Y(n_1762)
);

NAND4xp75_ASAP7_75t_L g1763 ( 
.A(n_1744),
.B(n_1726),
.C(n_1717),
.D(n_1725),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1746),
.B(n_1719),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1746),
.B(n_1719),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1748),
.B(n_1724),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1748),
.B(n_1724),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1761),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1761),
.Y(n_1769)
);

AOI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1752),
.A2(n_1728),
.B1(n_1725),
.B2(n_1736),
.Y(n_1770)
);

OA21x2_ASAP7_75t_L g1771 ( 
.A1(n_1752),
.A2(n_1732),
.B(n_1729),
.Y(n_1771)
);

INVx2_ASAP7_75t_L g1772 ( 
.A(n_1761),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1750),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1748),
.B(n_1679),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1750),
.Y(n_1775)
);

HB1xp67_ASAP7_75t_L g1776 ( 
.A(n_1760),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_L g1777 ( 
.A(n_1753),
.B(n_1679),
.Y(n_1777)
);

OAI21xp5_ASAP7_75t_L g1778 ( 
.A1(n_1744),
.A2(n_1729),
.B(n_1705),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1750),
.Y(n_1779)
);

AOI21xp5_ASAP7_75t_L g1780 ( 
.A1(n_1740),
.A2(n_1709),
.B(n_1711),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1750),
.Y(n_1781)
);

INVxp67_ASAP7_75t_L g1782 ( 
.A(n_1758),
.Y(n_1782)
);

OR2x2_ASAP7_75t_L g1783 ( 
.A(n_1776),
.B(n_1756),
.Y(n_1783)
);

AOI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1770),
.A2(n_1758),
.B1(n_1754),
.B2(n_1743),
.Y(n_1784)
);

INVx2_ASAP7_75t_SL g1785 ( 
.A(n_1768),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1776),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1764),
.B(n_1756),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1768),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1782),
.B(n_1749),
.Y(n_1789)
);

INVxp67_ASAP7_75t_SL g1790 ( 
.A(n_1771),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1769),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1769),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1772),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1778),
.B(n_1749),
.Y(n_1794)
);

NAND3xp33_ASAP7_75t_L g1795 ( 
.A(n_1790),
.B(n_1771),
.C(n_1741),
.Y(n_1795)
);

AOI22xp5_ASAP7_75t_L g1796 ( 
.A1(n_1790),
.A2(n_1754),
.B1(n_1753),
.B2(n_1747),
.Y(n_1796)
);

NOR3xp33_ASAP7_75t_SL g1797 ( 
.A(n_1786),
.B(n_1763),
.C(n_1765),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1789),
.B(n_1741),
.Y(n_1798)
);

NOR2xp33_ASAP7_75t_L g1799 ( 
.A(n_1783),
.B(n_1763),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1785),
.Y(n_1800)
);

OAI211xp5_ASAP7_75t_L g1801 ( 
.A1(n_1784),
.A2(n_1771),
.B(n_1740),
.C(n_1780),
.Y(n_1801)
);

OAI22xp5_ASAP7_75t_L g1802 ( 
.A1(n_1787),
.A2(n_1760),
.B1(n_1753),
.B2(n_1777),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_SL g1803 ( 
.A(n_1794),
.B(n_1760),
.Y(n_1803)
);

AOI221xp5_ASAP7_75t_L g1804 ( 
.A1(n_1794),
.A2(n_1781),
.B1(n_1779),
.B2(n_1775),
.C(n_1773),
.Y(n_1804)
);

AOI22xp33_ASAP7_75t_L g1805 ( 
.A1(n_1788),
.A2(n_1754),
.B1(n_1743),
.B2(n_1745),
.Y(n_1805)
);

NOR2x1_ASAP7_75t_L g1806 ( 
.A(n_1795),
.B(n_1772),
.Y(n_1806)
);

NOR2xp33_ASAP7_75t_L g1807 ( 
.A(n_1798),
.B(n_1742),
.Y(n_1807)
);

INVx2_ASAP7_75t_SL g1808 ( 
.A(n_1800),
.Y(n_1808)
);

O2A1O1Ixp33_ASAP7_75t_L g1809 ( 
.A1(n_1801),
.A2(n_1785),
.B(n_1792),
.C(n_1791),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_SL g1810 ( 
.A1(n_1799),
.A2(n_1737),
.B1(n_1802),
.B2(n_1749),
.Y(n_1810)
);

AOI211xp5_ASAP7_75t_L g1811 ( 
.A1(n_1803),
.A2(n_1766),
.B(n_1767),
.C(n_1737),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1796),
.Y(n_1812)
);

INVx1_ASAP7_75t_SL g1813 ( 
.A(n_1805),
.Y(n_1813)
);

INVx1_ASAP7_75t_SL g1814 ( 
.A(n_1806),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1810),
.B(n_1797),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1813),
.B(n_1804),
.Y(n_1816)
);

AND2x2_ASAP7_75t_SL g1817 ( 
.A(n_1807),
.B(n_1791),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_SL g1818 ( 
.A(n_1811),
.B(n_1737),
.Y(n_1818)
);

NOR2xp33_ASAP7_75t_L g1819 ( 
.A(n_1812),
.B(n_1793),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_SL g1820 ( 
.A(n_1808),
.B(n_1747),
.Y(n_1820)
);

XNOR2xp5_ASAP7_75t_L g1821 ( 
.A(n_1815),
.B(n_1742),
.Y(n_1821)
);

NOR2x1_ASAP7_75t_L g1822 ( 
.A(n_1814),
.B(n_1809),
.Y(n_1822)
);

AOI222xp33_ASAP7_75t_L g1823 ( 
.A1(n_1816),
.A2(n_1717),
.B1(n_1793),
.B2(n_1738),
.C1(n_1755),
.C2(n_1761),
.Y(n_1823)
);

HB1xp67_ASAP7_75t_L g1824 ( 
.A(n_1820),
.Y(n_1824)
);

OAI22xp5_ASAP7_75t_L g1825 ( 
.A1(n_1818),
.A2(n_1774),
.B1(n_1747),
.B2(n_1739),
.Y(n_1825)
);

INVx1_ASAP7_75t_SL g1826 ( 
.A(n_1817),
.Y(n_1826)
);

AO21x1_ASAP7_75t_L g1827 ( 
.A1(n_1824),
.A2(n_1819),
.B(n_1825),
.Y(n_1827)
);

NAND5xp2_ASAP7_75t_L g1828 ( 
.A(n_1823),
.B(n_1739),
.C(n_1743),
.D(n_1745),
.E(n_1759),
.Y(n_1828)
);

AOI21xp5_ASAP7_75t_SL g1829 ( 
.A1(n_1821),
.A2(n_1755),
.B(n_1738),
.Y(n_1829)
);

AOI22xp5_ASAP7_75t_L g1830 ( 
.A1(n_1827),
.A2(n_1826),
.B1(n_1822),
.B2(n_1739),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1830),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1831),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1831),
.B(n_1829),
.Y(n_1833)
);

OR2x2_ASAP7_75t_L g1834 ( 
.A(n_1833),
.B(n_1828),
.Y(n_1834)
);

OAI22x1_ASAP7_75t_L g1835 ( 
.A1(n_1832),
.A2(n_1755),
.B1(n_1738),
.B2(n_1757),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1835),
.B(n_1834),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1835),
.Y(n_1837)
);

OAI21xp5_ASAP7_75t_L g1838 ( 
.A1(n_1836),
.A2(n_1755),
.B(n_1738),
.Y(n_1838)
);

NOR2x1_ASAP7_75t_L g1839 ( 
.A(n_1838),
.B(n_1837),
.Y(n_1839)
);

OAI22xp5_ASAP7_75t_L g1840 ( 
.A1(n_1839),
.A2(n_1757),
.B1(n_1751),
.B2(n_1762),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1840),
.Y(n_1841)
);

AOI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1841),
.A2(n_1745),
.B1(n_1759),
.B2(n_1757),
.Y(n_1842)
);

AOI211xp5_ASAP7_75t_L g1843 ( 
.A1(n_1842),
.A2(n_1751),
.B(n_1759),
.C(n_1762),
.Y(n_1843)
);


endmodule