module fake_netlist_5_2589_n_2003 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_196, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_2003);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_196;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_2003;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_1960;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_1948;
wire n_1984;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_845;
wire n_663;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_901;
wire n_553;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1986;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1891;
wire n_1662;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_433;
wire n_314;
wire n_604;
wire n_368;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1406;
wire n_1279;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_1851;
wire n_758;
wire n_999;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_783;
wire n_555;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_681;
wire n_584;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1988;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_1999;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1995;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1969;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1990;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx2_ASAP7_75t_L g200 ( 
.A(n_37),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_114),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_95),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_96),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_7),
.Y(n_204)
);

BUFx10_ASAP7_75t_L g205 ( 
.A(n_172),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_54),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_22),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_26),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_52),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_60),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_8),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_19),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_46),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_142),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_70),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_115),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_51),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_0),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_91),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_109),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_131),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_151),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_88),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_99),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_66),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_176),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_135),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g228 ( 
.A(n_179),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_46),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_165),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_192),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_48),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_112),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_85),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_145),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_79),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_184),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_106),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_36),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_12),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_101),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_55),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_108),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_31),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_75),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_187),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_122),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_64),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_111),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g250 ( 
.A(n_62),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_143),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_104),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_23),
.Y(n_253)
);

INVxp67_ASAP7_75t_SL g254 ( 
.A(n_89),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_26),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_180),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_77),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_28),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_67),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_86),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_44),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_124),
.Y(n_262)
);

BUFx5_ASAP7_75t_L g263 ( 
.A(n_58),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_44),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_107),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_31),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_20),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_141),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_136),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_90),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_157),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_16),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_94),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_23),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_148),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_163),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_196),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_67),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_70),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_20),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_171),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_11),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_34),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_168),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_78),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_17),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_175),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_116),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_65),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_16),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_38),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_73),
.Y(n_292)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_49),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_173),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_190),
.Y(n_295)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_36),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_100),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_49),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_63),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_58),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_149),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_45),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_155),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_43),
.Y(n_304)
);

BUFx10_ASAP7_75t_L g305 ( 
.A(n_117),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_189),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_119),
.Y(n_307)
);

BUFx5_ASAP7_75t_L g308 ( 
.A(n_55),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_138),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_35),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_14),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_68),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_66),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_182),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_25),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_63),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_167),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_47),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_33),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_11),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_38),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_54),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_154),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_160),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_62),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_6),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_33),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_110),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_170),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_56),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_156),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_29),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_126),
.Y(n_333)
);

CKINVDCx14_ASAP7_75t_R g334 ( 
.A(n_161),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_193),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_24),
.Y(n_336)
);

BUFx5_ASAP7_75t_L g337 ( 
.A(n_146),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_93),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_19),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_40),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_32),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_39),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_42),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_9),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g345 ( 
.A(n_28),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_147),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_132),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g348 ( 
.A(n_7),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_12),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_127),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_188),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_80),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_4),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_68),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_74),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_43),
.Y(n_356)
);

INVx1_ASAP7_75t_SL g357 ( 
.A(n_29),
.Y(n_357)
);

INVx1_ASAP7_75t_SL g358 ( 
.A(n_183),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_134),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_139),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_103),
.Y(n_361)
);

BUFx10_ASAP7_75t_L g362 ( 
.A(n_158),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_174),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_87),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_14),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_50),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_65),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_130),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_197),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_137),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_191),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_113),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_74),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_15),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g375 ( 
.A(n_1),
.Y(n_375)
);

INVx1_ASAP7_75t_SL g376 ( 
.A(n_40),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_144),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_133),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_51),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_53),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_75),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_48),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_53),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_3),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_118),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_185),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_64),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_152),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_17),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_194),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_181),
.Y(n_391)
);

INVx2_ASAP7_75t_SL g392 ( 
.A(n_34),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_25),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_24),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_3),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_18),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g397 ( 
.A(n_76),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_60),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_18),
.Y(n_399)
);

INVxp67_ASAP7_75t_SL g400 ( 
.A(n_324),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_201),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_263),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_263),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_214),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_263),
.B(n_0),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_216),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_203),
.Y(n_407)
);

INVxp33_ASAP7_75t_SL g408 ( 
.A(n_292),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_219),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_263),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_227),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_263),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_228),
.B(n_202),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_352),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_370),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_377),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_221),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_222),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_263),
.Y(n_419)
);

INVx1_ASAP7_75t_SL g420 ( 
.A(n_293),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_263),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_263),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_223),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_293),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_378),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_308),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_308),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_308),
.B(n_1),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_224),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_228),
.B(n_2),
.Y(n_430)
);

INVxp33_ASAP7_75t_SL g431 ( 
.A(n_204),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_308),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_281),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_226),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_230),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_308),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_308),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_209),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_308),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_281),
.Y(n_440)
);

INVxp67_ASAP7_75t_SL g441 ( 
.A(n_324),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_308),
.B(n_2),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_236),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_218),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_260),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_237),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_218),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_218),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_334),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_238),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_243),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_218),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_246),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_249),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_252),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_256),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_218),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_265),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_356),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_268),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_269),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_200),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_270),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_200),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_209),
.Y(n_465)
);

INVxp33_ASAP7_75t_L g466 ( 
.A(n_213),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_213),
.Y(n_467)
);

INVxp33_ASAP7_75t_SL g468 ( 
.A(n_206),
.Y(n_468)
);

INVx1_ASAP7_75t_SL g469 ( 
.A(n_240),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_202),
.B(n_4),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_215),
.Y(n_471)
);

BUFx2_ASAP7_75t_L g472 ( 
.A(n_212),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_271),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_215),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_337),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_275),
.Y(n_476)
);

HB1xp67_ASAP7_75t_L g477 ( 
.A(n_356),
.Y(n_477)
);

INVxp33_ASAP7_75t_L g478 ( 
.A(n_217),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_276),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_217),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_277),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_284),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_285),
.Y(n_483)
);

HB1xp67_ASAP7_75t_L g484 ( 
.A(n_207),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_247),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_225),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_225),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_253),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_253),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_287),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_264),
.Y(n_491)
);

NOR2xp67_ASAP7_75t_L g492 ( 
.A(n_296),
.B(n_5),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_288),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_264),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_274),
.Y(n_495)
);

CKINVDCx16_ASAP7_75t_R g496 ( 
.A(n_205),
.Y(n_496)
);

CKINVDCx16_ASAP7_75t_R g497 ( 
.A(n_205),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_274),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_283),
.Y(n_499)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_208),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_444),
.Y(n_501)
);

INVx3_ASAP7_75t_L g502 ( 
.A(n_485),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_444),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_400),
.B(n_329),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_402),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_402),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_485),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_447),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_408),
.A2(n_420),
.B1(n_440),
.B2(n_433),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_403),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_450),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_447),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_441),
.B(n_329),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_448),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_485),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_448),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_485),
.Y(n_517)
);

AND2x4_ASAP7_75t_L g518 ( 
.A(n_452),
.B(n_351),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_413),
.B(n_351),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_430),
.B(n_452),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_459),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_457),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_457),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_403),
.B(n_295),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_465),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_407),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_410),
.Y(n_527)
);

AND2x4_ASAP7_75t_L g528 ( 
.A(n_410),
.B(n_361),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_412),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_412),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_419),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g532 ( 
.A(n_477),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_419),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_465),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_467),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_467),
.Y(n_536)
);

BUFx8_ASAP7_75t_L g537 ( 
.A(n_472),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_472),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_421),
.B(n_297),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_421),
.B(n_301),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_485),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_475),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_471),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_422),
.Y(n_544)
);

AND2x4_ASAP7_75t_L g545 ( 
.A(n_422),
.B(n_361),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_471),
.Y(n_546)
);

INVxp67_ASAP7_75t_L g547 ( 
.A(n_484),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_474),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_474),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_431),
.B(n_358),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_426),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_451),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_480),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_480),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_486),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_486),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_426),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_427),
.B(n_306),
.Y(n_558)
);

AND2x4_ASAP7_75t_L g559 ( 
.A(n_427),
.B(n_233),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_470),
.A2(n_399),
.B1(n_261),
.B2(n_341),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_432),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_475),
.Y(n_562)
);

CKINVDCx8_ASAP7_75t_R g563 ( 
.A(n_496),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_432),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_487),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_411),
.B(n_310),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_487),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_488),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_436),
.B(n_212),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_488),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_436),
.B(n_250),
.Y(n_571)
);

INVx6_ASAP7_75t_L g572 ( 
.A(n_496),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_491),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_491),
.Y(n_574)
);

AND2x2_ASAP7_75t_L g575 ( 
.A(n_437),
.B(n_250),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_437),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_439),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_439),
.Y(n_578)
);

HB1xp67_ASAP7_75t_L g579 ( 
.A(n_500),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_494),
.B(n_307),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_530),
.Y(n_581)
);

INVx6_ASAP7_75t_L g582 ( 
.A(n_518),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_505),
.Y(n_583)
);

BUFx10_ASAP7_75t_L g584 ( 
.A(n_550),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_504),
.B(n_462),
.Y(n_585)
);

INVxp67_ASAP7_75t_SL g586 ( 
.A(n_502),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_505),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_530),
.Y(n_588)
);

BUFx6f_ASAP7_75t_SL g589 ( 
.A(n_528),
.Y(n_589)
);

AND2x6_ASAP7_75t_L g590 ( 
.A(n_528),
.B(n_233),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_530),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_505),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_505),
.Y(n_593)
);

NOR3xp33_ASAP7_75t_L g594 ( 
.A(n_550),
.B(n_469),
.C(n_497),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_524),
.B(n_401),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_506),
.Y(n_596)
);

INVx2_ASAP7_75t_SL g597 ( 
.A(n_538),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_547),
.B(n_468),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_524),
.B(n_404),
.Y(n_599)
);

BUFx10_ASAP7_75t_L g600 ( 
.A(n_572),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_506),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_538),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_506),
.Y(n_603)
);

OR2x6_ASAP7_75t_L g604 ( 
.A(n_572),
.B(n_296),
.Y(n_604)
);

NAND3xp33_ASAP7_75t_L g605 ( 
.A(n_560),
.B(n_409),
.C(n_406),
.Y(n_605)
);

XNOR2xp5_ASAP7_75t_L g606 ( 
.A(n_566),
.B(n_414),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_506),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_510),
.Y(n_608)
);

INVx4_ASAP7_75t_L g609 ( 
.A(n_577),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_547),
.B(n_417),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_539),
.B(n_418),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_510),
.Y(n_612)
);

AOI22xp33_ASAP7_75t_SL g613 ( 
.A1(n_537),
.A2(n_445),
.B1(n_416),
.B2(n_425),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_539),
.B(n_423),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_507),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_510),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_510),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_540),
.B(n_429),
.Y(n_618)
);

CKINVDCx20_ASAP7_75t_R g619 ( 
.A(n_526),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_520),
.B(n_434),
.Y(n_620)
);

INVx4_ASAP7_75t_L g621 ( 
.A(n_577),
.Y(n_621)
);

BUFx10_ASAP7_75t_L g622 ( 
.A(n_572),
.Y(n_622)
);

OAI22xp33_ASAP7_75t_L g623 ( 
.A1(n_560),
.A2(n_336),
.B1(n_345),
.B2(n_272),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_504),
.B(n_462),
.Y(n_624)
);

AND2x6_ASAP7_75t_L g625 ( 
.A(n_528),
.B(n_359),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_520),
.B(n_435),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_L g627 ( 
.A1(n_528),
.A2(n_405),
.B1(n_442),
.B2(n_428),
.Y(n_627)
);

BUFx2_ASAP7_75t_L g628 ( 
.A(n_521),
.Y(n_628)
);

OAI22xp33_ASAP7_75t_L g629 ( 
.A1(n_579),
.A2(n_357),
.B1(n_375),
.B2(n_348),
.Y(n_629)
);

OR2x2_ASAP7_75t_L g630 ( 
.A(n_521),
.B(n_424),
.Y(n_630)
);

NOR2x1p5_ASAP7_75t_L g631 ( 
.A(n_511),
.B(n_552),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_527),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_540),
.B(n_443),
.Y(n_633)
);

BUFx4f_ASAP7_75t_L g634 ( 
.A(n_577),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_525),
.Y(n_635)
);

NAND3xp33_ASAP7_75t_L g636 ( 
.A(n_580),
.B(n_454),
.C(n_446),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_507),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_507),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_527),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_528),
.A2(n_392),
.B1(n_492),
.B2(n_289),
.Y(n_640)
);

BUFx2_ASAP7_75t_L g641 ( 
.A(n_532),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_545),
.A2(n_519),
.B1(n_571),
.B2(n_569),
.Y(n_642)
);

BUFx3_ASAP7_75t_L g643 ( 
.A(n_518),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_L g644 ( 
.A1(n_545),
.A2(n_392),
.B1(n_289),
.B2(n_299),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_563),
.B(n_456),
.Y(n_645)
);

BUFx10_ASAP7_75t_L g646 ( 
.A(n_572),
.Y(n_646)
);

OR2x2_ASAP7_75t_L g647 ( 
.A(n_532),
.B(n_460),
.Y(n_647)
);

INVxp67_ASAP7_75t_SL g648 ( 
.A(n_502),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_527),
.Y(n_649)
);

BUFx3_ASAP7_75t_L g650 ( 
.A(n_518),
.Y(n_650)
);

BUFx3_ASAP7_75t_L g651 ( 
.A(n_518),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_580),
.B(n_473),
.Y(n_652)
);

OR2x2_ASAP7_75t_L g653 ( 
.A(n_558),
.B(n_479),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_527),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_558),
.B(n_545),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_529),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_529),
.Y(n_657)
);

BUFx3_ASAP7_75t_L g658 ( 
.A(n_518),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_545),
.B(n_481),
.Y(n_659)
);

INVx6_ASAP7_75t_L g660 ( 
.A(n_545),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_529),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_529),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_531),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_519),
.A2(n_299),
.B1(n_302),
.B2(n_283),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_563),
.B(n_490),
.Y(n_665)
);

INVxp67_ASAP7_75t_SL g666 ( 
.A(n_502),
.Y(n_666)
);

INVx5_ASAP7_75t_L g667 ( 
.A(n_577),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_531),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_507),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_531),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_531),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_533),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_504),
.B(n_493),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_533),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_563),
.B(n_449),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_513),
.B(n_391),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_511),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_533),
.Y(n_678)
);

INVx6_ASAP7_75t_L g679 ( 
.A(n_569),
.Y(n_679)
);

BUFx3_ASAP7_75t_L g680 ( 
.A(n_569),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_513),
.B(n_397),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_513),
.B(n_571),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_519),
.Y(n_683)
);

BUFx2_ASAP7_75t_L g684 ( 
.A(n_537),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_571),
.B(n_309),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_575),
.B(n_314),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_575),
.B(n_317),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_533),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_507),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_544),
.Y(n_690)
);

AND2x6_ASAP7_75t_L g691 ( 
.A(n_559),
.B(n_359),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_544),
.Y(n_692)
);

INVxp67_ASAP7_75t_SL g693 ( 
.A(n_502),
.Y(n_693)
);

OR2x2_ASAP7_75t_L g694 ( 
.A(n_579),
.B(n_466),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_578),
.Y(n_695)
);

AND3x2_ASAP7_75t_L g696 ( 
.A(n_575),
.B(n_231),
.C(n_220),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_544),
.B(n_551),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_544),
.Y(n_698)
);

INVx3_ASAP7_75t_L g699 ( 
.A(n_507),
.Y(n_699)
);

NOR2x1p5_ASAP7_75t_L g700 ( 
.A(n_552),
.B(n_210),
.Y(n_700)
);

OR2x6_ASAP7_75t_L g701 ( 
.A(n_572),
.B(n_438),
.Y(n_701)
);

BUFx3_ASAP7_75t_L g702 ( 
.A(n_559),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_551),
.Y(n_703)
);

NAND2xp33_ASAP7_75t_L g704 ( 
.A(n_577),
.B(n_247),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_551),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_551),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_525),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_534),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_534),
.B(n_464),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_578),
.Y(n_710)
);

NAND3xp33_ASAP7_75t_L g711 ( 
.A(n_537),
.B(n_489),
.C(n_229),
.Y(n_711)
);

AND2x6_ASAP7_75t_L g712 ( 
.A(n_559),
.B(n_247),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_557),
.Y(n_713)
);

CKINVDCx20_ASAP7_75t_R g714 ( 
.A(n_526),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_557),
.Y(n_715)
);

INVx3_ASAP7_75t_L g716 ( 
.A(n_507),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_557),
.Y(n_717)
);

INVx3_ASAP7_75t_L g718 ( 
.A(n_507),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_537),
.B(n_453),
.Y(n_719)
);

NAND2xp33_ASAP7_75t_SL g720 ( 
.A(n_535),
.B(n_455),
.Y(n_720)
);

BUFx3_ASAP7_75t_L g721 ( 
.A(n_559),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_557),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_L g723 ( 
.A1(n_559),
.A2(n_564),
.B1(n_576),
.B2(n_561),
.Y(n_723)
);

BUFx2_ASAP7_75t_L g724 ( 
.A(n_537),
.Y(n_724)
);

INVxp67_ASAP7_75t_SL g725 ( 
.A(n_502),
.Y(n_725)
);

BUFx3_ASAP7_75t_L g726 ( 
.A(n_577),
.Y(n_726)
);

INVx4_ASAP7_75t_L g727 ( 
.A(n_577),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_561),
.B(n_323),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_561),
.B(n_331),
.Y(n_729)
);

INVxp67_ASAP7_75t_SL g730 ( 
.A(n_541),
.Y(n_730)
);

NAND2xp33_ASAP7_75t_L g731 ( 
.A(n_577),
.B(n_247),
.Y(n_731)
);

NOR2x1p5_ASAP7_75t_L g732 ( 
.A(n_535),
.B(n_211),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_572),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_679),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_655),
.B(n_247),
.Y(n_735)
);

CKINVDCx8_ASAP7_75t_R g736 ( 
.A(n_677),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_682),
.B(n_509),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_679),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_620),
.B(n_561),
.Y(n_739)
);

NAND2xp33_ASAP7_75t_L g740 ( 
.A(n_590),
.B(n_337),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_682),
.B(n_509),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_626),
.B(n_679),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_673),
.B(n_458),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_679),
.Y(n_744)
);

BUFx5_ASAP7_75t_L g745 ( 
.A(n_590),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_677),
.Y(n_746)
);

INVx4_ASAP7_75t_L g747 ( 
.A(n_660),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_680),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_680),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_642),
.B(n_347),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_652),
.B(n_564),
.Y(n_751)
);

INVxp67_ASAP7_75t_SL g752 ( 
.A(n_723),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_581),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_595),
.B(n_564),
.Y(n_754)
);

AOI22xp5_ASAP7_75t_L g755 ( 
.A1(n_683),
.A2(n_463),
.B1(n_476),
.B2(n_461),
.Y(n_755)
);

NOR2xp67_ASAP7_75t_L g756 ( 
.A(n_605),
.B(n_536),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_683),
.B(n_482),
.Y(n_757)
);

INVx1_ASAP7_75t_SL g758 ( 
.A(n_694),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_599),
.B(n_564),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_653),
.B(n_483),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_653),
.B(n_376),
.Y(n_761)
);

NOR2xp33_ASAP7_75t_L g762 ( 
.A(n_676),
.B(n_478),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_611),
.B(n_576),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_581),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_619),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_614),
.B(n_347),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_618),
.B(n_347),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_633),
.B(n_347),
.Y(n_768)
);

AOI22xp5_ASAP7_75t_L g769 ( 
.A1(n_720),
.A2(n_415),
.B1(n_254),
.B2(n_346),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_643),
.B(n_650),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_SL g771 ( 
.A(n_684),
.B(n_205),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_681),
.A2(n_386),
.B1(n_338),
.B2(n_350),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_597),
.B(n_536),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_588),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_585),
.B(n_576),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_702),
.Y(n_776)
);

NAND3xp33_ASAP7_75t_L g777 ( 
.A(n_598),
.B(n_239),
.C(n_232),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_643),
.B(n_347),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_597),
.B(n_543),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_591),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_702),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_585),
.B(n_576),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_732),
.Y(n_783)
);

NOR2xp67_ASAP7_75t_L g784 ( 
.A(n_636),
.B(n_543),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_624),
.B(n_578),
.Y(n_785)
);

INVx8_ASAP7_75t_L g786 ( 
.A(n_604),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_694),
.B(n_360),
.Y(n_787)
);

NOR2xp33_ASAP7_75t_L g788 ( 
.A(n_659),
.B(n_242),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_624),
.B(n_578),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_721),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_635),
.B(n_542),
.Y(n_791)
);

O2A1O1Ixp33_ASAP7_75t_L g792 ( 
.A1(n_591),
.A2(n_574),
.B(n_573),
.C(n_570),
.Y(n_792)
);

O2A1O1Ixp33_ASAP7_75t_L g793 ( 
.A1(n_685),
.A2(n_574),
.B(n_573),
.C(n_570),
.Y(n_793)
);

NOR3xp33_ASAP7_75t_L g794 ( 
.A(n_623),
.B(n_245),
.C(n_244),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_721),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_686),
.B(n_248),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_583),
.Y(n_797)
);

OAI22xp5_ASAP7_75t_L g798 ( 
.A1(n_627),
.A2(n_363),
.B1(n_335),
.B2(n_333),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_602),
.B(n_546),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_583),
.Y(n_800)
);

AOI22xp5_ASAP7_75t_L g801 ( 
.A1(n_660),
.A2(n_372),
.B1(n_364),
.B2(n_368),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_650),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_707),
.B(n_542),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_708),
.B(n_542),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_687),
.B(n_255),
.Y(n_805)
);

OR2x6_ASAP7_75t_L g806 ( 
.A(n_684),
.B(n_302),
.Y(n_806)
);

AOI22xp5_ASAP7_75t_L g807 ( 
.A1(n_660),
.A2(n_388),
.B1(n_369),
.B2(n_385),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_584),
.B(n_258),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_587),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_587),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_651),
.Y(n_811)
);

INVx3_ASAP7_75t_L g812 ( 
.A(n_651),
.Y(n_812)
);

INVx2_ASAP7_75t_SL g813 ( 
.A(n_647),
.Y(n_813)
);

O2A1O1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_704),
.A2(n_568),
.B(n_567),
.C(n_565),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_658),
.B(n_337),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_728),
.B(n_542),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_729),
.B(n_542),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_590),
.A2(n_320),
.B1(n_398),
.B2(n_393),
.Y(n_818)
);

INVx2_ASAP7_75t_SL g819 ( 
.A(n_647),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_592),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_586),
.B(n_562),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_584),
.B(n_259),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_584),
.B(n_546),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_648),
.B(n_562),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_666),
.B(n_562),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_592),
.Y(n_826)
);

BUFx6f_ASAP7_75t_SL g827 ( 
.A(n_701),
.Y(n_827)
);

OR2x2_ASAP7_75t_L g828 ( 
.A(n_630),
.B(n_566),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_733),
.B(n_305),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_660),
.A2(n_303),
.B1(n_390),
.B2(n_371),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_589),
.A2(n_303),
.B1(n_390),
.B2(n_371),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_658),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_693),
.B(n_562),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_593),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_725),
.B(n_562),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_709),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_619),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_730),
.B(n_503),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_709),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_726),
.B(n_503),
.Y(n_840)
);

OAI221xp5_ASAP7_75t_L g841 ( 
.A1(n_664),
.A2(n_393),
.B1(n_326),
.B2(n_327),
.C(n_332),
.Y(n_841)
);

BUFx6f_ASAP7_75t_L g842 ( 
.A(n_582),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_726),
.B(n_512),
.Y(n_843)
);

INVx8_ASAP7_75t_L g844 ( 
.A(n_604),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_628),
.B(n_548),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_582),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_615),
.B(n_512),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_733),
.B(n_305),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_615),
.B(n_514),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_593),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_596),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_615),
.B(n_514),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_596),
.Y(n_853)
);

HB1xp67_ASAP7_75t_L g854 ( 
.A(n_628),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_610),
.B(n_266),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_701),
.B(n_267),
.Y(n_856)
);

OAI22xp5_ASAP7_75t_L g857 ( 
.A1(n_604),
.A2(n_294),
.B1(n_220),
.B2(n_231),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_634),
.A2(n_517),
.B(n_515),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_582),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_582),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_641),
.Y(n_861)
);

AO22x2_ASAP7_75t_L g862 ( 
.A1(n_719),
.A2(n_566),
.B1(n_235),
.B2(n_234),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_607),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_601),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_637),
.B(n_516),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_601),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_600),
.B(n_337),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_600),
.B(n_337),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_603),
.Y(n_869)
);

BUFx5_ASAP7_75t_L g870 ( 
.A(n_590),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_603),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_701),
.B(n_278),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_637),
.B(n_516),
.Y(n_873)
);

AOI22xp33_ASAP7_75t_L g874 ( 
.A1(n_590),
.A2(n_320),
.B1(n_398),
.B2(n_389),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_637),
.B(n_522),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_L g876 ( 
.A1(n_590),
.A2(n_342),
.B1(n_326),
.B2(n_327),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_612),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_638),
.B(n_669),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_638),
.B(n_522),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_638),
.B(n_523),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_669),
.B(n_523),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_701),
.B(n_279),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_607),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_669),
.B(n_699),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_699),
.B(n_501),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_600),
.B(n_305),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_622),
.B(n_362),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_612),
.Y(n_888)
);

INVx8_ASAP7_75t_L g889 ( 
.A(n_604),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_622),
.B(n_646),
.Y(n_890)
);

NAND2xp33_ASAP7_75t_L g891 ( 
.A(n_590),
.B(n_337),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_699),
.B(n_501),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_716),
.B(n_501),
.Y(n_893)
);

INVxp67_ASAP7_75t_L g894 ( 
.A(n_641),
.Y(n_894)
);

AOI22xp33_ASAP7_75t_L g895 ( 
.A1(n_625),
.A2(n_349),
.B1(n_332),
.B2(n_340),
.Y(n_895)
);

INVx2_ASAP7_75t_SL g896 ( 
.A(n_630),
.Y(n_896)
);

NAND3xp33_ASAP7_75t_SL g897 ( 
.A(n_594),
.B(n_282),
.C(n_280),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_616),
.Y(n_898)
);

A2O1A1Ixp33_ASAP7_75t_L g899 ( 
.A1(n_640),
.A2(n_363),
.B(n_235),
.C(n_241),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_716),
.B(n_718),
.Y(n_900)
);

INVxp67_ASAP7_75t_L g901 ( 
.A(n_606),
.Y(n_901)
);

INVx3_ASAP7_75t_L g902 ( 
.A(n_589),
.Y(n_902)
);

AND2x6_ASAP7_75t_SL g903 ( 
.A(n_714),
.B(n_340),
.Y(n_903)
);

O2A1O1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_704),
.A2(n_568),
.B(n_567),
.C(n_565),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_742),
.A2(n_634),
.B(n_621),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_751),
.A2(n_634),
.B(n_621),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_762),
.B(n_724),
.Y(n_907)
);

AND2x4_ASAP7_75t_L g908 ( 
.A(n_748),
.B(n_711),
.Y(n_908)
);

O2A1O1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_798),
.A2(n_629),
.B(n_665),
.C(n_645),
.Y(n_909)
);

OAI22xp5_ASAP7_75t_L g910 ( 
.A1(n_752),
.A2(n_724),
.B1(n_589),
.B2(n_644),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_753),
.Y(n_911)
);

OAI21xp5_ASAP7_75t_L g912 ( 
.A1(n_754),
.A2(n_697),
.B(n_617),
.Y(n_912)
);

AOI21xp33_ASAP7_75t_L g913 ( 
.A1(n_761),
.A2(n_675),
.B(n_613),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_739),
.A2(n_817),
.B(n_816),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_842),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_758),
.B(n_608),
.Y(n_916)
);

BUFx4f_ASAP7_75t_L g917 ( 
.A(n_786),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_761),
.B(n_762),
.Y(n_918)
);

OAI22xp5_ASAP7_75t_L g919 ( 
.A1(n_759),
.A2(n_335),
.B1(n_234),
.B2(n_241),
.Y(n_919)
);

OAI21xp5_ASAP7_75t_L g920 ( 
.A1(n_763),
.A2(n_617),
.B(n_608),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_775),
.A2(n_621),
.B(n_609),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_745),
.B(n_622),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_753),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_764),
.Y(n_924)
);

BUFx12f_ASAP7_75t_L g925 ( 
.A(n_765),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_782),
.A2(n_727),
.B(n_609),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_743),
.B(n_632),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_785),
.A2(n_727),
.B(n_609),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_796),
.B(n_625),
.Y(n_929)
);

INVx4_ASAP7_75t_L g930 ( 
.A(n_842),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_764),
.Y(n_931)
);

A2O1A1Ixp33_ASAP7_75t_L g932 ( 
.A1(n_796),
.A2(n_353),
.B(n_389),
.C(n_342),
.Y(n_932)
);

NOR2xp67_ASAP7_75t_L g933 ( 
.A(n_755),
.B(n_606),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_789),
.A2(n_727),
.B(n_689),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_890),
.A2(n_689),
.B(n_667),
.Y(n_935)
);

BUFx2_ASAP7_75t_L g936 ( 
.A(n_854),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_774),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_890),
.A2(n_747),
.B(n_878),
.Y(n_938)
);

CKINVDCx14_ASAP7_75t_R g939 ( 
.A(n_837),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_805),
.B(n_625),
.Y(n_940)
);

INVx6_ASAP7_75t_L g941 ( 
.A(n_786),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_774),
.Y(n_942)
);

AOI22xp5_ASAP7_75t_L g943 ( 
.A1(n_743),
.A2(n_625),
.B1(n_691),
.B2(n_700),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_SL g944 ( 
.A(n_745),
.B(n_646),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_842),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_747),
.A2(n_689),
.B(n_667),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_780),
.Y(n_947)
);

AOI21x1_ASAP7_75t_L g948 ( 
.A1(n_867),
.A2(n_639),
.B(n_632),
.Y(n_948)
);

INVx4_ASAP7_75t_L g949 ( 
.A(n_842),
.Y(n_949)
);

OAI21xp5_ASAP7_75t_L g950 ( 
.A1(n_735),
.A2(n_750),
.B(n_884),
.Y(n_950)
);

NOR2xp67_ASAP7_75t_L g951 ( 
.A(n_777),
.B(n_548),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_780),
.Y(n_952)
);

NOR3xp33_ASAP7_75t_L g953 ( 
.A(n_760),
.B(n_257),
.C(n_251),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_900),
.A2(n_689),
.B(n_667),
.Y(n_954)
);

INVxp67_ASAP7_75t_L g955 ( 
.A(n_861),
.Y(n_955)
);

NOR2x1_ASAP7_75t_L g956 ( 
.A(n_897),
.B(n_631),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_813),
.B(n_639),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_805),
.B(n_625),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_797),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_749),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_770),
.A2(n_689),
.B(n_667),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_745),
.B(n_646),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_770),
.A2(n_667),
.B(n_731),
.Y(n_963)
);

A2O1A1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_788),
.A2(n_251),
.B(n_333),
.C(n_257),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_788),
.B(n_625),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_773),
.B(n_625),
.Y(n_966)
);

NAND3xp33_ASAP7_75t_SL g967 ( 
.A(n_855),
.B(n_822),
.C(n_808),
.Y(n_967)
);

AO21x1_ASAP7_75t_L g968 ( 
.A1(n_750),
.A2(n_273),
.B(n_262),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_821),
.A2(n_731),
.B(n_718),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_776),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_819),
.B(n_654),
.Y(n_971)
);

AOI21x1_ASAP7_75t_L g972 ( 
.A1(n_867),
.A2(n_656),
.B(n_654),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_779),
.B(n_656),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_737),
.B(n_741),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_824),
.A2(n_718),
.B(n_716),
.Y(n_975)
);

OAI21xp5_ASAP7_75t_L g976 ( 
.A1(n_735),
.A2(n_662),
.B(n_661),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_845),
.B(n_799),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_781),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_797),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_836),
.B(n_839),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_902),
.Y(n_981)
);

OAI21xp5_ASAP7_75t_L g982 ( 
.A1(n_815),
.A2(n_662),
.B(n_661),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_823),
.B(n_722),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_R g984 ( 
.A(n_746),
.B(n_714),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_812),
.B(n_668),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_812),
.B(n_668),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_734),
.B(n_722),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_825),
.A2(n_835),
.B(n_833),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_896),
.B(n_670),
.Y(n_989)
);

OAI21xp5_ASAP7_75t_L g990 ( 
.A1(n_815),
.A2(n_672),
.B(n_670),
.Y(n_990)
);

NAND2xp33_ASAP7_75t_L g991 ( 
.A(n_745),
.B(n_691),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_SL g992 ( 
.A(n_745),
.B(n_616),
.Y(n_992)
);

BUFx2_ASAP7_75t_L g993 ( 
.A(n_894),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_800),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_738),
.B(n_672),
.Y(n_995)
);

AOI21xp33_ASAP7_75t_L g996 ( 
.A1(n_855),
.A2(n_760),
.B(n_808),
.Y(n_996)
);

INVx3_ASAP7_75t_L g997 ( 
.A(n_846),
.Y(n_997)
);

INVx3_ASAP7_75t_L g998 ( 
.A(n_859),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_860),
.A2(n_657),
.B(n_649),
.Y(n_999)
);

INVx4_ASAP7_75t_L g1000 ( 
.A(n_902),
.Y(n_1000)
);

O2A1O1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_899),
.A2(n_703),
.B(n_715),
.C(n_713),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_744),
.B(n_674),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_840),
.A2(n_657),
.B(n_649),
.Y(n_1003)
);

NAND2x1_ASAP7_75t_L g1004 ( 
.A(n_800),
.B(n_691),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_790),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_786),
.Y(n_1006)
);

AND2x2_ASAP7_75t_SL g1007 ( 
.A(n_771),
.B(n_262),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_822),
.B(n_549),
.Y(n_1008)
);

NAND2xp33_ASAP7_75t_L g1009 ( 
.A(n_745),
.B(n_691),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_901),
.Y(n_1010)
);

AOI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_756),
.A2(n_691),
.B1(n_712),
.B2(n_713),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_843),
.A2(n_671),
.B(n_663),
.Y(n_1012)
);

INVxp67_ASAP7_75t_L g1013 ( 
.A(n_856),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_868),
.A2(n_671),
.B(n_663),
.Y(n_1014)
);

INVx1_ASAP7_75t_SL g1015 ( 
.A(n_828),
.Y(n_1015)
);

O2A1O1Ixp33_ASAP7_75t_SL g1016 ( 
.A1(n_766),
.A2(n_273),
.B(n_328),
.C(n_294),
.Y(n_1016)
);

OAI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_793),
.A2(n_678),
.B(n_674),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_795),
.B(n_678),
.Y(n_1018)
);

OAI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_885),
.A2(n_692),
.B(n_688),
.Y(n_1019)
);

A2O1A1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_841),
.A2(n_349),
.B(n_353),
.C(n_328),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_868),
.A2(n_717),
.B(n_690),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_757),
.B(n_549),
.Y(n_1022)
);

AND2x4_ASAP7_75t_L g1023 ( 
.A(n_783),
.B(n_696),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_802),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_811),
.Y(n_1025)
);

OAI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_892),
.A2(n_688),
.B(n_715),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_832),
.Y(n_1027)
);

AO22x1_ASAP7_75t_L g1028 ( 
.A1(n_794),
.A2(n_291),
.B1(n_286),
.B2(n_290),
.Y(n_1028)
);

BUFx6f_ASAP7_75t_L g1029 ( 
.A(n_844),
.Y(n_1029)
);

INVx2_ASAP7_75t_SL g1030 ( 
.A(n_787),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_856),
.B(n_553),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_784),
.B(n_692),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_740),
.A2(n_717),
.B(n_690),
.Y(n_1033)
);

INVx1_ASAP7_75t_SL g1034 ( 
.A(n_903),
.Y(n_1034)
);

OAI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_818),
.A2(n_698),
.B1(n_706),
.B2(n_705),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_809),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_872),
.B(n_553),
.Y(n_1037)
);

NOR3xp33_ASAP7_75t_L g1038 ( 
.A(n_872),
.B(n_554),
.C(n_555),
.Y(n_1038)
);

BUFx8_ASAP7_75t_L g1039 ( 
.A(n_827),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_838),
.B(n_698),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_809),
.Y(n_1041)
);

CKINVDCx14_ASAP7_75t_R g1042 ( 
.A(n_769),
.Y(n_1042)
);

O2A1O1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_792),
.A2(n_706),
.B(n_705),
.C(n_703),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_863),
.B(n_695),
.Y(n_1044)
);

INVx4_ASAP7_75t_L g1045 ( 
.A(n_844),
.Y(n_1045)
);

INVxp67_ASAP7_75t_L g1046 ( 
.A(n_882),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_893),
.A2(n_710),
.B(n_695),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_883),
.B(n_710),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_810),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_891),
.A2(n_515),
.B(n_517),
.Y(n_1050)
);

OAI22xp5_ASAP7_75t_L g1051 ( 
.A1(n_818),
.A2(n_554),
.B1(n_555),
.B2(n_556),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_810),
.Y(n_1052)
);

A2O1A1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_882),
.A2(n_556),
.B(n_508),
.C(n_298),
.Y(n_1053)
);

OAI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_820),
.A2(n_691),
.B(n_712),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_847),
.A2(n_517),
.B(n_515),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_820),
.Y(n_1056)
);

AO21x1_ASAP7_75t_L g1057 ( 
.A1(n_766),
.A2(n_508),
.B(n_495),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_826),
.Y(n_1058)
);

HB1xp67_ASAP7_75t_L g1059 ( 
.A(n_806),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_834),
.Y(n_1060)
);

OR2x6_ASAP7_75t_SL g1061 ( 
.A(n_857),
.B(n_300),
.Y(n_1061)
);

BUFx6f_ASAP7_75t_L g1062 ( 
.A(n_844),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_829),
.B(n_304),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_806),
.B(n_494),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_849),
.A2(n_517),
.B(n_515),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_834),
.Y(n_1066)
);

A2O1A1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_874),
.A2(n_498),
.B(n_495),
.C(n_499),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_852),
.A2(n_515),
.B(n_517),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_850),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_848),
.B(n_311),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_865),
.A2(n_515),
.B(n_517),
.Y(n_1071)
);

OAI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_850),
.A2(n_691),
.B(n_712),
.Y(n_1072)
);

INVxp67_ASAP7_75t_L g1073 ( 
.A(n_806),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_873),
.A2(n_517),
.B(n_515),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_851),
.B(n_712),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_851),
.B(n_712),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_889),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_889),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_853),
.B(n_712),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_853),
.Y(n_1080)
);

AND2x2_ASAP7_75t_L g1081 ( 
.A(n_862),
.B(n_498),
.Y(n_1081)
);

OAI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_864),
.A2(n_869),
.B(n_866),
.Y(n_1082)
);

OAI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_864),
.A2(n_712),
.B(n_508),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_866),
.B(n_541),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_869),
.B(n_541),
.Y(n_1085)
);

AOI22xp33_ASAP7_75t_L g1086 ( 
.A1(n_874),
.A2(n_337),
.B1(n_362),
.B2(n_312),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_862),
.B(n_499),
.Y(n_1087)
);

O2A1O1Ixp33_ASAP7_75t_L g1088 ( 
.A1(n_778),
.A2(n_464),
.B(n_541),
.C(n_362),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_875),
.A2(n_517),
.B(n_515),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_SL g1090 ( 
.A(n_870),
.B(n_337),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_772),
.B(n_313),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_871),
.Y(n_1092)
);

A2O1A1Ixp33_ASAP7_75t_SL g1093 ( 
.A1(n_918),
.A2(n_904),
.B(n_814),
.C(n_831),
.Y(n_1093)
);

NOR2xp67_ASAP7_75t_SL g1094 ( 
.A(n_1006),
.B(n_886),
.Y(n_1094)
);

AOI21x1_ASAP7_75t_L g1095 ( 
.A1(n_938),
.A2(n_905),
.B(n_914),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_918),
.B(n_887),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_911),
.Y(n_1097)
);

OAI21xp33_ASAP7_75t_L g1098 ( 
.A1(n_996),
.A2(n_862),
.B(n_895),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_929),
.A2(n_778),
.B(n_767),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_977),
.B(n_876),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_974),
.B(n_1008),
.Y(n_1101)
);

BUFx3_ASAP7_75t_L g1102 ( 
.A(n_936),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_974),
.B(n_801),
.Y(n_1103)
);

AND2x2_ASAP7_75t_L g1104 ( 
.A(n_907),
.B(n_767),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_931),
.Y(n_1105)
);

INVx2_ASAP7_75t_SL g1106 ( 
.A(n_993),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_1013),
.B(n_807),
.Y(n_1107)
);

HB1xp67_ASAP7_75t_L g1108 ( 
.A(n_955),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_940),
.A2(n_768),
.B(n_880),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_909),
.A2(n_768),
.B(n_830),
.C(n_889),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_1031),
.B(n_876),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_927),
.B(n_895),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_958),
.A2(n_881),
.B(n_879),
.Y(n_1113)
);

NAND2x1p5_ASAP7_75t_L g1114 ( 
.A(n_1045),
.B(n_871),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_1013),
.B(n_791),
.Y(n_1115)
);

OAI21xp33_ASAP7_75t_L g1116 ( 
.A1(n_1091),
.A2(n_374),
.B(n_316),
.Y(n_1116)
);

O2A1O1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_967),
.A2(n_953),
.B(n_913),
.C(n_932),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_927),
.B(n_877),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_1046),
.A2(n_804),
.B1(n_803),
.B2(n_877),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1037),
.B(n_888),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_983),
.B(n_888),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1041),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_1046),
.B(n_898),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_967),
.B(n_955),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_991),
.A2(n_858),
.B(n_898),
.Y(n_1125)
);

INVx1_ASAP7_75t_SL g1126 ( 
.A(n_1015),
.Y(n_1126)
);

NAND2x1p5_ASAP7_75t_L g1127 ( 
.A(n_1045),
.B(n_870),
.Y(n_1127)
);

BUFx8_ASAP7_75t_L g1128 ( 
.A(n_925),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_966),
.A2(n_870),
.B1(n_366),
.B2(n_396),
.Y(n_1129)
);

NOR2x1_ASAP7_75t_L g1130 ( 
.A(n_1000),
.B(n_541),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_1041),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_1064),
.B(n_315),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_916),
.B(n_973),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_916),
.B(n_870),
.Y(n_1134)
);

BUFx2_ASAP7_75t_SL g1135 ( 
.A(n_1006),
.Y(n_1135)
);

BUFx3_ASAP7_75t_L g1136 ( 
.A(n_1039),
.Y(n_1136)
);

INVxp67_ASAP7_75t_L g1137 ( 
.A(n_1022),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_923),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_984),
.Y(n_1139)
);

AND2x2_ASAP7_75t_SL g1140 ( 
.A(n_1007),
.B(n_5),
.Y(n_1140)
);

O2A1O1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_953),
.A2(n_318),
.B(n_319),
.C(n_321),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1009),
.A2(n_870),
.B(n_395),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_980),
.B(n_957),
.Y(n_1143)
);

O2A1O1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_932),
.A2(n_322),
.B(n_325),
.C(n_330),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_924),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_SL g1146 ( 
.A(n_1007),
.B(n_1030),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_937),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_947),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_965),
.A2(n_870),
.B(n_394),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_SL g1150 ( 
.A(n_908),
.B(n_339),
.Y(n_1150)
);

AOI21xp5_ASAP7_75t_L g1151 ( 
.A1(n_950),
.A2(n_387),
.B(n_384),
.Y(n_1151)
);

AOI22xp33_ASAP7_75t_L g1152 ( 
.A1(n_1091),
.A2(n_383),
.B1(n_382),
.B2(n_381),
.Y(n_1152)
);

NOR2xp67_ASAP7_75t_L g1153 ( 
.A(n_1010),
.B(n_81),
.Y(n_1153)
);

AOI22xp33_ASAP7_75t_L g1154 ( 
.A1(n_1038),
.A2(n_380),
.B1(n_379),
.B2(n_373),
.Y(n_1154)
);

A2O1A1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_1063),
.A2(n_367),
.B(n_365),
.C(n_355),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_908),
.B(n_354),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_R g1157 ( 
.A(n_939),
.B(n_344),
.Y(n_1157)
);

OR2x6_ASAP7_75t_L g1158 ( 
.A(n_941),
.B(n_83),
.Y(n_1158)
);

A2O1A1Ixp33_ASAP7_75t_L g1159 ( 
.A1(n_1063),
.A2(n_343),
.B(n_8),
.C(n_9),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_988),
.A2(n_84),
.B(n_198),
.Y(n_1160)
);

NAND2xp33_ASAP7_75t_R g1161 ( 
.A(n_984),
.B(n_82),
.Y(n_1161)
);

OAI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_920),
.A2(n_199),
.B(n_195),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_957),
.B(n_6),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_942),
.Y(n_1164)
);

NOR2x1_ASAP7_75t_SL g1165 ( 
.A(n_915),
.B(n_186),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_906),
.A2(n_944),
.B(n_922),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_971),
.B(n_10),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_922),
.A2(n_128),
.B(n_177),
.Y(n_1168)
);

AND2x2_ASAP7_75t_L g1169 ( 
.A(n_1081),
.B(n_10),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_971),
.B(n_13),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_981),
.B(n_178),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_944),
.A2(n_125),
.B(n_166),
.Y(n_1172)
);

A2O1A1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_1070),
.A2(n_13),
.B(n_15),
.C(n_21),
.Y(n_1173)
);

AOI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1070),
.A2(n_169),
.B1(n_164),
.B2(n_162),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_962),
.A2(n_159),
.B(n_153),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_962),
.A2(n_150),
.B(n_140),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_1042),
.B(n_21),
.Y(n_1177)
);

INVx3_ASAP7_75t_L g1178 ( 
.A(n_915),
.Y(n_1178)
);

AND2x2_ASAP7_75t_L g1179 ( 
.A(n_1087),
.B(n_22),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_L g1180 ( 
.A(n_1073),
.B(n_27),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_981),
.B(n_129),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_989),
.B(n_27),
.Y(n_1182)
);

NOR2xp67_ASAP7_75t_SL g1183 ( 
.A(n_1006),
.B(n_1029),
.Y(n_1183)
);

O2A1O1Ixp5_ASAP7_75t_L g1184 ( 
.A1(n_1090),
.A2(n_123),
.B(n_121),
.C(n_120),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_952),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_981),
.B(n_105),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_989),
.B(n_30),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_934),
.A2(n_98),
.B(n_97),
.Y(n_1188)
);

A2O1A1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_1053),
.A2(n_30),
.B(n_32),
.C(n_35),
.Y(n_1189)
);

AOI21xp33_ASAP7_75t_L g1190 ( 
.A1(n_910),
.A2(n_37),
.B(n_39),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1038),
.B(n_41),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_981),
.B(n_102),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_1073),
.B(n_41),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_921),
.A2(n_92),
.B(n_45),
.Y(n_1194)
);

BUFx3_ASAP7_75t_L g1195 ( 
.A(n_1039),
.Y(n_1195)
);

O2A1O1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_964),
.A2(n_42),
.B(n_47),
.C(n_50),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_L g1197 ( 
.A(n_960),
.B(n_52),
.Y(n_1197)
);

BUFx6f_ASAP7_75t_L g1198 ( 
.A(n_1029),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_SL g1199 ( 
.A(n_1029),
.B(n_56),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_926),
.A2(n_57),
.B(n_59),
.Y(n_1200)
);

INVx5_ASAP7_75t_L g1201 ( 
.A(n_915),
.Y(n_1201)
);

O2A1O1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_919),
.A2(n_57),
.B(n_59),
.C(n_61),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_970),
.B(n_61),
.Y(n_1203)
);

AOI22x1_ASAP7_75t_L g1204 ( 
.A1(n_969),
.A2(n_69),
.B1(n_71),
.B2(n_72),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1059),
.B(n_69),
.Y(n_1205)
);

NAND2x1p5_ASAP7_75t_L g1206 ( 
.A(n_1029),
.B(n_71),
.Y(n_1206)
);

BUFx6f_ASAP7_75t_L g1207 ( 
.A(n_1062),
.Y(n_1207)
);

BUFx6f_ASAP7_75t_L g1208 ( 
.A(n_1062),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_928),
.A2(n_73),
.B(n_1019),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_1062),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1040),
.A2(n_992),
.B(n_985),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1026),
.A2(n_912),
.B(n_1033),
.Y(n_1212)
);

INVx5_ASAP7_75t_L g1213 ( 
.A(n_915),
.Y(n_1213)
);

NOR2xp67_ASAP7_75t_SL g1214 ( 
.A(n_1062),
.B(n_1077),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_978),
.B(n_1005),
.Y(n_1215)
);

OA21x2_ASAP7_75t_L g1216 ( 
.A1(n_1017),
.A2(n_976),
.B(n_982),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1056),
.Y(n_1217)
);

OR2x2_ASAP7_75t_L g1218 ( 
.A(n_933),
.B(n_1024),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_SL g1219 ( 
.A(n_1077),
.B(n_1078),
.Y(n_1219)
);

AOI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1090),
.A2(n_972),
.B(n_948),
.Y(n_1220)
);

INVx2_ASAP7_75t_L g1221 ( 
.A(n_959),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_R g1222 ( 
.A(n_917),
.B(n_1077),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1058),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_L g1224 ( 
.A(n_1025),
.B(n_1027),
.Y(n_1224)
);

AOI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_951),
.A2(n_956),
.B1(n_943),
.B2(n_941),
.Y(n_1225)
);

INVx6_ASAP7_75t_L g1226 ( 
.A(n_1077),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_979),
.B(n_994),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_L g1228 ( 
.A(n_1061),
.B(n_1028),
.Y(n_1228)
);

AOI22x1_ASAP7_75t_L g1229 ( 
.A1(n_963),
.A2(n_975),
.B1(n_1052),
.B2(n_1066),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_SL g1230 ( 
.A(n_917),
.B(n_1034),
.Y(n_1230)
);

NOR2xp67_ASAP7_75t_SL g1231 ( 
.A(n_1078),
.B(n_941),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_986),
.A2(n_992),
.B(n_1032),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1023),
.B(n_1078),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1047),
.A2(n_1021),
.B(n_1014),
.Y(n_1234)
);

NAND2xp33_ASAP7_75t_SL g1235 ( 
.A(n_1078),
.B(n_1000),
.Y(n_1235)
);

BUFx2_ASAP7_75t_L g1236 ( 
.A(n_945),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_997),
.A2(n_998),
.B1(n_945),
.B2(n_1018),
.Y(n_1237)
);

O2A1O1Ixp33_ASAP7_75t_L g1238 ( 
.A1(n_1020),
.A2(n_1051),
.B(n_1016),
.C(n_1067),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1036),
.B(n_1049),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1080),
.B(n_1092),
.Y(n_1240)
);

O2A1O1Ixp33_ASAP7_75t_L g1241 ( 
.A1(n_1020),
.A2(n_1016),
.B(n_1067),
.C(n_1043),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_SL g1242 ( 
.A(n_945),
.B(n_997),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1060),
.B(n_1069),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_987),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_995),
.Y(n_1245)
);

A2O1A1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_1001),
.A2(n_1011),
.B(n_990),
.C(n_1054),
.Y(n_1246)
);

BUFx6f_ASAP7_75t_L g1247 ( 
.A(n_945),
.Y(n_1247)
);

OAI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1002),
.A2(n_1044),
.B1(n_1048),
.B2(n_930),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_SL g1249 ( 
.A(n_930),
.B(n_949),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1082),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1212),
.A2(n_1004),
.B(n_946),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1125),
.A2(n_1012),
.B(n_1003),
.Y(n_1252)
);

CKINVDCx16_ASAP7_75t_R g1253 ( 
.A(n_1157),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_SL g1254 ( 
.A(n_1101),
.B(n_949),
.Y(n_1254)
);

AND2x4_ASAP7_75t_L g1255 ( 
.A(n_1233),
.B(n_1072),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1133),
.B(n_1086),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1212),
.A2(n_1211),
.B(n_1113),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1113),
.A2(n_1099),
.B(n_1134),
.Y(n_1258)
);

AO31x2_ASAP7_75t_L g1259 ( 
.A1(n_1209),
.A2(n_1057),
.A3(n_968),
.B(n_1035),
.Y(n_1259)
);

AO31x2_ASAP7_75t_L g1260 ( 
.A1(n_1209),
.A2(n_935),
.A3(n_961),
.B(n_999),
.Y(n_1260)
);

INVx2_ASAP7_75t_SL g1261 ( 
.A(n_1102),
.Y(n_1261)
);

O2A1O1Ixp33_ASAP7_75t_L g1262 ( 
.A1(n_1096),
.A2(n_1117),
.B(n_1159),
.C(n_1190),
.Y(n_1262)
);

INVx1_ASAP7_75t_SL g1263 ( 
.A(n_1126),
.Y(n_1263)
);

INVx3_ASAP7_75t_L g1264 ( 
.A(n_1198),
.Y(n_1264)
);

AO31x2_ASAP7_75t_L g1265 ( 
.A1(n_1234),
.A2(n_1089),
.A3(n_1074),
.B(n_1055),
.Y(n_1265)
);

AO31x2_ASAP7_75t_L g1266 ( 
.A1(n_1234),
.A2(n_1065),
.A3(n_1068),
.B(n_1071),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1143),
.B(n_1086),
.Y(n_1267)
);

HB1xp67_ASAP7_75t_L g1268 ( 
.A(n_1106),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1099),
.A2(n_954),
.B(n_1083),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1125),
.A2(n_1050),
.B(n_1084),
.Y(n_1270)
);

INVx8_ASAP7_75t_L g1271 ( 
.A(n_1201),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1229),
.A2(n_1085),
.B(n_1076),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1223),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1221),
.Y(n_1274)
);

O2A1O1Ixp33_ASAP7_75t_L g1275 ( 
.A1(n_1173),
.A2(n_1088),
.B(n_1075),
.C(n_1079),
.Y(n_1275)
);

AOI21xp33_ASAP7_75t_L g1276 ( 
.A1(n_1098),
.A2(n_1103),
.B(n_1124),
.Y(n_1276)
);

OAI221xp5_ASAP7_75t_L g1277 ( 
.A1(n_1152),
.A2(n_1116),
.B1(n_1150),
.B2(n_1156),
.C(n_1155),
.Y(n_1277)
);

HB1xp67_ASAP7_75t_L g1278 ( 
.A(n_1108),
.Y(n_1278)
);

AO31x2_ASAP7_75t_L g1279 ( 
.A1(n_1246),
.A2(n_1166),
.A3(n_1109),
.B(n_1149),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1097),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1105),
.Y(n_1281)
);

NAND3xp33_ASAP7_75t_L g1282 ( 
.A(n_1191),
.B(n_1141),
.C(n_1189),
.Y(n_1282)
);

INVx3_ASAP7_75t_L g1283 ( 
.A(n_1198),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1111),
.B(n_1137),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1109),
.A2(n_1166),
.B(n_1118),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1232),
.A2(n_1149),
.B(n_1216),
.Y(n_1286)
);

OA21x2_ASAP7_75t_L g1287 ( 
.A1(n_1232),
.A2(n_1162),
.B(n_1095),
.Y(n_1287)
);

AOI21xp5_ASAP7_75t_L g1288 ( 
.A1(n_1216),
.A2(n_1110),
.B(n_1120),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1244),
.B(n_1245),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1142),
.A2(n_1112),
.B(n_1248),
.Y(n_1290)
);

AO31x2_ASAP7_75t_L g1291 ( 
.A1(n_1194),
.A2(n_1200),
.A3(n_1250),
.B(n_1119),
.Y(n_1291)
);

NOR4xp25_ASAP7_75t_L g1292 ( 
.A(n_1202),
.B(n_1196),
.C(n_1167),
.D(n_1170),
.Y(n_1292)
);

AO31x2_ASAP7_75t_L g1293 ( 
.A1(n_1194),
.A2(n_1200),
.A3(n_1160),
.B(n_1237),
.Y(n_1293)
);

CKINVDCx16_ASAP7_75t_R g1294 ( 
.A(n_1136),
.Y(n_1294)
);

AO221x1_ASAP7_75t_L g1295 ( 
.A1(n_1129),
.A2(n_1247),
.B1(n_1178),
.B2(n_1198),
.C(n_1207),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_1148),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1215),
.Y(n_1297)
);

INVx2_ASAP7_75t_L g1298 ( 
.A(n_1138),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_1107),
.B(n_1218),
.Y(n_1299)
);

INVx5_ASAP7_75t_L g1300 ( 
.A(n_1158),
.Y(n_1300)
);

NAND3xp33_ASAP7_75t_SL g1301 ( 
.A(n_1177),
.B(n_1154),
.C(n_1228),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1115),
.B(n_1123),
.Y(n_1302)
);

O2A1O1Ixp33_ASAP7_75t_SL g1303 ( 
.A1(n_1093),
.A2(n_1192),
.B(n_1181),
.C(n_1171),
.Y(n_1303)
);

AO32x2_ASAP7_75t_L g1304 ( 
.A1(n_1204),
.A2(n_1140),
.A3(n_1241),
.B1(n_1238),
.B2(n_1144),
.Y(n_1304)
);

AO32x2_ASAP7_75t_L g1305 ( 
.A1(n_1163),
.A2(n_1187),
.A3(n_1182),
.B1(n_1151),
.B2(n_1104),
.Y(n_1305)
);

A2O1A1Ixp33_ASAP7_75t_L g1306 ( 
.A1(n_1151),
.A2(n_1225),
.B(n_1100),
.C(n_1146),
.Y(n_1306)
);

A2O1A1Ixp33_ASAP7_75t_L g1307 ( 
.A1(n_1224),
.A2(n_1160),
.B(n_1197),
.C(n_1175),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1145),
.Y(n_1308)
);

AOI221x1_ASAP7_75t_L g1309 ( 
.A1(n_1188),
.A2(n_1172),
.B1(n_1168),
.B2(n_1175),
.C(n_1176),
.Y(n_1309)
);

OAI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1142),
.A2(n_1188),
.B(n_1176),
.Y(n_1310)
);

OAI21xp33_ASAP7_75t_SL g1311 ( 
.A1(n_1158),
.A2(n_1203),
.B(n_1243),
.Y(n_1311)
);

O2A1O1Ixp33_ASAP7_75t_SL g1312 ( 
.A1(n_1186),
.A2(n_1242),
.B(n_1199),
.C(n_1172),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1121),
.A2(n_1235),
.B(n_1168),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1169),
.B(n_1179),
.Y(n_1314)
);

OAI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1184),
.A2(n_1220),
.B(n_1240),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1127),
.A2(n_1130),
.B(n_1114),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1127),
.A2(n_1114),
.B(n_1239),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1201),
.A2(n_1213),
.B(n_1249),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1201),
.A2(n_1213),
.B(n_1227),
.Y(n_1319)
);

AOI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1094),
.A2(n_1185),
.B(n_1219),
.Y(n_1320)
);

AOI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1147),
.A2(n_1164),
.B(n_1131),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1178),
.A2(n_1122),
.B(n_1206),
.Y(n_1322)
);

INVxp67_ASAP7_75t_L g1323 ( 
.A(n_1205),
.Y(n_1323)
);

OAI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1174),
.A2(n_1193),
.B(n_1180),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1201),
.A2(n_1213),
.B(n_1165),
.Y(n_1325)
);

BUFx6f_ASAP7_75t_L g1326 ( 
.A(n_1207),
.Y(n_1326)
);

OA21x2_ASAP7_75t_L g1327 ( 
.A1(n_1236),
.A2(n_1132),
.B(n_1153),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_SL g1328 ( 
.A(n_1139),
.B(n_1222),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1206),
.A2(n_1183),
.B(n_1214),
.Y(n_1329)
);

AO31x2_ASAP7_75t_L g1330 ( 
.A1(n_1247),
.A2(n_1231),
.A3(n_1161),
.B(n_1135),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_SL g1331 ( 
.A1(n_1207),
.A2(n_1208),
.B(n_1210),
.Y(n_1331)
);

INVx6_ASAP7_75t_L g1332 ( 
.A(n_1128),
.Y(n_1332)
);

AO31x2_ASAP7_75t_L g1333 ( 
.A1(n_1247),
.A2(n_1226),
.A3(n_1208),
.B(n_1210),
.Y(n_1333)
);

AO32x2_ASAP7_75t_L g1334 ( 
.A1(n_1226),
.A2(n_1208),
.A3(n_1210),
.B1(n_1230),
.B2(n_1195),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_SL g1335 ( 
.A(n_1128),
.B(n_1226),
.Y(n_1335)
);

AND2x2_ASAP7_75t_SL g1336 ( 
.A(n_1140),
.B(n_1007),
.Y(n_1336)
);

AOI221x1_ASAP7_75t_L g1337 ( 
.A1(n_1190),
.A2(n_996),
.B1(n_953),
.B2(n_967),
.C(n_1098),
.Y(n_1337)
);

AO31x2_ASAP7_75t_L g1338 ( 
.A1(n_1209),
.A2(n_1212),
.A3(n_1234),
.B(n_1246),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1132),
.B(n_974),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1217),
.Y(n_1340)
);

OAI22x1_ASAP7_75t_L g1341 ( 
.A1(n_1096),
.A2(n_918),
.B1(n_1228),
.B2(n_1046),
.Y(n_1341)
);

NAND2xp33_ASAP7_75t_L g1342 ( 
.A(n_1222),
.B(n_1112),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1125),
.A2(n_1229),
.B(n_1220),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1221),
.Y(n_1344)
);

AND2x4_ASAP7_75t_L g1345 ( 
.A(n_1233),
.B(n_1045),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_SL g1346 ( 
.A1(n_1162),
.A2(n_890),
.B(n_1110),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1221),
.Y(n_1347)
);

BUFx12f_ASAP7_75t_L g1348 ( 
.A(n_1128),
.Y(n_1348)
);

INVx4_ASAP7_75t_L g1349 ( 
.A(n_1198),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1217),
.Y(n_1350)
);

AO31x2_ASAP7_75t_L g1351 ( 
.A1(n_1209),
.A2(n_1212),
.A3(n_1234),
.B(n_1246),
.Y(n_1351)
);

AOI21xp5_ASAP7_75t_L g1352 ( 
.A1(n_1212),
.A2(n_1009),
.B(n_991),
.Y(n_1352)
);

AOI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1140),
.A2(n_918),
.B1(n_974),
.B2(n_967),
.Y(n_1353)
);

CKINVDCx20_ASAP7_75t_R g1354 ( 
.A(n_1128),
.Y(n_1354)
);

INVx2_ASAP7_75t_L g1355 ( 
.A(n_1221),
.Y(n_1355)
);

AOI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1140),
.A2(n_918),
.B1(n_974),
.B2(n_967),
.Y(n_1356)
);

O2A1O1Ixp5_ASAP7_75t_L g1357 ( 
.A1(n_1209),
.A2(n_996),
.B(n_918),
.C(n_1096),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1125),
.A2(n_1229),
.B(n_1220),
.Y(n_1358)
);

A2O1A1Ixp33_ASAP7_75t_L g1359 ( 
.A1(n_1117),
.A2(n_918),
.B(n_996),
.C(n_1096),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1212),
.A2(n_1009),
.B(n_991),
.Y(n_1360)
);

O2A1O1Ixp5_ASAP7_75t_SL g1361 ( 
.A1(n_1190),
.A2(n_996),
.B(n_798),
.C(n_766),
.Y(n_1361)
);

INVx1_ASAP7_75t_SL g1362 ( 
.A(n_1126),
.Y(n_1362)
);

BUFx6f_ASAP7_75t_L g1363 ( 
.A(n_1198),
.Y(n_1363)
);

AOI21xp33_ASAP7_75t_L g1364 ( 
.A1(n_1117),
.A2(n_918),
.B(n_996),
.Y(n_1364)
);

AOI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1140),
.A2(n_918),
.B1(n_996),
.B2(n_967),
.Y(n_1365)
);

OR2x6_ASAP7_75t_L g1366 ( 
.A(n_1158),
.B(n_1135),
.Y(n_1366)
);

AOI221x1_ASAP7_75t_L g1367 ( 
.A1(n_1190),
.A2(n_996),
.B1(n_953),
.B2(n_967),
.C(n_1098),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1125),
.A2(n_1229),
.B(n_1220),
.Y(n_1368)
);

NOR2x1_ASAP7_75t_L g1369 ( 
.A(n_1101),
.B(n_967),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1101),
.B(n_918),
.Y(n_1370)
);

NOR2xp67_ASAP7_75t_SL g1371 ( 
.A(n_1135),
.B(n_736),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1125),
.A2(n_1229),
.B(n_1220),
.Y(n_1372)
);

O2A1O1Ixp33_ASAP7_75t_SL g1373 ( 
.A1(n_1110),
.A2(n_996),
.B(n_967),
.C(n_1190),
.Y(n_1373)
);

BUFx2_ASAP7_75t_L g1374 ( 
.A(n_1102),
.Y(n_1374)
);

AO31x2_ASAP7_75t_L g1375 ( 
.A1(n_1209),
.A2(n_1212),
.A3(n_1234),
.B(n_1246),
.Y(n_1375)
);

INVx3_ASAP7_75t_L g1376 ( 
.A(n_1198),
.Y(n_1376)
);

INVx1_ASAP7_75t_SL g1377 ( 
.A(n_1126),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1221),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1221),
.Y(n_1379)
);

AOI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1140),
.A2(n_918),
.B1(n_974),
.B2(n_967),
.Y(n_1380)
);

OA21x2_ASAP7_75t_L g1381 ( 
.A1(n_1209),
.A2(n_1212),
.B(n_1099),
.Y(n_1381)
);

INVx2_ASAP7_75t_L g1382 ( 
.A(n_1221),
.Y(n_1382)
);

A2O1A1Ixp33_ASAP7_75t_L g1383 ( 
.A1(n_1117),
.A2(n_918),
.B(n_996),
.C(n_1096),
.Y(n_1383)
);

BUFx6f_ASAP7_75t_SL g1384 ( 
.A(n_1136),
.Y(n_1384)
);

AO31x2_ASAP7_75t_L g1385 ( 
.A1(n_1209),
.A2(n_1212),
.A3(n_1234),
.B(n_1246),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1125),
.A2(n_1229),
.B(n_1220),
.Y(n_1386)
);

OAI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1112),
.A2(n_918),
.B1(n_1101),
.B2(n_1143),
.Y(n_1387)
);

OAI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1246),
.A2(n_1117),
.B(n_918),
.Y(n_1388)
);

BUFx6f_ASAP7_75t_L g1389 ( 
.A(n_1198),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_SL g1390 ( 
.A1(n_1165),
.A2(n_1162),
.B(n_1168),
.Y(n_1390)
);

AO31x2_ASAP7_75t_L g1391 ( 
.A1(n_1209),
.A2(n_1212),
.A3(n_1234),
.B(n_1246),
.Y(n_1391)
);

BUFx2_ASAP7_75t_R g1392 ( 
.A(n_1139),
.Y(n_1392)
);

AO31x2_ASAP7_75t_L g1393 ( 
.A1(n_1209),
.A2(n_1212),
.A3(n_1234),
.B(n_1246),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_L g1394 ( 
.A(n_1096),
.B(n_918),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1221),
.Y(n_1395)
);

AO31x2_ASAP7_75t_L g1396 ( 
.A1(n_1209),
.A2(n_1212),
.A3(n_1234),
.B(n_1246),
.Y(n_1396)
);

AO22x1_ASAP7_75t_L g1397 ( 
.A1(n_1177),
.A2(n_918),
.B1(n_677),
.B2(n_537),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_SL g1398 ( 
.A(n_1101),
.B(n_996),
.Y(n_1398)
);

AO31x2_ASAP7_75t_L g1399 ( 
.A1(n_1209),
.A2(n_1212),
.A3(n_1234),
.B(n_1246),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1101),
.B(n_918),
.Y(n_1400)
);

A2O1A1Ixp33_ASAP7_75t_L g1401 ( 
.A1(n_1117),
.A2(n_918),
.B(n_996),
.C(n_1096),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1217),
.Y(n_1402)
);

BUFx3_ASAP7_75t_L g1403 ( 
.A(n_1102),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1221),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1212),
.A2(n_1009),
.B(n_991),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1125),
.A2(n_1229),
.B(n_1220),
.Y(n_1406)
);

OA21x2_ASAP7_75t_L g1407 ( 
.A1(n_1209),
.A2(n_1212),
.B(n_1099),
.Y(n_1407)
);

INVx4_ASAP7_75t_L g1408 ( 
.A(n_1198),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1217),
.Y(n_1409)
);

NOR2xp33_ASAP7_75t_L g1410 ( 
.A(n_1096),
.B(n_918),
.Y(n_1410)
);

CKINVDCx11_ASAP7_75t_R g1411 ( 
.A(n_1348),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1394),
.A2(n_1410),
.B1(n_1336),
.B2(n_1276),
.Y(n_1412)
);

BUFx3_ASAP7_75t_L g1413 ( 
.A(n_1403),
.Y(n_1413)
);

OAI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1353),
.A2(n_1356),
.B1(n_1380),
.B2(n_1400),
.Y(n_1414)
);

INVx2_ASAP7_75t_SL g1415 ( 
.A(n_1374),
.Y(n_1415)
);

INVx6_ASAP7_75t_L g1416 ( 
.A(n_1271),
.Y(n_1416)
);

INVxp67_ASAP7_75t_L g1417 ( 
.A(n_1278),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1339),
.B(n_1299),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_SL g1419 ( 
.A1(n_1277),
.A2(n_1324),
.B1(n_1300),
.B2(n_1388),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1276),
.A2(n_1364),
.B1(n_1365),
.B2(n_1388),
.Y(n_1420)
);

BUFx2_ASAP7_75t_SL g1421 ( 
.A(n_1261),
.Y(n_1421)
);

HB1xp67_ASAP7_75t_L g1422 ( 
.A(n_1263),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1364),
.A2(n_1324),
.B1(n_1380),
.B2(n_1356),
.Y(n_1423)
);

AOI22xp5_ASAP7_75t_SL g1424 ( 
.A1(n_1397),
.A2(n_1341),
.B1(n_1314),
.B2(n_1302),
.Y(n_1424)
);

INVx6_ASAP7_75t_L g1425 ( 
.A(n_1271),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1353),
.A2(n_1301),
.B1(n_1282),
.B2(n_1398),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1282),
.A2(n_1387),
.B1(n_1370),
.B2(n_1369),
.Y(n_1427)
);

BUFx4_ASAP7_75t_R g1428 ( 
.A(n_1300),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_SL g1429 ( 
.A1(n_1300),
.A2(n_1390),
.B1(n_1387),
.B2(n_1311),
.Y(n_1429)
);

INVx1_ASAP7_75t_SL g1430 ( 
.A(n_1263),
.Y(n_1430)
);

CKINVDCx11_ASAP7_75t_R g1431 ( 
.A(n_1354),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_1253),
.Y(n_1432)
);

CKINVDCx11_ASAP7_75t_R g1433 ( 
.A(n_1294),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1296),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1369),
.A2(n_1256),
.B1(n_1267),
.B2(n_1284),
.Y(n_1435)
);

CKINVDCx11_ASAP7_75t_R g1436 ( 
.A(n_1362),
.Y(n_1436)
);

INVx8_ASAP7_75t_L g1437 ( 
.A(n_1271),
.Y(n_1437)
);

OAI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1359),
.A2(n_1401),
.B1(n_1383),
.B2(n_1289),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1321),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1273),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1297),
.A2(n_1342),
.B1(n_1289),
.B2(n_1255),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1281),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1340),
.Y(n_1443)
);

BUFx2_ASAP7_75t_SL g1444 ( 
.A(n_1384),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_SL g1445 ( 
.A1(n_1311),
.A2(n_1295),
.B1(n_1366),
.B2(n_1332),
.Y(n_1445)
);

BUFx2_ASAP7_75t_L g1446 ( 
.A(n_1268),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1255),
.A2(n_1323),
.B1(n_1407),
.B2(n_1381),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1381),
.A2(n_1407),
.B1(n_1366),
.B2(n_1350),
.Y(n_1448)
);

OAI22xp5_ASAP7_75t_SL g1449 ( 
.A1(n_1332),
.A2(n_1366),
.B1(n_1362),
.B2(n_1377),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_1384),
.Y(n_1450)
);

INVx1_ASAP7_75t_SL g1451 ( 
.A(n_1377),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1402),
.Y(n_1452)
);

BUFx12f_ASAP7_75t_L g1453 ( 
.A(n_1326),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1409),
.A2(n_1395),
.B1(n_1274),
.B2(n_1379),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1298),
.Y(n_1455)
);

BUFx6f_ASAP7_75t_L g1456 ( 
.A(n_1326),
.Y(n_1456)
);

AOI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1308),
.A2(n_1347),
.B1(n_1344),
.B2(n_1378),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1355),
.A2(n_1382),
.B1(n_1404),
.B2(n_1290),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_SL g1459 ( 
.A1(n_1310),
.A2(n_1327),
.B1(n_1262),
.B2(n_1367),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_L g1460 ( 
.A1(n_1254),
.A2(n_1288),
.B1(n_1337),
.B2(n_1335),
.Y(n_1460)
);

INVx3_ASAP7_75t_L g1461 ( 
.A(n_1349),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_1392),
.Y(n_1462)
);

BUFx4f_ASAP7_75t_SL g1463 ( 
.A(n_1328),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1357),
.A2(n_1287),
.B1(n_1257),
.B2(n_1345),
.Y(n_1464)
);

CKINVDCx11_ASAP7_75t_R g1465 ( 
.A(n_1326),
.Y(n_1465)
);

INVxp67_ASAP7_75t_SL g1466 ( 
.A(n_1329),
.Y(n_1466)
);

BUFx12f_ASAP7_75t_L g1467 ( 
.A(n_1363),
.Y(n_1467)
);

INVx2_ASAP7_75t_SL g1468 ( 
.A(n_1363),
.Y(n_1468)
);

INVx3_ASAP7_75t_SL g1469 ( 
.A(n_1363),
.Y(n_1469)
);

CKINVDCx20_ASAP7_75t_R g1470 ( 
.A(n_1389),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1307),
.A2(n_1306),
.B1(n_1346),
.B2(n_1405),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1338),
.Y(n_1472)
);

INVx6_ASAP7_75t_L g1473 ( 
.A(n_1349),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1373),
.B(n_1292),
.Y(n_1474)
);

BUFx6f_ASAP7_75t_L g1475 ( 
.A(n_1389),
.Y(n_1475)
);

OAI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1309),
.A2(n_1313),
.B1(n_1320),
.B2(n_1408),
.Y(n_1476)
);

INVx6_ASAP7_75t_L g1477 ( 
.A(n_1408),
.Y(n_1477)
);

AOI22xp33_ASAP7_75t_L g1478 ( 
.A1(n_1287),
.A2(n_1285),
.B1(n_1258),
.B2(n_1292),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1351),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1334),
.Y(n_1480)
);

OAI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1361),
.A2(n_1275),
.B(n_1360),
.Y(n_1481)
);

BUFx3_ASAP7_75t_L g1482 ( 
.A(n_1389),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1304),
.A2(n_1315),
.B1(n_1286),
.B2(n_1352),
.Y(n_1483)
);

CKINVDCx11_ASAP7_75t_R g1484 ( 
.A(n_1371),
.Y(n_1484)
);

CKINVDCx20_ASAP7_75t_R g1485 ( 
.A(n_1264),
.Y(n_1485)
);

BUFx4f_ASAP7_75t_SL g1486 ( 
.A(n_1264),
.Y(n_1486)
);

CKINVDCx14_ASAP7_75t_R g1487 ( 
.A(n_1283),
.Y(n_1487)
);

CKINVDCx11_ASAP7_75t_R g1488 ( 
.A(n_1331),
.Y(n_1488)
);

NAND2x1p5_ASAP7_75t_L g1489 ( 
.A(n_1322),
.B(n_1316),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_1283),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_SL g1491 ( 
.A1(n_1304),
.A2(n_1325),
.B1(n_1315),
.B2(n_1269),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1351),
.B(n_1391),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1251),
.A2(n_1376),
.B1(n_1305),
.B2(n_1319),
.Y(n_1493)
);

BUFx12f_ASAP7_75t_L g1494 ( 
.A(n_1330),
.Y(n_1494)
);

INVx4_ASAP7_75t_L g1495 ( 
.A(n_1376),
.Y(n_1495)
);

INVx6_ASAP7_75t_L g1496 ( 
.A(n_1330),
.Y(n_1496)
);

BUFx4f_ASAP7_75t_SL g1497 ( 
.A(n_1333),
.Y(n_1497)
);

BUFx2_ASAP7_75t_L g1498 ( 
.A(n_1333),
.Y(n_1498)
);

CKINVDCx10_ASAP7_75t_R g1499 ( 
.A(n_1305),
.Y(n_1499)
);

INVx6_ASAP7_75t_L g1500 ( 
.A(n_1318),
.Y(n_1500)
);

CKINVDCx11_ASAP7_75t_R g1501 ( 
.A(n_1305),
.Y(n_1501)
);

OAI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1303),
.A2(n_1312),
.B1(n_1385),
.B2(n_1375),
.Y(n_1502)
);

AOI22xp33_ASAP7_75t_L g1503 ( 
.A1(n_1270),
.A2(n_1358),
.B1(n_1386),
.B2(n_1372),
.Y(n_1503)
);

NAND2x1p5_ASAP7_75t_L g1504 ( 
.A(n_1317),
.B(n_1343),
.Y(n_1504)
);

CKINVDCx20_ASAP7_75t_R g1505 ( 
.A(n_1375),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_L g1506 ( 
.A1(n_1368),
.A2(n_1406),
.B1(n_1252),
.B2(n_1272),
.Y(n_1506)
);

BUFx2_ASAP7_75t_L g1507 ( 
.A(n_1385),
.Y(n_1507)
);

INVxp67_ASAP7_75t_SL g1508 ( 
.A(n_1385),
.Y(n_1508)
);

BUFx2_ASAP7_75t_SL g1509 ( 
.A(n_1293),
.Y(n_1509)
);

BUFx6f_ASAP7_75t_L g1510 ( 
.A(n_1279),
.Y(n_1510)
);

INVx4_ASAP7_75t_L g1511 ( 
.A(n_1293),
.Y(n_1511)
);

OAI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1391),
.A2(n_1399),
.B1(n_1396),
.B2(n_1393),
.Y(n_1512)
);

NAND2xp5_ASAP7_75t_L g1513 ( 
.A(n_1393),
.B(n_1399),
.Y(n_1513)
);

INVx6_ASAP7_75t_L g1514 ( 
.A(n_1293),
.Y(n_1514)
);

BUFx12f_ASAP7_75t_L g1515 ( 
.A(n_1259),
.Y(n_1515)
);

OAI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1393),
.A2(n_1399),
.B1(n_1396),
.B2(n_1291),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_1291),
.Y(n_1517)
);

INVx3_ASAP7_75t_SL g1518 ( 
.A(n_1259),
.Y(n_1518)
);

CKINVDCx11_ASAP7_75t_R g1519 ( 
.A(n_1259),
.Y(n_1519)
);

BUFx10_ASAP7_75t_L g1520 ( 
.A(n_1260),
.Y(n_1520)
);

OAI21xp33_ASAP7_75t_L g1521 ( 
.A1(n_1279),
.A2(n_1265),
.B(n_1266),
.Y(n_1521)
);

CKINVDCx6p67_ASAP7_75t_R g1522 ( 
.A(n_1260),
.Y(n_1522)
);

INVx6_ASAP7_75t_L g1523 ( 
.A(n_1279),
.Y(n_1523)
);

BUFx8_ASAP7_75t_L g1524 ( 
.A(n_1260),
.Y(n_1524)
);

OAI22xp33_ASAP7_75t_R g1525 ( 
.A1(n_1265),
.A2(n_1394),
.B1(n_1410),
.B2(n_828),
.Y(n_1525)
);

OAI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1265),
.A2(n_1410),
.B1(n_1394),
.B2(n_1365),
.Y(n_1526)
);

CKINVDCx20_ASAP7_75t_R g1527 ( 
.A(n_1266),
.Y(n_1527)
);

INVx2_ASAP7_75t_SL g1528 ( 
.A(n_1403),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1280),
.Y(n_1529)
);

OAI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1353),
.A2(n_1356),
.B1(n_1380),
.B2(n_1394),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1394),
.A2(n_1410),
.B1(n_918),
.B2(n_1336),
.Y(n_1531)
);

OAI22xp33_ASAP7_75t_L g1532 ( 
.A1(n_1353),
.A2(n_1356),
.B1(n_1380),
.B2(n_1394),
.Y(n_1532)
);

CKINVDCx11_ASAP7_75t_R g1533 ( 
.A(n_1348),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1394),
.B(n_1410),
.Y(n_1534)
);

CKINVDCx20_ASAP7_75t_R g1535 ( 
.A(n_1354),
.Y(n_1535)
);

OAI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1394),
.A2(n_1410),
.B1(n_1365),
.B2(n_918),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1280),
.Y(n_1537)
);

BUFx12f_ASAP7_75t_L g1538 ( 
.A(n_1348),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1394),
.B(n_1410),
.Y(n_1539)
);

OAI22xp5_ASAP7_75t_L g1540 ( 
.A1(n_1394),
.A2(n_1410),
.B1(n_1365),
.B2(n_918),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1280),
.Y(n_1541)
);

CKINVDCx11_ASAP7_75t_R g1542 ( 
.A(n_1348),
.Y(n_1542)
);

BUFx2_ASAP7_75t_SL g1543 ( 
.A(n_1403),
.Y(n_1543)
);

OAI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1353),
.A2(n_1356),
.B1(n_1380),
.B2(n_1394),
.Y(n_1544)
);

BUFx6f_ASAP7_75t_L g1545 ( 
.A(n_1271),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1280),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1280),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1280),
.Y(n_1548)
);

BUFx2_ASAP7_75t_L g1549 ( 
.A(n_1374),
.Y(n_1549)
);

BUFx4f_ASAP7_75t_SL g1550 ( 
.A(n_1348),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1280),
.Y(n_1551)
);

BUFx3_ASAP7_75t_L g1552 ( 
.A(n_1403),
.Y(n_1552)
);

INVx3_ASAP7_75t_L g1553 ( 
.A(n_1271),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1280),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1280),
.Y(n_1555)
);

INVx2_ASAP7_75t_L g1556 ( 
.A(n_1439),
.Y(n_1556)
);

CKINVDCx20_ASAP7_75t_R g1557 ( 
.A(n_1431),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1472),
.Y(n_1558)
);

INVx3_ASAP7_75t_L g1559 ( 
.A(n_1496),
.Y(n_1559)
);

INVx4_ASAP7_75t_L g1560 ( 
.A(n_1428),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1439),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1440),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1536),
.A2(n_1540),
.B1(n_1419),
.B2(n_1530),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_1422),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1442),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1534),
.B(n_1539),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1418),
.B(n_1531),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1531),
.B(n_1412),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1412),
.B(n_1427),
.Y(n_1569)
);

BUFx6f_ASAP7_75t_L g1570 ( 
.A(n_1488),
.Y(n_1570)
);

AND2x4_ASAP7_75t_L g1571 ( 
.A(n_1442),
.B(n_1443),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1479),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1443),
.Y(n_1573)
);

AOI22xp33_ASAP7_75t_L g1574 ( 
.A1(n_1532),
.A2(n_1544),
.B1(n_1423),
.B2(n_1426),
.Y(n_1574)
);

NOR2xp33_ASAP7_75t_L g1575 ( 
.A(n_1436),
.B(n_1463),
.Y(n_1575)
);

AO21x2_ASAP7_75t_L g1576 ( 
.A1(n_1481),
.A2(n_1476),
.B(n_1471),
.Y(n_1576)
);

CKINVDCx6p67_ASAP7_75t_R g1577 ( 
.A(n_1431),
.Y(n_1577)
);

INVx2_ASAP7_75t_SL g1578 ( 
.A(n_1416),
.Y(n_1578)
);

OAI21x1_ASAP7_75t_L g1579 ( 
.A1(n_1504),
.A2(n_1506),
.B(n_1503),
.Y(n_1579)
);

CKINVDCx12_ASAP7_75t_R g1580 ( 
.A(n_1449),
.Y(n_1580)
);

INVx3_ASAP7_75t_L g1581 ( 
.A(n_1496),
.Y(n_1581)
);

INVx3_ASAP7_75t_L g1582 ( 
.A(n_1496),
.Y(n_1582)
);

INVx2_ASAP7_75t_SL g1583 ( 
.A(n_1416),
.Y(n_1583)
);

OR2x6_ASAP7_75t_L g1584 ( 
.A(n_1494),
.B(n_1509),
.Y(n_1584)
);

NOR2xp33_ASAP7_75t_SL g1585 ( 
.A(n_1462),
.B(n_1432),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1427),
.B(n_1435),
.Y(n_1586)
);

OAI21x1_ASAP7_75t_L g1587 ( 
.A1(n_1504),
.A2(n_1506),
.B(n_1503),
.Y(n_1587)
);

OAI21xp33_ASAP7_75t_SL g1588 ( 
.A1(n_1420),
.A2(n_1426),
.B(n_1474),
.Y(n_1588)
);

INVx3_ASAP7_75t_L g1589 ( 
.A(n_1494),
.Y(n_1589)
);

BUFx2_ASAP7_75t_L g1590 ( 
.A(n_1498),
.Y(n_1590)
);

NAND2xp33_ASAP7_75t_R g1591 ( 
.A(n_1450),
.B(n_1549),
.Y(n_1591)
);

NOR2xp33_ASAP7_75t_L g1592 ( 
.A(n_1430),
.B(n_1451),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1452),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1434),
.Y(n_1594)
);

NOR2xp67_ASAP7_75t_SL g1595 ( 
.A(n_1444),
.B(n_1543),
.Y(n_1595)
);

INVx3_ASAP7_75t_L g1596 ( 
.A(n_1497),
.Y(n_1596)
);

A2O1A1Ixp33_ASAP7_75t_L g1597 ( 
.A1(n_1424),
.A2(n_1420),
.B(n_1438),
.C(n_1429),
.Y(n_1597)
);

INVx3_ASAP7_75t_L g1598 ( 
.A(n_1489),
.Y(n_1598)
);

BUFx2_ASAP7_75t_L g1599 ( 
.A(n_1480),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1537),
.Y(n_1600)
);

OAI21x1_ASAP7_75t_L g1601 ( 
.A1(n_1502),
.A2(n_1478),
.B(n_1464),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1435),
.B(n_1414),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1541),
.Y(n_1603)
);

BUFx6f_ASAP7_75t_L g1604 ( 
.A(n_1545),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1507),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1492),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1501),
.B(n_1505),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1513),
.B(n_1512),
.Y(n_1608)
);

AOI21x1_ASAP7_75t_L g1609 ( 
.A1(n_1516),
.A2(n_1526),
.B(n_1554),
.Y(n_1609)
);

HB1xp67_ASAP7_75t_L g1610 ( 
.A(n_1417),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1517),
.B(n_1518),
.Y(n_1611)
);

OA21x2_ASAP7_75t_L g1612 ( 
.A1(n_1483),
.A2(n_1478),
.B(n_1521),
.Y(n_1612)
);

AOI22xp33_ASAP7_75t_L g1613 ( 
.A1(n_1525),
.A2(n_1441),
.B1(n_1519),
.B2(n_1445),
.Y(n_1613)
);

OAI21x1_ASAP7_75t_L g1614 ( 
.A1(n_1464),
.A2(n_1483),
.B(n_1493),
.Y(n_1614)
);

OA21x2_ASAP7_75t_L g1615 ( 
.A1(n_1493),
.A2(n_1448),
.B(n_1508),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1529),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1518),
.B(n_1447),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1441),
.A2(n_1527),
.B1(n_1484),
.B2(n_1459),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1447),
.B(n_1448),
.Y(n_1619)
);

INVxp67_ASAP7_75t_L g1620 ( 
.A(n_1446),
.Y(n_1620)
);

BUFx3_ASAP7_75t_L g1621 ( 
.A(n_1413),
.Y(n_1621)
);

INVxp67_ASAP7_75t_L g1622 ( 
.A(n_1415),
.Y(n_1622)
);

OAI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1460),
.A2(n_1485),
.B1(n_1487),
.B2(n_1454),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1515),
.B(n_1511),
.Y(n_1624)
);

AO21x1_ASAP7_75t_L g1625 ( 
.A1(n_1511),
.A2(n_1466),
.B(n_1499),
.Y(n_1625)
);

OR2x6_ASAP7_75t_L g1626 ( 
.A(n_1523),
.B(n_1514),
.Y(n_1626)
);

OAI21x1_ASAP7_75t_L g1627 ( 
.A1(n_1458),
.A2(n_1454),
.B(n_1457),
.Y(n_1627)
);

INVx4_ASAP7_75t_L g1628 ( 
.A(n_1428),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1514),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_1546),
.Y(n_1630)
);

INVxp67_ASAP7_75t_L g1631 ( 
.A(n_1421),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1514),
.Y(n_1632)
);

BUFx2_ASAP7_75t_L g1633 ( 
.A(n_1524),
.Y(n_1633)
);

OAI21x1_ASAP7_75t_SL g1634 ( 
.A1(n_1458),
.A2(n_1457),
.B(n_1551),
.Y(n_1634)
);

OAI21x1_ASAP7_75t_L g1635 ( 
.A1(n_1547),
.A2(n_1555),
.B(n_1548),
.Y(n_1635)
);

BUFx2_ASAP7_75t_L g1636 ( 
.A(n_1524),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1510),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1524),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1522),
.Y(n_1639)
);

HB1xp67_ASAP7_75t_L g1640 ( 
.A(n_1487),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_L g1641 ( 
.A(n_1528),
.B(n_1413),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1455),
.Y(n_1642)
);

BUFx12f_ASAP7_75t_L g1643 ( 
.A(n_1411),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1552),
.B(n_1490),
.Y(n_1644)
);

INVx4_ASAP7_75t_L g1645 ( 
.A(n_1437),
.Y(n_1645)
);

OAI21x1_ASAP7_75t_L g1646 ( 
.A1(n_1553),
.A2(n_1520),
.B(n_1491),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1500),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1500),
.Y(n_1648)
);

INVxp67_ASAP7_75t_L g1649 ( 
.A(n_1552),
.Y(n_1649)
);

OAI21x1_ASAP7_75t_L g1650 ( 
.A1(n_1553),
.A2(n_1461),
.B(n_1437),
.Y(n_1650)
);

AND2x4_ASAP7_75t_L g1651 ( 
.A(n_1545),
.B(n_1495),
.Y(n_1651)
);

OR2x2_ASAP7_75t_L g1652 ( 
.A(n_1469),
.B(n_1461),
.Y(n_1652)
);

OAI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1470),
.A2(n_1486),
.B1(n_1425),
.B2(n_1416),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1456),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1475),
.Y(n_1655)
);

O2A1O1Ixp33_ASAP7_75t_SL g1656 ( 
.A1(n_1597),
.A2(n_1468),
.B(n_1437),
.C(n_1535),
.Y(n_1656)
);

OAI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1563),
.A2(n_1482),
.B(n_1433),
.Y(n_1657)
);

AO32x2_ASAP7_75t_L g1658 ( 
.A1(n_1623),
.A2(n_1465),
.A3(n_1453),
.B1(n_1467),
.B2(n_1425),
.Y(n_1658)
);

NAND3xp33_ASAP7_75t_L g1659 ( 
.A(n_1574),
.B(n_1545),
.C(n_1533),
.Y(n_1659)
);

OAI21xp5_ASAP7_75t_L g1660 ( 
.A1(n_1588),
.A2(n_1477),
.B(n_1473),
.Y(n_1660)
);

NAND4xp25_ASAP7_75t_L g1661 ( 
.A(n_1566),
.B(n_1550),
.C(n_1542),
.D(n_1538),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1607),
.B(n_1453),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1564),
.B(n_1473),
.Y(n_1663)
);

A2O1A1Ixp33_ASAP7_75t_L g1664 ( 
.A1(n_1602),
.A2(n_1613),
.B(n_1607),
.C(n_1569),
.Y(n_1664)
);

NOR2xp33_ASAP7_75t_L g1665 ( 
.A(n_1586),
.B(n_1568),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1573),
.Y(n_1666)
);

OAI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1618),
.A2(n_1477),
.B(n_1467),
.Y(n_1667)
);

AOI21xp5_ASAP7_75t_L g1668 ( 
.A1(n_1576),
.A2(n_1538),
.B(n_1626),
.Y(n_1668)
);

INVxp67_ASAP7_75t_L g1669 ( 
.A(n_1592),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1630),
.B(n_1610),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1619),
.B(n_1611),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1571),
.B(n_1567),
.Y(n_1672)
);

OAI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1601),
.A2(n_1627),
.B(n_1631),
.Y(n_1673)
);

AOI21xp5_ASAP7_75t_L g1674 ( 
.A1(n_1576),
.A2(n_1626),
.B(n_1584),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1619),
.B(n_1611),
.Y(n_1675)
);

NAND2xp33_ASAP7_75t_R g1676 ( 
.A(n_1633),
.B(n_1636),
.Y(n_1676)
);

OAI21xp5_ASAP7_75t_L g1677 ( 
.A1(n_1647),
.A2(n_1648),
.B(n_1609),
.Y(n_1677)
);

O2A1O1Ixp33_ASAP7_75t_SL g1678 ( 
.A1(n_1638),
.A2(n_1653),
.B(n_1639),
.C(n_1596),
.Y(n_1678)
);

OR2x2_ASAP7_75t_L g1679 ( 
.A(n_1608),
.B(n_1617),
.Y(n_1679)
);

OAI21xp5_ASAP7_75t_L g1680 ( 
.A1(n_1647),
.A2(n_1648),
.B(n_1614),
.Y(n_1680)
);

OAI211xp5_ASAP7_75t_L g1681 ( 
.A1(n_1620),
.A2(n_1622),
.B(n_1560),
.C(n_1628),
.Y(n_1681)
);

INVx5_ASAP7_75t_SL g1682 ( 
.A(n_1577),
.Y(n_1682)
);

NOR2x1_ASAP7_75t_SL g1683 ( 
.A(n_1584),
.B(n_1626),
.Y(n_1683)
);

NOR3xp33_ASAP7_75t_SL g1684 ( 
.A(n_1591),
.B(n_1575),
.C(n_1641),
.Y(n_1684)
);

AND2x4_ASAP7_75t_L g1685 ( 
.A(n_1589),
.B(n_1638),
.Y(n_1685)
);

OA21x2_ASAP7_75t_L g1686 ( 
.A1(n_1614),
.A2(n_1579),
.B(n_1587),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1642),
.B(n_1616),
.Y(n_1687)
);

AOI22xp33_ASAP7_75t_L g1688 ( 
.A1(n_1625),
.A2(n_1576),
.B1(n_1628),
.B2(n_1560),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1608),
.B(n_1606),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1606),
.B(n_1617),
.Y(n_1690)
);

NOR2xp33_ASAP7_75t_L g1691 ( 
.A(n_1580),
.B(n_1560),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1593),
.B(n_1612),
.Y(n_1692)
);

OAI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1628),
.A2(n_1570),
.B1(n_1649),
.B2(n_1640),
.Y(n_1693)
);

A2O1A1Ixp33_ASAP7_75t_L g1694 ( 
.A1(n_1633),
.A2(n_1636),
.B(n_1595),
.C(n_1646),
.Y(n_1694)
);

AND2x4_ASAP7_75t_L g1695 ( 
.A(n_1589),
.B(n_1639),
.Y(n_1695)
);

INVxp67_ASAP7_75t_L g1696 ( 
.A(n_1621),
.Y(n_1696)
);

CKINVDCx20_ASAP7_75t_R g1697 ( 
.A(n_1557),
.Y(n_1697)
);

A2O1A1Ixp33_ASAP7_75t_L g1698 ( 
.A1(n_1595),
.A2(n_1646),
.B(n_1596),
.C(n_1625),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1612),
.B(n_1573),
.Y(n_1699)
);

OAI21xp5_ASAP7_75t_L g1700 ( 
.A1(n_1635),
.A2(n_1644),
.B(n_1650),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1612),
.B(n_1624),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1562),
.B(n_1565),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1642),
.B(n_1594),
.Y(n_1703)
);

BUFx6f_ASAP7_75t_L g1704 ( 
.A(n_1570),
.Y(n_1704)
);

AND2x6_ASAP7_75t_L g1705 ( 
.A(n_1559),
.B(n_1581),
.Y(n_1705)
);

AOI211xp5_ASAP7_75t_L g1706 ( 
.A1(n_1570),
.A2(n_1580),
.B(n_1652),
.C(n_1624),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1612),
.B(n_1556),
.Y(n_1707)
);

AOI21xp5_ASAP7_75t_L g1708 ( 
.A1(n_1626),
.A2(n_1584),
.B(n_1615),
.Y(n_1708)
);

A2O1A1Ixp33_ASAP7_75t_L g1709 ( 
.A1(n_1570),
.A2(n_1590),
.B(n_1605),
.C(n_1650),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1561),
.B(n_1637),
.Y(n_1710)
);

OAI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1570),
.A2(n_1557),
.B1(n_1577),
.B2(n_1578),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1654),
.B(n_1655),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1635),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1600),
.B(n_1603),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1689),
.B(n_1599),
.Y(n_1715)
);

BUFx2_ASAP7_75t_L g1716 ( 
.A(n_1699),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1689),
.B(n_1599),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1690),
.B(n_1665),
.Y(n_1718)
);

AOI22xp33_ASAP7_75t_L g1719 ( 
.A1(n_1665),
.A2(n_1643),
.B1(n_1634),
.B2(n_1615),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1701),
.B(n_1615),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1690),
.B(n_1671),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1707),
.Y(n_1722)
);

HB1xp67_ASAP7_75t_L g1723 ( 
.A(n_1692),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1692),
.B(n_1686),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1679),
.B(n_1590),
.Y(n_1725)
);

AOI22xp33_ASAP7_75t_L g1726 ( 
.A1(n_1659),
.A2(n_1643),
.B1(n_1615),
.B2(n_1585),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1666),
.Y(n_1727)
);

BUFx2_ASAP7_75t_L g1728 ( 
.A(n_1700),
.Y(n_1728)
);

AOI22xp33_ASAP7_75t_SL g1729 ( 
.A1(n_1657),
.A2(n_1581),
.B1(n_1559),
.B2(n_1582),
.Y(n_1729)
);

BUFx2_ASAP7_75t_L g1730 ( 
.A(n_1680),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_SL g1731 ( 
.A(n_1706),
.B(n_1598),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1675),
.B(n_1558),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1675),
.B(n_1558),
.Y(n_1733)
);

INVx5_ASAP7_75t_L g1734 ( 
.A(n_1705),
.Y(n_1734)
);

AOI22xp5_ASAP7_75t_L g1735 ( 
.A1(n_1664),
.A2(n_1578),
.B1(n_1583),
.B2(n_1645),
.Y(n_1735)
);

HB1xp67_ASAP7_75t_L g1736 ( 
.A(n_1713),
.Y(n_1736)
);

OAI221xp5_ASAP7_75t_L g1737 ( 
.A1(n_1664),
.A2(n_1583),
.B1(n_1632),
.B2(n_1629),
.C(n_1645),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1672),
.B(n_1572),
.Y(n_1738)
);

BUFx2_ASAP7_75t_L g1739 ( 
.A(n_1673),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1710),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1670),
.B(n_1708),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1687),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1702),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1742),
.B(n_1718),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1736),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1736),
.Y(n_1746)
);

AOI221xp5_ASAP7_75t_L g1747 ( 
.A1(n_1737),
.A2(n_1656),
.B1(n_1669),
.B2(n_1678),
.C(n_1668),
.Y(n_1747)
);

INVx5_ASAP7_75t_L g1748 ( 
.A(n_1734),
.Y(n_1748)
);

AOI22xp33_ASAP7_75t_L g1749 ( 
.A1(n_1739),
.A2(n_1726),
.B1(n_1729),
.B2(n_1728),
.Y(n_1749)
);

NAND3xp33_ASAP7_75t_L g1750 ( 
.A(n_1735),
.B(n_1684),
.C(n_1698),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1727),
.Y(n_1751)
);

HB1xp67_ASAP7_75t_L g1752 ( 
.A(n_1725),
.Y(n_1752)
);

HB1xp67_ASAP7_75t_L g1753 ( 
.A(n_1725),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1723),
.B(n_1674),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1727),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1742),
.B(n_1718),
.Y(n_1756)
);

AND2x4_ASAP7_75t_L g1757 ( 
.A(n_1734),
.B(n_1683),
.Y(n_1757)
);

INVxp67_ASAP7_75t_L g1758 ( 
.A(n_1741),
.Y(n_1758)
);

OR2x2_ASAP7_75t_L g1759 ( 
.A(n_1723),
.B(n_1694),
.Y(n_1759)
);

OAI22xp5_ASAP7_75t_L g1760 ( 
.A1(n_1735),
.A2(n_1688),
.B1(n_1667),
.B2(n_1697),
.Y(n_1760)
);

BUFx2_ASAP7_75t_L g1761 ( 
.A(n_1734),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1716),
.B(n_1685),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1741),
.B(n_1712),
.Y(n_1763)
);

OR2x2_ASAP7_75t_L g1764 ( 
.A(n_1741),
.B(n_1694),
.Y(n_1764)
);

HB1xp67_ASAP7_75t_L g1765 ( 
.A(n_1715),
.Y(n_1765)
);

INVxp67_ASAP7_75t_SL g1766 ( 
.A(n_1724),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1732),
.B(n_1733),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1720),
.B(n_1695),
.Y(n_1768)
);

INVx3_ASAP7_75t_L g1769 ( 
.A(n_1722),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_L g1770 ( 
.A(n_1732),
.B(n_1677),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1733),
.B(n_1709),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1720),
.B(n_1695),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1738),
.B(n_1709),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1721),
.B(n_1703),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1738),
.B(n_1714),
.Y(n_1775)
);

HB1xp67_ASAP7_75t_L g1776 ( 
.A(n_1715),
.Y(n_1776)
);

INVx1_ASAP7_75t_SL g1777 ( 
.A(n_1764),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1768),
.B(n_1720),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1758),
.B(n_1730),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1769),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1768),
.B(n_1739),
.Y(n_1781)
);

HB1xp67_ASAP7_75t_L g1782 ( 
.A(n_1752),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1758),
.B(n_1770),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1770),
.B(n_1728),
.Y(n_1784)
);

NAND3xp33_ASAP7_75t_L g1785 ( 
.A(n_1750),
.B(n_1728),
.C(n_1739),
.Y(n_1785)
);

NAND4xp25_ASAP7_75t_L g1786 ( 
.A(n_1750),
.B(n_1726),
.C(n_1719),
.D(n_1737),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1769),
.Y(n_1787)
);

NOR2xp33_ASAP7_75t_L g1788 ( 
.A(n_1774),
.B(n_1661),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1772),
.B(n_1730),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1772),
.B(n_1730),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1769),
.Y(n_1791)
);

INVx2_ASAP7_75t_SL g1792 ( 
.A(n_1762),
.Y(n_1792)
);

INVxp67_ASAP7_75t_L g1793 ( 
.A(n_1771),
.Y(n_1793)
);

INVx2_ASAP7_75t_SL g1794 ( 
.A(n_1762),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1773),
.B(n_1724),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1773),
.B(n_1724),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1745),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1771),
.B(n_1743),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1745),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1744),
.B(n_1756),
.Y(n_1800)
);

OR2x2_ASAP7_75t_L g1801 ( 
.A(n_1754),
.B(n_1717),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1746),
.Y(n_1802)
);

OR2x2_ASAP7_75t_L g1803 ( 
.A(n_1754),
.B(n_1717),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1746),
.Y(n_1804)
);

AND2x4_ASAP7_75t_L g1805 ( 
.A(n_1748),
.B(n_1734),
.Y(n_1805)
);

AOI22xp5_ASAP7_75t_L g1806 ( 
.A1(n_1760),
.A2(n_1656),
.B1(n_1688),
.B2(n_1729),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1744),
.B(n_1743),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1751),
.Y(n_1808)
);

OR2x2_ASAP7_75t_L g1809 ( 
.A(n_1759),
.B(n_1740),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1769),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1751),
.Y(n_1811)
);

OR2x2_ASAP7_75t_L g1812 ( 
.A(n_1759),
.B(n_1738),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1755),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1755),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1793),
.B(n_1763),
.Y(n_1815)
);

INVx1_ASAP7_75t_SL g1816 ( 
.A(n_1777),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1789),
.B(n_1764),
.Y(n_1817)
);

NOR3xp33_ASAP7_75t_L g1818 ( 
.A(n_1785),
.B(n_1760),
.C(n_1747),
.Y(n_1818)
);

NAND3xp33_ASAP7_75t_L g1819 ( 
.A(n_1785),
.B(n_1749),
.C(n_1747),
.Y(n_1819)
);

AND4x1_ASAP7_75t_L g1820 ( 
.A(n_1806),
.B(n_1691),
.C(n_1698),
.D(n_1660),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1789),
.B(n_1766),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1797),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1797),
.Y(n_1823)
);

OR2x2_ASAP7_75t_L g1824 ( 
.A(n_1812),
.B(n_1763),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1799),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1777),
.B(n_1756),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1790),
.B(n_1766),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1799),
.Y(n_1828)
);

NOR2xp33_ASAP7_75t_L g1829 ( 
.A(n_1788),
.B(n_1697),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1802),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1802),
.Y(n_1831)
);

NOR2xp33_ASAP7_75t_L g1832 ( 
.A(n_1786),
.B(n_1682),
.Y(n_1832)
);

INVxp67_ASAP7_75t_L g1833 ( 
.A(n_1782),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1780),
.Y(n_1834)
);

INVx2_ASAP7_75t_L g1835 ( 
.A(n_1780),
.Y(n_1835)
);

NOR2x1p5_ASAP7_75t_L g1836 ( 
.A(n_1786),
.B(n_1704),
.Y(n_1836)
);

NAND2x1p5_ASAP7_75t_L g1837 ( 
.A(n_1805),
.B(n_1748),
.Y(n_1837)
);

AO22x1_ASAP7_75t_L g1838 ( 
.A1(n_1805),
.A2(n_1748),
.B1(n_1711),
.B2(n_1704),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1780),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1790),
.B(n_1757),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1804),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1804),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1787),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1781),
.B(n_1757),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1787),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1808),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1781),
.B(n_1757),
.Y(n_1847)
);

AOI211xp5_ASAP7_75t_L g1848 ( 
.A1(n_1806),
.A2(n_1678),
.B(n_1691),
.C(n_1731),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1792),
.B(n_1757),
.Y(n_1849)
);

AND2x2_ASAP7_75t_L g1850 ( 
.A(n_1792),
.B(n_1761),
.Y(n_1850)
);

INVx2_ASAP7_75t_L g1851 ( 
.A(n_1787),
.Y(n_1851)
);

AND2x4_ASAP7_75t_L g1852 ( 
.A(n_1805),
.B(n_1748),
.Y(n_1852)
);

INVx1_ASAP7_75t_SL g1853 ( 
.A(n_1812),
.Y(n_1853)
);

NOR2xp33_ASAP7_75t_L g1854 ( 
.A(n_1784),
.B(n_1682),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1783),
.B(n_1765),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1808),
.Y(n_1856)
);

AND2x4_ASAP7_75t_L g1857 ( 
.A(n_1805),
.B(n_1748),
.Y(n_1857)
);

OR2x2_ASAP7_75t_L g1858 ( 
.A(n_1795),
.B(n_1753),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1811),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1783),
.B(n_1776),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1834),
.Y(n_1861)
);

OR2x2_ASAP7_75t_L g1862 ( 
.A(n_1816),
.B(n_1795),
.Y(n_1862)
);

OR2x2_ASAP7_75t_L g1863 ( 
.A(n_1853),
.B(n_1796),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1822),
.Y(n_1864)
);

INVx1_ASAP7_75t_SL g1865 ( 
.A(n_1837),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1822),
.Y(n_1866)
);

BUFx2_ASAP7_75t_L g1867 ( 
.A(n_1837),
.Y(n_1867)
);

OR2x2_ASAP7_75t_L g1868 ( 
.A(n_1824),
.B(n_1796),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1823),
.Y(n_1869)
);

AOI22xp33_ASAP7_75t_L g1870 ( 
.A1(n_1818),
.A2(n_1819),
.B1(n_1836),
.B2(n_1832),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1824),
.B(n_1784),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1836),
.B(n_1798),
.Y(n_1872)
);

HB1xp67_ASAP7_75t_L g1873 ( 
.A(n_1833),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1817),
.B(n_1852),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1823),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1825),
.Y(n_1876)
);

INVx2_ASAP7_75t_L g1877 ( 
.A(n_1834),
.Y(n_1877)
);

HB1xp67_ASAP7_75t_L g1878 ( 
.A(n_1817),
.Y(n_1878)
);

AND2x4_ASAP7_75t_L g1879 ( 
.A(n_1852),
.B(n_1748),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1825),
.Y(n_1880)
);

HB1xp67_ASAP7_75t_L g1881 ( 
.A(n_1826),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1834),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1852),
.B(n_1794),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_L g1884 ( 
.A(n_1819),
.B(n_1798),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1848),
.B(n_1800),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_SL g1886 ( 
.A(n_1848),
.B(n_1748),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1828),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1852),
.B(n_1794),
.Y(n_1888)
);

OR2x2_ASAP7_75t_L g1889 ( 
.A(n_1858),
.B(n_1779),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1828),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1815),
.B(n_1800),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1830),
.Y(n_1892)
);

HB1xp67_ASAP7_75t_L g1893 ( 
.A(n_1830),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1831),
.Y(n_1894)
);

OR2x2_ASAP7_75t_L g1895 ( 
.A(n_1858),
.B(n_1779),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1857),
.B(n_1778),
.Y(n_1896)
);

AND2x4_ASAP7_75t_L g1897 ( 
.A(n_1857),
.B(n_1840),
.Y(n_1897)
);

INVx1_ASAP7_75t_SL g1898 ( 
.A(n_1874),
.Y(n_1898)
);

NOR2xp33_ASAP7_75t_L g1899 ( 
.A(n_1870),
.B(n_1829),
.Y(n_1899)
);

AOI32xp33_ASAP7_75t_L g1900 ( 
.A1(n_1885),
.A2(n_1850),
.A3(n_1854),
.B1(n_1820),
.B2(n_1857),
.Y(n_1900)
);

AOI211xp5_ASAP7_75t_L g1901 ( 
.A1(n_1886),
.A2(n_1838),
.B(n_1857),
.C(n_1820),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1884),
.B(n_1855),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1897),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1893),
.Y(n_1904)
);

NOR3xp33_ASAP7_75t_L g1905 ( 
.A(n_1873),
.B(n_1838),
.C(n_1860),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1864),
.Y(n_1906)
);

OAI22xp5_ASAP7_75t_L g1907 ( 
.A1(n_1878),
.A2(n_1837),
.B1(n_1731),
.B2(n_1719),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1864),
.Y(n_1908)
);

OR2x2_ASAP7_75t_L g1909 ( 
.A(n_1862),
.B(n_1872),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1881),
.B(n_1821),
.Y(n_1910)
);

INVxp67_ASAP7_75t_SL g1911 ( 
.A(n_1861),
.Y(n_1911)
);

OR2x2_ASAP7_75t_L g1912 ( 
.A(n_1862),
.B(n_1801),
.Y(n_1912)
);

OAI22xp5_ASAP7_75t_L g1913 ( 
.A1(n_1897),
.A2(n_1863),
.B1(n_1891),
.B2(n_1867),
.Y(n_1913)
);

NOR2xp33_ASAP7_75t_R g1914 ( 
.A(n_1867),
.B(n_1676),
.Y(n_1914)
);

NOR2xp33_ASAP7_75t_L g1915 ( 
.A(n_1874),
.B(n_1682),
.Y(n_1915)
);

AND2x2_ASAP7_75t_L g1916 ( 
.A(n_1897),
.B(n_1840),
.Y(n_1916)
);

AOI22xp5_ASAP7_75t_L g1917 ( 
.A1(n_1897),
.A2(n_1676),
.B1(n_1849),
.B2(n_1850),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1866),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1866),
.Y(n_1919)
);

INVx2_ASAP7_75t_SL g1920 ( 
.A(n_1883),
.Y(n_1920)
);

NAND2x1p5_ASAP7_75t_L g1921 ( 
.A(n_1865),
.B(n_1704),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1869),
.Y(n_1922)
);

INVx1_ASAP7_75t_SL g1923 ( 
.A(n_1883),
.Y(n_1923)
);

OAI221xp5_ASAP7_75t_SL g1924 ( 
.A1(n_1863),
.A2(n_1681),
.B1(n_1827),
.B2(n_1821),
.C(n_1831),
.Y(n_1924)
);

INVxp67_ASAP7_75t_SL g1925 ( 
.A(n_1901),
.Y(n_1925)
);

OAI21xp33_ASAP7_75t_L g1926 ( 
.A1(n_1899),
.A2(n_1888),
.B(n_1889),
.Y(n_1926)
);

AOI22xp5_ASAP7_75t_L g1927 ( 
.A1(n_1899),
.A2(n_1905),
.B1(n_1898),
.B2(n_1907),
.Y(n_1927)
);

AOI22xp5_ASAP7_75t_L g1928 ( 
.A1(n_1905),
.A2(n_1888),
.B1(n_1879),
.B2(n_1865),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1911),
.Y(n_1929)
);

OAI211xp5_ASAP7_75t_L g1930 ( 
.A1(n_1900),
.A2(n_1924),
.B(n_1902),
.C(n_1904),
.Y(n_1930)
);

OAI31xp33_ASAP7_75t_L g1931 ( 
.A1(n_1924),
.A2(n_1879),
.A3(n_1895),
.B(n_1889),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1916),
.Y(n_1932)
);

AND2x4_ASAP7_75t_L g1933 ( 
.A(n_1903),
.B(n_1896),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1911),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1906),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1908),
.Y(n_1936)
);

OAI221xp5_ASAP7_75t_L g1937 ( 
.A1(n_1917),
.A2(n_1895),
.B1(n_1871),
.B2(n_1868),
.C(n_1896),
.Y(n_1937)
);

OAI21xp5_ASAP7_75t_L g1938 ( 
.A1(n_1913),
.A2(n_1879),
.B(n_1871),
.Y(n_1938)
);

NOR2xp33_ASAP7_75t_L g1939 ( 
.A(n_1915),
.B(n_1879),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1918),
.Y(n_1940)
);

O2A1O1Ixp33_ASAP7_75t_L g1941 ( 
.A1(n_1909),
.A2(n_1894),
.B(n_1892),
.C(n_1890),
.Y(n_1941)
);

AOI22xp5_ASAP7_75t_L g1942 ( 
.A1(n_1923),
.A2(n_1849),
.B1(n_1847),
.B2(n_1844),
.Y(n_1942)
);

HB1xp67_ASAP7_75t_L g1943 ( 
.A(n_1920),
.Y(n_1943)
);

OR2x2_ASAP7_75t_L g1944 ( 
.A(n_1910),
.B(n_1868),
.Y(n_1944)
);

INVxp67_ASAP7_75t_L g1945 ( 
.A(n_1912),
.Y(n_1945)
);

O2A1O1Ixp5_ASAP7_75t_L g1946 ( 
.A1(n_1919),
.A2(n_1894),
.B(n_1892),
.C(n_1890),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1929),
.Y(n_1947)
);

HB1xp67_ASAP7_75t_L g1948 ( 
.A(n_1934),
.Y(n_1948)
);

OAI222xp33_ASAP7_75t_L g1949 ( 
.A1(n_1927),
.A2(n_1921),
.B1(n_1922),
.B2(n_1914),
.C1(n_1887),
.C2(n_1875),
.Y(n_1949)
);

OR2x2_ASAP7_75t_L g1950 ( 
.A(n_1944),
.B(n_1945),
.Y(n_1950)
);

AOI21xp33_ASAP7_75t_SL g1951 ( 
.A1(n_1931),
.A2(n_1921),
.B(n_1875),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1946),
.Y(n_1952)
);

AOI221xp5_ASAP7_75t_L g1953 ( 
.A1(n_1925),
.A2(n_1887),
.B1(n_1869),
.B2(n_1880),
.C(n_1876),
.Y(n_1953)
);

XOR2x2_ASAP7_75t_L g1954 ( 
.A(n_1928),
.B(n_1662),
.Y(n_1954)
);

OA21x2_ASAP7_75t_SL g1955 ( 
.A1(n_1933),
.A2(n_1807),
.B(n_1775),
.Y(n_1955)
);

AOI22xp5_ASAP7_75t_L g1956 ( 
.A1(n_1930),
.A2(n_1880),
.B1(n_1876),
.B2(n_1761),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1946),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1943),
.Y(n_1958)
);

NOR3xp33_ASAP7_75t_L g1959 ( 
.A(n_1951),
.B(n_1930),
.C(n_1939),
.Y(n_1959)
);

OR2x2_ASAP7_75t_L g1960 ( 
.A(n_1958),
.B(n_1932),
.Y(n_1960)
);

HB1xp67_ASAP7_75t_L g1961 ( 
.A(n_1948),
.Y(n_1961)
);

OAI211xp5_ASAP7_75t_L g1962 ( 
.A1(n_1952),
.A2(n_1938),
.B(n_1941),
.C(n_1926),
.Y(n_1962)
);

INVx1_ASAP7_75t_SL g1963 ( 
.A(n_1950),
.Y(n_1963)
);

OAI21xp33_ASAP7_75t_L g1964 ( 
.A1(n_1954),
.A2(n_1942),
.B(n_1933),
.Y(n_1964)
);

NOR2x1_ASAP7_75t_SL g1965 ( 
.A(n_1947),
.B(n_1935),
.Y(n_1965)
);

AOI22xp5_ASAP7_75t_L g1966 ( 
.A1(n_1957),
.A2(n_1937),
.B1(n_1940),
.B2(n_1936),
.Y(n_1966)
);

OR2x2_ASAP7_75t_L g1967 ( 
.A(n_1956),
.B(n_1827),
.Y(n_1967)
);

O2A1O1Ixp33_ASAP7_75t_L g1968 ( 
.A1(n_1949),
.A2(n_1941),
.B(n_1882),
.C(n_1877),
.Y(n_1968)
);

AOI21xp33_ASAP7_75t_SL g1969 ( 
.A1(n_1959),
.A2(n_1955),
.B(n_1953),
.Y(n_1969)
);

AOI322xp5_ASAP7_75t_L g1970 ( 
.A1(n_1964),
.A2(n_1953),
.A3(n_1842),
.B1(n_1841),
.B2(n_1861),
.C1(n_1882),
.C2(n_1877),
.Y(n_1970)
);

NAND3xp33_ASAP7_75t_L g1971 ( 
.A(n_1962),
.B(n_1877),
.C(n_1861),
.Y(n_1971)
);

AOI32xp33_ASAP7_75t_L g1972 ( 
.A1(n_1963),
.A2(n_1882),
.A3(n_1847),
.B1(n_1844),
.B2(n_1841),
.Y(n_1972)
);

AOI21xp33_ASAP7_75t_L g1973 ( 
.A1(n_1968),
.A2(n_1842),
.B(n_1835),
.Y(n_1973)
);

NOR2x1_ASAP7_75t_L g1974 ( 
.A(n_1960),
.B(n_1846),
.Y(n_1974)
);

AOI211xp5_ASAP7_75t_SL g1975 ( 
.A1(n_1973),
.A2(n_1961),
.B(n_1966),
.C(n_1967),
.Y(n_1975)
);

INVx2_ASAP7_75t_SL g1976 ( 
.A(n_1974),
.Y(n_1976)
);

AOI221xp5_ASAP7_75t_SL g1977 ( 
.A1(n_1969),
.A2(n_1965),
.B1(n_1859),
.B2(n_1856),
.C(n_1846),
.Y(n_1977)
);

AOI221xp5_ASAP7_75t_L g1978 ( 
.A1(n_1971),
.A2(n_1859),
.B1(n_1856),
.B2(n_1835),
.C(n_1845),
.Y(n_1978)
);

NOR3xp33_ASAP7_75t_L g1979 ( 
.A(n_1972),
.B(n_1693),
.C(n_1645),
.Y(n_1979)
);

AOI221xp5_ASAP7_75t_L g1980 ( 
.A1(n_1970),
.A2(n_1845),
.B1(n_1835),
.B2(n_1851),
.C(n_1839),
.Y(n_1980)
);

OAI22xp5_ASAP7_75t_L g1981 ( 
.A1(n_1969),
.A2(n_1809),
.B1(n_1801),
.B2(n_1803),
.Y(n_1981)
);

BUFx6f_ASAP7_75t_L g1982 ( 
.A(n_1976),
.Y(n_1982)
);

NAND4xp75_ASAP7_75t_L g1983 ( 
.A(n_1977),
.B(n_1845),
.C(n_1851),
.D(n_1843),
.Y(n_1983)
);

NAND4xp75_ASAP7_75t_L g1984 ( 
.A(n_1978),
.B(n_1843),
.C(n_1839),
.D(n_1663),
.Y(n_1984)
);

NOR4xp75_ASAP7_75t_L g1985 ( 
.A(n_1981),
.B(n_1807),
.C(n_1767),
.D(n_1775),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1979),
.Y(n_1986)
);

OAI22xp5_ASAP7_75t_L g1987 ( 
.A1(n_1980),
.A2(n_1809),
.B1(n_1803),
.B2(n_1791),
.Y(n_1987)
);

XNOR2xp5_ASAP7_75t_L g1988 ( 
.A(n_1986),
.B(n_1975),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1982),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1984),
.Y(n_1990)
);

INVx1_ASAP7_75t_SL g1991 ( 
.A(n_1989),
.Y(n_1991)
);

CKINVDCx20_ASAP7_75t_R g1992 ( 
.A(n_1991),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1992),
.Y(n_1993)
);

OAI22xp5_ASAP7_75t_SL g1994 ( 
.A1(n_1992),
.A2(n_1988),
.B1(n_1990),
.B2(n_1987),
.Y(n_1994)
);

INVx2_ASAP7_75t_L g1995 ( 
.A(n_1993),
.Y(n_1995)
);

INVx2_ASAP7_75t_L g1996 ( 
.A(n_1994),
.Y(n_1996)
);

OAI21xp33_ASAP7_75t_L g1997 ( 
.A1(n_1996),
.A2(n_1985),
.B(n_1983),
.Y(n_1997)
);

OAI21x1_ASAP7_75t_L g1998 ( 
.A1(n_1995),
.A2(n_1810),
.B(n_1791),
.Y(n_1998)
);

OA21x2_ASAP7_75t_L g1999 ( 
.A1(n_1997),
.A2(n_1810),
.B(n_1791),
.Y(n_1999)
);

AOI22xp5_ASAP7_75t_L g2000 ( 
.A1(n_1999),
.A2(n_1998),
.B1(n_1704),
.B2(n_1810),
.Y(n_2000)
);

CKINVDCx20_ASAP7_75t_R g2001 ( 
.A(n_2000),
.Y(n_2001)
);

OAI221xp5_ASAP7_75t_R g2002 ( 
.A1(n_2001),
.A2(n_1814),
.B1(n_1811),
.B2(n_1813),
.C(n_1658),
.Y(n_2002)
);

AOI211xp5_ASAP7_75t_L g2003 ( 
.A1(n_2002),
.A2(n_1604),
.B(n_1696),
.C(n_1651),
.Y(n_2003)
);


endmodule