module fake_jpeg_30677_n_447 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_447);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_447;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx16f_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_14),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_11),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_48),
.B(n_66),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_50),
.Y(n_105)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_45),
.Y(n_51)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_52),
.Y(n_132)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_53),
.Y(n_135)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_54),
.Y(n_99)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_55),
.Y(n_142)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_21),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_57),
.B(n_58),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_29),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_60),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_30),
.B(n_0),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_75),
.Y(n_94)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_63),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_64),
.Y(n_141)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_22),
.B(n_0),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_16),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_16),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_29),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g121 ( 
.A(n_69),
.Y(n_121)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_71),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_72),
.Y(n_131)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_74),
.Y(n_143)
);

OR2x2_ASAP7_75t_SL g75 ( 
.A(n_42),
.B(n_0),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_18),
.Y(n_77)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_77),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_29),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_78),
.B(n_79),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_42),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_19),
.Y(n_80)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_18),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_24),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_27),
.Y(n_83)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_83),
.Y(n_145)
);

CKINVDCx9p33_ASAP7_75t_R g84 ( 
.A(n_41),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_84),
.Y(n_96)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_17),
.Y(n_85)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_28),
.B(n_1),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_86),
.B(n_91),
.Y(n_126)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

BUFx4f_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_17),
.Y(n_89)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_90),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_35),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_92),
.B(n_41),
.Y(n_127)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_20),
.Y(n_93)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_84),
.A2(n_37),
.B1(n_35),
.B2(n_27),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_103),
.A2(n_114),
.B1(n_130),
.B2(n_92),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_93),
.A2(n_37),
.B1(n_35),
.B2(n_27),
.Y(n_114)
);

OAI22xp33_ASAP7_75t_L g116 ( 
.A1(n_65),
.A2(n_20),
.B1(n_37),
.B2(n_40),
.Y(n_116)
);

OA22x2_ASAP7_75t_L g177 ( 
.A1(n_116),
.A2(n_81),
.B1(n_77),
.B2(n_74),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_75),
.B(n_44),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_123),
.B(n_140),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_127),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_64),
.A2(n_20),
.B1(n_47),
.B2(n_31),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_88),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_133),
.B(n_138),
.Y(n_147)
);

AO22x1_ASAP7_75t_SL g136 ( 
.A1(n_52),
.A2(n_20),
.B1(n_47),
.B2(n_31),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_136),
.B(n_72),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_50),
.A2(n_22),
.B1(n_44),
.B2(n_39),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_137),
.A2(n_36),
.B1(n_25),
.B2(n_26),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_69),
.B(n_33),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_49),
.B(n_33),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_139),
.B(n_49),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_53),
.B(n_34),
.Y(n_140)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_97),
.Y(n_148)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_148),
.Y(n_197)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_108),
.Y(n_149)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_149),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_94),
.B(n_55),
.C(n_63),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_150),
.B(n_156),
.C(n_158),
.Y(n_200)
);

A2O1A1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_94),
.A2(n_88),
.B(n_46),
.C(n_40),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_151),
.B(n_152),
.Y(n_208)
);

A2O1A1Ixp33_ASAP7_75t_L g152 ( 
.A1(n_118),
.A2(n_46),
.B(n_23),
.C(n_92),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_119),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_153),
.B(n_164),
.Y(n_199)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_128),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_154),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_105),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_155),
.Y(n_195)
);

AND2x2_ASAP7_75t_SL g156 ( 
.A(n_95),
.B(n_87),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_157),
.A2(n_162),
.B1(n_178),
.B2(n_141),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_109),
.B(n_76),
.C(n_82),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_102),
.B(n_60),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_159),
.Y(n_225)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_99),
.Y(n_160)
);

INVx4_ASAP7_75t_L g231 ( 
.A(n_160),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_105),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_161),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_32),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_163),
.B(n_166),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_117),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_144),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_165),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_136),
.B(n_32),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_112),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_167),
.Y(n_203)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_110),
.Y(n_168)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_168),
.Y(n_213)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_100),
.Y(n_169)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_169),
.Y(n_215)
);

OA22x2_ASAP7_75t_L g221 ( 
.A1(n_170),
.A2(n_177),
.B1(n_192),
.B2(n_145),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_103),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_171),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_113),
.Y(n_172)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_172),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_101),
.Y(n_173)
);

BUFx2_ASAP7_75t_SL g211 ( 
.A(n_173),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_126),
.B(n_26),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_174),
.B(n_184),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_113),
.Y(n_175)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_175),
.Y(n_222)
);

INVx6_ASAP7_75t_SL g176 ( 
.A(n_121),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_176),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_96),
.A2(n_83),
.B1(n_25),
.B2(n_39),
.Y(n_178)
);

INVx8_ASAP7_75t_L g179 ( 
.A(n_98),
.Y(n_179)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_179),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_114),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_180),
.Y(n_219)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_128),
.Y(n_181)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_181),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_183),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_104),
.B(n_106),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_107),
.B(n_36),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_185),
.B(n_187),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_112),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_186),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_121),
.B(n_34),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_116),
.B(n_68),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_188),
.B(n_190),
.Y(n_229)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_124),
.Y(n_189)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_189),
.Y(n_234)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_124),
.Y(n_190)
);

AOI21xp33_ASAP7_75t_SL g191 ( 
.A1(n_130),
.A2(n_71),
.B(n_67),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_134),
.C(n_111),
.Y(n_202)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_125),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_120),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_193),
.Y(n_209)
);

INVx11_ASAP7_75t_L g194 ( 
.A(n_122),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_194),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_180),
.A2(n_134),
.B1(n_111),
.B2(n_143),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_198),
.A2(n_212),
.B1(n_223),
.B2(n_6),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_201),
.B(n_202),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_166),
.A2(n_120),
.B(n_132),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_206),
.A2(n_193),
.B(n_154),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_162),
.A2(n_143),
.B1(n_115),
.B2(n_131),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_150),
.B(n_142),
.C(n_135),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_218),
.B(n_226),
.C(n_228),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_221),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_177),
.A2(n_131),
.B1(n_115),
.B2(n_145),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_158),
.B(n_98),
.C(n_141),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_182),
.B(n_122),
.C(n_2),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_229),
.A2(n_188),
.B1(n_177),
.B2(n_184),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_236),
.A2(n_238),
.B1(n_239),
.B2(n_256),
.Y(n_279)
);

OAI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_221),
.A2(n_152),
.B1(n_157),
.B2(n_151),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_229),
.A2(n_177),
.B1(n_185),
.B2(n_163),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_220),
.B(n_187),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_240),
.B(n_242),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_220),
.B(n_148),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_214),
.B(n_147),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_243),
.B(n_253),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_208),
.A2(n_156),
.B1(n_159),
.B2(n_169),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_244),
.A2(n_245),
.B1(n_247),
.B2(n_252),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_208),
.A2(n_156),
.B1(n_159),
.B2(n_160),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_200),
.B(n_218),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_246),
.B(n_228),
.C(n_205),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_221),
.A2(n_192),
.B1(n_146),
.B2(n_190),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_199),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_248),
.B(n_257),
.Y(n_289)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_227),
.Y(n_249)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_249),
.Y(n_300)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_197),
.Y(n_250)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_250),
.Y(n_274)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_197),
.Y(n_251)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_251),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_221),
.A2(n_189),
.B1(n_149),
.B2(n_155),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_199),
.B(n_174),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_214),
.B(n_168),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_254),
.B(n_265),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g295 ( 
.A1(n_255),
.A2(n_258),
.B(n_204),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_219),
.A2(n_175),
.B1(n_172),
.B2(n_161),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_211),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_206),
.A2(n_176),
.B(n_181),
.Y(n_258)
);

O2A1O1Ixp33_ASAP7_75t_L g259 ( 
.A1(n_219),
.A2(n_173),
.B(n_194),
.C(n_179),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_259),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_195),
.Y(n_260)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_260),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_195),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_261),
.Y(n_280)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_213),
.Y(n_262)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_262),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_225),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_263),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_L g264 ( 
.A1(n_223),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_264),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_216),
.B(n_3),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_224),
.B(n_3),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_270),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_267),
.A2(n_271),
.B1(n_203),
.B2(n_207),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_216),
.B(n_6),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_268),
.B(n_272),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_226),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_202),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_200),
.B(n_7),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_248),
.B(n_235),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_282),
.B(n_290),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_283),
.A2(n_285),
.B1(n_287),
.B2(n_302),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_241),
.A2(n_205),
.B1(n_212),
.B2(n_235),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_286),
.B(n_305),
.C(n_272),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_241),
.A2(n_236),
.B1(n_239),
.B2(n_267),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_243),
.B(n_196),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_290),
.B(n_294),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_246),
.B(n_213),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_SL g330 ( 
.A(n_293),
.B(n_215),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_242),
.B(n_196),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_295),
.A2(n_301),
.B(n_247),
.Y(n_307)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_250),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_297),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_261),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_298),
.Y(n_316)
);

XOR2x2_ASAP7_75t_L g299 ( 
.A(n_269),
.B(n_237),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_299),
.B(n_7),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_258),
.A2(n_234),
.B(n_198),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_269),
.A2(n_233),
.B1(n_230),
.B2(n_234),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_269),
.A2(n_230),
.B1(n_222),
.B2(n_217),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_303),
.B(n_306),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_237),
.B(n_232),
.C(n_209),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_255),
.A2(n_222),
.B1(n_217),
.B2(n_215),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_307),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_308),
.B(n_311),
.C(n_321),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_SL g309 ( 
.A(n_299),
.B(n_271),
.C(n_263),
.Y(n_309)
);

NOR2x1_ASAP7_75t_L g336 ( 
.A(n_309),
.B(n_283),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_295),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_310),
.B(n_326),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_240),
.C(n_254),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_281),
.Y(n_312)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_312),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_282),
.B(n_253),
.Y(n_313)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_313),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_289),
.B(n_268),
.Y(n_314)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_314),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_288),
.A2(n_252),
.B(n_259),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_317),
.A2(n_277),
.B(n_297),
.Y(n_359)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_280),
.Y(n_318)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_318),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_289),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_319),
.Y(n_345)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_281),
.Y(n_320)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_320),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_293),
.B(n_245),
.Y(n_321)
);

A2O1A1Ixp33_ASAP7_75t_L g322 ( 
.A1(n_294),
.A2(n_265),
.B(n_244),
.C(n_251),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_322),
.B(n_324),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_278),
.B(n_257),
.Y(n_323)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_323),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_305),
.B(n_262),
.C(n_232),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_275),
.B(n_231),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_325),
.B(n_274),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_273),
.B(n_256),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_329),
.B(n_277),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_330),
.B(n_331),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_286),
.B(n_204),
.C(n_249),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_304),
.A2(n_210),
.B1(n_260),
.B2(n_231),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_333),
.A2(n_328),
.B1(n_306),
.B2(n_329),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_273),
.B(n_227),
.C(n_260),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_334),
.B(n_335),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_336),
.B(n_317),
.Y(n_368)
);

OAI22x1_ASAP7_75t_SL g340 ( 
.A1(n_309),
.A2(n_276),
.B1(n_301),
.B2(n_287),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_340),
.A2(n_341),
.B1(n_342),
.B2(n_348),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_319),
.A2(n_279),
.B1(n_296),
.B2(n_275),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_332),
.A2(n_304),
.B1(n_276),
.B2(n_302),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_343),
.B(n_349),
.Y(n_363)
);

MAJx2_ASAP7_75t_L g344 ( 
.A(n_311),
.B(n_291),
.C(n_284),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_344),
.B(n_354),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_332),
.A2(n_279),
.B1(n_303),
.B2(n_285),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_307),
.A2(n_310),
.B1(n_328),
.B2(n_321),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_330),
.B(n_291),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_355),
.A2(n_333),
.B1(n_322),
.B2(n_327),
.Y(n_370)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_357),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_359),
.B(n_292),
.Y(n_379)
);

BUFx24_ASAP7_75t_SL g361 ( 
.A(n_346),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_361),
.B(n_379),
.Y(n_383)
);

XOR2x2_ASAP7_75t_L g365 ( 
.A(n_340),
.B(n_335),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_365),
.B(n_367),
.Y(n_397)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_347),
.Y(n_366)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_366),
.Y(n_395)
);

MAJx2_ASAP7_75t_L g367 ( 
.A(n_353),
.B(n_308),
.C(n_315),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_368),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_351),
.B(n_284),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_369),
.B(n_378),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_370),
.A2(n_339),
.B1(n_320),
.B2(n_312),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_353),
.B(n_324),
.C(n_331),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_371),
.B(n_373),
.C(n_375),
.Y(n_385)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_347),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_372),
.B(n_380),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_356),
.B(n_334),
.C(n_315),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_345),
.B(n_316),
.Y(n_374)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_374),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_356),
.B(n_316),
.C(n_318),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_357),
.Y(n_376)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_376),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_337),
.B(n_292),
.C(n_274),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_359),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g381 ( 
.A(n_360),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_381),
.B(n_300),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_363),
.A2(n_348),
.B1(n_342),
.B2(n_349),
.Y(n_384)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_384),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g387 ( 
.A1(n_363),
.A2(n_336),
.B1(n_338),
.B2(n_352),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_387),
.B(n_390),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_370),
.A2(n_338),
.B1(n_358),
.B2(n_350),
.Y(n_390)
);

AOI221xp5_ASAP7_75t_L g391 ( 
.A1(n_366),
.A2(n_355),
.B1(n_339),
.B2(n_344),
.C(n_350),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_391),
.A2(n_365),
.B1(n_362),
.B2(n_280),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_392),
.B(n_393),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_374),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_SL g407 ( 
.A(n_396),
.B(n_377),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_364),
.A2(n_337),
.B1(n_354),
.B2(n_298),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_398),
.A2(n_378),
.B1(n_380),
.B2(n_372),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_385),
.B(n_371),
.C(n_367),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_402),
.B(n_404),
.C(n_408),
.Y(n_414)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_382),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_403),
.B(n_392),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_385),
.B(n_375),
.C(n_373),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_405),
.B(n_407),
.Y(n_421)
);

AOI211xp5_ASAP7_75t_L g406 ( 
.A1(n_388),
.A2(n_382),
.B(n_376),
.C(n_362),
.Y(n_406)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_406),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_398),
.B(n_377),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_397),
.B(n_396),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_409),
.B(n_410),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_397),
.B(n_8),
.C(n_9),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_411),
.B(n_389),
.C(n_386),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_399),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_412),
.B(n_416),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_401),
.A2(n_383),
.B1(n_388),
.B2(n_393),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_406),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_417),
.B(n_419),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_402),
.A2(n_409),
.B(n_394),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_418),
.A2(n_404),
.B(n_411),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_405),
.A2(n_395),
.B1(n_389),
.B2(n_386),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_420),
.A2(n_422),
.B1(n_10),
.B2(n_12),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_421),
.B(n_400),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_423),
.B(n_425),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_421),
.B(n_407),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_426),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_413),
.B(n_408),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_427),
.B(n_431),
.Y(n_435)
);

AOI21xp33_ASAP7_75t_L g429 ( 
.A1(n_415),
.A2(n_8),
.B(n_10),
.Y(n_429)
);

OAI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_429),
.A2(n_424),
.B(n_430),
.Y(n_436)
);

OR2x2_ASAP7_75t_L g430 ( 
.A(n_420),
.B(n_8),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_SL g433 ( 
.A1(n_430),
.A2(n_412),
.B(n_422),
.Y(n_433)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_433),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_436),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_428),
.B(n_414),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_437),
.B(n_427),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_432),
.B(n_414),
.C(n_423),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_440),
.B(n_441),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_439),
.B(n_435),
.C(n_434),
.Y(n_442)
);

A2O1A1O1Ixp25_ASAP7_75t_L g444 ( 
.A1(n_442),
.A2(n_438),
.B(n_433),
.C(n_425),
.D(n_13),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_444),
.A2(n_443),
.B(n_10),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_445),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_446),
.B(n_12),
.Y(n_447)
);


endmodule