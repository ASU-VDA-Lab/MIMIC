module fake_jpeg_13323_n_107 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_107);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_107;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_106;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_29),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_23),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_24),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_42),
.Y(n_45)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_42),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_47),
.A2(n_42),
.B1(n_44),
.B2(n_39),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_48),
.B(n_51),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_43),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_2),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_36),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_41),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_56),
.B(n_57),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_41),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_43),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_58),
.B(n_62),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_61),
.A2(n_42),
.B(n_54),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_35),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_73),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_40),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_71),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_3),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_61),
.A2(n_38),
.B1(n_5),
.B2(n_6),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_74),
.A2(n_79),
.B1(n_15),
.B2(n_16),
.Y(n_89)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_65),
.A2(n_38),
.B1(n_6),
.B2(n_7),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_76),
.B(n_12),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_53),
.B(n_4),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_78),
.Y(n_84)
);

AO22x2_ASAP7_75t_L g78 ( 
.A1(n_65),
.A2(n_20),
.B1(n_33),
.B2(n_10),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_63),
.A2(n_4),
.B1(n_7),
.B2(n_11),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_66),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_81),
.B(n_87),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_85),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_63),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_13),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_14),
.Y(n_88)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_89),
.Y(n_97)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_90),
.B(n_82),
.C(n_84),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_78),
.C(n_21),
.Y(n_100)
);

AOI322xp5_ASAP7_75t_L g98 ( 
.A1(n_97),
.A2(n_88),
.A3(n_90),
.B1(n_78),
.B2(n_80),
.C1(n_25),
.C2(n_26),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_100),
.C(n_94),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_95),
.B(n_17),
.Y(n_99)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_99),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_95),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_102),
.Y(n_104)
);

OAI21x1_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_92),
.B(n_96),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_105),
.A2(n_18),
.B1(n_22),
.B2(n_27),
.Y(n_106)
);

NOR3xp33_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_30),
.C(n_32),
.Y(n_107)
);


endmodule