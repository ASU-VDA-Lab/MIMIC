module fake_netlist_6_1469_n_1801 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1801);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1801;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_1796;
wire n_170;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_297;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1774;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1475;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_162;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1721;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_130),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_3),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_118),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_7),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_160),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_58),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_64),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_81),
.Y(n_168)
);

INVx2_ASAP7_75t_SL g169 ( 
.A(n_58),
.Y(n_169)
);

INVx4_ASAP7_75t_R g170 ( 
.A(n_148),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_89),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_138),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_145),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_19),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_8),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_61),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_137),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_101),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_15),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_48),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_30),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_22),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_15),
.Y(n_183)
);

BUFx10_ASAP7_75t_L g184 ( 
.A(n_127),
.Y(n_184)
);

BUFx10_ASAP7_75t_L g185 ( 
.A(n_80),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_56),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_9),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_72),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_131),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_55),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_6),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_87),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_116),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_7),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_158),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_83),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_54),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_10),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_155),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_17),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_106),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_76),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_29),
.Y(n_203)
);

BUFx10_ASAP7_75t_L g204 ( 
.A(n_129),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_67),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_43),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_79),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_82),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_120),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_111),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_159),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_32),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_109),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_56),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_33),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_49),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_5),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_110),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_25),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_107),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_94),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_113),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_135),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_86),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_121),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_75),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_49),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_17),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_31),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_66),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_157),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_25),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_78),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_151),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_132),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_97),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_9),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_142),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_68),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_140),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_62),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_44),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_14),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_123),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_2),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_41),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_23),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_47),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_69),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_96),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_2),
.Y(n_251)
);

BUFx10_ASAP7_75t_L g252 ( 
.A(n_28),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_12),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_39),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_112),
.Y(n_255)
);

BUFx8_ASAP7_75t_SL g256 ( 
.A(n_122),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_156),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_32),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_100),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_50),
.Y(n_260)
);

BUFx5_ASAP7_75t_L g261 ( 
.A(n_98),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_51),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_139),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_143),
.Y(n_264)
);

BUFx10_ASAP7_75t_L g265 ( 
.A(n_6),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_117),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_73),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_16),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_104),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_21),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_99),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_43),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_13),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_103),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_144),
.Y(n_275)
);

BUFx3_ASAP7_75t_L g276 ( 
.A(n_26),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_114),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_42),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_45),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_45),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_57),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_20),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_14),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_124),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_84),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_105),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_153),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_28),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_134),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_95),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_16),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_27),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_29),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_13),
.Y(n_294)
);

INVx2_ASAP7_75t_SL g295 ( 
.A(n_92),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_39),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_37),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_44),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_26),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_19),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_115),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_108),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_54),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_146),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_93),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_24),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_3),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_23),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_57),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_24),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_88),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_10),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_18),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_53),
.Y(n_314)
);

BUFx5_ASAP7_75t_L g315 ( 
.A(n_126),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_1),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_60),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_8),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_1),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_174),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_R g321 ( 
.A(n_163),
.B(n_102),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_174),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_174),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_258),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_174),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_174),
.Y(n_326)
);

INVxp67_ASAP7_75t_SL g327 ( 
.A(n_191),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_261),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_261),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_257),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_191),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_227),
.Y(n_332)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_221),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_175),
.B(n_187),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_256),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_196),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_199),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_168),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_227),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_293),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_293),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_201),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_193),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_261),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_261),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_165),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_209),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_228),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_211),
.Y(n_349)
);

NOR2xp67_ASAP7_75t_L g350 ( 
.A(n_169),
.B(n_0),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_261),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_312),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_312),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_202),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_215),
.Y(n_355)
);

BUFx6f_ASAP7_75t_SL g356 ( 
.A(n_184),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_261),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_215),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_237),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_213),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_218),
.Y(n_361)
);

INVxp33_ASAP7_75t_SL g362 ( 
.A(n_166),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_237),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_184),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_207),
.Y(n_365)
);

NOR2xp67_ASAP7_75t_L g366 ( 
.A(n_169),
.B(n_0),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_253),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_223),
.Y(n_368)
);

NOR2xp67_ASAP7_75t_L g369 ( 
.A(n_294),
.B(n_4),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_224),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_184),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_172),
.B(n_295),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_226),
.Y(n_373)
);

INVxp67_ASAP7_75t_SL g374 ( 
.A(n_253),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_276),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_241),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_264),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_230),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_231),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_276),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_162),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_172),
.B(n_4),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_164),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_186),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_234),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_190),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_225),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_185),
.Y(n_388)
);

BUFx2_ASAP7_75t_L g389 ( 
.A(n_166),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_236),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_238),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_239),
.Y(n_392)
);

INVxp33_ASAP7_75t_SL g393 ( 
.A(n_179),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_240),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_197),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_372),
.B(n_295),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_387),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_320),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_320),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_382),
.B(n_322),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_322),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_367),
.B(n_173),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_323),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_333),
.B(n_220),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_387),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_323),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_336),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_374),
.B(n_173),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_325),
.B(n_161),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_325),
.B(n_161),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_387),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_389),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_326),
.Y(n_413)
);

OR2x6_ASAP7_75t_L g414 ( 
.A(n_350),
.B(n_294),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_326),
.B(n_346),
.Y(n_415)
);

AND2x2_ASAP7_75t_L g416 ( 
.A(n_346),
.B(n_250),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_387),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_381),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_381),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_346),
.B(n_167),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_383),
.Y(n_421)
);

INVx5_ASAP7_75t_L g422 ( 
.A(n_387),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_327),
.B(n_167),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_327),
.B(n_171),
.Y(n_424)
);

INVx6_ASAP7_75t_L g425 ( 
.A(n_387),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_337),
.B(n_235),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_328),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_334),
.A2(n_262),
.B1(n_316),
.B2(n_273),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_328),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_383),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_328),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_355),
.B(n_171),
.Y(n_432)
);

AND2x4_ASAP7_75t_L g433 ( 
.A(n_329),
.B(n_250),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_SL g434 ( 
.A(n_364),
.B(n_252),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_384),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_362),
.B(n_274),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_384),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_329),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_329),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_386),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_386),
.Y(n_441)
);

BUFx2_ASAP7_75t_L g442 ( 
.A(n_324),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_364),
.B(n_252),
.Y(n_443)
);

CKINVDCx8_ASAP7_75t_R g444 ( 
.A(n_371),
.Y(n_444)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_371),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_395),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_395),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_388),
.B(n_185),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_344),
.Y(n_449)
);

AND2x4_ASAP7_75t_SL g450 ( 
.A(n_385),
.B(n_185),
.Y(n_450)
);

BUFx2_ASAP7_75t_L g451 ( 
.A(n_389),
.Y(n_451)
);

INVx4_ASAP7_75t_L g452 ( 
.A(n_344),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_331),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_344),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_345),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_331),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_345),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g458 ( 
.A(n_342),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g459 ( 
.A(n_350),
.Y(n_459)
);

INVx4_ASAP7_75t_L g460 ( 
.A(n_345),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_351),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_332),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_351),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_351),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_332),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_388),
.B(n_204),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_357),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_426),
.B(n_347),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_442),
.Y(n_469)
);

OR2x6_ASAP7_75t_L g470 ( 
.A(n_414),
.B(n_274),
.Y(n_470)
);

OR2x6_ASAP7_75t_L g471 ( 
.A(n_414),
.B(n_277),
.Y(n_471)
);

NAND2xp33_ASAP7_75t_SL g472 ( 
.A(n_448),
.B(n_356),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g473 ( 
.A(n_433),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_404),
.B(n_349),
.Y(n_474)
);

AND3x2_ASAP7_75t_L g475 ( 
.A(n_434),
.B(n_183),
.C(n_277),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_452),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_452),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_452),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_429),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_396),
.B(n_360),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_460),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_460),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_429),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_404),
.B(n_361),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_460),
.Y(n_485)
);

NAND3xp33_ASAP7_75t_L g486 ( 
.A(n_396),
.B(n_369),
.C(n_366),
.Y(n_486)
);

INVx3_ASAP7_75t_L g487 ( 
.A(n_460),
.Y(n_487)
);

INVx1_ASAP7_75t_SL g488 ( 
.A(n_442),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_433),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_434),
.B(n_368),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_429),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_431),
.Y(n_492)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_402),
.B(n_355),
.Y(n_493)
);

AOI22xp33_ASAP7_75t_L g494 ( 
.A1(n_402),
.A2(n_330),
.B1(n_348),
.B2(n_366),
.Y(n_494)
);

OAI21xp33_ASAP7_75t_SL g495 ( 
.A1(n_400),
.A2(n_369),
.B(n_359),
.Y(n_495)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_427),
.Y(n_496)
);

OR2x6_ASAP7_75t_L g497 ( 
.A(n_414),
.B(n_301),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_433),
.Y(n_498)
);

INVx1_ASAP7_75t_SL g499 ( 
.A(n_451),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_433),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_459),
.B(n_370),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_444),
.Y(n_502)
);

AOI22xp33_ASAP7_75t_L g503 ( 
.A1(n_402),
.A2(n_330),
.B1(n_393),
.B2(n_232),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_433),
.Y(n_504)
);

BUFx10_ASAP7_75t_L g505 ( 
.A(n_407),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_459),
.B(n_373),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_431),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_436),
.B(n_378),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_436),
.B(n_379),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_408),
.B(n_358),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_400),
.B(n_390),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_408),
.B(n_358),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_431),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_443),
.B(n_394),
.Y(n_514)
);

BUFx2_ASAP7_75t_L g515 ( 
.A(n_451),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_398),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_439),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_443),
.B(n_321),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_408),
.B(n_359),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_398),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_423),
.B(n_391),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_427),
.Y(n_522)
);

BUFx3_ASAP7_75t_L g523 ( 
.A(n_415),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_420),
.B(n_330),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_427),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_439),
.Y(n_526)
);

INVx1_ASAP7_75t_SL g527 ( 
.A(n_450),
.Y(n_527)
);

NAND3xp33_ASAP7_75t_L g528 ( 
.A(n_416),
.B(n_424),
.C(n_423),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_439),
.Y(n_529)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_415),
.Y(n_530)
);

INVx2_ASAP7_75t_SL g531 ( 
.A(n_414),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_399),
.Y(n_532)
);

BUFx4f_ASAP7_75t_L g533 ( 
.A(n_427),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_420),
.B(n_244),
.Y(n_534)
);

NAND3xp33_ASAP7_75t_L g535 ( 
.A(n_416),
.B(n_301),
.C(n_177),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_399),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_416),
.B(n_424),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_401),
.Y(n_538)
);

BUFx4f_ASAP7_75t_L g539 ( 
.A(n_427),
.Y(n_539)
);

OR2x2_ASAP7_75t_L g540 ( 
.A(n_412),
.B(n_363),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_458),
.B(n_392),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_458),
.Y(n_542)
);

INVxp67_ASAP7_75t_SL g543 ( 
.A(n_427),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_449),
.Y(n_544)
);

OR2x2_ASAP7_75t_L g545 ( 
.A(n_412),
.B(n_363),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_401),
.Y(n_546)
);

OR2x2_ASAP7_75t_L g547 ( 
.A(n_409),
.B(n_375),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_409),
.B(n_249),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_449),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_466),
.B(n_335),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_403),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_449),
.Y(n_552)
);

AO22x2_ASAP7_75t_L g553 ( 
.A1(n_432),
.A2(n_198),
.B1(n_254),
.B2(n_318),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_403),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_427),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_406),
.Y(n_556)
);

INVx1_ASAP7_75t_SL g557 ( 
.A(n_450),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_461),
.Y(n_558)
);

CKINVDCx6p67_ASAP7_75t_R g559 ( 
.A(n_445),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_461),
.Y(n_560)
);

INVx1_ASAP7_75t_SL g561 ( 
.A(n_450),
.Y(n_561)
);

NAND3xp33_ASAP7_75t_SL g562 ( 
.A(n_444),
.B(n_291),
.C(n_280),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_438),
.Y(n_563)
);

BUFx2_ASAP7_75t_L g564 ( 
.A(n_414),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_406),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_461),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_410),
.B(n_255),
.Y(n_567)
);

NOR3xp33_ASAP7_75t_L g568 ( 
.A(n_428),
.B(n_214),
.C(n_206),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_467),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_438),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_410),
.B(n_267),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_467),
.Y(n_572)
);

INVx4_ASAP7_75t_L g573 ( 
.A(n_438),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_413),
.Y(n_574)
);

NAND3xp33_ASAP7_75t_L g575 ( 
.A(n_432),
.B(n_188),
.C(n_176),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_453),
.B(n_456),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_444),
.B(n_204),
.Y(n_577)
);

INVx1_ASAP7_75t_SL g578 ( 
.A(n_445),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_467),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_425),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_413),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_454),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_438),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_414),
.B(n_269),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_418),
.B(n_356),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_454),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_438),
.B(n_271),
.Y(n_587)
);

OR2x6_ASAP7_75t_L g588 ( 
.A(n_418),
.B(n_195),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_454),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_438),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_419),
.B(n_356),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_419),
.B(n_356),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_421),
.B(n_375),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_454),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_438),
.B(n_205),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_455),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_425),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_421),
.B(n_204),
.Y(n_598)
);

OR2x2_ASAP7_75t_L g599 ( 
.A(n_430),
.B(n_380),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_455),
.B(n_208),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_455),
.B(n_210),
.Y(n_601)
);

NAND3xp33_ASAP7_75t_L g602 ( 
.A(n_430),
.B(n_233),
.C(n_222),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_457),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_435),
.B(n_178),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_435),
.B(n_380),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_455),
.B(n_259),
.Y(n_606)
);

INVx4_ASAP7_75t_L g607 ( 
.A(n_455),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_437),
.B(n_338),
.Y(n_608)
);

INVx4_ASAP7_75t_L g609 ( 
.A(n_455),
.Y(n_609)
);

INVx5_ASAP7_75t_L g610 ( 
.A(n_455),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_457),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_463),
.B(n_263),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_457),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_437),
.B(n_178),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_457),
.Y(n_615)
);

AOI22xp33_ASAP7_75t_L g616 ( 
.A1(n_440),
.A2(n_303),
.B1(n_281),
.B2(n_260),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_464),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_528),
.B(n_225),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_473),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_511),
.B(n_189),
.Y(n_620)
);

OR2x6_ASAP7_75t_L g621 ( 
.A(n_542),
.B(n_428),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_480),
.B(n_189),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_528),
.B(n_487),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_523),
.B(n_463),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_576),
.B(n_440),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_473),
.Y(n_626)
);

NOR3xp33_ASAP7_75t_L g627 ( 
.A(n_562),
.B(n_446),
.C(n_441),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_484),
.B(n_192),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_487),
.B(n_225),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_523),
.B(n_463),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_499),
.B(n_493),
.Y(n_631)
);

HB1xp67_ASAP7_75t_L g632 ( 
.A(n_499),
.Y(n_632)
);

BUFx6f_ASAP7_75t_L g633 ( 
.A(n_498),
.Y(n_633)
);

INVxp67_ASAP7_75t_L g634 ( 
.A(n_469),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_530),
.A2(n_248),
.B1(n_217),
.B2(n_243),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_489),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_530),
.B(n_463),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_521),
.B(n_192),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_537),
.B(n_463),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_489),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_500),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_500),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_504),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_504),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_487),
.B(n_463),
.Y(n_645)
);

BUFx3_ASAP7_75t_L g646 ( 
.A(n_542),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_516),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_493),
.B(n_343),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_468),
.B(n_463),
.Y(n_649)
);

NAND3xp33_ASAP7_75t_L g650 ( 
.A(n_486),
.B(n_509),
.C(n_508),
.Y(n_650)
);

NOR3xp33_ASAP7_75t_L g651 ( 
.A(n_518),
.B(n_446),
.C(n_441),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_576),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_516),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_476),
.B(n_464),
.Y(n_654)
);

AND2x4_ASAP7_75t_SL g655 ( 
.A(n_505),
.B(n_354),
.Y(n_655)
);

INVxp67_ASAP7_75t_L g656 ( 
.A(n_515),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_599),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_476),
.B(n_464),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_477),
.B(n_464),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_540),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_477),
.B(n_397),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_478),
.B(n_397),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_478),
.B(n_397),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_599),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_531),
.B(n_225),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_524),
.B(n_474),
.Y(n_666)
);

NAND2xp33_ASAP7_75t_L g667 ( 
.A(n_531),
.B(n_534),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_501),
.B(n_506),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_510),
.B(n_365),
.Y(n_669)
);

AOI21xp5_ASAP7_75t_L g670 ( 
.A1(n_587),
.A2(n_422),
.B(n_405),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_486),
.B(n_564),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_520),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_564),
.B(n_284),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_481),
.B(n_411),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_540),
.B(n_545),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_520),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_532),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_481),
.B(n_225),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_532),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_536),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_536),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_482),
.B(n_261),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_482),
.B(n_411),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_510),
.B(n_447),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_L g685 ( 
.A1(n_553),
.A2(n_245),
.B1(n_288),
.B2(n_296),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_538),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_L g687 ( 
.A1(n_553),
.A2(n_310),
.B1(n_314),
.B2(n_308),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_485),
.B(n_548),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_SL g689 ( 
.A(n_505),
.B(n_376),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_545),
.B(n_284),
.Y(n_690)
);

BUFx3_ASAP7_75t_L g691 ( 
.A(n_505),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_485),
.B(n_567),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_571),
.B(n_411),
.Y(n_693)
);

NAND3xp33_ASAP7_75t_L g694 ( 
.A(n_503),
.B(n_494),
.C(n_495),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_538),
.Y(n_695)
);

INVxp67_ASAP7_75t_L g696 ( 
.A(n_515),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_547),
.B(n_285),
.Y(n_697)
);

O2A1O1Ixp33_ASAP7_75t_L g698 ( 
.A1(n_495),
.A2(n_447),
.B(n_462),
.C(n_456),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_547),
.B(n_417),
.Y(n_699)
);

OR2x2_ASAP7_75t_L g700 ( 
.A(n_488),
.B(n_334),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_546),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_546),
.Y(n_702)
);

INVxp33_ASAP7_75t_L g703 ( 
.A(n_608),
.Y(n_703)
);

OAI22xp33_ASAP7_75t_L g704 ( 
.A1(n_470),
.A2(n_377),
.B1(n_266),
.B2(n_275),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_490),
.B(n_285),
.Y(n_705)
);

INVx2_ASAP7_75t_SL g706 ( 
.A(n_512),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_512),
.B(n_417),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_519),
.B(n_252),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_551),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_519),
.A2(n_286),
.B1(n_287),
.B2(n_289),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_551),
.Y(n_711)
);

HB1xp67_ASAP7_75t_L g712 ( 
.A(n_588),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_554),
.B(n_417),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_554),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_475),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_556),
.B(n_290),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_584),
.B(n_286),
.Y(n_717)
);

BUFx5_ASAP7_75t_L g718 ( 
.A(n_582),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_556),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_514),
.B(n_287),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_565),
.B(n_302),
.Y(n_721)
);

NAND2xp33_ASAP7_75t_L g722 ( 
.A(n_565),
.B(n_261),
.Y(n_722)
);

AOI21xp5_ASAP7_75t_L g723 ( 
.A1(n_543),
.A2(n_539),
.B(n_533),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_574),
.B(n_581),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_574),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_581),
.B(n_315),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_582),
.B(n_453),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_580),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_577),
.B(n_604),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_586),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_586),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_611),
.B(n_462),
.Y(n_732)
);

NOR2xp67_ASAP7_75t_L g733 ( 
.A(n_550),
.B(n_465),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_479),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_472),
.A2(n_289),
.B1(n_304),
.B2(n_305),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_611),
.B(n_315),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_613),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_613),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_615),
.B(n_465),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_615),
.Y(n_740)
);

AOI22xp5_ASAP7_75t_L g741 ( 
.A1(n_470),
.A2(n_304),
.B1(n_305),
.B2(n_311),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_585),
.B(n_311),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_496),
.B(n_522),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_593),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_614),
.B(n_317),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_479),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_483),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_575),
.B(n_317),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_L g749 ( 
.A1(n_553),
.A2(n_292),
.B1(n_309),
.B2(n_315),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_505),
.B(n_265),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_563),
.B(n_315),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_496),
.B(n_315),
.Y(n_752)
);

AND2x6_ASAP7_75t_SL g753 ( 
.A(n_588),
.B(n_339),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_496),
.B(n_315),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_522),
.B(n_315),
.Y(n_755)
);

INVxp67_ASAP7_75t_L g756 ( 
.A(n_605),
.Y(n_756)
);

BUFx6f_ASAP7_75t_L g757 ( 
.A(n_580),
.Y(n_757)
);

NAND2xp33_ASAP7_75t_SL g758 ( 
.A(n_502),
.B(n_179),
.Y(n_758)
);

INVx4_ASAP7_75t_L g759 ( 
.A(n_563),
.Y(n_759)
);

INVx4_ASAP7_75t_L g760 ( 
.A(n_563),
.Y(n_760)
);

O2A1O1Ixp33_ASAP7_75t_L g761 ( 
.A1(n_575),
.A2(n_353),
.B(n_352),
.C(n_341),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_591),
.B(n_194),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_553),
.A2(n_315),
.B1(n_180),
.B2(n_181),
.Y(n_763)
);

BUFx2_ASAP7_75t_L g764 ( 
.A(n_578),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_592),
.B(n_200),
.Y(n_765)
);

AND2x6_ASAP7_75t_SL g766 ( 
.A(n_588),
.B(n_339),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_589),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_568),
.A2(n_278),
.B1(n_180),
.B2(n_182),
.Y(n_768)
);

AOI22xp5_ASAP7_75t_SL g769 ( 
.A1(n_502),
.A2(n_319),
.B1(n_313),
.B2(n_307),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_597),
.Y(n_770)
);

INVx4_ASAP7_75t_L g771 ( 
.A(n_563),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_589),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_578),
.B(n_265),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_483),
.Y(n_774)
);

BUFx5_ASAP7_75t_L g775 ( 
.A(n_597),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_491),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_598),
.B(n_203),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_522),
.B(n_425),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_491),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_525),
.B(n_425),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_492),
.Y(n_781)
);

AND2x6_ASAP7_75t_L g782 ( 
.A(n_525),
.B(n_555),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_492),
.Y(n_783)
);

INVx4_ASAP7_75t_L g784 ( 
.A(n_563),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_507),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_525),
.B(n_425),
.Y(n_786)
);

OAI21xp5_ASAP7_75t_L g787 ( 
.A1(n_623),
.A2(n_533),
.B(n_539),
.Y(n_787)
);

OAI21xp5_ASAP7_75t_L g788 ( 
.A1(n_623),
.A2(n_533),
.B(n_539),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_668),
.B(n_470),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_668),
.B(n_470),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_650),
.A2(n_497),
.B1(n_470),
.B2(n_471),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_636),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_723),
.A2(n_639),
.B(n_645),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_633),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_631),
.B(n_527),
.Y(n_795)
);

INVx4_ASAP7_75t_L g796 ( 
.A(n_633),
.Y(n_796)
);

AOI22xp5_ASAP7_75t_L g797 ( 
.A1(n_666),
.A2(n_471),
.B1(n_497),
.B2(n_541),
.Y(n_797)
);

AND2x6_ASAP7_75t_SL g798 ( 
.A(n_621),
.B(n_588),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_666),
.B(n_622),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_703),
.B(n_557),
.Y(n_800)
);

AOI21x1_ASAP7_75t_L g801 ( 
.A1(n_629),
.A2(n_595),
.B(n_600),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_622),
.B(n_756),
.Y(n_802)
);

INVx1_ASAP7_75t_SL g803 ( 
.A(n_632),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_641),
.Y(n_804)
);

NOR2xp67_ASAP7_75t_L g805 ( 
.A(n_634),
.B(n_535),
.Y(n_805)
);

AOI21x1_ASAP7_75t_L g806 ( 
.A1(n_629),
.A2(n_601),
.B(n_606),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_744),
.B(n_471),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_641),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_649),
.A2(n_573),
.B(n_609),
.Y(n_809)
);

OAI22xp5_ASAP7_75t_L g810 ( 
.A1(n_688),
.A2(n_471),
.B1(n_497),
.B2(n_561),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_624),
.A2(n_573),
.B(n_609),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_620),
.B(n_471),
.Y(n_812)
);

O2A1O1Ixp33_ASAP7_75t_SL g813 ( 
.A1(n_618),
.A2(n_535),
.B(n_612),
.C(n_602),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_630),
.A2(n_573),
.B(n_609),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_620),
.A2(n_729),
.B1(n_671),
.B2(n_619),
.Y(n_815)
);

OR2x6_ASAP7_75t_L g816 ( 
.A(n_764),
.B(n_497),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_692),
.B(n_497),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_637),
.A2(n_607),
.B(n_583),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_693),
.A2(n_607),
.B(n_583),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_707),
.A2(n_607),
.B(n_583),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_633),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_675),
.B(n_559),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_697),
.B(n_588),
.Y(n_823)
);

OAI21xp5_ASAP7_75t_L g824 ( 
.A1(n_618),
.A2(n_555),
.B(n_570),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_697),
.B(n_555),
.Y(n_825)
);

OAI21xp5_ASAP7_75t_L g826 ( 
.A1(n_682),
.A2(n_570),
.B(n_596),
.Y(n_826)
);

AOI22xp5_ASAP7_75t_L g827 ( 
.A1(n_729),
.A2(n_570),
.B1(n_596),
.B2(n_559),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_647),
.Y(n_828)
);

AOI21x1_ASAP7_75t_L g829 ( 
.A1(n_682),
.A2(n_579),
.B(n_544),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_647),
.Y(n_830)
);

INVx2_ASAP7_75t_SL g831 ( 
.A(n_648),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_675),
.B(n_596),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_759),
.A2(n_583),
.B(n_590),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_676),
.B(n_594),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_653),
.Y(n_835)
);

BUFx3_ASAP7_75t_L g836 ( 
.A(n_646),
.Y(n_836)
);

HB1xp67_ASAP7_75t_L g837 ( 
.A(n_656),
.Y(n_837)
);

INVx4_ASAP7_75t_L g838 ( 
.A(n_633),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_759),
.A2(n_583),
.B(n_590),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_733),
.B(n_590),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_640),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_642),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_680),
.B(n_594),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_660),
.B(n_616),
.Y(n_844)
);

CKINVDCx20_ASAP7_75t_R g845 ( 
.A(n_655),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_708),
.B(n_669),
.Y(n_846)
);

OAI321xp33_ASAP7_75t_L g847 ( 
.A1(n_749),
.A2(n_602),
.A3(n_340),
.B1(n_353),
.B2(n_352),
.C(n_341),
.Y(n_847)
);

AOI22xp33_ASAP7_75t_L g848 ( 
.A1(n_763),
.A2(n_265),
.B1(n_181),
.B2(n_300),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_701),
.B(n_603),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_709),
.B(n_603),
.Y(n_850)
);

INVxp67_ASAP7_75t_L g851 ( 
.A(n_773),
.Y(n_851)
);

OAI22xp5_ASAP7_75t_L g852 ( 
.A1(n_694),
.A2(n_590),
.B1(n_617),
.B2(n_526),
.Y(n_852)
);

INVxp67_ASAP7_75t_L g853 ( 
.A(n_690),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_760),
.A2(n_590),
.B(n_610),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_711),
.B(n_617),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_714),
.B(n_507),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_725),
.B(n_513),
.Y(n_857)
);

AND2x4_ASAP7_75t_L g858 ( 
.A(n_625),
.B(n_513),
.Y(n_858)
);

NOR2xp67_ASAP7_75t_L g859 ( 
.A(n_696),
.B(n_517),
.Y(n_859)
);

INVx1_ASAP7_75t_SL g860 ( 
.A(n_646),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_760),
.A2(n_610),
.B(n_422),
.Y(n_861)
);

INVx2_ASAP7_75t_SL g862 ( 
.A(n_684),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_718),
.B(n_517),
.Y(n_863)
);

O2A1O1Ixp5_ASAP7_75t_L g864 ( 
.A1(n_665),
.A2(n_558),
.B(n_579),
.C(n_572),
.Y(n_864)
);

HB1xp67_ASAP7_75t_L g865 ( 
.A(n_706),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_771),
.A2(n_610),
.B(n_422),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_653),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_771),
.A2(n_610),
.B(n_422),
.Y(n_868)
);

INVx2_ASAP7_75t_SL g869 ( 
.A(n_684),
.Y(n_869)
);

AOI21x1_ASAP7_75t_L g870 ( 
.A1(n_654),
.A2(n_549),
.B(n_572),
.Y(n_870)
);

BUFx2_ASAP7_75t_L g871 ( 
.A(n_700),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_784),
.A2(n_610),
.B(n_422),
.Y(n_872)
);

A2O1A1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_687),
.A2(n_298),
.B(n_278),
.C(n_279),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_672),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_784),
.A2(n_610),
.B(n_422),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_699),
.B(n_526),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_625),
.B(n_529),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_724),
.B(n_529),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_652),
.B(n_544),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_658),
.A2(n_422),
.B(n_569),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_659),
.A2(n_569),
.B(n_566),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_672),
.B(n_549),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_690),
.B(n_340),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_743),
.A2(n_566),
.B(n_560),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_677),
.B(n_552),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_718),
.B(n_552),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_677),
.B(n_679),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_679),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_638),
.B(n_657),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_681),
.B(n_558),
.Y(n_890)
);

AOI21x1_ASAP7_75t_L g891 ( 
.A1(n_661),
.A2(n_560),
.B(n_357),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_667),
.A2(n_357),
.B(n_170),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_681),
.B(n_212),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_686),
.B(n_216),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_664),
.B(n_219),
.Y(n_895)
);

NOR2x1_ASAP7_75t_R g896 ( 
.A(n_691),
.B(n_182),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_686),
.Y(n_897)
);

OAI21xp33_ASAP7_75t_L g898 ( 
.A1(n_768),
.A2(n_319),
.B(n_313),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_643),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_695),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_628),
.B(n_229),
.Y(n_901)
);

BUFx4f_ASAP7_75t_L g902 ( 
.A(n_655),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_695),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_702),
.B(n_242),
.Y(n_904)
);

HB1xp67_ASAP7_75t_L g905 ( 
.A(n_712),
.Y(n_905)
);

INVx2_ASAP7_75t_SL g906 ( 
.A(n_750),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_702),
.B(n_246),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_719),
.B(n_247),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_719),
.B(n_251),
.Y(n_909)
);

BUFx6f_ASAP7_75t_L g910 ( 
.A(n_728),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_644),
.B(n_268),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_651),
.B(n_270),
.Y(n_912)
);

OAI21xp5_ASAP7_75t_L g913 ( 
.A1(n_662),
.A2(n_272),
.B(n_306),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_734),
.Y(n_914)
);

AND2x4_ASAP7_75t_L g915 ( 
.A(n_626),
.B(n_63),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_730),
.Y(n_916)
);

NAND2xp33_ASAP7_75t_L g917 ( 
.A(n_782),
.B(n_307),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_691),
.B(n_297),
.Y(n_918)
);

AOI21x1_ASAP7_75t_L g919 ( 
.A1(n_663),
.A2(n_59),
.B(n_154),
.Y(n_919)
);

INVx11_ASAP7_75t_L g920 ( 
.A(n_782),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_728),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_674),
.A2(n_299),
.B(n_297),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_731),
.Y(n_923)
);

NOR2xp67_ASAP7_75t_L g924 ( 
.A(n_715),
.B(n_128),
.Y(n_924)
);

INVx2_ASAP7_75t_SL g925 ( 
.A(n_757),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_748),
.B(n_283),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_737),
.B(n_283),
.Y(n_927)
);

INVxp33_ASAP7_75t_SL g928 ( 
.A(n_689),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_705),
.B(n_282),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_718),
.B(n_282),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_683),
.A2(n_279),
.B(n_152),
.Y(n_931)
);

AOI21xp33_ASAP7_75t_L g932 ( 
.A1(n_705),
.A2(n_5),
.B(n_11),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_738),
.B(n_11),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_740),
.B(n_12),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_716),
.B(n_721),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_745),
.B(n_18),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_713),
.Y(n_937)
);

AND2x2_ASAP7_75t_L g938 ( 
.A(n_777),
.B(n_20),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_745),
.B(n_720),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_720),
.B(n_21),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_727),
.B(n_22),
.Y(n_941)
);

HB1xp67_ASAP7_75t_L g942 ( 
.A(n_627),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_767),
.Y(n_943)
);

NAND2x1p5_ASAP7_75t_L g944 ( 
.A(n_757),
.B(n_150),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_777),
.B(n_27),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_732),
.B(n_30),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_734),
.Y(n_947)
);

OAI21xp5_ASAP7_75t_L g948 ( 
.A1(n_665),
.A2(n_149),
.B(n_147),
.Y(n_948)
);

OAI21xp5_ASAP7_75t_L g949 ( 
.A1(n_678),
.A2(n_141),
.B(n_136),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_769),
.B(n_31),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_778),
.A2(n_133),
.B(n_125),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_739),
.B(n_33),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_698),
.B(n_34),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_772),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_718),
.B(n_34),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_780),
.A2(n_119),
.B(n_91),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_786),
.A2(n_90),
.B(n_85),
.Y(n_957)
);

AND2x6_ASAP7_75t_SL g958 ( 
.A(n_621),
.B(n_35),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_746),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_746),
.Y(n_960)
);

OAI21xp5_ASAP7_75t_L g961 ( 
.A1(n_678),
.A2(n_77),
.B(n_74),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_670),
.A2(n_71),
.B(n_70),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_718),
.B(n_65),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_747),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_718),
.B(n_35),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_752),
.A2(n_36),
.B(n_37),
.Y(n_966)
);

INVx3_ASAP7_75t_L g967 ( 
.A(n_757),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_747),
.Y(n_968)
);

A2O1A1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_687),
.A2(n_36),
.B(n_38),
.C(n_40),
.Y(n_969)
);

AOI22xp5_ASAP7_75t_L g970 ( 
.A1(n_717),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_774),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_774),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_704),
.B(n_42),
.Y(n_973)
);

AND2x4_ASAP7_75t_L g974 ( 
.A(n_836),
.B(n_673),
.Y(n_974)
);

O2A1O1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_939),
.A2(n_742),
.B(n_762),
.C(n_765),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_799),
.B(n_635),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_802),
.B(n_758),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_793),
.A2(n_770),
.B(n_757),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_853),
.B(n_741),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_929),
.B(n_621),
.Y(n_980)
);

OAI21xp5_ASAP7_75t_L g981 ( 
.A1(n_832),
.A2(n_726),
.B(n_736),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_794),
.Y(n_982)
);

INVx4_ASAP7_75t_L g983 ( 
.A(n_794),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_883),
.B(n_749),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_937),
.B(n_635),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_804),
.Y(n_986)
);

O2A1O1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_929),
.A2(n_726),
.B(n_763),
.C(n_736),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_815),
.B(n_710),
.Y(n_988)
);

NAND2xp33_ASAP7_75t_SL g989 ( 
.A(n_936),
.B(n_685),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_822),
.B(n_735),
.Y(n_990)
);

NAND3xp33_ASAP7_75t_SL g991 ( 
.A(n_926),
.B(n_768),
.C(n_685),
.Y(n_991)
);

OAI22xp33_ASAP7_75t_L g992 ( 
.A1(n_940),
.A2(n_754),
.B1(n_755),
.B2(n_770),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_795),
.B(n_785),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_873),
.A2(n_785),
.B1(n_783),
.B2(n_781),
.Y(n_994)
);

BUFx2_ASAP7_75t_L g995 ( 
.A(n_803),
.Y(n_995)
);

OR2x6_ASAP7_75t_L g996 ( 
.A(n_816),
.B(n_770),
.Y(n_996)
);

O2A1O1Ixp5_ASAP7_75t_SL g997 ( 
.A1(n_932),
.A2(n_751),
.B(n_722),
.C(n_753),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_822),
.B(n_766),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_851),
.B(n_770),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_804),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_832),
.B(n_783),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_809),
.A2(n_751),
.B(n_781),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_828),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_935),
.A2(n_779),
.B(n_776),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_819),
.A2(n_779),
.B(n_776),
.Y(n_1005)
);

AOI22xp33_ASAP7_75t_L g1006 ( 
.A1(n_938),
.A2(n_782),
.B1(n_775),
.B2(n_761),
.Y(n_1006)
);

HB1xp67_ASAP7_75t_L g1007 ( 
.A(n_837),
.Y(n_1007)
);

BUFx6f_ASAP7_75t_L g1008 ( 
.A(n_794),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_820),
.A2(n_775),
.B(n_782),
.Y(n_1009)
);

BUFx2_ASAP7_75t_L g1010 ( 
.A(n_871),
.Y(n_1010)
);

NAND2x1p5_ASAP7_75t_L g1011 ( 
.A(n_796),
.B(n_775),
.Y(n_1011)
);

BUFx6f_ASAP7_75t_L g1012 ( 
.A(n_794),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_845),
.Y(n_1013)
);

O2A1O1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_973),
.A2(n_46),
.B(n_47),
.C(n_48),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_846),
.B(n_46),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_889),
.B(n_841),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_817),
.A2(n_775),
.B(n_51),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_889),
.B(n_775),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_910),
.Y(n_1019)
);

INVx3_ASAP7_75t_L g1020 ( 
.A(n_910),
.Y(n_1020)
);

A2O1A1Ixp33_ASAP7_75t_L g1021 ( 
.A1(n_945),
.A2(n_775),
.B(n_52),
.C(n_53),
.Y(n_1021)
);

BUFx12f_ASAP7_75t_L g1022 ( 
.A(n_831),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_844),
.B(n_50),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_842),
.B(n_52),
.Y(n_1024)
);

CKINVDCx20_ASAP7_75t_R g1025 ( 
.A(n_845),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_787),
.A2(n_55),
.B(n_788),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_899),
.B(n_916),
.Y(n_1027)
);

O2A1O1Ixp33_ASAP7_75t_SL g1028 ( 
.A1(n_963),
.A2(n_969),
.B(n_812),
.C(n_823),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_923),
.B(n_789),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_897),
.B(n_790),
.Y(n_1030)
);

BUFx2_ASAP7_75t_L g1031 ( 
.A(n_837),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_910),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_SL g1033 ( 
.A(n_797),
.B(n_928),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_897),
.B(n_942),
.Y(n_1034)
);

INVx3_ASAP7_75t_L g1035 ( 
.A(n_910),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_873),
.A2(n_969),
.B1(n_848),
.B2(n_973),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_830),
.B(n_835),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_830),
.B(n_835),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_792),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_800),
.B(n_928),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_918),
.B(n_895),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_862),
.B(n_869),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_808),
.Y(n_1043)
);

INVxp67_ASAP7_75t_L g1044 ( 
.A(n_942),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_867),
.Y(n_1045)
);

A2O1A1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_901),
.A2(n_807),
.B(n_805),
.C(n_847),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_874),
.B(n_888),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_874),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_SL g1049 ( 
.A(n_902),
.B(n_800),
.Y(n_1049)
);

AND2x4_ASAP7_75t_L g1050 ( 
.A(n_836),
.B(n_862),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_888),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_900),
.Y(n_1052)
);

A2O1A1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_901),
.A2(n_791),
.B(n_913),
.C(n_953),
.Y(n_1053)
);

NOR3xp33_ASAP7_75t_SL g1054 ( 
.A(n_898),
.B(n_895),
.C(n_912),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_900),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_903),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_SL g1057 ( 
.A(n_902),
.B(n_860),
.Y(n_1057)
);

OAI22x1_ASAP7_75t_L g1058 ( 
.A1(n_950),
.A2(n_905),
.B1(n_906),
.B2(n_970),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_903),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_914),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_865),
.B(n_905),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_811),
.A2(n_814),
.B(n_818),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_816),
.B(n_859),
.Y(n_1063)
);

INVx1_ASAP7_75t_SL g1064 ( 
.A(n_865),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_798),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_887),
.B(n_825),
.Y(n_1066)
);

O2A1O1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_933),
.A2(n_934),
.B(n_952),
.C(n_941),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_914),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_878),
.B(n_876),
.Y(n_1069)
);

INVx4_ASAP7_75t_L g1070 ( 
.A(n_921),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_840),
.A2(n_892),
.B(n_886),
.Y(n_1071)
);

NAND2x1p5_ASAP7_75t_L g1072 ( 
.A(n_796),
.B(n_838),
.Y(n_1072)
);

HB1xp67_ASAP7_75t_L g1073 ( 
.A(n_816),
.Y(n_1073)
);

INVxp67_ASAP7_75t_SL g1074 ( 
.A(n_921),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_810),
.B(n_858),
.Y(n_1075)
);

AOI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_915),
.A2(n_858),
.B1(n_911),
.B2(n_930),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_947),
.B(n_879),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_921),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_947),
.B(n_858),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_840),
.A2(n_886),
.B(n_863),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_863),
.A2(n_839),
.B(n_833),
.Y(n_1081)
);

O2A1O1Ixp5_ASAP7_75t_L g1082 ( 
.A1(n_930),
.A2(n_946),
.B(n_965),
.C(n_955),
.Y(n_1082)
);

OAI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_920),
.A2(n_915),
.B1(n_877),
.B2(n_796),
.Y(n_1083)
);

CKINVDCx5p33_ASAP7_75t_R g1084 ( 
.A(n_958),
.Y(n_1084)
);

O2A1O1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_927),
.A2(n_894),
.B(n_904),
.C(n_907),
.Y(n_1085)
);

CKINVDCx20_ASAP7_75t_R g1086 ( 
.A(n_893),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_959),
.Y(n_1087)
);

AOI221xp5_ASAP7_75t_SL g1088 ( 
.A1(n_922),
.A2(n_908),
.B1(n_909),
.B2(n_917),
.C(n_966),
.Y(n_1088)
);

OAI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_915),
.A2(n_838),
.B1(n_954),
.B2(n_943),
.Y(n_1089)
);

NOR3xp33_ASAP7_75t_SL g1090 ( 
.A(n_963),
.B(n_948),
.C(n_961),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_SL g1091 ( 
.A(n_838),
.B(n_921),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_824),
.A2(n_813),
.B(n_852),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_829),
.A2(n_870),
.B(n_891),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_896),
.B(n_821),
.Y(n_1094)
);

O2A1O1Ixp33_ASAP7_75t_SL g1095 ( 
.A1(n_949),
.A2(n_857),
.B(n_856),
.C(n_849),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_827),
.A2(n_931),
.B(n_917),
.C(n_924),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_884),
.A2(n_881),
.B(n_864),
.Y(n_1097)
);

NAND2x1p5_ASAP7_75t_L g1098 ( 
.A(n_967),
.B(n_925),
.Y(n_1098)
);

OR2x2_ASAP7_75t_L g1099 ( 
.A(n_834),
.B(n_850),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_960),
.Y(n_1100)
);

AOI22xp33_ASAP7_75t_L g1101 ( 
.A1(n_964),
.A2(n_972),
.B1(n_971),
.B2(n_968),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_967),
.Y(n_1102)
);

OAI22xp5_ASAP7_75t_L g1103 ( 
.A1(n_925),
.A2(n_944),
.B1(n_855),
.B2(n_843),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_R g1104 ( 
.A(n_919),
.B(n_801),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_944),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_SL g1106 ( 
.A(n_882),
.B(n_885),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_890),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_806),
.Y(n_1108)
);

BUFx6f_ASAP7_75t_L g1109 ( 
.A(n_962),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_813),
.B(n_826),
.Y(n_1110)
);

BUFx12f_ASAP7_75t_L g1111 ( 
.A(n_951),
.Y(n_1111)
);

A2O1A1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_880),
.A2(n_957),
.B(n_956),
.C(n_854),
.Y(n_1112)
);

O2A1O1Ixp5_ASAP7_75t_SL g1113 ( 
.A1(n_861),
.A2(n_866),
.B(n_868),
.C(n_872),
.Y(n_1113)
);

CKINVDCx8_ASAP7_75t_R g1114 ( 
.A(n_875),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_939),
.B(n_802),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_799),
.B(n_802),
.Y(n_1116)
);

BUFx8_ASAP7_75t_L g1117 ( 
.A(n_871),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_793),
.A2(n_723),
.B(n_487),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_799),
.B(n_802),
.Y(n_1119)
);

OR2x2_ASAP7_75t_L g1120 ( 
.A(n_871),
.B(n_700),
.Y(n_1120)
);

OAI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_1116),
.A2(n_1119),
.B1(n_1053),
.B2(n_990),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_1116),
.A2(n_1119),
.B1(n_976),
.B2(n_984),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1115),
.B(n_993),
.Y(n_1123)
);

O2A1O1Ixp5_ASAP7_75t_L g1124 ( 
.A1(n_980),
.A2(n_988),
.B(n_1026),
.C(n_989),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_1041),
.B(n_1040),
.Y(n_1125)
);

O2A1O1Ixp5_ASAP7_75t_L g1126 ( 
.A1(n_1082),
.A2(n_1112),
.B(n_1036),
.C(n_1096),
.Y(n_1126)
);

OAI21xp5_ASAP7_75t_SL g1127 ( 
.A1(n_998),
.A2(n_991),
.B(n_1036),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_977),
.B(n_1120),
.Y(n_1128)
);

BUFx10_ASAP7_75t_L g1129 ( 
.A(n_1094),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1118),
.A2(n_978),
.B(n_1092),
.Y(n_1130)
);

AO31x2_ASAP7_75t_L g1131 ( 
.A1(n_1108),
.A2(n_1103),
.A3(n_1071),
.B(n_994),
.Y(n_1131)
);

OR2x2_ASAP7_75t_L g1132 ( 
.A(n_1010),
.B(n_995),
.Y(n_1132)
);

INVx4_ASAP7_75t_L g1133 ( 
.A(n_982),
.Y(n_1133)
);

AND2x4_ASAP7_75t_L g1134 ( 
.A(n_1063),
.B(n_1050),
.Y(n_1134)
);

INVxp67_ASAP7_75t_L g1135 ( 
.A(n_1031),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_SL g1136 ( 
.A1(n_1029),
.A2(n_1030),
.B(n_1089),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1066),
.A2(n_1069),
.B(n_1062),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_982),
.Y(n_1138)
);

AO21x2_ASAP7_75t_L g1139 ( 
.A1(n_1104),
.A2(n_1110),
.B(n_1028),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1066),
.A2(n_1069),
.B(n_1095),
.Y(n_1140)
);

AO31x2_ASAP7_75t_L g1141 ( 
.A1(n_1103),
.A2(n_994),
.A3(n_1046),
.B(n_1017),
.Y(n_1141)
);

OAI21xp33_ASAP7_75t_L g1142 ( 
.A1(n_1054),
.A2(n_1016),
.B(n_1049),
.Y(n_1142)
);

BUFx3_ASAP7_75t_L g1143 ( 
.A(n_1022),
.Y(n_1143)
);

AO31x2_ASAP7_75t_L g1144 ( 
.A1(n_1081),
.A2(n_1089),
.A3(n_1058),
.B(n_1021),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1037),
.Y(n_1145)
);

OAI21x1_ASAP7_75t_L g1146 ( 
.A1(n_1093),
.A2(n_1097),
.B(n_1002),
.Y(n_1146)
);

AO21x1_ASAP7_75t_L g1147 ( 
.A1(n_1067),
.A2(n_1075),
.B(n_1033),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_1063),
.B(n_1050),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_984),
.B(n_1023),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1015),
.B(n_1044),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_1009),
.A2(n_1005),
.B(n_1113),
.Y(n_1151)
);

INVx2_ASAP7_75t_SL g1152 ( 
.A(n_1117),
.Y(n_1152)
);

OR2x2_ASAP7_75t_L g1153 ( 
.A(n_1064),
.B(n_1007),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1018),
.A2(n_1085),
.B(n_1109),
.Y(n_1154)
);

A2O1A1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_975),
.A2(n_1090),
.B(n_987),
.C(n_1076),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_1034),
.B(n_985),
.Y(n_1156)
);

OAI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_1027),
.A2(n_1006),
.B1(n_996),
.B2(n_979),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1107),
.B(n_1099),
.Y(n_1158)
);

AO31x2_ASAP7_75t_L g1159 ( 
.A1(n_1080),
.A2(n_1001),
.A3(n_1004),
.B(n_1083),
.Y(n_1159)
);

INVx3_ASAP7_75t_L g1160 ( 
.A(n_1072),
.Y(n_1160)
);

INVx3_ASAP7_75t_SL g1161 ( 
.A(n_1013),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1011),
.A2(n_981),
.B(n_1038),
.Y(n_1162)
);

AOI221x1_ASAP7_75t_L g1163 ( 
.A1(n_981),
.A2(n_1083),
.B1(n_1001),
.B2(n_1109),
.C(n_1024),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_1011),
.A2(n_1038),
.B(n_1047),
.Y(n_1164)
);

AOI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_1086),
.A2(n_974),
.B1(n_999),
.B2(n_1057),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1000),
.Y(n_1166)
);

A2O1A1Ixp33_ASAP7_75t_L g1167 ( 
.A1(n_1014),
.A2(n_1088),
.B(n_1043),
.C(n_1039),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1109),
.A2(n_992),
.B(n_1106),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1003),
.Y(n_1169)
);

O2A1O1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_1073),
.A2(n_1042),
.B(n_1061),
.C(n_974),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_SL g1171 ( 
.A1(n_1077),
.A2(n_1079),
.B(n_1087),
.Y(n_1171)
);

INVxp67_ASAP7_75t_SL g1172 ( 
.A(n_1079),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1100),
.B(n_1102),
.Y(n_1173)
);

BUFx6f_ASAP7_75t_L g1174 ( 
.A(n_982),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1091),
.A2(n_1074),
.B(n_996),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_996),
.A2(n_1072),
.B(n_1105),
.Y(n_1176)
);

AO221x2_ASAP7_75t_L g1177 ( 
.A1(n_997),
.A2(n_1059),
.B1(n_986),
.B2(n_1051),
.C(n_1048),
.Y(n_1177)
);

AO21x1_ASAP7_75t_L g1178 ( 
.A1(n_1052),
.A2(n_1055),
.B(n_1098),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_L g1179 ( 
.A1(n_1101),
.A2(n_1098),
.B(n_1068),
.Y(n_1179)
);

AO32x2_ASAP7_75t_L g1180 ( 
.A1(n_983),
.A2(n_1070),
.A3(n_1111),
.B1(n_1114),
.B2(n_1105),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1060),
.A2(n_1056),
.B(n_1045),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1105),
.A2(n_1035),
.B(n_1020),
.Y(n_1182)
);

AND2x6_ASAP7_75t_SL g1183 ( 
.A(n_1117),
.B(n_1084),
.Y(n_1183)
);

AOI22xp33_ASAP7_75t_L g1184 ( 
.A1(n_1065),
.A2(n_1008),
.B1(n_1012),
.B2(n_1019),
.Y(n_1184)
);

O2A1O1Ixp33_ASAP7_75t_SL g1185 ( 
.A1(n_1008),
.A2(n_1012),
.B(n_1019),
.C(n_1032),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1032),
.A2(n_1078),
.B(n_1025),
.Y(n_1186)
);

AOI22xp33_ASAP7_75t_L g1187 ( 
.A1(n_1032),
.A2(n_991),
.B1(n_929),
.B2(n_668),
.Y(n_1187)
);

OR2x2_ASAP7_75t_L g1188 ( 
.A(n_1078),
.B(n_1120),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_SL g1189 ( 
.A(n_1078),
.B(n_1040),
.Y(n_1189)
);

INVx5_ASAP7_75t_L g1190 ( 
.A(n_982),
.Y(n_1190)
);

A2O1A1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_1053),
.A2(n_668),
.B(n_939),
.C(n_799),
.Y(n_1191)
);

BUFx3_ASAP7_75t_L g1192 ( 
.A(n_995),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1037),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_SL g1194 ( 
.A(n_1040),
.B(n_928),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1116),
.B(n_1119),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1118),
.A2(n_793),
.B(n_723),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1118),
.A2(n_793),
.B(n_723),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_1040),
.B(n_928),
.Y(n_1198)
);

AND2x4_ASAP7_75t_L g1199 ( 
.A(n_1063),
.B(n_1050),
.Y(n_1199)
);

AOI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_980),
.A2(n_929),
.B1(n_991),
.B2(n_668),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1037),
.Y(n_1201)
);

NOR3xp33_ASAP7_75t_L g1202 ( 
.A(n_980),
.B(n_668),
.C(n_929),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1118),
.A2(n_793),
.B(n_723),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1093),
.A2(n_1118),
.B(n_1081),
.Y(n_1204)
);

INVx3_ASAP7_75t_L g1205 ( 
.A(n_1072),
.Y(n_1205)
);

OA22x2_ASAP7_75t_L g1206 ( 
.A1(n_1084),
.A2(n_428),
.B1(n_334),
.B2(n_475),
.Y(n_1206)
);

O2A1O1Ixp5_ASAP7_75t_SL g1207 ( 
.A1(n_1036),
.A2(n_932),
.B(n_939),
.C(n_973),
.Y(n_1207)
);

AO32x2_ASAP7_75t_L g1208 ( 
.A1(n_1036),
.A2(n_994),
.A3(n_1089),
.B1(n_1103),
.B2(n_810),
.Y(n_1208)
);

AOI221x1_ASAP7_75t_L g1209 ( 
.A1(n_1053),
.A2(n_1036),
.B1(n_1026),
.B2(n_939),
.C(n_989),
.Y(n_1209)
);

OAI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1053),
.A2(n_799),
.B(n_939),
.Y(n_1210)
);

OR2x2_ASAP7_75t_L g1211 ( 
.A(n_1120),
.B(n_1116),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_L g1212 ( 
.A(n_1040),
.B(n_703),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1093),
.A2(n_1118),
.B(n_1081),
.Y(n_1213)
);

BUFx6f_ASAP7_75t_L g1214 ( 
.A(n_982),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1093),
.A2(n_1118),
.B(n_1081),
.Y(n_1215)
);

OR2x2_ASAP7_75t_L g1216 ( 
.A(n_1120),
.B(n_1116),
.Y(n_1216)
);

OAI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1053),
.A2(n_799),
.B(n_939),
.Y(n_1217)
);

AOI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1092),
.A2(n_1071),
.B(n_1103),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_1013),
.Y(n_1219)
);

OAI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1093),
.A2(n_1118),
.B(n_1081),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1118),
.A2(n_793),
.B(n_723),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_1013),
.Y(n_1222)
);

AOI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_980),
.A2(n_929),
.B1(n_991),
.B2(n_668),
.Y(n_1223)
);

OA21x2_ASAP7_75t_L g1224 ( 
.A1(n_1082),
.A2(n_1092),
.B(n_1026),
.Y(n_1224)
);

BUFx6f_ASAP7_75t_L g1225 ( 
.A(n_982),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1118),
.A2(n_793),
.B(n_723),
.Y(n_1226)
);

BUFx2_ASAP7_75t_L g1227 ( 
.A(n_995),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1093),
.A2(n_1118),
.B(n_1081),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1037),
.Y(n_1229)
);

INVx2_ASAP7_75t_SL g1230 ( 
.A(n_995),
.Y(n_1230)
);

AOI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_980),
.A2(n_929),
.B1(n_991),
.B2(n_668),
.Y(n_1231)
);

CKINVDCx20_ASAP7_75t_R g1232 ( 
.A(n_1025),
.Y(n_1232)
);

INVx1_ASAP7_75t_SL g1233 ( 
.A(n_995),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1118),
.A2(n_793),
.B(n_723),
.Y(n_1234)
);

AO31x2_ASAP7_75t_L g1235 ( 
.A1(n_1053),
.A2(n_1026),
.A3(n_1092),
.B(n_1108),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1037),
.Y(n_1236)
);

OR2x2_ASAP7_75t_L g1237 ( 
.A(n_1120),
.B(n_1116),
.Y(n_1237)
);

O2A1O1Ixp33_ASAP7_75t_SL g1238 ( 
.A1(n_1053),
.A2(n_939),
.B(n_799),
.C(n_1046),
.Y(n_1238)
);

AO31x2_ASAP7_75t_L g1239 ( 
.A1(n_1053),
.A2(n_1026),
.A3(n_1092),
.B(n_1108),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1093),
.A2(n_1118),
.B(n_1081),
.Y(n_1240)
);

OR2x2_ASAP7_75t_L g1241 ( 
.A(n_1120),
.B(n_1116),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1041),
.B(n_631),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1040),
.B(n_928),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1118),
.A2(n_793),
.B(n_723),
.Y(n_1244)
);

BUFx6f_ASAP7_75t_L g1245 ( 
.A(n_982),
.Y(n_1245)
);

A2O1A1Ixp33_ASAP7_75t_L g1246 ( 
.A1(n_1053),
.A2(n_668),
.B(n_939),
.C(n_799),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1041),
.B(n_631),
.Y(n_1247)
);

A2O1A1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_1053),
.A2(n_668),
.B(n_939),
.C(n_799),
.Y(n_1248)
);

OR2x2_ASAP7_75t_L g1249 ( 
.A(n_1120),
.B(n_1116),
.Y(n_1249)
);

O2A1O1Ixp33_ASAP7_75t_SL g1250 ( 
.A1(n_1053),
.A2(n_939),
.B(n_799),
.C(n_1046),
.Y(n_1250)
);

OA21x2_ASAP7_75t_L g1251 ( 
.A1(n_1082),
.A2(n_1092),
.B(n_1026),
.Y(n_1251)
);

BUFx6f_ASAP7_75t_L g1252 ( 
.A(n_982),
.Y(n_1252)
);

AOI22xp5_ASAP7_75t_L g1253 ( 
.A1(n_980),
.A2(n_668),
.B1(n_622),
.B2(n_990),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1037),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1116),
.B(n_1119),
.Y(n_1255)
);

AO31x2_ASAP7_75t_L g1256 ( 
.A1(n_1053),
.A2(n_1026),
.A3(n_1092),
.B(n_1108),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_L g1257 ( 
.A1(n_1093),
.A2(n_1118),
.B(n_1081),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1116),
.B(n_1119),
.Y(n_1258)
);

BUFx2_ASAP7_75t_L g1259 ( 
.A(n_995),
.Y(n_1259)
);

A2O1A1Ixp33_ASAP7_75t_L g1260 ( 
.A1(n_1053),
.A2(n_668),
.B(n_939),
.C(n_799),
.Y(n_1260)
);

OA21x2_ASAP7_75t_L g1261 ( 
.A1(n_1082),
.A2(n_1092),
.B(n_1026),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1037),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1037),
.Y(n_1263)
);

OR2x6_ASAP7_75t_L g1264 ( 
.A(n_995),
.B(n_996),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1118),
.A2(n_793),
.B(n_723),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1093),
.A2(n_1118),
.B(n_1081),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1041),
.B(n_631),
.Y(n_1267)
);

AOI22xp5_ASAP7_75t_SL g1268 ( 
.A1(n_980),
.A2(n_928),
.B1(n_668),
.B2(n_334),
.Y(n_1268)
);

A2O1A1Ixp33_ASAP7_75t_L g1269 ( 
.A1(n_1053),
.A2(n_668),
.B(n_939),
.C(n_799),
.Y(n_1269)
);

BUFx3_ASAP7_75t_L g1270 ( 
.A(n_995),
.Y(n_1270)
);

INVx6_ASAP7_75t_L g1271 ( 
.A(n_1190),
.Y(n_1271)
);

AOI22xp33_ASAP7_75t_L g1272 ( 
.A1(n_1202),
.A2(n_1253),
.B1(n_1200),
.B2(n_1223),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1166),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1200),
.A2(n_1223),
.B1(n_1231),
.B2(n_1121),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1169),
.Y(n_1275)
);

INVxp67_ASAP7_75t_L g1276 ( 
.A(n_1153),
.Y(n_1276)
);

BUFx6f_ASAP7_75t_SL g1277 ( 
.A(n_1192),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1122),
.B(n_1195),
.Y(n_1278)
);

BUFx8_ASAP7_75t_SL g1279 ( 
.A(n_1232),
.Y(n_1279)
);

INVx1_ASAP7_75t_SL g1280 ( 
.A(n_1132),
.Y(n_1280)
);

AOI22xp33_ASAP7_75t_SL g1281 ( 
.A1(n_1268),
.A2(n_1206),
.B1(n_1128),
.B2(n_1212),
.Y(n_1281)
);

BUFx3_ASAP7_75t_L g1282 ( 
.A(n_1270),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1123),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1181),
.Y(n_1284)
);

AOI22xp5_ASAP7_75t_L g1285 ( 
.A1(n_1231),
.A2(n_1127),
.B1(n_1194),
.B2(n_1243),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1255),
.B(n_1258),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1158),
.Y(n_1287)
);

CKINVDCx11_ASAP7_75t_R g1288 ( 
.A(n_1183),
.Y(n_1288)
);

BUFx12f_ASAP7_75t_L g1289 ( 
.A(n_1219),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1177),
.Y(n_1290)
);

INVx2_ASAP7_75t_SL g1291 ( 
.A(n_1227),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1147),
.A2(n_1142),
.B1(n_1210),
.B2(n_1217),
.Y(n_1292)
);

BUFx8_ASAP7_75t_SL g1293 ( 
.A(n_1222),
.Y(n_1293)
);

BUFx10_ASAP7_75t_L g1294 ( 
.A(n_1230),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1125),
.A2(n_1187),
.B1(n_1157),
.B2(n_1247),
.Y(n_1295)
);

INVx5_ASAP7_75t_L g1296 ( 
.A(n_1190),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_SL g1297 ( 
.A1(n_1242),
.A2(n_1267),
.B1(n_1149),
.B2(n_1172),
.Y(n_1297)
);

BUFx12f_ASAP7_75t_L g1298 ( 
.A(n_1129),
.Y(n_1298)
);

INVx6_ASAP7_75t_L g1299 ( 
.A(n_1134),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_SL g1300 ( 
.A1(n_1150),
.A2(n_1173),
.B1(n_1134),
.B2(n_1199),
.Y(n_1300)
);

BUFx6f_ASAP7_75t_SL g1301 ( 
.A(n_1152),
.Y(n_1301)
);

INVx6_ASAP7_75t_L g1302 ( 
.A(n_1148),
.Y(n_1302)
);

BUFx12f_ASAP7_75t_L g1303 ( 
.A(n_1259),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1156),
.B(n_1191),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1177),
.Y(n_1305)
);

INVx1_ASAP7_75t_SL g1306 ( 
.A(n_1233),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1198),
.A2(n_1241),
.B1(n_1216),
.B2(n_1237),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_SL g1308 ( 
.A1(n_1148),
.A2(n_1199),
.B1(n_1211),
.B2(n_1249),
.Y(n_1308)
);

BUFx8_ASAP7_75t_L g1309 ( 
.A(n_1188),
.Y(n_1309)
);

BUFx2_ASAP7_75t_L g1310 ( 
.A(n_1264),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1269),
.A2(n_1248),
.B1(n_1246),
.B2(n_1260),
.Y(n_1311)
);

BUFx3_ASAP7_75t_L g1312 ( 
.A(n_1143),
.Y(n_1312)
);

CKINVDCx20_ASAP7_75t_R g1313 ( 
.A(n_1161),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1171),
.Y(n_1314)
);

INVx8_ASAP7_75t_L g1315 ( 
.A(n_1264),
.Y(n_1315)
);

BUFx2_ASAP7_75t_L g1316 ( 
.A(n_1135),
.Y(n_1316)
);

OAI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1165),
.A2(n_1155),
.B1(n_1201),
.B2(n_1193),
.Y(n_1317)
);

CKINVDCx11_ASAP7_75t_R g1318 ( 
.A(n_1138),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_1165),
.Y(n_1319)
);

BUFx2_ASAP7_75t_SL g1320 ( 
.A(n_1138),
.Y(n_1320)
);

BUFx12f_ASAP7_75t_L g1321 ( 
.A(n_1138),
.Y(n_1321)
);

BUFx2_ASAP7_75t_SL g1322 ( 
.A(n_1174),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_SL g1323 ( 
.A1(n_1136),
.A2(n_1139),
.B1(n_1224),
.B2(n_1261),
.Y(n_1323)
);

OAI22xp5_ASAP7_75t_L g1324 ( 
.A1(n_1145),
.A2(n_1193),
.B1(n_1229),
.B2(n_1236),
.Y(n_1324)
);

BUFx3_ASAP7_75t_L g1325 ( 
.A(n_1174),
.Y(n_1325)
);

INVx4_ASAP7_75t_L g1326 ( 
.A(n_1174),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1196),
.A2(n_1197),
.B(n_1234),
.Y(n_1327)
);

BUFx6f_ASAP7_75t_L g1328 ( 
.A(n_1214),
.Y(n_1328)
);

INVx2_ASAP7_75t_SL g1329 ( 
.A(n_1214),
.Y(n_1329)
);

INVx2_ASAP7_75t_SL g1330 ( 
.A(n_1214),
.Y(n_1330)
);

INVx6_ASAP7_75t_L g1331 ( 
.A(n_1133),
.Y(n_1331)
);

INVx6_ASAP7_75t_L g1332 ( 
.A(n_1133),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1189),
.A2(n_1168),
.B1(n_1154),
.B2(n_1139),
.Y(n_1333)
);

AOI22xp33_ASAP7_75t_L g1334 ( 
.A1(n_1186),
.A2(n_1178),
.B1(n_1201),
.B2(n_1254),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_SL g1335 ( 
.A1(n_1224),
.A2(n_1251),
.B1(n_1261),
.B2(n_1209),
.Y(n_1335)
);

OAI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1163),
.A2(n_1176),
.B1(n_1175),
.B2(n_1262),
.Y(n_1336)
);

BUFx8_ASAP7_75t_SL g1337 ( 
.A(n_1225),
.Y(n_1337)
);

BUFx10_ASAP7_75t_L g1338 ( 
.A(n_1225),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1254),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_SL g1340 ( 
.A1(n_1251),
.A2(n_1205),
.B1(n_1160),
.B2(n_1207),
.Y(n_1340)
);

OR2x6_ASAP7_75t_L g1341 ( 
.A(n_1170),
.B(n_1179),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1263),
.A2(n_1137),
.B1(n_1184),
.B2(n_1205),
.Y(n_1342)
);

INVx1_ASAP7_75t_SL g1343 ( 
.A(n_1225),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1263),
.A2(n_1140),
.B1(n_1162),
.B2(n_1130),
.Y(n_1344)
);

OAI22xp5_ASAP7_75t_L g1345 ( 
.A1(n_1167),
.A2(n_1208),
.B1(n_1238),
.B2(n_1250),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1180),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1180),
.Y(n_1347)
);

INVx4_ASAP7_75t_L g1348 ( 
.A(n_1245),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1203),
.A2(n_1244),
.B1(n_1265),
.B2(n_1226),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1235),
.B(n_1256),
.Y(n_1350)
);

OAI21xp5_ASAP7_75t_SL g1351 ( 
.A1(n_1218),
.A2(n_1221),
.B(n_1124),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1185),
.Y(n_1352)
);

CKINVDCx11_ASAP7_75t_R g1353 ( 
.A(n_1245),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1245),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1182),
.A2(n_1252),
.B1(n_1164),
.B2(n_1266),
.Y(n_1355)
);

INVx1_ASAP7_75t_SL g1356 ( 
.A(n_1252),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1144),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1141),
.B(n_1208),
.Y(n_1358)
);

AND2x4_ASAP7_75t_L g1359 ( 
.A(n_1141),
.B(n_1256),
.Y(n_1359)
);

CKINVDCx6p67_ASAP7_75t_R g1360 ( 
.A(n_1208),
.Y(n_1360)
);

CKINVDCx5p33_ASAP7_75t_R g1361 ( 
.A(n_1126),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1204),
.A2(n_1220),
.B1(n_1240),
.B2(n_1228),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1235),
.B(n_1256),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1141),
.A2(n_1239),
.B1(n_1235),
.B2(n_1131),
.Y(n_1364)
);

BUFx2_ASAP7_75t_L g1365 ( 
.A(n_1239),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_SL g1366 ( 
.A1(n_1151),
.A2(n_1213),
.B1(n_1215),
.B2(n_1257),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1146),
.A2(n_1202),
.B1(n_980),
.B2(n_668),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1159),
.A2(n_1202),
.B1(n_980),
.B2(n_668),
.Y(n_1368)
);

BUFx12f_ASAP7_75t_L g1369 ( 
.A(n_1159),
.Y(n_1369)
);

BUFx3_ASAP7_75t_L g1370 ( 
.A(n_1192),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_1219),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1166),
.Y(n_1372)
);

AOI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1202),
.A2(n_1253),
.B1(n_980),
.B2(n_668),
.Y(n_1373)
);

CKINVDCx20_ASAP7_75t_R g1374 ( 
.A(n_1232),
.Y(n_1374)
);

AOI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1202),
.A2(n_1253),
.B1(n_980),
.B2(n_668),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1253),
.A2(n_1255),
.B1(n_1258),
.B2(n_1195),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_SL g1377 ( 
.A1(n_1268),
.A2(n_434),
.B1(n_443),
.B2(n_928),
.Y(n_1377)
);

BUFx2_ASAP7_75t_L g1378 ( 
.A(n_1192),
.Y(n_1378)
);

BUFx2_ASAP7_75t_L g1379 ( 
.A(n_1192),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1166),
.Y(n_1380)
);

BUFx2_ASAP7_75t_L g1381 ( 
.A(n_1192),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1166),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_1219),
.Y(n_1383)
);

OAI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1253),
.A2(n_1255),
.B1(n_1258),
.B2(n_1195),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_SL g1385 ( 
.A1(n_1268),
.A2(n_980),
.B1(n_928),
.B2(n_434),
.Y(n_1385)
);

BUFx6f_ASAP7_75t_L g1386 ( 
.A(n_1190),
.Y(n_1386)
);

CKINVDCx11_ASAP7_75t_R g1387 ( 
.A(n_1183),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1121),
.B(n_1122),
.Y(n_1388)
);

INVx6_ASAP7_75t_L g1389 ( 
.A(n_1190),
.Y(n_1389)
);

INVx1_ASAP7_75t_SL g1390 ( 
.A(n_1153),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1202),
.A2(n_980),
.B1(n_668),
.B2(n_991),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1202),
.A2(n_980),
.B1(n_668),
.B2(n_991),
.Y(n_1392)
);

INVx6_ASAP7_75t_L g1393 ( 
.A(n_1190),
.Y(n_1393)
);

BUFx2_ASAP7_75t_SL g1394 ( 
.A(n_1192),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1327),
.A2(n_1362),
.B(n_1349),
.Y(n_1395)
);

AND2x4_ASAP7_75t_L g1396 ( 
.A(n_1314),
.B(n_1359),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1360),
.B(n_1358),
.Y(n_1397)
);

AO21x2_ASAP7_75t_L g1398 ( 
.A1(n_1327),
.A2(n_1351),
.B(n_1336),
.Y(n_1398)
);

NOR2xp33_ASAP7_75t_L g1399 ( 
.A(n_1319),
.B(n_1373),
.Y(n_1399)
);

BUFx2_ASAP7_75t_L g1400 ( 
.A(n_1346),
.Y(n_1400)
);

HB1xp67_ASAP7_75t_L g1401 ( 
.A(n_1390),
.Y(n_1401)
);

INVx6_ASAP7_75t_L g1402 ( 
.A(n_1296),
.Y(n_1402)
);

BUFx12f_ASAP7_75t_L g1403 ( 
.A(n_1288),
.Y(n_1403)
);

BUFx6f_ASAP7_75t_L g1404 ( 
.A(n_1369),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1357),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1274),
.B(n_1290),
.Y(n_1406)
);

OAI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1375),
.A2(n_1392),
.B(n_1391),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1278),
.B(n_1376),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1284),
.Y(n_1409)
);

AOI22xp33_ASAP7_75t_SL g1410 ( 
.A1(n_1311),
.A2(n_1388),
.B1(n_1361),
.B2(n_1345),
.Y(n_1410)
);

AO21x2_ASAP7_75t_L g1411 ( 
.A1(n_1350),
.A2(n_1363),
.B(n_1388),
.Y(n_1411)
);

AOI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1377),
.A2(n_1272),
.B1(n_1385),
.B2(n_1285),
.Y(n_1412)
);

INVxp67_ASAP7_75t_L g1413 ( 
.A(n_1316),
.Y(n_1413)
);

INVx2_ASAP7_75t_L g1414 ( 
.A(n_1350),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_1293),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1365),
.Y(n_1416)
);

INVx2_ASAP7_75t_SL g1417 ( 
.A(n_1315),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1344),
.A2(n_1363),
.B(n_1364),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_1279),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1390),
.Y(n_1420)
);

OA21x2_ASAP7_75t_L g1421 ( 
.A1(n_1292),
.A2(n_1368),
.B(n_1333),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1339),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1347),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1364),
.A2(n_1311),
.B(n_1355),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1324),
.Y(n_1425)
);

BUFx2_ASAP7_75t_L g1426 ( 
.A(n_1341),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1324),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1377),
.A2(n_1281),
.B1(n_1308),
.B2(n_1295),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1341),
.Y(n_1429)
);

BUFx2_ASAP7_75t_L g1430 ( 
.A(n_1341),
.Y(n_1430)
);

BUFx3_ASAP7_75t_L g1431 ( 
.A(n_1315),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1278),
.Y(n_1432)
);

HB1xp67_ASAP7_75t_L g1433 ( 
.A(n_1280),
.Y(n_1433)
);

HB1xp67_ASAP7_75t_L g1434 ( 
.A(n_1280),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1304),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1376),
.B(n_1384),
.Y(n_1436)
);

HB1xp67_ASAP7_75t_L g1437 ( 
.A(n_1276),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1304),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1305),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1345),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1323),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1323),
.Y(n_1442)
);

OR2x6_ASAP7_75t_L g1443 ( 
.A(n_1315),
.B(n_1317),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_1371),
.Y(n_1444)
);

INVx2_ASAP7_75t_SL g1445 ( 
.A(n_1271),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1384),
.B(n_1286),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1317),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1335),
.Y(n_1448)
);

INVx4_ASAP7_75t_L g1449 ( 
.A(n_1296),
.Y(n_1449)
);

AOI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1286),
.A2(n_1335),
.B(n_1366),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1273),
.Y(n_1451)
);

BUFx3_ASAP7_75t_L g1452 ( 
.A(n_1309),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1275),
.Y(n_1453)
);

AOI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1352),
.A2(n_1283),
.B(n_1380),
.Y(n_1454)
);

INVxp67_ASAP7_75t_L g1455 ( 
.A(n_1306),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1372),
.Y(n_1456)
);

BUFx2_ASAP7_75t_L g1457 ( 
.A(n_1309),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1382),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1340),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1334),
.Y(n_1460)
);

OAI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1342),
.A2(n_1367),
.B(n_1354),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1297),
.A2(n_1300),
.B1(n_1310),
.B2(n_1307),
.Y(n_1462)
);

OAI21x1_ASAP7_75t_L g1463 ( 
.A1(n_1287),
.A2(n_1297),
.B(n_1296),
.Y(n_1463)
);

OA21x2_ASAP7_75t_L g1464 ( 
.A1(n_1343),
.A2(n_1356),
.B(n_1329),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1389),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_1383),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1393),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1393),
.Y(n_1468)
);

INVx2_ASAP7_75t_SL g1469 ( 
.A(n_1331),
.Y(n_1469)
);

O2A1O1Ixp33_ASAP7_75t_SL g1470 ( 
.A1(n_1343),
.A2(n_1356),
.B(n_1330),
.C(n_1313),
.Y(n_1470)
);

AOI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1306),
.A2(n_1302),
.B1(n_1299),
.B2(n_1291),
.Y(n_1471)
);

OAI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1320),
.A2(n_1322),
.B(n_1338),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1386),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1299),
.B(n_1302),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1397),
.B(n_1381),
.Y(n_1475)
);

INVx2_ASAP7_75t_SL g1476 ( 
.A(n_1452),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1397),
.B(n_1378),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1433),
.B(n_1379),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1434),
.B(n_1401),
.Y(n_1479)
);

OAI21xp5_ASAP7_75t_L g1480 ( 
.A1(n_1407),
.A2(n_1374),
.B(n_1282),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1420),
.B(n_1394),
.Y(n_1481)
);

A2O1A1Ixp33_ASAP7_75t_L g1482 ( 
.A1(n_1412),
.A2(n_1386),
.B(n_1370),
.C(n_1325),
.Y(n_1482)
);

O2A1O1Ixp33_ASAP7_75t_SL g1483 ( 
.A1(n_1412),
.A2(n_1387),
.B(n_1337),
.C(n_1353),
.Y(n_1483)
);

NAND2xp33_ASAP7_75t_SL g1484 ( 
.A(n_1428),
.B(n_1277),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1422),
.Y(n_1485)
);

OR2x2_ASAP7_75t_L g1486 ( 
.A(n_1437),
.B(n_1312),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1446),
.B(n_1299),
.Y(n_1487)
);

NAND2x1_ASAP7_75t_L g1488 ( 
.A(n_1402),
.B(n_1443),
.Y(n_1488)
);

INVx3_ASAP7_75t_L g1489 ( 
.A(n_1464),
.Y(n_1489)
);

A2O1A1Ixp33_ASAP7_75t_L g1490 ( 
.A1(n_1407),
.A2(n_1328),
.B(n_1318),
.C(n_1277),
.Y(n_1490)
);

OAI21xp5_ASAP7_75t_L g1491 ( 
.A1(n_1399),
.A2(n_1326),
.B(n_1348),
.Y(n_1491)
);

HB1xp67_ASAP7_75t_L g1492 ( 
.A(n_1464),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1406),
.B(n_1294),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1405),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1471),
.B(n_1303),
.Y(n_1495)
);

NAND3xp33_ASAP7_75t_L g1496 ( 
.A(n_1410),
.B(n_1348),
.C(n_1298),
.Y(n_1496)
);

AND2x4_ASAP7_75t_L g1497 ( 
.A(n_1396),
.B(n_1321),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_SL g1498 ( 
.A(n_1415),
.B(n_1289),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1446),
.B(n_1331),
.Y(n_1499)
);

OAI22xp5_ASAP7_75t_L g1500 ( 
.A1(n_1462),
.A2(n_1301),
.B1(n_1332),
.B2(n_1436),
.Y(n_1500)
);

AOI211xp5_ASAP7_75t_L g1501 ( 
.A1(n_1436),
.A2(n_1332),
.B(n_1408),
.C(n_1470),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1408),
.B(n_1332),
.Y(n_1502)
);

AOI221xp5_ASAP7_75t_SL g1503 ( 
.A1(n_1439),
.A2(n_1459),
.B1(n_1455),
.B2(n_1447),
.C(n_1450),
.Y(n_1503)
);

A2O1A1Ixp33_ASAP7_75t_L g1504 ( 
.A1(n_1463),
.A2(n_1447),
.B(n_1424),
.C(n_1450),
.Y(n_1504)
);

OA21x2_ASAP7_75t_L g1505 ( 
.A1(n_1418),
.A2(n_1424),
.B(n_1395),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1443),
.A2(n_1413),
.B1(n_1457),
.B2(n_1452),
.Y(n_1506)
);

O2A1O1Ixp33_ASAP7_75t_L g1507 ( 
.A1(n_1460),
.A2(n_1432),
.B(n_1439),
.C(n_1459),
.Y(n_1507)
);

AO21x2_ASAP7_75t_L g1508 ( 
.A1(n_1454),
.A2(n_1395),
.B(n_1398),
.Y(n_1508)
);

AOI21xp5_ASAP7_75t_L g1509 ( 
.A1(n_1398),
.A2(n_1395),
.B(n_1432),
.Y(n_1509)
);

A2O1A1Ixp33_ASAP7_75t_L g1510 ( 
.A1(n_1463),
.A2(n_1424),
.B(n_1460),
.C(n_1418),
.Y(n_1510)
);

INVxp67_ASAP7_75t_L g1511 ( 
.A(n_1464),
.Y(n_1511)
);

AND2x2_ASAP7_75t_SL g1512 ( 
.A(n_1426),
.B(n_1430),
.Y(n_1512)
);

OAI21xp5_ASAP7_75t_L g1513 ( 
.A1(n_1461),
.A2(n_1463),
.B(n_1421),
.Y(n_1513)
);

INVx2_ASAP7_75t_SL g1514 ( 
.A(n_1452),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1456),
.B(n_1458),
.Y(n_1515)
);

AOI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1421),
.A2(n_1457),
.B1(n_1417),
.B2(n_1474),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1409),
.Y(n_1517)
);

OR2x6_ASAP7_75t_L g1518 ( 
.A(n_1426),
.B(n_1430),
.Y(n_1518)
);

OAI211xp5_ASAP7_75t_L g1519 ( 
.A1(n_1421),
.A2(n_1442),
.B(n_1441),
.C(n_1448),
.Y(n_1519)
);

NOR2xp33_ASAP7_75t_L g1520 ( 
.A(n_1435),
.B(n_1438),
.Y(n_1520)
);

BUFx4f_ASAP7_75t_SL g1521 ( 
.A(n_1403),
.Y(n_1521)
);

OA21x2_ASAP7_75t_L g1522 ( 
.A1(n_1418),
.A2(n_1442),
.B(n_1441),
.Y(n_1522)
);

A2O1A1Ixp33_ASAP7_75t_L g1523 ( 
.A1(n_1461),
.A2(n_1440),
.B(n_1427),
.C(n_1425),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1451),
.B(n_1453),
.Y(n_1524)
);

OR2x6_ASAP7_75t_L g1525 ( 
.A(n_1429),
.B(n_1404),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1522),
.B(n_1448),
.Y(n_1526)
);

OR2x2_ASAP7_75t_L g1527 ( 
.A(n_1522),
.B(n_1429),
.Y(n_1527)
);

INVx3_ASAP7_75t_L g1528 ( 
.A(n_1489),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1485),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1520),
.B(n_1411),
.Y(n_1530)
);

AND2x4_ASAP7_75t_L g1531 ( 
.A(n_1517),
.B(n_1429),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1522),
.B(n_1505),
.Y(n_1532)
);

BUFx2_ASAP7_75t_L g1533 ( 
.A(n_1525),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1492),
.B(n_1400),
.Y(n_1534)
);

BUFx2_ASAP7_75t_L g1535 ( 
.A(n_1525),
.Y(n_1535)
);

BUFx2_ASAP7_75t_L g1536 ( 
.A(n_1525),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1520),
.B(n_1411),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1505),
.B(n_1398),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1494),
.Y(n_1539)
);

OR2x2_ASAP7_75t_L g1540 ( 
.A(n_1492),
.B(n_1400),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1505),
.B(n_1398),
.Y(n_1541)
);

INVxp67_ASAP7_75t_SL g1542 ( 
.A(n_1511),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1523),
.B(n_1411),
.Y(n_1543)
);

BUFx2_ASAP7_75t_L g1544 ( 
.A(n_1518),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1523),
.B(n_1425),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1513),
.B(n_1414),
.Y(n_1546)
);

OR2x2_ASAP7_75t_L g1547 ( 
.A(n_1510),
.B(n_1423),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1510),
.B(n_1416),
.Y(n_1548)
);

BUFx3_ASAP7_75t_L g1549 ( 
.A(n_1488),
.Y(n_1549)
);

INVxp67_ASAP7_75t_SL g1550 ( 
.A(n_1507),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1484),
.A2(n_1421),
.B1(n_1403),
.B2(n_1440),
.Y(n_1551)
);

CKINVDCx5p33_ASAP7_75t_R g1552 ( 
.A(n_1521),
.Y(n_1552)
);

AOI22xp33_ASAP7_75t_L g1553 ( 
.A1(n_1484),
.A2(n_1403),
.B1(n_1461),
.B2(n_1431),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1504),
.B(n_1414),
.Y(n_1554)
);

INVxp67_ASAP7_75t_SL g1555 ( 
.A(n_1507),
.Y(n_1555)
);

NOR2x1_ASAP7_75t_L g1556 ( 
.A(n_1549),
.B(n_1519),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1532),
.B(n_1504),
.Y(n_1557)
);

OAI33xp33_ASAP7_75t_L g1558 ( 
.A1(n_1545),
.A2(n_1499),
.A3(n_1500),
.B1(n_1502),
.B2(n_1478),
.B3(n_1487),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1526),
.B(n_1509),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1532),
.B(n_1508),
.Y(n_1560)
);

INVx3_ASAP7_75t_L g1561 ( 
.A(n_1528),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1534),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1530),
.B(n_1524),
.Y(n_1563)
);

OAI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1555),
.A2(n_1482),
.B1(n_1501),
.B2(n_1490),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1532),
.B(n_1516),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1538),
.B(n_1515),
.Y(n_1566)
);

INVxp67_ASAP7_75t_SL g1567 ( 
.A(n_1542),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1527),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1527),
.Y(n_1569)
);

INVx1_ASAP7_75t_SL g1570 ( 
.A(n_1540),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_L g1571 ( 
.A1(n_1551),
.A2(n_1480),
.B1(n_1496),
.B2(n_1521),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1529),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1541),
.B(n_1518),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1528),
.Y(n_1574)
);

BUFx2_ASAP7_75t_L g1575 ( 
.A(n_1542),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1539),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1530),
.B(n_1503),
.Y(n_1577)
);

BUFx3_ASAP7_75t_L g1578 ( 
.A(n_1549),
.Y(n_1578)
);

OAI31xp33_ASAP7_75t_L g1579 ( 
.A1(n_1551),
.A2(n_1482),
.A3(n_1490),
.B(n_1483),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1529),
.Y(n_1580)
);

NOR2x1_ASAP7_75t_SL g1581 ( 
.A(n_1548),
.B(n_1404),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1554),
.B(n_1512),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1537),
.B(n_1479),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1554),
.B(n_1512),
.Y(n_1584)
);

NOR2xp67_ASAP7_75t_L g1585 ( 
.A(n_1557),
.B(n_1526),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1572),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1577),
.B(n_1546),
.Y(n_1587)
);

AND2x4_ASAP7_75t_SL g1588 ( 
.A(n_1582),
.B(n_1404),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1573),
.B(n_1544),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1577),
.B(n_1537),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1573),
.B(n_1544),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1577),
.B(n_1547),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1573),
.B(n_1549),
.Y(n_1593)
);

OR2x2_ASAP7_75t_L g1594 ( 
.A(n_1563),
.B(n_1547),
.Y(n_1594)
);

INVxp67_ASAP7_75t_L g1595 ( 
.A(n_1583),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1578),
.B(n_1533),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1573),
.B(n_1533),
.Y(n_1597)
);

AND2x4_ASAP7_75t_L g1598 ( 
.A(n_1578),
.B(n_1535),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1563),
.B(n_1547),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1582),
.B(n_1535),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1582),
.B(n_1536),
.Y(n_1601)
);

AND2x4_ASAP7_75t_L g1602 ( 
.A(n_1578),
.B(n_1536),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1572),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1582),
.B(n_1546),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1583),
.B(n_1546),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1584),
.B(n_1554),
.Y(n_1606)
);

INVx1_ASAP7_75t_SL g1607 ( 
.A(n_1578),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1584),
.B(n_1531),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1563),
.B(n_1543),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1572),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1580),
.Y(n_1611)
);

NAND2x1_ASAP7_75t_L g1612 ( 
.A(n_1556),
.B(n_1548),
.Y(n_1612)
);

NOR2x1_ASAP7_75t_L g1613 ( 
.A(n_1556),
.B(n_1578),
.Y(n_1613)
);

OR2x2_ASAP7_75t_L g1614 ( 
.A(n_1583),
.B(n_1543),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1580),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1557),
.B(n_1550),
.Y(n_1616)
);

INVx2_ASAP7_75t_SL g1617 ( 
.A(n_1576),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1562),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1584),
.B(n_1531),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1580),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1584),
.B(n_1565),
.Y(n_1621)
);

INVx1_ASAP7_75t_SL g1622 ( 
.A(n_1556),
.Y(n_1622)
);

INVx2_ASAP7_75t_SL g1623 ( 
.A(n_1613),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1586),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1616),
.B(n_1587),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1592),
.B(n_1559),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1586),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1592),
.B(n_1565),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_SL g1629 ( 
.A(n_1613),
.B(n_1579),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1594),
.B(n_1559),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1621),
.B(n_1565),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1618),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1595),
.B(n_1565),
.Y(n_1633)
);

AOI21xp5_ASAP7_75t_L g1634 ( 
.A1(n_1612),
.A2(n_1564),
.B(n_1579),
.Y(n_1634)
);

INVxp67_ASAP7_75t_L g1635 ( 
.A(n_1612),
.Y(n_1635)
);

OR2x2_ASAP7_75t_L g1636 ( 
.A(n_1594),
.B(n_1559),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1603),
.Y(n_1637)
);

INVx1_ASAP7_75t_SL g1638 ( 
.A(n_1622),
.Y(n_1638)
);

BUFx3_ASAP7_75t_L g1639 ( 
.A(n_1588),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1603),
.Y(n_1640)
);

AO21x2_ASAP7_75t_L g1641 ( 
.A1(n_1585),
.A2(n_1557),
.B(n_1560),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1610),
.Y(n_1642)
);

INVx2_ASAP7_75t_SL g1643 ( 
.A(n_1588),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_R g1644 ( 
.A(n_1621),
.B(n_1476),
.Y(n_1644)
);

AND2x4_ASAP7_75t_L g1645 ( 
.A(n_1588),
.B(n_1581),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1599),
.B(n_1559),
.Y(n_1646)
);

INVx2_ASAP7_75t_SL g1647 ( 
.A(n_1596),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1599),
.B(n_1570),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1610),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1617),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1606),
.B(n_1557),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1611),
.Y(n_1652)
);

OR2x2_ASAP7_75t_L g1653 ( 
.A(n_1590),
.B(n_1570),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1590),
.B(n_1550),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1606),
.B(n_1581),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1611),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1604),
.B(n_1593),
.Y(n_1657)
);

INVx2_ASAP7_75t_SL g1658 ( 
.A(n_1596),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1615),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1604),
.B(n_1581),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1617),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1615),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1620),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1593),
.B(n_1566),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1620),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1634),
.B(n_1638),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1627),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1629),
.B(n_1600),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1628),
.B(n_1609),
.Y(n_1669)
);

HB1xp67_ASAP7_75t_L g1670 ( 
.A(n_1632),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1627),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1654),
.B(n_1609),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1625),
.B(n_1600),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1637),
.Y(n_1674)
);

OR2x6_ASAP7_75t_L g1675 ( 
.A(n_1635),
.B(n_1623),
.Y(n_1675)
);

BUFx2_ASAP7_75t_L g1676 ( 
.A(n_1639),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1657),
.B(n_1601),
.Y(n_1677)
);

OAI22xp33_ASAP7_75t_L g1678 ( 
.A1(n_1643),
.A2(n_1564),
.B1(n_1555),
.B2(n_1585),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1657),
.B(n_1596),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1626),
.B(n_1614),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1651),
.B(n_1655),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1641),
.Y(n_1682)
);

AOI22xp33_ASAP7_75t_L g1683 ( 
.A1(n_1639),
.A2(n_1571),
.B1(n_1579),
.B2(n_1558),
.Y(n_1683)
);

OAI211xp5_ASAP7_75t_L g1684 ( 
.A1(n_1623),
.A2(n_1571),
.B(n_1564),
.C(n_1553),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_SL g1685 ( 
.A(n_1643),
.B(n_1558),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1651),
.B(n_1596),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1637),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1640),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1655),
.B(n_1598),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1664),
.B(n_1601),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1626),
.B(n_1614),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1645),
.B(n_1598),
.Y(n_1692)
);

AND4x1_ASAP7_75t_L g1693 ( 
.A(n_1660),
.B(n_1498),
.C(n_1491),
.D(n_1553),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1640),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1645),
.B(n_1598),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1664),
.B(n_1631),
.Y(n_1696)
);

OAI21xp5_ASAP7_75t_L g1697 ( 
.A1(n_1647),
.A2(n_1602),
.B(n_1598),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1645),
.B(n_1602),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1631),
.B(n_1607),
.Y(n_1699)
);

AOI22xp33_ASAP7_75t_L g1700 ( 
.A1(n_1647),
.A2(n_1602),
.B1(n_1589),
.B2(n_1591),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1633),
.B(n_1597),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1668),
.B(n_1648),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1676),
.Y(n_1703)
);

OAI22xp5_ASAP7_75t_L g1704 ( 
.A1(n_1683),
.A2(n_1658),
.B1(n_1660),
.B2(n_1602),
.Y(n_1704)
);

OAI22xp33_ASAP7_75t_SL g1705 ( 
.A1(n_1685),
.A2(n_1658),
.B1(n_1648),
.B2(n_1653),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1667),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1666),
.B(n_1589),
.Y(n_1707)
);

NAND2x1p5_ASAP7_75t_L g1708 ( 
.A(n_1693),
.B(n_1575),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1679),
.B(n_1591),
.Y(n_1709)
);

AOI22xp33_ASAP7_75t_L g1710 ( 
.A1(n_1685),
.A2(n_1641),
.B1(n_1495),
.B2(n_1493),
.Y(n_1710)
);

OAI221xp5_ASAP7_75t_L g1711 ( 
.A1(n_1684),
.A2(n_1646),
.B1(n_1636),
.B2(n_1630),
.C(n_1653),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1670),
.B(n_1641),
.Y(n_1712)
);

AOI211xp5_ASAP7_75t_L g1713 ( 
.A1(n_1678),
.A2(n_1483),
.B(n_1646),
.C(n_1636),
.Y(n_1713)
);

INVx1_ASAP7_75t_SL g1714 ( 
.A(n_1676),
.Y(n_1714)
);

NOR3xp33_ASAP7_75t_SL g1715 ( 
.A(n_1697),
.B(n_1552),
.C(n_1419),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1677),
.B(n_1597),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1667),
.Y(n_1717)
);

AOI221xp5_ASAP7_75t_L g1718 ( 
.A1(n_1700),
.A2(n_1630),
.B1(n_1560),
.B2(n_1662),
.C(n_1663),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1671),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1679),
.B(n_1650),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1693),
.B(n_1444),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1671),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1674),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1686),
.B(n_1605),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1674),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1687),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1687),
.Y(n_1727)
);

OAI221xp5_ASAP7_75t_L g1728 ( 
.A1(n_1710),
.A2(n_1708),
.B1(n_1713),
.B2(n_1705),
.C(n_1704),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_SL g1729 ( 
.A(n_1714),
.B(n_1466),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1703),
.B(n_1673),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1703),
.Y(n_1731)
);

OAI221xp5_ASAP7_75t_L g1732 ( 
.A1(n_1710),
.A2(n_1708),
.B1(n_1718),
.B2(n_1715),
.C(n_1721),
.Y(n_1732)
);

OAI221xp5_ASAP7_75t_L g1733 ( 
.A1(n_1715),
.A2(n_1699),
.B1(n_1701),
.B2(n_1675),
.C(n_1672),
.Y(n_1733)
);

AOI221xp5_ASAP7_75t_L g1734 ( 
.A1(n_1711),
.A2(n_1682),
.B1(n_1694),
.B2(n_1688),
.C(n_1696),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1709),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1707),
.B(n_1681),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1702),
.B(n_1688),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1720),
.B(n_1692),
.Y(n_1738)
);

XOR2x2_ASAP7_75t_L g1739 ( 
.A(n_1721),
.B(n_1690),
.Y(n_1739)
);

O2A1O1Ixp5_ASAP7_75t_L g1740 ( 
.A1(n_1712),
.A2(n_1682),
.B(n_1695),
.C(n_1698),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1716),
.B(n_1672),
.Y(n_1741)
);

INVx2_ASAP7_75t_L g1742 ( 
.A(n_1720),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1724),
.B(n_1692),
.Y(n_1743)
);

OAI21xp33_ASAP7_75t_L g1744 ( 
.A1(n_1706),
.A2(n_1686),
.B(n_1695),
.Y(n_1744)
);

OAI22xp33_ASAP7_75t_L g1745 ( 
.A1(n_1717),
.A2(n_1675),
.B1(n_1682),
.B2(n_1669),
.Y(n_1745)
);

INVxp67_ASAP7_75t_L g1746 ( 
.A(n_1719),
.Y(n_1746)
);

NOR2xp33_ASAP7_75t_L g1747 ( 
.A(n_1729),
.B(n_1698),
.Y(n_1747)
);

XOR2x2_ASAP7_75t_L g1748 ( 
.A(n_1739),
.B(n_1514),
.Y(n_1748)
);

HB1xp67_ASAP7_75t_L g1749 ( 
.A(n_1738),
.Y(n_1749)
);

NOR3xp33_ASAP7_75t_L g1750 ( 
.A(n_1728),
.B(n_1723),
.C(n_1722),
.Y(n_1750)
);

XNOR2xp5_ASAP7_75t_L g1751 ( 
.A(n_1733),
.B(n_1506),
.Y(n_1751)
);

AOI221xp5_ASAP7_75t_L g1752 ( 
.A1(n_1734),
.A2(n_1727),
.B1(n_1726),
.B2(n_1725),
.C(n_1694),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1742),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1731),
.Y(n_1754)
);

AOI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1729),
.A2(n_1675),
.B1(n_1689),
.B2(n_1681),
.Y(n_1755)
);

OAI21xp33_ASAP7_75t_SL g1756 ( 
.A1(n_1732),
.A2(n_1675),
.B(n_1689),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1735),
.B(n_1675),
.Y(n_1757)
);

INVx1_ASAP7_75t_SL g1758 ( 
.A(n_1730),
.Y(n_1758)
);

AOI221xp5_ASAP7_75t_L g1759 ( 
.A1(n_1750),
.A2(n_1745),
.B1(n_1740),
.B2(n_1744),
.C(n_1730),
.Y(n_1759)
);

OAI31xp33_ASAP7_75t_L g1760 ( 
.A1(n_1758),
.A2(n_1746),
.A3(n_1737),
.B(n_1741),
.Y(n_1760)
);

INVx2_ASAP7_75t_SL g1761 ( 
.A(n_1749),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1747),
.B(n_1743),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1754),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1753),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_SL g1765 ( 
.A(n_1755),
.B(n_1736),
.Y(n_1765)
);

AOI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1756),
.A2(n_1737),
.B1(n_1669),
.B2(n_1680),
.Y(n_1766)
);

OR2x2_ASAP7_75t_L g1767 ( 
.A(n_1758),
.B(n_1680),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1757),
.Y(n_1768)
);

OAI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1751),
.A2(n_1691),
.B1(n_1650),
.B2(n_1661),
.Y(n_1769)
);

AOI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1759),
.A2(n_1748),
.B1(n_1752),
.B2(n_1691),
.Y(n_1770)
);

OAI21xp5_ASAP7_75t_SL g1771 ( 
.A1(n_1760),
.A2(n_1481),
.B(n_1486),
.Y(n_1771)
);

AOI221xp5_ASAP7_75t_L g1772 ( 
.A1(n_1760),
.A2(n_1567),
.B1(n_1575),
.B2(n_1665),
.C(n_1659),
.Y(n_1772)
);

NAND4xp75_ASAP7_75t_L g1773 ( 
.A(n_1761),
.B(n_1661),
.C(n_1642),
.D(n_1665),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1767),
.Y(n_1774)
);

AO221x1_ASAP7_75t_L g1775 ( 
.A1(n_1774),
.A2(n_1769),
.B1(n_1764),
.B2(n_1768),
.C(n_1763),
.Y(n_1775)
);

XOR2x2_ASAP7_75t_L g1776 ( 
.A(n_1770),
.B(n_1765),
.Y(n_1776)
);

AOI222xp33_ASAP7_75t_L g1777 ( 
.A1(n_1772),
.A2(n_1771),
.B1(n_1762),
.B2(n_1766),
.C1(n_1773),
.C2(n_1567),
.Y(n_1777)
);

AOI22xp5_ASAP7_75t_L g1778 ( 
.A1(n_1770),
.A2(n_1659),
.B1(n_1642),
.B2(n_1652),
.Y(n_1778)
);

AOI22xp33_ASAP7_75t_L g1779 ( 
.A1(n_1770),
.A2(n_1404),
.B1(n_1649),
.B2(n_1624),
.Y(n_1779)
);

A2O1A1Ixp33_ASAP7_75t_L g1780 ( 
.A1(n_1770),
.A2(n_1575),
.B(n_1656),
.C(n_1560),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1775),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1777),
.B(n_1776),
.Y(n_1782)
);

AOI211x1_ASAP7_75t_L g1783 ( 
.A1(n_1780),
.A2(n_1644),
.B(n_1560),
.C(n_1619),
.Y(n_1783)
);

NAND4xp75_ASAP7_75t_L g1784 ( 
.A(n_1778),
.B(n_1417),
.C(n_1469),
.D(n_1445),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1779),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1785),
.Y(n_1786)
);

AOI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1781),
.A2(n_1570),
.B1(n_1477),
.B2(n_1475),
.Y(n_1787)
);

OAI21xp5_ASAP7_75t_L g1788 ( 
.A1(n_1782),
.A2(n_1784),
.B(n_1783),
.Y(n_1788)
);

XNOR2x1_ASAP7_75t_L g1789 ( 
.A(n_1786),
.B(n_1497),
.Y(n_1789)
);

OAI22x1_ASAP7_75t_L g1790 ( 
.A1(n_1789),
.A2(n_1787),
.B1(n_1788),
.B2(n_1644),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1790),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1790),
.B(n_1608),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1792),
.Y(n_1793)
);

OAI22xp5_ASAP7_75t_SL g1794 ( 
.A1(n_1791),
.A2(n_1469),
.B1(n_1445),
.B2(n_1402),
.Y(n_1794)
);

OAI21xp5_ASAP7_75t_L g1795 ( 
.A1(n_1793),
.A2(n_1619),
.B(n_1608),
.Y(n_1795)
);

AOI21xp5_ASAP7_75t_L g1796 ( 
.A1(n_1794),
.A2(n_1569),
.B(n_1568),
.Y(n_1796)
);

OAI22xp5_ASAP7_75t_L g1797 ( 
.A1(n_1795),
.A2(n_1796),
.B1(n_1569),
.B2(n_1568),
.Y(n_1797)
);

AOI22x1_ASAP7_75t_L g1798 ( 
.A1(n_1797),
.A2(n_1449),
.B1(n_1473),
.B2(n_1468),
.Y(n_1798)
);

AOI21xp33_ASAP7_75t_L g1799 ( 
.A1(n_1798),
.A2(n_1569),
.B(n_1473),
.Y(n_1799)
);

AOI221xp5_ASAP7_75t_L g1800 ( 
.A1(n_1799),
.A2(n_1569),
.B1(n_1568),
.B2(n_1574),
.C(n_1561),
.Y(n_1800)
);

AOI211xp5_ASAP7_75t_L g1801 ( 
.A1(n_1800),
.A2(n_1472),
.B(n_1465),
.C(n_1467),
.Y(n_1801)
);


endmodule