module fake_ariane_1215_n_1860 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_172, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1860);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1860;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1733;
wire n_1524;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1288;
wire n_1201;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_236;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_76),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_4),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_136),
.Y(n_176)
);

BUFx8_ASAP7_75t_SL g177 ( 
.A(n_150),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_37),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_29),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_156),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_134),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_92),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_71),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_19),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_119),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_51),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_145),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_51),
.Y(n_188)
);

BUFx10_ASAP7_75t_L g189 ( 
.A(n_37),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_30),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_101),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_59),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_155),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_130),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_53),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_62),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_131),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_4),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_110),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_157),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_151),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_87),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_52),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_91),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_33),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_100),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_173),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_154),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_138),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_75),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_106),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_153),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_54),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_94),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_49),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_3),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_103),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_126),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_27),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_109),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_171),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_116),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_133),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_141),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_28),
.Y(n_225)
);

BUFx5_ASAP7_75t_L g226 ( 
.A(n_148),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_66),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_44),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_123),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_26),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_45),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_97),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_108),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_69),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_16),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_61),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_16),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_172),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_58),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_83),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_58),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_86),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_28),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_90),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_120),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_79),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_144),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_78),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_0),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_98),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_36),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_52),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_46),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_73),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_49),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_38),
.Y(n_256)
);

INVxp67_ASAP7_75t_SL g257 ( 
.A(n_56),
.Y(n_257)
);

BUFx10_ASAP7_75t_L g258 ( 
.A(n_43),
.Y(n_258)
);

INVxp67_ASAP7_75t_SL g259 ( 
.A(n_36),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_128),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_127),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_146),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_95),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_12),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_20),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_121),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_46),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_124),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_20),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_113),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_139),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_125),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_166),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_158),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_54),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_118),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_99),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_143),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_59),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_104),
.Y(n_280)
);

BUFx10_ASAP7_75t_L g281 ( 
.A(n_149),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_0),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_132),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_163),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_22),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_105),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_140),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_25),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_30),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_167),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_169),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_70),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_129),
.Y(n_293)
);

CKINVDCx12_ASAP7_75t_R g294 ( 
.A(n_25),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_42),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_74),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_89),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_10),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_26),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_96),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_65),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_102),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_43),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_39),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_88),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_39),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_115),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_5),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_47),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_1),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_63),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_112),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_107),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_67),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_40),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_29),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_53),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_165),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_3),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_147),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_23),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_80),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_84),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_164),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_31),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_18),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_81),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_33),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_10),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_57),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_45),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_18),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_85),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_27),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_122),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_19),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_22),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_56),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_34),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_23),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_82),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_160),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_31),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_177),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_216),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_319),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_302),
.B(n_1),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_178),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_267),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_178),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_210),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_178),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_316),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_246),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_178),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_312),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_219),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_225),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_178),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_192),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_319),
.B(n_2),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_230),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_192),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_207),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_241),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_207),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_215),
.Y(n_367)
);

INVxp67_ASAP7_75t_SL g368 ( 
.A(n_190),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_228),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_243),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_220),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_265),
.Y(n_372)
);

INVxp67_ASAP7_75t_SL g373 ( 
.A(n_195),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_189),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_176),
.B(n_2),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_220),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_221),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_249),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_221),
.Y(n_379)
);

INVxp33_ASAP7_75t_SL g380 ( 
.A(n_175),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_251),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_270),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_270),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_253),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_183),
.B(n_5),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_300),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_189),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_300),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_198),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_291),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_231),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_237),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_264),
.Y(n_393)
);

INVxp67_ASAP7_75t_SL g394 ( 
.A(n_239),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_235),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_269),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_252),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_279),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_255),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_275),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_288),
.Y(n_401)
);

INVxp67_ASAP7_75t_SL g402 ( 
.A(n_304),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_315),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_282),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_232),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_317),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_256),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_285),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_321),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_185),
.B(n_6),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_289),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_193),
.B(n_6),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_329),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_197),
.B(n_7),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_331),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_337),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_295),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_298),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_200),
.B(n_7),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_340),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_201),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_206),
.B(n_8),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_299),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_294),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_175),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_208),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_309),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_211),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_303),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_421),
.B(n_281),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g431 ( 
.A(n_421),
.B(n_281),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_348),
.Y(n_432)
);

HB1xp67_ASAP7_75t_L g433 ( 
.A(n_372),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_348),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_426),
.B(n_222),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_350),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_350),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_352),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_352),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_355),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_355),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_359),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_426),
.B(n_224),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_359),
.Y(n_444)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_364),
.Y(n_445)
);

AND3x2_ASAP7_75t_L g446 ( 
.A(n_374),
.B(n_259),
.C(n_257),
.Y(n_446)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_428),
.B(n_281),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_345),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_364),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_366),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_366),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_371),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_371),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_376),
.Y(n_454)
);

BUFx6f_ASAP7_75t_L g455 ( 
.A(n_376),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_428),
.B(n_377),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_377),
.B(n_227),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_379),
.Y(n_458)
);

AND2x4_ASAP7_75t_L g459 ( 
.A(n_379),
.B(n_191),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_382),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_382),
.Y(n_461)
);

INVxp33_ASAP7_75t_SL g462 ( 
.A(n_344),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_346),
.B(n_273),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_383),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_383),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_386),
.Y(n_466)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_367),
.A2(n_328),
.B1(n_188),
.B2(n_339),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_386),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_347),
.B(n_191),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_388),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_388),
.B(n_233),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_360),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_360),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_363),
.Y(n_474)
);

INVx5_ASAP7_75t_L g475 ( 
.A(n_405),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_363),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_375),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_410),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_389),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g480 ( 
.A(n_368),
.B(n_273),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_389),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_391),
.Y(n_482)
);

AND2x4_ASAP7_75t_L g483 ( 
.A(n_373),
.B(n_296),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_391),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_354),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_392),
.Y(n_486)
);

AND2x4_ASAP7_75t_L g487 ( 
.A(n_394),
.B(n_296),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_392),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_402),
.B(n_234),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_399),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_399),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_400),
.Y(n_492)
);

INVx3_ASAP7_75t_L g493 ( 
.A(n_400),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_401),
.B(n_189),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_401),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_403),
.Y(n_496)
);

INVx3_ASAP7_75t_L g497 ( 
.A(n_403),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_406),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_406),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_409),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_409),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_413),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_413),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_415),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_415),
.B(n_258),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_416),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_430),
.B(n_431),
.Y(n_507)
);

BUFx3_ASAP7_75t_L g508 ( 
.A(n_458),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_432),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_467),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_475),
.B(n_390),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_475),
.B(n_357),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_445),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_437),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_430),
.B(n_416),
.Y(n_515)
);

INVx6_ASAP7_75t_L g516 ( 
.A(n_475),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_445),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_432),
.Y(n_518)
);

INVxp33_ASAP7_75t_L g519 ( 
.A(n_433),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_430),
.B(n_405),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_432),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_434),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_445),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_475),
.B(n_358),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_475),
.B(n_362),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_437),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_437),
.Y(n_527)
);

INVxp67_ASAP7_75t_SL g528 ( 
.A(n_456),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_445),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_434),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_434),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_438),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_438),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_437),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_431),
.A2(n_380),
.B1(n_365),
.B2(n_396),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_L g536 ( 
.A1(n_469),
.A2(n_414),
.B1(n_412),
.B2(n_385),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_437),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_438),
.Y(n_538)
);

BUFx2_ASAP7_75t_L g539 ( 
.A(n_433),
.Y(n_539)
);

AND2x6_ASAP7_75t_L g540 ( 
.A(n_431),
.B(n_261),
.Y(n_540)
);

NAND3xp33_ASAP7_75t_L g541 ( 
.A(n_469),
.B(n_378),
.C(n_370),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_475),
.B(n_381),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_439),
.Y(n_543)
);

BUFx3_ASAP7_75t_L g544 ( 
.A(n_458),
.Y(n_544)
);

NOR2x1p5_ASAP7_75t_L g545 ( 
.A(n_494),
.B(n_349),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_447),
.B(n_384),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_SL g547 ( 
.A(n_462),
.B(n_353),
.Y(n_547)
);

AND3x2_ASAP7_75t_L g548 ( 
.A(n_448),
.B(n_387),
.C(n_424),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_447),
.B(n_393),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_439),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_445),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_439),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_445),
.Y(n_553)
);

AND2x2_ASAP7_75t_SL g554 ( 
.A(n_447),
.B(n_419),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_440),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_467),
.Y(n_556)
);

NAND2xp33_ASAP7_75t_SL g557 ( 
.A(n_494),
.B(n_398),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_475),
.B(n_404),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_478),
.B(n_408),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_440),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_458),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_494),
.A2(n_429),
.B1(n_411),
.B2(n_423),
.Y(n_562)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_485),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_440),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_478),
.B(n_417),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_505),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_478),
.B(n_418),
.Y(n_567)
);

INVxp67_ASAP7_75t_SL g568 ( 
.A(n_456),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_475),
.B(n_425),
.Y(n_569)
);

AND3x2_ASAP7_75t_L g570 ( 
.A(n_448),
.B(n_361),
.C(n_422),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_444),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_L g572 ( 
.A1(n_480),
.A2(n_487),
.B1(n_483),
.B2(n_505),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_441),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_444),
.Y(n_574)
);

AND3x1_ASAP7_75t_L g575 ( 
.A(n_505),
.B(n_484),
.C(n_479),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_445),
.Y(n_576)
);

INVx2_ASAP7_75t_SL g577 ( 
.A(n_463),
.Y(n_577)
);

BUFx3_ASAP7_75t_L g578 ( 
.A(n_458),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_499),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_441),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_480),
.B(n_483),
.Y(n_581)
);

INVx4_ASAP7_75t_L g582 ( 
.A(n_477),
.Y(n_582)
);

AND2x2_ASAP7_75t_SL g583 ( 
.A(n_477),
.B(n_242),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_444),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_477),
.B(n_420),
.Y(n_585)
);

INVxp67_ASAP7_75t_L g586 ( 
.A(n_485),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_445),
.Y(n_587)
);

BUFx10_ASAP7_75t_L g588 ( 
.A(n_480),
.Y(n_588)
);

AND2x6_ASAP7_75t_L g589 ( 
.A(n_477),
.B(n_261),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_445),
.Y(n_590)
);

AND2x6_ASAP7_75t_L g591 ( 
.A(n_477),
.B(n_261),
.Y(n_591)
);

INVx1_ASAP7_75t_SL g592 ( 
.A(n_463),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_477),
.B(n_420),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_L g594 ( 
.A1(n_477),
.A2(n_306),
.B1(n_203),
.B2(n_213),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_444),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_480),
.B(n_483),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_441),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_442),
.Y(n_598)
);

INVxp33_ASAP7_75t_L g599 ( 
.A(n_463),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_480),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_477),
.B(n_351),
.Y(n_601)
);

OR2x6_ASAP7_75t_L g602 ( 
.A(n_480),
.B(n_244),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_444),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_442),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_444),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_450),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_450),
.Y(n_607)
);

BUFx10_ASAP7_75t_L g608 ( 
.A(n_483),
.Y(n_608)
);

INVx4_ASAP7_75t_L g609 ( 
.A(n_481),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_483),
.B(n_174),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g611 ( 
.A1(n_483),
.A2(n_258),
.B1(n_278),
.B2(n_250),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_487),
.B(n_174),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_487),
.B(n_266),
.Y(n_613)
);

AOI22xp5_ASAP7_75t_L g614 ( 
.A1(n_487),
.A2(n_343),
.B1(n_186),
.B2(n_184),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_442),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_450),
.Y(n_616)
);

INVx4_ASAP7_75t_L g617 ( 
.A(n_481),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_L g618 ( 
.A1(n_489),
.A2(n_179),
.B1(n_188),
.B2(n_203),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_449),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_449),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_487),
.B(n_274),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_487),
.B(n_180),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_450),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_449),
.Y(n_624)
);

BUFx4f_ASAP7_75t_L g625 ( 
.A(n_476),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_449),
.Y(n_626)
);

INVx4_ASAP7_75t_L g627 ( 
.A(n_481),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_499),
.B(n_180),
.Y(n_628)
);

AOI22xp33_ASAP7_75t_L g629 ( 
.A1(n_499),
.A2(n_501),
.B1(n_459),
.B2(n_472),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_449),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_449),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_453),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_499),
.B(n_181),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_450),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_450),
.Y(n_635)
);

AND3x1_ASAP7_75t_L g636 ( 
.A(n_506),
.B(n_258),
.C(n_205),
.Y(n_636)
);

INVx4_ASAP7_75t_L g637 ( 
.A(n_481),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_453),
.Y(n_638)
);

BUFx10_ASAP7_75t_L g639 ( 
.A(n_446),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_501),
.B(n_356),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_450),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_453),
.Y(n_642)
);

INVx3_ASAP7_75t_L g643 ( 
.A(n_450),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g644 ( 
.A(n_501),
.Y(n_644)
);

BUFx2_ASAP7_75t_L g645 ( 
.A(n_446),
.Y(n_645)
);

INVx5_ASAP7_75t_L g646 ( 
.A(n_436),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_450),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_501),
.B(n_181),
.Y(n_648)
);

OR2x6_ASAP7_75t_L g649 ( 
.A(n_435),
.B(n_247),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_462),
.B(n_182),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_481),
.B(n_182),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g652 ( 
.A(n_481),
.B(n_248),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_451),
.Y(n_653)
);

BUFx3_ASAP7_75t_L g654 ( 
.A(n_482),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_588),
.Y(n_655)
);

OAI221xp5_ASAP7_75t_L g656 ( 
.A1(n_536),
.A2(n_443),
.B1(n_435),
.B2(n_310),
.C(n_325),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_619),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_588),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_528),
.B(n_482),
.Y(n_659)
);

INVx2_ASAP7_75t_SL g660 ( 
.A(n_639),
.Y(n_660)
);

AND2x4_ASAP7_75t_L g661 ( 
.A(n_566),
.B(n_479),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_619),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_514),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_620),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_568),
.B(n_482),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_620),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_559),
.B(n_482),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_599),
.B(n_482),
.Y(n_668)
);

O2A1O1Ixp33_ASAP7_75t_L g669 ( 
.A1(n_507),
.A2(n_482),
.B(n_486),
.C(n_493),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_639),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_577),
.B(n_486),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_546),
.B(n_486),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_588),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_592),
.B(n_479),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_563),
.Y(n_675)
);

O2A1O1Ixp33_ASAP7_75t_L g676 ( 
.A1(n_566),
.A2(n_486),
.B(n_493),
.C(n_495),
.Y(n_676)
);

OR2x2_ASAP7_75t_L g677 ( 
.A(n_539),
.B(n_519),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_577),
.B(n_486),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_554),
.B(n_486),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_554),
.B(n_493),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_608),
.B(n_493),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_549),
.B(n_493),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_583),
.A2(n_488),
.B1(n_504),
.B2(n_498),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_624),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_572),
.B(n_493),
.Y(n_685)
);

NAND3xp33_ASAP7_75t_L g686 ( 
.A(n_565),
.B(n_443),
.C(n_484),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_515),
.B(n_495),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_515),
.B(n_600),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_624),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_626),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_539),
.B(n_484),
.Y(n_691)
);

OAI22xp5_ASAP7_75t_L g692 ( 
.A1(n_583),
.A2(n_575),
.B1(n_600),
.B2(n_567),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_626),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_585),
.B(n_495),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_608),
.B(n_495),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_630),
.Y(n_696)
);

OAI22xp5_ASAP7_75t_L g697 ( 
.A1(n_602),
.A2(n_495),
.B1(n_497),
.B2(n_506),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_630),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_540),
.B(n_495),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_631),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_608),
.B(n_497),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_631),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_540),
.B(n_497),
.Y(n_703)
);

AOI22xp5_ASAP7_75t_L g704 ( 
.A1(n_540),
.A2(n_459),
.B1(n_492),
.B2(n_503),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_609),
.B(n_497),
.Y(n_705)
);

NOR3xp33_ASAP7_75t_L g706 ( 
.A(n_586),
.B(n_497),
.C(n_205),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_639),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_526),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_632),
.Y(n_709)
);

AND2x4_ASAP7_75t_L g710 ( 
.A(n_545),
.B(n_490),
.Y(n_710)
);

AOI22xp33_ASAP7_75t_L g711 ( 
.A1(n_649),
.A2(n_498),
.B1(n_504),
.B2(n_488),
.Y(n_711)
);

OR2x2_ASAP7_75t_L g712 ( 
.A(n_520),
.B(n_490),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_632),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_609),
.B(n_490),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_527),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_638),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_540),
.B(n_491),
.Y(n_717)
);

A2O1A1Ixp33_ASAP7_75t_L g718 ( 
.A1(n_581),
.A2(n_468),
.B(n_465),
.C(n_453),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_645),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_540),
.A2(n_459),
.B1(n_496),
.B2(n_503),
.Y(n_720)
);

AOI22xp5_ASAP7_75t_L g721 ( 
.A1(n_649),
.A2(n_459),
.B1(n_496),
.B2(n_503),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_596),
.B(n_491),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_613),
.B(n_491),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_621),
.B(n_492),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_609),
.B(n_492),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_649),
.B(n_496),
.Y(n_726)
);

NAND2xp33_ASAP7_75t_L g727 ( 
.A(n_523),
.B(n_553),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_527),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_523),
.Y(n_729)
);

NAND2xp33_ASAP7_75t_L g730 ( 
.A(n_523),
.B(n_500),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_649),
.B(n_500),
.Y(n_731)
);

CKINVDCx14_ASAP7_75t_R g732 ( 
.A(n_557),
.Y(n_732)
);

CKINVDCx11_ASAP7_75t_R g733 ( 
.A(n_510),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_617),
.B(n_500),
.Y(n_734)
);

INVx2_ASAP7_75t_SL g735 ( 
.A(n_645),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_629),
.B(n_502),
.Y(n_736)
);

BUFx6f_ASAP7_75t_L g737 ( 
.A(n_523),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_617),
.B(n_502),
.Y(n_738)
);

INVxp67_ASAP7_75t_L g739 ( 
.A(n_640),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_601),
.B(n_502),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_541),
.B(n_506),
.Y(n_741)
);

INVx4_ASAP7_75t_L g742 ( 
.A(n_579),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_617),
.B(n_459),
.Y(n_743)
);

AND2x4_ASAP7_75t_L g744 ( 
.A(n_602),
.B(n_459),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_562),
.B(n_535),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_627),
.B(n_453),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_534),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_627),
.B(n_453),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_610),
.B(n_612),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_627),
.B(n_465),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_637),
.B(n_465),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_L g752 ( 
.A(n_622),
.B(n_465),
.Y(n_752)
);

BUFx6f_ASAP7_75t_SL g753 ( 
.A(n_602),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_534),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_637),
.B(n_465),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_509),
.Y(n_756)
);

OAI22xp33_ASAP7_75t_L g757 ( 
.A1(n_602),
.A2(n_614),
.B1(n_618),
.B2(n_556),
.Y(n_757)
);

INVxp67_ASAP7_75t_L g758 ( 
.A(n_547),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_537),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_637),
.B(n_465),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_571),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_582),
.B(n_468),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_593),
.B(n_468),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_582),
.B(n_468),
.Y(n_764)
);

AOI22xp5_ASAP7_75t_L g765 ( 
.A1(n_557),
.A2(n_504),
.B1(n_498),
.B2(n_488),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_571),
.Y(n_766)
);

AO22x2_ASAP7_75t_L g767 ( 
.A1(n_510),
.A2(n_460),
.B1(n_472),
.B2(n_473),
.Y(n_767)
);

AO22x2_ASAP7_75t_L g768 ( 
.A1(n_556),
.A2(n_460),
.B1(n_472),
.B2(n_473),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_638),
.Y(n_769)
);

OR2x2_ASAP7_75t_L g770 ( 
.A(n_594),
.B(n_488),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_512),
.A2(n_504),
.B(n_498),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_642),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_518),
.Y(n_773)
);

BUFx3_ASAP7_75t_L g774 ( 
.A(n_508),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_518),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_574),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_582),
.B(n_654),
.Y(n_777)
);

BUFx8_ASAP7_75t_L g778 ( 
.A(n_548),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_642),
.B(n_468),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_521),
.Y(n_780)
);

OR2x2_ASAP7_75t_L g781 ( 
.A(n_650),
.B(n_457),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_654),
.B(n_460),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_521),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_SL g784 ( 
.A(n_523),
.B(n_451),
.Y(n_784)
);

BUFx5_ASAP7_75t_L g785 ( 
.A(n_589),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_611),
.B(n_369),
.Y(n_786)
);

INVx1_ASAP7_75t_SL g787 ( 
.A(n_628),
.Y(n_787)
);

O2A1O1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_522),
.A2(n_473),
.B(n_474),
.C(n_471),
.Y(n_788)
);

INVxp67_ASAP7_75t_L g789 ( 
.A(n_636),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_574),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_584),
.Y(n_791)
);

OR2x2_ASAP7_75t_L g792 ( 
.A(n_633),
.B(n_457),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_553),
.B(n_451),
.Y(n_793)
);

OAI22xp5_ASAP7_75t_L g794 ( 
.A1(n_644),
.A2(n_310),
.B1(n_338),
.B2(n_339),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_584),
.Y(n_795)
);

NOR2xp33_ASAP7_75t_L g796 ( 
.A(n_644),
.B(n_471),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_508),
.B(n_544),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_544),
.B(n_561),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_561),
.B(n_474),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_522),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_530),
.A2(n_454),
.B1(n_464),
.B2(n_466),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_553),
.B(n_451),
.Y(n_802)
);

INVxp67_ASAP7_75t_L g803 ( 
.A(n_652),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_578),
.B(n_454),
.Y(n_804)
);

INVx3_ASAP7_75t_L g805 ( 
.A(n_578),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_553),
.B(n_451),
.Y(n_806)
);

INVx2_ASAP7_75t_SL g807 ( 
.A(n_570),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_595),
.B(n_454),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_530),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_531),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_595),
.B(n_454),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_603),
.B(n_464),
.Y(n_812)
);

OAI22xp5_ASAP7_75t_L g813 ( 
.A1(n_651),
.A2(n_213),
.B1(n_179),
.B2(n_306),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_603),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_587),
.B(n_451),
.Y(n_815)
);

O2A1O1Ixp33_ASAP7_75t_L g816 ( 
.A1(n_656),
.A2(n_648),
.B(n_564),
.C(n_598),
.Y(n_816)
);

OAI21xp33_ASAP7_75t_L g817 ( 
.A1(n_803),
.A2(n_325),
.B(n_308),
.Y(n_817)
);

O2A1O1Ixp33_ASAP7_75t_L g818 ( 
.A1(n_679),
.A2(n_604),
.B(n_555),
.C(n_560),
.Y(n_818)
);

OAI22xp5_ASAP7_75t_L g819 ( 
.A1(n_680),
.A2(n_538),
.B1(n_564),
.B2(n_573),
.Y(n_819)
);

NAND2xp33_ASAP7_75t_L g820 ( 
.A(n_655),
.B(n_587),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_672),
.B(n_531),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_746),
.A2(n_525),
.B(n_524),
.Y(n_822)
);

OAI21xp5_ASAP7_75t_L g823 ( 
.A1(n_762),
.A2(n_625),
.B(n_533),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_756),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_672),
.B(n_532),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_L g826 ( 
.A(n_739),
.B(n_395),
.Y(n_826)
);

OAI22xp5_ASAP7_75t_L g827 ( 
.A1(n_667),
.A2(n_543),
.B1(n_532),
.B2(n_533),
.Y(n_827)
);

BUFx4f_ASAP7_75t_L g828 ( 
.A(n_677),
.Y(n_828)
);

O2A1O1Ixp33_ASAP7_75t_L g829 ( 
.A1(n_688),
.A2(n_543),
.B(n_580),
.C(n_538),
.Y(n_829)
);

AOI21xp5_ASAP7_75t_L g830 ( 
.A1(n_738),
.A2(n_558),
.B(n_542),
.Y(n_830)
);

HB1xp67_ASAP7_75t_L g831 ( 
.A(n_675),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_705),
.A2(n_625),
.B(n_569),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_705),
.A2(n_625),
.B(n_605),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_655),
.B(n_511),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_682),
.B(n_550),
.Y(n_835)
);

AOI22xp33_ASAP7_75t_L g836 ( 
.A1(n_767),
.A2(n_397),
.B1(n_427),
.B2(n_407),
.Y(n_836)
);

INVx4_ASAP7_75t_L g837 ( 
.A(n_655),
.Y(n_837)
);

AOI21xp33_ASAP7_75t_L g838 ( 
.A1(n_757),
.A2(n_552),
.B(n_550),
.Y(n_838)
);

A2O1A1Ixp33_ASAP7_75t_L g839 ( 
.A1(n_741),
.A2(n_682),
.B(n_749),
.C(n_668),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_694),
.A2(n_605),
.B(n_517),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_780),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_745),
.B(n_552),
.Y(n_842)
);

INVx2_ASAP7_75t_SL g843 ( 
.A(n_719),
.Y(n_843)
);

OR2x6_ASAP7_75t_L g844 ( 
.A(n_767),
.B(n_464),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_792),
.B(n_756),
.Y(n_845)
);

A2O1A1Ixp33_ASAP7_75t_L g846 ( 
.A1(n_741),
.A2(n_597),
.B(n_555),
.C(n_560),
.Y(n_846)
);

INVx4_ASAP7_75t_L g847 ( 
.A(n_655),
.Y(n_847)
);

CKINVDCx8_ASAP7_75t_R g848 ( 
.A(n_710),
.Y(n_848)
);

A2O1A1Ixp33_ASAP7_75t_L g849 ( 
.A1(n_749),
.A2(n_598),
.B(n_573),
.C(n_580),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_758),
.B(n_597),
.Y(n_850)
);

OAI22xp5_ASAP7_75t_L g851 ( 
.A1(n_783),
.A2(n_604),
.B1(n_615),
.B2(n_513),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_673),
.B(n_587),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_787),
.B(n_615),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_673),
.B(n_587),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_673),
.B(n_587),
.Y(n_855)
);

AOI21xp5_ASAP7_75t_L g856 ( 
.A1(n_748),
.A2(n_517),
.B(n_513),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_748),
.A2(n_751),
.B(n_750),
.Y(n_857)
);

INVxp67_ASAP7_75t_L g858 ( 
.A(n_691),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_SL g859 ( 
.A(n_753),
.B(n_308),
.Y(n_859)
);

INVx4_ASAP7_75t_L g860 ( 
.A(n_673),
.Y(n_860)
);

INVx4_ASAP7_75t_L g861 ( 
.A(n_753),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_744),
.B(n_513),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_674),
.B(n_464),
.Y(n_863)
);

BUFx3_ASAP7_75t_L g864 ( 
.A(n_778),
.Y(n_864)
);

INVx4_ASAP7_75t_L g865 ( 
.A(n_774),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_750),
.A2(n_653),
.B(n_647),
.Y(n_866)
);

OAI21xp5_ASAP7_75t_L g867 ( 
.A1(n_762),
.A2(n_764),
.B(n_669),
.Y(n_867)
);

AOI21x1_ASAP7_75t_L g868 ( 
.A1(n_784),
.A2(n_616),
.B(n_606),
.Y(n_868)
);

A2O1A1Ixp33_ASAP7_75t_L g869 ( 
.A1(n_668),
.A2(n_653),
.B(n_647),
.C(n_517),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_773),
.B(n_529),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_751),
.A2(n_653),
.B(n_647),
.Y(n_871)
);

OAI321xp33_ASAP7_75t_L g872 ( 
.A1(n_757),
.A2(n_341),
.A3(n_333),
.B1(n_313),
.B2(n_287),
.C(n_286),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_755),
.A2(n_551),
.B(n_643),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_735),
.B(n_529),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_755),
.A2(n_551),
.B(n_643),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_744),
.B(n_529),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_773),
.B(n_551),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_760),
.A2(n_623),
.B(n_643),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_775),
.B(n_576),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_781),
.B(n_576),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_658),
.B(n_576),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_760),
.A2(n_623),
.B(n_641),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_800),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_714),
.A2(n_623),
.B(n_641),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_714),
.A2(n_641),
.B(n_590),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_809),
.Y(n_886)
);

NOR3xp33_ASAP7_75t_L g887 ( 
.A(n_789),
.B(n_332),
.C(n_334),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_775),
.B(n_590),
.Y(n_888)
);

CKINVDCx8_ASAP7_75t_R g889 ( 
.A(n_710),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_810),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_657),
.Y(n_891)
);

AOI22xp5_ASAP7_75t_L g892 ( 
.A1(n_732),
.A2(n_589),
.B1(n_591),
.B2(n_590),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_764),
.A2(n_635),
.B(n_634),
.Y(n_893)
);

O2A1O1Ixp5_ASAP7_75t_L g894 ( 
.A1(n_740),
.A2(n_606),
.B(n_635),
.C(n_634),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_725),
.A2(n_616),
.B(n_607),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_662),
.Y(n_896)
);

AOI22xp5_ASAP7_75t_L g897 ( 
.A1(n_732),
.A2(n_591),
.B1(n_589),
.B2(n_607),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_740),
.B(n_589),
.Y(n_898)
);

OAI22xp5_ASAP7_75t_L g899 ( 
.A1(n_743),
.A2(n_516),
.B1(n_326),
.B2(n_328),
.Y(n_899)
);

AO21x1_ASAP7_75t_L g900 ( 
.A1(n_692),
.A2(n_322),
.B(n_280),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_725),
.A2(n_646),
.B(n_516),
.Y(n_901)
);

BUFx3_ASAP7_75t_L g902 ( 
.A(n_778),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_687),
.B(n_796),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_734),
.A2(n_646),
.B(n_516),
.Y(n_904)
);

OAI22xp5_ASAP7_75t_L g905 ( 
.A1(n_721),
.A2(n_516),
.B1(n_326),
.B2(n_330),
.Y(n_905)
);

AOI22xp5_ASAP7_75t_L g906 ( 
.A1(n_767),
.A2(n_589),
.B1(n_591),
.B2(n_214),
.Y(n_906)
);

A2O1A1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_796),
.A2(n_276),
.B(n_284),
.C(n_283),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_664),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_734),
.A2(n_646),
.B(n_342),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_666),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_659),
.A2(n_646),
.B(n_342),
.Y(n_911)
);

BUFx6f_ASAP7_75t_L g912 ( 
.A(n_774),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_723),
.B(n_591),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_729),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_665),
.A2(n_646),
.B(n_335),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_684),
.Y(n_916)
);

AO21x1_ASAP7_75t_L g917 ( 
.A1(n_771),
.A2(n_591),
.B(n_226),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_663),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_763),
.A2(n_214),
.B(n_212),
.Y(n_919)
);

OR2x2_ASAP7_75t_L g920 ( 
.A(n_786),
.B(n_330),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_729),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_777),
.A2(n_212),
.B(n_209),
.Y(n_922)
);

OR2x6_ASAP7_75t_L g923 ( 
.A(n_768),
.B(n_476),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_724),
.B(n_451),
.Y(n_924)
);

INVx1_ASAP7_75t_SL g925 ( 
.A(n_733),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_689),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_661),
.B(n_451),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_777),
.A2(n_209),
.B(n_202),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_690),
.Y(n_929)
);

INVxp67_ASAP7_75t_L g930 ( 
.A(n_768),
.Y(n_930)
);

OAI22xp5_ASAP7_75t_L g931 ( 
.A1(n_782),
.A2(n_332),
.B1(n_334),
.B2(n_336),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_779),
.A2(n_202),
.B(n_199),
.Y(n_932)
);

OAI21xp33_ASAP7_75t_L g933 ( 
.A1(n_813),
.A2(n_336),
.B(n_338),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_661),
.B(n_452),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_727),
.A2(n_199),
.B(n_196),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_808),
.A2(n_196),
.B(n_194),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_658),
.B(n_187),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_811),
.A2(n_204),
.B(n_187),
.Y(n_938)
);

AOI33xp33_ASAP7_75t_L g939 ( 
.A1(n_807),
.A2(n_8),
.A3(n_9),
.B1(n_11),
.B2(n_12),
.B3(n_13),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_660),
.B(n_476),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_SL g941 ( 
.A(n_670),
.B(n_194),
.Y(n_941)
);

INVx3_ASAP7_75t_L g942 ( 
.A(n_742),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_685),
.B(n_452),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_693),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_696),
.Y(n_945)
);

OAI321xp33_ASAP7_75t_L g946 ( 
.A1(n_686),
.A2(n_476),
.A3(n_470),
.B1(n_466),
.B2(n_461),
.C(n_455),
.Y(n_946)
);

A2O1A1Ixp33_ASAP7_75t_L g947 ( 
.A1(n_676),
.A2(n_470),
.B(n_466),
.C(n_461),
.Y(n_947)
);

A2O1A1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_752),
.A2(n_470),
.B(n_466),
.C(n_461),
.Y(n_948)
);

NOR2x1p5_ASAP7_75t_L g949 ( 
.A(n_712),
.B(n_204),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_768),
.B(n_476),
.Y(n_950)
);

O2A1O1Ixp33_ASAP7_75t_L g951 ( 
.A1(n_718),
.A2(n_9),
.B(n_11),
.C(n_13),
.Y(n_951)
);

HB1xp67_ASAP7_75t_L g952 ( 
.A(n_707),
.Y(n_952)
);

OAI21xp5_ASAP7_75t_L g953 ( 
.A1(n_718),
.A2(n_307),
.B(n_311),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_698),
.Y(n_954)
);

OAI21xp5_ASAP7_75t_L g955 ( 
.A1(n_752),
.A2(n_307),
.B(n_311),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_700),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_722),
.B(n_702),
.Y(n_957)
);

NOR2x1p5_ASAP7_75t_SL g958 ( 
.A(n_785),
.B(n_226),
.Y(n_958)
);

NOR3xp33_ASAP7_75t_L g959 ( 
.A(n_706),
.B(n_314),
.C(n_335),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_681),
.B(n_314),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_681),
.B(n_695),
.Y(n_961)
);

OAI21xp5_ASAP7_75t_L g962 ( 
.A1(n_709),
.A2(n_318),
.B(n_320),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_812),
.A2(n_318),
.B(n_320),
.Y(n_963)
);

O2A1O1Ixp33_ASAP7_75t_L g964 ( 
.A1(n_671),
.A2(n_14),
.B(n_15),
.C(n_17),
.Y(n_964)
);

BUFx2_ASAP7_75t_L g965 ( 
.A(n_726),
.Y(n_965)
);

A2O1A1Ixp33_ASAP7_75t_L g966 ( 
.A1(n_731),
.A2(n_452),
.B(n_470),
.C(n_466),
.Y(n_966)
);

AOI22xp5_ASAP7_75t_L g967 ( 
.A1(n_695),
.A2(n_323),
.B1(n_327),
.B2(n_324),
.Y(n_967)
);

OAI21xp5_ASAP7_75t_L g968 ( 
.A1(n_713),
.A2(n_323),
.B(n_324),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_701),
.A2(n_327),
.B(n_217),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_716),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_701),
.A2(n_271),
.B(n_223),
.Y(n_971)
);

OAI21xp5_ASAP7_75t_L g972 ( 
.A1(n_769),
.A2(n_272),
.B(n_229),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_772),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_L g974 ( 
.A(n_805),
.B(n_476),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_805),
.B(n_476),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_678),
.B(n_455),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_708),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_711),
.B(n_455),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_711),
.B(n_455),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_736),
.B(n_455),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_715),
.B(n_455),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_728),
.Y(n_982)
);

AOI21x1_ASAP7_75t_L g983 ( 
.A1(n_793),
.A2(n_436),
.B(n_470),
.Y(n_983)
);

O2A1O1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_697),
.A2(n_14),
.B(n_15),
.C(n_17),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_794),
.B(n_476),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_797),
.A2(n_277),
.B(n_236),
.Y(n_986)
);

BUFx6f_ASAP7_75t_L g987 ( 
.A(n_729),
.Y(n_987)
);

INVxp67_ASAP7_75t_L g988 ( 
.A(n_765),
.Y(n_988)
);

OR2x2_ASAP7_75t_L g989 ( 
.A(n_747),
.B(n_476),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_798),
.A2(n_290),
.B(n_238),
.Y(n_990)
);

AO21x1_ASAP7_75t_L g991 ( 
.A1(n_804),
.A2(n_226),
.B(n_466),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_799),
.A2(n_292),
.B(n_240),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_754),
.B(n_470),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_759),
.Y(n_994)
);

BUFx2_ASAP7_75t_L g995 ( 
.A(n_742),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_761),
.Y(n_996)
);

NOR3xp33_ASAP7_75t_L g997 ( 
.A(n_826),
.B(n_788),
.C(n_730),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_842),
.A2(n_770),
.B1(n_804),
.B2(n_704),
.Y(n_998)
);

AOI21xp5_ASAP7_75t_L g999 ( 
.A1(n_821),
.A2(n_815),
.B(n_806),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_841),
.Y(n_1000)
);

INVx2_ASAP7_75t_L g1001 ( 
.A(n_824),
.Y(n_1001)
);

INVxp67_ASAP7_75t_L g1002 ( 
.A(n_965),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_853),
.B(n_683),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_831),
.B(n_766),
.Y(n_1004)
);

AOI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_821),
.A2(n_815),
.B(n_806),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_845),
.B(n_683),
.Y(n_1006)
);

A2O1A1Ixp33_ASAP7_75t_L g1007 ( 
.A1(n_839),
.A2(n_720),
.B(n_717),
.C(n_703),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_845),
.B(n_776),
.Y(n_1008)
);

INVx1_ASAP7_75t_SL g1009 ( 
.A(n_843),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_912),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_825),
.A2(n_802),
.B(n_729),
.Y(n_1011)
);

INVx1_ASAP7_75t_SL g1012 ( 
.A(n_920),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_912),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_883),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_886),
.Y(n_1015)
);

NOR2xp33_ASAP7_75t_L g1016 ( 
.A(n_828),
.B(n_814),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_858),
.B(n_790),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_828),
.B(n_737),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_903),
.A2(n_737),
.B1(n_795),
.B2(n_791),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_912),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_850),
.B(n_801),
.Y(n_1021)
);

NOR2xp33_ASAP7_75t_SL g1022 ( 
.A(n_848),
.B(n_699),
.Y(n_1022)
);

BUFx3_ASAP7_75t_L g1023 ( 
.A(n_864),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_890),
.Y(n_1024)
);

CKINVDCx20_ASAP7_75t_R g1025 ( 
.A(n_902),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_918),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_825),
.A2(n_802),
.B(n_737),
.Y(n_1027)
);

A2O1A1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_838),
.A2(n_801),
.B(n_737),
.C(n_466),
.Y(n_1028)
);

INVxp67_ASAP7_75t_L g1029 ( 
.A(n_859),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_903),
.B(n_470),
.Y(n_1030)
);

OR2x6_ASAP7_75t_L g1031 ( 
.A(n_844),
.B(n_455),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_891),
.Y(n_1032)
);

OAI22xp33_ASAP7_75t_L g1033 ( 
.A1(n_923),
.A2(n_452),
.B1(n_470),
.B2(n_466),
.Y(n_1033)
);

INVx1_ASAP7_75t_SL g1034 ( 
.A(n_925),
.Y(n_1034)
);

AND2x4_ASAP7_75t_L g1035 ( 
.A(n_861),
.B(n_452),
.Y(n_1035)
);

AOI22xp33_ASAP7_75t_L g1036 ( 
.A1(n_844),
.A2(n_470),
.B1(n_466),
.B2(n_461),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_835),
.A2(n_461),
.B(n_455),
.Y(n_1037)
);

OAI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_898),
.A2(n_894),
.B(n_857),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_827),
.A2(n_461),
.B(n_452),
.Y(n_1039)
);

INVx4_ASAP7_75t_L g1040 ( 
.A(n_865),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_837),
.Y(n_1041)
);

CKINVDCx11_ASAP7_75t_R g1042 ( 
.A(n_889),
.Y(n_1042)
);

BUFx2_ASAP7_75t_L g1043 ( 
.A(n_861),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_896),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_863),
.B(n_461),
.Y(n_1045)
);

O2A1O1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_838),
.A2(n_21),
.B(n_24),
.C(n_32),
.Y(n_1046)
);

AOI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_941),
.A2(n_988),
.B1(n_949),
.B2(n_844),
.Y(n_1047)
);

O2A1O1Ixp5_ASAP7_75t_L g1048 ( 
.A1(n_991),
.A2(n_785),
.B(n_452),
.C(n_436),
.Y(n_1048)
);

AOI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_960),
.A2(n_785),
.B1(n_263),
.B2(n_305),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_837),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_931),
.B(n_21),
.Y(n_1051)
);

INVx1_ASAP7_75t_SL g1052 ( 
.A(n_952),
.Y(n_1052)
);

OAI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_898),
.A2(n_262),
.B(n_245),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_836),
.B(n_923),
.Y(n_1054)
);

O2A1O1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_849),
.A2(n_24),
.B(n_32),
.C(n_34),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_908),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_880),
.B(n_785),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_865),
.B(n_872),
.Y(n_1058)
);

OAI22xp5_ASAP7_75t_L g1059 ( 
.A1(n_957),
.A2(n_268),
.B1(n_301),
.B2(n_297),
.Y(n_1059)
);

INVx4_ASAP7_75t_L g1060 ( 
.A(n_847),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_817),
.B(n_218),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_SL g1062 ( 
.A(n_995),
.B(n_260),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_910),
.Y(n_1063)
);

BUFx2_ASAP7_75t_L g1064 ( 
.A(n_950),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_957),
.B(n_35),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_916),
.B(n_35),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_926),
.B(n_40),
.Y(n_1067)
);

INVx4_ASAP7_75t_L g1068 ( 
.A(n_847),
.Y(n_1068)
);

INVx2_ASAP7_75t_SL g1069 ( 
.A(n_940),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_923),
.B(n_41),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_SL g1071 ( 
.A(n_961),
.B(n_254),
.Y(n_1071)
);

AND2x2_ASAP7_75t_L g1072 ( 
.A(n_930),
.B(n_41),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_929),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_860),
.B(n_436),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_868),
.A2(n_226),
.B(n_436),
.Y(n_1075)
);

INVx4_ASAP7_75t_L g1076 ( 
.A(n_860),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_914),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_914),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_R g1079 ( 
.A(n_914),
.B(n_921),
.Y(n_1079)
);

AOI21x1_ASAP7_75t_L g1080 ( 
.A1(n_917),
.A2(n_436),
.B(n_226),
.Y(n_1080)
);

AOI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_955),
.A2(n_436),
.B1(n_226),
.B2(n_261),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_944),
.Y(n_1082)
);

INVx3_ASAP7_75t_L g1083 ( 
.A(n_921),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_972),
.B(n_436),
.Y(n_1084)
);

BUFx6f_ASAP7_75t_L g1085 ( 
.A(n_921),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_945),
.B(n_954),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_956),
.B(n_42),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_970),
.B(n_47),
.Y(n_1088)
);

AOI22xp33_ASAP7_75t_L g1089 ( 
.A1(n_933),
.A2(n_293),
.B1(n_226),
.B2(n_55),
.Y(n_1089)
);

AND2x4_ASAP7_75t_L g1090 ( 
.A(n_862),
.B(n_48),
.Y(n_1090)
);

OAI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_819),
.A2(n_846),
.B1(n_973),
.B2(n_934),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_977),
.Y(n_1092)
);

BUFx2_ASAP7_75t_L g1093 ( 
.A(n_940),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_R g1094 ( 
.A(n_987),
.B(n_117),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_830),
.A2(n_293),
.B(n_226),
.Y(n_1095)
);

INVx4_ASAP7_75t_L g1096 ( 
.A(n_987),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_822),
.A2(n_946),
.B(n_840),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_962),
.B(n_50),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_994),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_996),
.Y(n_1100)
);

INVxp67_ASAP7_75t_L g1101 ( 
.A(n_874),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_987),
.Y(n_1102)
);

A2O1A1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_818),
.A2(n_293),
.B(n_55),
.C(n_57),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_942),
.Y(n_1104)
);

BUFx3_ASAP7_75t_L g1105 ( 
.A(n_982),
.Y(n_1105)
);

OAI22xp5_ASAP7_75t_SL g1106 ( 
.A1(n_906),
.A2(n_50),
.B1(n_60),
.B2(n_64),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_L g1107 ( 
.A(n_876),
.B(n_60),
.Y(n_1107)
);

INVxp67_ASAP7_75t_L g1108 ( 
.A(n_927),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_SL g1109 ( 
.A(n_887),
.B(n_68),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_968),
.B(n_927),
.Y(n_1110)
);

INVxp67_ASAP7_75t_L g1111 ( 
.A(n_934),
.Y(n_1111)
);

A2O1A1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_816),
.A2(n_72),
.B(n_77),
.C(n_93),
.Y(n_1112)
);

BUFx3_ASAP7_75t_L g1113 ( 
.A(n_942),
.Y(n_1113)
);

O2A1O1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_984),
.A2(n_111),
.B(n_114),
.C(n_135),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_937),
.B(n_137),
.Y(n_1115)
);

BUFx6f_ASAP7_75t_L g1116 ( 
.A(n_989),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_959),
.B(n_142),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_967),
.B(n_152),
.Y(n_1118)
);

O2A1O1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_907),
.A2(n_159),
.B(n_161),
.C(n_162),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_870),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_820),
.A2(n_168),
.B(n_170),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_905),
.B(n_953),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_892),
.B(n_829),
.Y(n_1123)
);

OAI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_851),
.A2(n_924),
.B1(n_879),
.B2(n_870),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_SL g1125 ( 
.A(n_900),
.B(n_935),
.Y(n_1125)
);

INVx3_ASAP7_75t_L g1126 ( 
.A(n_985),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_877),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_924),
.B(n_939),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_852),
.Y(n_1129)
);

O2A1O1Ixp5_ASAP7_75t_L g1130 ( 
.A1(n_867),
.A2(n_869),
.B(n_948),
.C(n_966),
.Y(n_1130)
);

INVxp67_ASAP7_75t_L g1131 ( 
.A(n_978),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_SL g1132 ( 
.A(n_899),
.B(n_969),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_R g1133 ( 
.A(n_978),
.B(n_979),
.Y(n_1133)
);

O2A1O1Ixp5_ASAP7_75t_L g1134 ( 
.A1(n_834),
.A2(n_947),
.B(n_855),
.C(n_854),
.Y(n_1134)
);

AOI21x1_ASAP7_75t_L g1135 ( 
.A1(n_983),
.A2(n_943),
.B(n_980),
.Y(n_1135)
);

NOR3xp33_ASAP7_75t_SL g1136 ( 
.A(n_932),
.B(n_919),
.C(n_964),
.Y(n_1136)
);

O2A1O1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_951),
.A2(n_888),
.B(n_879),
.C(n_877),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_833),
.A2(n_895),
.B(n_882),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_922),
.B(n_928),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_856),
.A2(n_873),
.B(n_866),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_871),
.A2(n_875),
.B(n_878),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_888),
.B(n_980),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_881),
.B(n_938),
.Y(n_1143)
);

AOI21x1_ASAP7_75t_L g1144 ( 
.A1(n_943),
.A2(n_911),
.B(n_915),
.Y(n_1144)
);

AOI22xp33_ASAP7_75t_L g1145 ( 
.A1(n_979),
.A2(n_913),
.B1(n_936),
.B2(n_963),
.Y(n_1145)
);

INVx1_ASAP7_75t_SL g1146 ( 
.A(n_981),
.Y(n_1146)
);

BUFx3_ASAP7_75t_L g1147 ( 
.A(n_1023),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1142),
.A2(n_823),
.B(n_976),
.Y(n_1148)
);

OAI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1122),
.A2(n_913),
.B(n_832),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_L g1150 ( 
.A1(n_1075),
.A2(n_893),
.B(n_885),
.Y(n_1150)
);

INVx4_ASAP7_75t_L g1151 ( 
.A(n_1042),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_1138),
.A2(n_884),
.B(n_981),
.Y(n_1152)
);

BUFx2_ASAP7_75t_L g1153 ( 
.A(n_1102),
.Y(n_1153)
);

AO31x2_ASAP7_75t_L g1154 ( 
.A1(n_1028),
.A2(n_976),
.A3(n_993),
.B(n_974),
.Y(n_1154)
);

BUFx8_ASAP7_75t_L g1155 ( 
.A(n_1043),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1138),
.A2(n_993),
.B(n_901),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1097),
.A2(n_975),
.B(n_904),
.Y(n_1157)
);

NAND2xp33_ASAP7_75t_SL g1158 ( 
.A(n_1051),
.B(n_1040),
.Y(n_1158)
);

AOI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_998),
.A2(n_1106),
.B1(n_1003),
.B2(n_1047),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1000),
.Y(n_1160)
);

INVxp67_ASAP7_75t_L g1161 ( 
.A(n_1004),
.Y(n_1161)
);

INVx1_ASAP7_75t_SL g1162 ( 
.A(n_1052),
.Y(n_1162)
);

AO31x2_ASAP7_75t_L g1163 ( 
.A1(n_1037),
.A2(n_992),
.A3(n_986),
.B(n_990),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1012),
.B(n_971),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1097),
.A2(n_1124),
.B(n_1123),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1014),
.Y(n_1166)
);

O2A1O1Ixp33_ASAP7_75t_SL g1167 ( 
.A1(n_1110),
.A2(n_909),
.B(n_897),
.C(n_958),
.Y(n_1167)
);

CKINVDCx20_ASAP7_75t_R g1168 ( 
.A(n_1025),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1140),
.A2(n_1141),
.B(n_1091),
.Y(n_1169)
);

INVxp67_ASAP7_75t_SL g1170 ( 
.A(n_1002),
.Y(n_1170)
);

OR2x2_ASAP7_75t_L g1171 ( 
.A(n_1002),
.B(n_1009),
.Y(n_1171)
);

OAI21xp33_ASAP7_75t_L g1172 ( 
.A1(n_1098),
.A2(n_997),
.B(n_1103),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1015),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1140),
.A2(n_1141),
.B(n_1030),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1011),
.A2(n_1027),
.B(n_1037),
.Y(n_1175)
);

NAND3xp33_ASAP7_75t_L g1176 ( 
.A(n_1046),
.B(n_1055),
.C(n_1114),
.Y(n_1176)
);

NOR2xp33_ASAP7_75t_L g1177 ( 
.A(n_1101),
.B(n_1034),
.Y(n_1177)
);

INVx1_ASAP7_75t_SL g1178 ( 
.A(n_1010),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1011),
.A2(n_1027),
.B(n_999),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_999),
.A2(n_1005),
.B(n_1038),
.Y(n_1180)
);

A2O1A1Ixp33_ASAP7_75t_L g1181 ( 
.A1(n_1061),
.A2(n_1114),
.B(n_1115),
.C(n_1046),
.Y(n_1181)
);

BUFx2_ASAP7_75t_L g1182 ( 
.A(n_1079),
.Y(n_1182)
);

OAI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1134),
.A2(n_1130),
.B(n_1005),
.Y(n_1183)
);

AO21x1_ASAP7_75t_L g1184 ( 
.A1(n_1055),
.A2(n_1125),
.B(n_1033),
.Y(n_1184)
);

AO22x2_ASAP7_75t_L g1185 ( 
.A1(n_1054),
.A2(n_1070),
.B1(n_1126),
.B2(n_1131),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_1006),
.B(n_1021),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1080),
.A2(n_1095),
.B(n_1135),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1016),
.B(n_1086),
.Y(n_1188)
);

OAI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1065),
.A2(n_1128),
.B1(n_1031),
.B2(n_1108),
.Y(n_1189)
);

O2A1O1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1112),
.A2(n_1109),
.B(n_1132),
.C(n_1117),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1144),
.A2(n_1048),
.B(n_1039),
.Y(n_1191)
);

BUFx2_ASAP7_75t_L g1192 ( 
.A(n_1010),
.Y(n_1192)
);

BUFx6f_ASAP7_75t_L g1193 ( 
.A(n_1010),
.Y(n_1193)
);

AO32x2_ASAP7_75t_L g1194 ( 
.A1(n_1019),
.A2(n_1069),
.A3(n_1059),
.B1(n_1096),
.B2(n_1133),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1031),
.A2(n_1108),
.B1(n_1111),
.B2(n_1049),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1039),
.A2(n_1084),
.B(n_1137),
.Y(n_1196)
);

CKINVDCx11_ASAP7_75t_R g1197 ( 
.A(n_1013),
.Y(n_1197)
);

INVx2_ASAP7_75t_SL g1198 ( 
.A(n_1013),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1024),
.B(n_1032),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1044),
.B(n_1056),
.Y(n_1200)
);

AOI221xp5_ASAP7_75t_SL g1201 ( 
.A1(n_1107),
.A2(n_1067),
.B1(n_1087),
.B2(n_1088),
.C(n_1066),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1063),
.Y(n_1202)
);

NOR2xp33_ASAP7_75t_L g1203 ( 
.A(n_1029),
.B(n_1090),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1048),
.A2(n_1130),
.B(n_1134),
.Y(n_1204)
);

A2O1A1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1081),
.A2(n_1137),
.B(n_1119),
.C(n_1089),
.Y(n_1205)
);

INVx6_ASAP7_75t_L g1206 ( 
.A(n_1013),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1057),
.A2(n_1007),
.B(n_1120),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1073),
.Y(n_1208)
);

NAND2xp33_ASAP7_75t_SL g1209 ( 
.A(n_1040),
.B(n_1104),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1082),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1127),
.A2(n_1121),
.B(n_1045),
.Y(n_1211)
);

OAI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1031),
.A2(n_1111),
.B1(n_1145),
.B2(n_1036),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1099),
.Y(n_1213)
);

OAI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1053),
.A2(n_1143),
.B(n_1017),
.Y(n_1214)
);

INVx3_ASAP7_75t_L g1215 ( 
.A(n_1096),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1100),
.Y(n_1216)
);

OA21x2_ASAP7_75t_L g1217 ( 
.A1(n_1131),
.A2(n_1121),
.B(n_1136),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1026),
.Y(n_1218)
);

BUFx3_ASAP7_75t_L g1219 ( 
.A(n_1020),
.Y(n_1219)
);

OAI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1058),
.A2(n_1071),
.B(n_1118),
.Y(n_1220)
);

OAI22x1_ASAP7_75t_L g1221 ( 
.A1(n_1090),
.A2(n_1072),
.B1(n_1064),
.B2(n_1018),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1008),
.B(n_1105),
.Y(n_1222)
);

NOR2xp67_ASAP7_75t_L g1223 ( 
.A(n_1083),
.B(n_1041),
.Y(n_1223)
);

BUFx2_ASAP7_75t_SL g1224 ( 
.A(n_1020),
.Y(n_1224)
);

HB1xp67_ASAP7_75t_L g1225 ( 
.A(n_1093),
.Y(n_1225)
);

AO22x1_ASAP7_75t_L g1226 ( 
.A1(n_1035),
.A2(n_1020),
.B1(n_1113),
.B2(n_1092),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1074),
.A2(n_1139),
.B(n_1146),
.Y(n_1227)
);

AO21x1_ASAP7_75t_L g1228 ( 
.A1(n_1119),
.A2(n_1035),
.B(n_1022),
.Y(n_1228)
);

AOI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1116),
.A2(n_1062),
.B1(n_1104),
.B2(n_1129),
.Y(n_1229)
);

BUFx2_ASAP7_75t_L g1230 ( 
.A(n_1077),
.Y(n_1230)
);

INVxp67_ASAP7_75t_SL g1231 ( 
.A(n_1116),
.Y(n_1231)
);

AND2x4_ASAP7_75t_L g1232 ( 
.A(n_1060),
.B(n_1068),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1104),
.A2(n_1041),
.B(n_1050),
.Y(n_1233)
);

INVx3_ASAP7_75t_L g1234 ( 
.A(n_1077),
.Y(n_1234)
);

NAND3xp33_ASAP7_75t_L g1235 ( 
.A(n_1129),
.B(n_1116),
.C(n_1077),
.Y(n_1235)
);

OR2x2_ASAP7_75t_L g1236 ( 
.A(n_1083),
.B(n_1050),
.Y(n_1236)
);

AOI221x1_ASAP7_75t_L g1237 ( 
.A1(n_1129),
.A2(n_1078),
.B1(n_1085),
.B2(n_1076),
.C(n_1094),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1078),
.A2(n_1085),
.B(n_821),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1078),
.A2(n_825),
.B(n_821),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1085),
.A2(n_825),
.B(n_821),
.Y(n_1240)
);

HB1xp67_ASAP7_75t_L g1241 ( 
.A(n_1052),
.Y(n_1241)
);

O2A1O1Ixp33_ASAP7_75t_SL g1242 ( 
.A1(n_1110),
.A2(n_839),
.B(n_1122),
.C(n_1098),
.Y(n_1242)
);

BUFx2_ASAP7_75t_L g1243 ( 
.A(n_1102),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1122),
.A2(n_842),
.B(n_739),
.Y(n_1244)
);

AOI221xp5_ASAP7_75t_SL g1245 ( 
.A1(n_1055),
.A2(n_656),
.B1(n_757),
.B2(n_933),
.C(n_1051),
.Y(n_1245)
);

AOI21x1_ASAP7_75t_L g1246 ( 
.A1(n_1080),
.A2(n_1144),
.B(n_1097),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_998),
.A2(n_842),
.B1(n_839),
.B2(n_739),
.Y(n_1247)
);

AO31x2_ASAP7_75t_L g1248 ( 
.A1(n_1028),
.A2(n_991),
.A3(n_917),
.B(n_1037),
.Y(n_1248)
);

OAI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1075),
.A2(n_1138),
.B(n_1080),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1001),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1142),
.A2(n_825),
.B(n_821),
.Y(n_1251)
);

A2O1A1Ixp33_ASAP7_75t_SL g1252 ( 
.A1(n_1143),
.A2(n_559),
.B(n_997),
.C(n_536),
.Y(n_1252)
);

O2A1O1Ixp33_ASAP7_75t_SL g1253 ( 
.A1(n_1110),
.A2(n_839),
.B(n_1122),
.C(n_1098),
.Y(n_1253)
);

OR2x6_ASAP7_75t_L g1254 ( 
.A(n_1023),
.B(n_861),
.Y(n_1254)
);

BUFx2_ASAP7_75t_L g1255 ( 
.A(n_1102),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1000),
.Y(n_1256)
);

INVx1_ASAP7_75t_SL g1257 ( 
.A(n_1042),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1000),
.Y(n_1258)
);

AOI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_998),
.A2(n_757),
.B1(n_842),
.B2(n_745),
.Y(n_1259)
);

O2A1O1Ixp33_ASAP7_75t_SL g1260 ( 
.A1(n_1110),
.A2(n_839),
.B(n_1122),
.C(n_1098),
.Y(n_1260)
);

A2O1A1Ixp33_ASAP7_75t_L g1261 ( 
.A1(n_998),
.A2(n_842),
.B(n_739),
.C(n_839),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1000),
.Y(n_1262)
);

A2O1A1Ixp33_ASAP7_75t_L g1263 ( 
.A1(n_998),
.A2(n_842),
.B(n_739),
.C(n_839),
.Y(n_1263)
);

NOR2xp67_ASAP7_75t_SL g1264 ( 
.A(n_1023),
.B(n_563),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1000),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1012),
.B(n_739),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1142),
.A2(n_825),
.B(n_821),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1142),
.A2(n_825),
.B(n_821),
.Y(n_1268)
);

AO31x2_ASAP7_75t_L g1269 ( 
.A1(n_1028),
.A2(n_991),
.A3(n_917),
.B(n_1037),
.Y(n_1269)
);

OAI21xp5_ASAP7_75t_SL g1270 ( 
.A1(n_1051),
.A2(n_745),
.B(n_757),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1012),
.B(n_739),
.Y(n_1271)
);

AOI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1142),
.A2(n_825),
.B(n_821),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1142),
.A2(n_825),
.B(n_821),
.Y(n_1273)
);

A2O1A1Ixp33_ASAP7_75t_L g1274 ( 
.A1(n_998),
.A2(n_842),
.B(n_739),
.C(n_839),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1000),
.Y(n_1275)
);

AO32x2_ASAP7_75t_L g1276 ( 
.A1(n_1106),
.A2(n_1091),
.A3(n_1124),
.B1(n_998),
.B2(n_1019),
.Y(n_1276)
);

NAND3x1_ASAP7_75t_L g1277 ( 
.A(n_1047),
.B(n_1051),
.C(n_745),
.Y(n_1277)
);

AOI221x1_ASAP7_75t_L g1278 ( 
.A1(n_1106),
.A2(n_997),
.B1(n_1103),
.B2(n_767),
.C(n_768),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1012),
.B(n_739),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1012),
.B(n_739),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1012),
.B(n_739),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_SL g1282 ( 
.A(n_1025),
.B(n_586),
.Y(n_1282)
);

INVxp67_ASAP7_75t_L g1283 ( 
.A(n_1004),
.Y(n_1283)
);

OAI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1122),
.A2(n_842),
.B(n_739),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1012),
.B(n_739),
.Y(n_1285)
);

NAND2xp33_ASAP7_75t_L g1286 ( 
.A(n_997),
.B(n_655),
.Y(n_1286)
);

O2A1O1Ixp33_ASAP7_75t_L g1287 ( 
.A1(n_1122),
.A2(n_739),
.B(n_745),
.C(n_839),
.Y(n_1287)
);

NOR2xp33_ASAP7_75t_SL g1288 ( 
.A(n_1025),
.B(n_586),
.Y(n_1288)
);

CKINVDCx11_ASAP7_75t_R g1289 ( 
.A(n_1025),
.Y(n_1289)
);

BUFx2_ASAP7_75t_L g1290 ( 
.A(n_1102),
.Y(n_1290)
);

A2O1A1Ixp33_ASAP7_75t_L g1291 ( 
.A1(n_998),
.A2(n_842),
.B(n_739),
.C(n_839),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1001),
.Y(n_1292)
);

INVx2_ASAP7_75t_L g1293 ( 
.A(n_1001),
.Y(n_1293)
);

OR2x6_ASAP7_75t_L g1294 ( 
.A(n_1023),
.B(n_861),
.Y(n_1294)
);

AOI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1142),
.A2(n_825),
.B(n_821),
.Y(n_1295)
);

OR2x6_ASAP7_75t_L g1296 ( 
.A(n_1023),
.B(n_861),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1012),
.B(n_739),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1142),
.A2(n_825),
.B(n_821),
.Y(n_1298)
);

A2O1A1Ixp33_ASAP7_75t_L g1299 ( 
.A1(n_998),
.A2(n_842),
.B(n_739),
.C(n_839),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1000),
.Y(n_1300)
);

AO22x1_ASAP7_75t_L g1301 ( 
.A1(n_1054),
.A2(n_485),
.B1(n_745),
.B2(n_354),
.Y(n_1301)
);

INVxp67_ASAP7_75t_L g1302 ( 
.A(n_1004),
.Y(n_1302)
);

AO31x2_ASAP7_75t_L g1303 ( 
.A1(n_1028),
.A2(n_991),
.A3(n_917),
.B(n_1037),
.Y(n_1303)
);

NAND2x1p5_ASAP7_75t_L g1304 ( 
.A(n_1182),
.B(n_1219),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1199),
.Y(n_1305)
);

BUFx6f_ASAP7_75t_L g1306 ( 
.A(n_1197),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1237),
.B(n_1231),
.Y(n_1307)
);

AOI22xp33_ASAP7_75t_L g1308 ( 
.A1(n_1259),
.A2(n_1159),
.B1(n_1247),
.B2(n_1176),
.Y(n_1308)
);

BUFx2_ASAP7_75t_L g1309 ( 
.A(n_1155),
.Y(n_1309)
);

AOI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1259),
.A2(n_1270),
.B1(n_1159),
.B2(n_1277),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_SL g1311 ( 
.A1(n_1176),
.A2(n_1185),
.B1(n_1278),
.B2(n_1244),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1172),
.A2(n_1284),
.B1(n_1184),
.B2(n_1203),
.Y(n_1312)
);

INVx6_ASAP7_75t_L g1313 ( 
.A(n_1155),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_SL g1314 ( 
.A1(n_1185),
.A2(n_1189),
.B1(n_1212),
.B2(n_1214),
.Y(n_1314)
);

CKINVDCx20_ASAP7_75t_R g1315 ( 
.A(n_1289),
.Y(n_1315)
);

BUFx10_ASAP7_75t_L g1316 ( 
.A(n_1177),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1188),
.B(n_1161),
.Y(n_1317)
);

OAI22xp5_ASAP7_75t_L g1318 ( 
.A1(n_1261),
.A2(n_1263),
.B1(n_1291),
.B2(n_1274),
.Y(n_1318)
);

INVx8_ASAP7_75t_L g1319 ( 
.A(n_1168),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1200),
.Y(n_1320)
);

INVx2_ASAP7_75t_SL g1321 ( 
.A(n_1147),
.Y(n_1321)
);

BUFx2_ASAP7_75t_SL g1322 ( 
.A(n_1151),
.Y(n_1322)
);

AOI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1282),
.A2(n_1288),
.B1(n_1283),
.B2(n_1302),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1172),
.A2(n_1221),
.B1(n_1186),
.B2(n_1158),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_1257),
.Y(n_1325)
);

INVx2_ASAP7_75t_SL g1326 ( 
.A(n_1153),
.Y(n_1326)
);

INVx3_ASAP7_75t_L g1327 ( 
.A(n_1193),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1299),
.A2(n_1181),
.B1(n_1287),
.B2(n_1165),
.Y(n_1328)
);

BUFx12f_ASAP7_75t_L g1329 ( 
.A(n_1151),
.Y(n_1329)
);

BUFx8_ASAP7_75t_SL g1330 ( 
.A(n_1243),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1160),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1205),
.A2(n_1170),
.B1(n_1279),
.B2(n_1285),
.Y(n_1332)
);

CKINVDCx20_ASAP7_75t_R g1333 ( 
.A(n_1255),
.Y(n_1333)
);

BUFx3_ASAP7_75t_L g1334 ( 
.A(n_1290),
.Y(n_1334)
);

INVx6_ASAP7_75t_L g1335 ( 
.A(n_1254),
.Y(n_1335)
);

OAI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1266),
.A2(n_1271),
.B1(n_1280),
.B2(n_1281),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1220),
.A2(n_1228),
.B1(n_1222),
.B2(n_1216),
.Y(n_1337)
);

INVx6_ASAP7_75t_L g1338 ( 
.A(n_1254),
.Y(n_1338)
);

OAI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1297),
.A2(n_1164),
.B1(n_1171),
.B2(n_1195),
.Y(n_1339)
);

INVx6_ASAP7_75t_L g1340 ( 
.A(n_1294),
.Y(n_1340)
);

OAI21xp5_ASAP7_75t_SL g1341 ( 
.A1(n_1183),
.A2(n_1190),
.B(n_1169),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1166),
.Y(n_1342)
);

CKINVDCx11_ASAP7_75t_R g1343 ( 
.A(n_1294),
.Y(n_1343)
);

CKINVDCx11_ASAP7_75t_R g1344 ( 
.A(n_1296),
.Y(n_1344)
);

BUFx12f_ASAP7_75t_L g1345 ( 
.A(n_1296),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1173),
.Y(n_1346)
);

OAI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1251),
.A2(n_1268),
.B1(n_1267),
.B2(n_1272),
.Y(n_1347)
);

BUFx3_ASAP7_75t_L g1348 ( 
.A(n_1206),
.Y(n_1348)
);

BUFx2_ASAP7_75t_L g1349 ( 
.A(n_1225),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1213),
.A2(n_1208),
.B1(n_1265),
.B2(n_1275),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1202),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1210),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1256),
.Y(n_1353)
);

BUFx2_ASAP7_75t_L g1354 ( 
.A(n_1193),
.Y(n_1354)
);

BUFx10_ASAP7_75t_L g1355 ( 
.A(n_1206),
.Y(n_1355)
);

BUFx3_ASAP7_75t_L g1356 ( 
.A(n_1192),
.Y(n_1356)
);

BUFx4f_ASAP7_75t_SL g1357 ( 
.A(n_1162),
.Y(n_1357)
);

OAI22xp5_ASAP7_75t_SL g1358 ( 
.A1(n_1301),
.A2(n_1229),
.B1(n_1241),
.B2(n_1300),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1258),
.Y(n_1359)
);

OAI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1276),
.A2(n_1262),
.B1(n_1245),
.B2(n_1229),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_SL g1361 ( 
.A1(n_1276),
.A2(n_1217),
.B1(n_1298),
.B2(n_1295),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1273),
.A2(n_1240),
.B1(n_1239),
.B2(n_1217),
.Y(n_1362)
);

CKINVDCx11_ASAP7_75t_R g1363 ( 
.A(n_1230),
.Y(n_1363)
);

OAI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1276),
.A2(n_1252),
.B1(n_1207),
.B2(n_1196),
.Y(n_1364)
);

BUFx12f_ASAP7_75t_L g1365 ( 
.A(n_1198),
.Y(n_1365)
);

BUFx2_ASAP7_75t_L g1366 ( 
.A(n_1234),
.Y(n_1366)
);

BUFx4_ASAP7_75t_R g1367 ( 
.A(n_1226),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1218),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_SL g1369 ( 
.A1(n_1286),
.A2(n_1201),
.B1(n_1149),
.B2(n_1194),
.Y(n_1369)
);

OAI21xp5_ASAP7_75t_SL g1370 ( 
.A1(n_1180),
.A2(n_1232),
.B(n_1179),
.Y(n_1370)
);

OAI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1236),
.A2(n_1227),
.B1(n_1223),
.B2(n_1148),
.Y(n_1371)
);

INVx6_ASAP7_75t_L g1372 ( 
.A(n_1232),
.Y(n_1372)
);

CKINVDCx6p67_ASAP7_75t_R g1373 ( 
.A(n_1224),
.Y(n_1373)
);

OAI22xp33_ASAP7_75t_SL g1374 ( 
.A1(n_1250),
.A2(n_1293),
.B1(n_1292),
.B2(n_1178),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1264),
.B(n_1234),
.Y(n_1375)
);

BUFx10_ASAP7_75t_L g1376 ( 
.A(n_1209),
.Y(n_1376)
);

BUFx2_ASAP7_75t_L g1377 ( 
.A(n_1215),
.Y(n_1377)
);

CKINVDCx11_ASAP7_75t_R g1378 ( 
.A(n_1223),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1215),
.A2(n_1238),
.B1(n_1211),
.B2(n_1235),
.Y(n_1379)
);

BUFx12f_ASAP7_75t_L g1380 ( 
.A(n_1235),
.Y(n_1380)
);

CKINVDCx20_ASAP7_75t_R g1381 ( 
.A(n_1233),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_SL g1382 ( 
.A(n_1157),
.B(n_1175),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1204),
.A2(n_1253),
.B1(n_1242),
.B2(n_1260),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1194),
.A2(n_1174),
.B1(n_1156),
.B2(n_1152),
.Y(n_1384)
);

BUFx3_ASAP7_75t_L g1385 ( 
.A(n_1154),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1194),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1150),
.A2(n_1191),
.B1(n_1187),
.B2(n_1249),
.Y(n_1387)
);

AOI22xp33_ASAP7_75t_L g1388 ( 
.A1(n_1167),
.A2(n_1248),
.B1(n_1269),
.B2(n_1303),
.Y(n_1388)
);

CKINVDCx11_ASAP7_75t_R g1389 ( 
.A(n_1163),
.Y(n_1389)
);

INVxp67_ASAP7_75t_SL g1390 ( 
.A(n_1246),
.Y(n_1390)
);

INVx5_ASAP7_75t_L g1391 ( 
.A(n_1269),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_L g1392 ( 
.A1(n_1303),
.A2(n_1259),
.B1(n_767),
.B2(n_768),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1199),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1259),
.A2(n_767),
.B1(n_768),
.B2(n_844),
.Y(n_1394)
);

INVx2_ASAP7_75t_SL g1395 ( 
.A(n_1147),
.Y(n_1395)
);

OAI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1259),
.A2(n_1261),
.B1(n_1274),
.B2(n_1263),
.Y(n_1396)
);

BUFx4f_ASAP7_75t_SL g1397 ( 
.A(n_1168),
.Y(n_1397)
);

BUFx6f_ASAP7_75t_SL g1398 ( 
.A(n_1151),
.Y(n_1398)
);

CKINVDCx6p67_ASAP7_75t_R g1399 ( 
.A(n_1289),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1199),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1199),
.Y(n_1401)
);

BUFx6f_ASAP7_75t_L g1402 ( 
.A(n_1197),
.Y(n_1402)
);

OAI22xp5_ASAP7_75t_L g1403 ( 
.A1(n_1259),
.A2(n_1261),
.B1(n_1274),
.B2(n_1263),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1199),
.Y(n_1404)
);

INVx6_ASAP7_75t_L g1405 ( 
.A(n_1155),
.Y(n_1405)
);

BUFx3_ASAP7_75t_L g1406 ( 
.A(n_1182),
.Y(n_1406)
);

BUFx8_ASAP7_75t_L g1407 ( 
.A(n_1153),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_1289),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1199),
.Y(n_1409)
);

OAI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1259),
.A2(n_1261),
.B1(n_1274),
.B2(n_1263),
.Y(n_1410)
);

BUFx3_ASAP7_75t_L g1411 ( 
.A(n_1182),
.Y(n_1411)
);

BUFx2_ASAP7_75t_SL g1412 ( 
.A(n_1168),
.Y(n_1412)
);

AND2x4_ASAP7_75t_SL g1413 ( 
.A(n_1254),
.B(n_1294),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1259),
.A2(n_767),
.B1(n_768),
.B2(n_844),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1199),
.Y(n_1415)
);

BUFx6f_ASAP7_75t_L g1416 ( 
.A(n_1197),
.Y(n_1416)
);

INVx1_ASAP7_75t_SL g1417 ( 
.A(n_1162),
.Y(n_1417)
);

OAI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1259),
.A2(n_1261),
.B1(n_1274),
.B2(n_1263),
.Y(n_1418)
);

BUFx2_ASAP7_75t_L g1419 ( 
.A(n_1155),
.Y(n_1419)
);

INVx4_ASAP7_75t_L g1420 ( 
.A(n_1197),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1259),
.A2(n_1261),
.B1(n_1274),
.B2(n_1263),
.Y(n_1421)
);

INVx1_ASAP7_75t_SL g1422 ( 
.A(n_1162),
.Y(n_1422)
);

INVx4_ASAP7_75t_L g1423 ( 
.A(n_1197),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_SL g1424 ( 
.A1(n_1247),
.A2(n_768),
.B1(n_767),
.B2(n_844),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1199),
.Y(n_1425)
);

OAI22xp5_ASAP7_75t_L g1426 ( 
.A1(n_1259),
.A2(n_1261),
.B1(n_1274),
.B2(n_1263),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1259),
.A2(n_767),
.B1(n_768),
.B2(n_844),
.Y(n_1427)
);

INVx4_ASAP7_75t_L g1428 ( 
.A(n_1367),
.Y(n_1428)
);

BUFx6f_ASAP7_75t_L g1429 ( 
.A(n_1391),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1317),
.B(n_1305),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1331),
.Y(n_1431)
);

OAI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1362),
.A2(n_1382),
.B(n_1384),
.Y(n_1432)
);

BUFx3_ASAP7_75t_L g1433 ( 
.A(n_1307),
.Y(n_1433)
);

BUFx3_ASAP7_75t_L g1434 ( 
.A(n_1307),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1342),
.Y(n_1435)
);

AOI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1382),
.A2(n_1347),
.B(n_1328),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1386),
.B(n_1346),
.Y(n_1437)
);

NAND2x1p5_ASAP7_75t_L g1438 ( 
.A(n_1391),
.B(n_1310),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1351),
.Y(n_1439)
);

NOR2xp33_ASAP7_75t_L g1440 ( 
.A(n_1397),
.B(n_1357),
.Y(n_1440)
);

INVx1_ASAP7_75t_SL g1441 ( 
.A(n_1357),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1352),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_1408),
.Y(n_1443)
);

BUFx12f_ASAP7_75t_L g1444 ( 
.A(n_1343),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1353),
.Y(n_1445)
);

OA21x2_ASAP7_75t_L g1446 ( 
.A1(n_1341),
.A2(n_1384),
.B(n_1388),
.Y(n_1446)
);

CKINVDCx8_ASAP7_75t_R g1447 ( 
.A(n_1412),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1359),
.B(n_1385),
.Y(n_1448)
);

INVx2_ASAP7_75t_SL g1449 ( 
.A(n_1335),
.Y(n_1449)
);

AO21x2_ASAP7_75t_L g1450 ( 
.A1(n_1364),
.A2(n_1360),
.B(n_1339),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1368),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1390),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1390),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1308),
.B(n_1350),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1370),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1350),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1379),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1320),
.Y(n_1458)
);

AND2x4_ASAP7_75t_L g1459 ( 
.A(n_1388),
.B(n_1356),
.Y(n_1459)
);

OA21x2_ASAP7_75t_L g1460 ( 
.A1(n_1387),
.A2(n_1337),
.B(n_1383),
.Y(n_1460)
);

INVx3_ASAP7_75t_L g1461 ( 
.A(n_1389),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1393),
.Y(n_1462)
);

INVx3_ASAP7_75t_L g1463 ( 
.A(n_1389),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1308),
.B(n_1361),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1400),
.Y(n_1465)
);

OAI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1396),
.A2(n_1421),
.B(n_1426),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1401),
.Y(n_1467)
);

AND2x2_ASAP7_75t_L g1468 ( 
.A(n_1361),
.B(n_1314),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1404),
.Y(n_1469)
);

INVx3_ASAP7_75t_L g1470 ( 
.A(n_1376),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1409),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1415),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1425),
.B(n_1332),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1360),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1371),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1314),
.B(n_1392),
.Y(n_1476)
);

OAI21x1_ASAP7_75t_L g1477 ( 
.A1(n_1387),
.A2(n_1383),
.B(n_1318),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_1399),
.Y(n_1478)
);

AOI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1403),
.A2(n_1410),
.B(n_1418),
.Y(n_1479)
);

OAI21x1_ASAP7_75t_L g1480 ( 
.A1(n_1337),
.A2(n_1324),
.B(n_1312),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1371),
.Y(n_1481)
);

INVx4_ASAP7_75t_L g1482 ( 
.A(n_1367),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1424),
.A2(n_1427),
.B1(n_1414),
.B2(n_1394),
.Y(n_1483)
);

HB1xp67_ASAP7_75t_L g1484 ( 
.A(n_1349),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1381),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1366),
.Y(n_1486)
);

OAI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1324),
.A2(n_1312),
.B(n_1327),
.Y(n_1487)
);

BUFx3_ASAP7_75t_L g1488 ( 
.A(n_1380),
.Y(n_1488)
);

OAI21x1_ASAP7_75t_L g1489 ( 
.A1(n_1392),
.A2(n_1304),
.B(n_1375),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1354),
.Y(n_1490)
);

INVx3_ASAP7_75t_L g1491 ( 
.A(n_1376),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1369),
.Y(n_1492)
);

INVx8_ASAP7_75t_L g1493 ( 
.A(n_1345),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1336),
.B(n_1339),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1311),
.Y(n_1495)
);

HB1xp67_ASAP7_75t_L g1496 ( 
.A(n_1377),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1311),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1424),
.B(n_1427),
.Y(n_1498)
);

OA21x2_ASAP7_75t_L g1499 ( 
.A1(n_1394),
.A2(n_1414),
.B(n_1323),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1374),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1358),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1417),
.B(n_1422),
.Y(n_1502)
);

AO21x1_ASAP7_75t_SL g1503 ( 
.A1(n_1378),
.A2(n_1372),
.B(n_1373),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1334),
.B(n_1411),
.Y(n_1504)
);

INVx2_ASAP7_75t_SL g1505 ( 
.A(n_1338),
.Y(n_1505)
);

AO21x1_ASAP7_75t_SL g1506 ( 
.A1(n_1372),
.A2(n_1344),
.B(n_1343),
.Y(n_1506)
);

INVx2_ASAP7_75t_SL g1507 ( 
.A(n_1340),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1413),
.B(n_1334),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1406),
.Y(n_1509)
);

AOI21x1_ASAP7_75t_L g1510 ( 
.A1(n_1326),
.A2(n_1309),
.B(n_1419),
.Y(n_1510)
);

INVx2_ASAP7_75t_SL g1511 ( 
.A(n_1411),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1511),
.B(n_1316),
.Y(n_1512)
);

OR2x6_ASAP7_75t_L g1513 ( 
.A(n_1428),
.B(n_1306),
.Y(n_1513)
);

OR2x2_ASAP7_75t_L g1514 ( 
.A(n_1484),
.B(n_1423),
.Y(n_1514)
);

AND2x4_ASAP7_75t_L g1515 ( 
.A(n_1433),
.B(n_1306),
.Y(n_1515)
);

A2O1A1Ixp33_ASAP7_75t_L g1516 ( 
.A1(n_1479),
.A2(n_1306),
.B(n_1416),
.C(n_1402),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1451),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1511),
.B(n_1316),
.Y(n_1518)
);

OAI21xp5_ASAP7_75t_L g1519 ( 
.A1(n_1466),
.A2(n_1395),
.B(n_1321),
.Y(n_1519)
);

AOI221xp5_ASAP7_75t_L g1520 ( 
.A1(n_1494),
.A2(n_1398),
.B1(n_1325),
.B2(n_1319),
.C(n_1416),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1476),
.A2(n_1344),
.B1(n_1416),
.B2(n_1402),
.Y(n_1521)
);

O2A1O1Ixp33_ASAP7_75t_L g1522 ( 
.A1(n_1455),
.A2(n_1348),
.B(n_1333),
.C(n_1315),
.Y(n_1522)
);

OA21x2_ASAP7_75t_L g1523 ( 
.A1(n_1432),
.A2(n_1363),
.B(n_1365),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1485),
.B(n_1416),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1430),
.B(n_1363),
.Y(n_1525)
);

BUFx6f_ASAP7_75t_L g1526 ( 
.A(n_1503),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1485),
.B(n_1402),
.Y(n_1527)
);

OR2x2_ASAP7_75t_L g1528 ( 
.A(n_1431),
.B(n_1423),
.Y(n_1528)
);

A2O1A1Ixp33_ASAP7_75t_L g1529 ( 
.A1(n_1468),
.A2(n_1402),
.B(n_1322),
.C(n_1319),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1504),
.B(n_1420),
.Y(n_1530)
);

BUFx12f_ASAP7_75t_L g1531 ( 
.A(n_1478),
.Y(n_1531)
);

BUFx6f_ASAP7_75t_L g1532 ( 
.A(n_1503),
.Y(n_1532)
);

O2A1O1Ixp33_ASAP7_75t_L g1533 ( 
.A1(n_1455),
.A2(n_1398),
.B(n_1330),
.C(n_1407),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1431),
.B(n_1420),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1435),
.B(n_1319),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1496),
.B(n_1313),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1435),
.B(n_1330),
.Y(n_1537)
);

AO21x2_ASAP7_75t_L g1538 ( 
.A1(n_1450),
.A2(n_1355),
.B(n_1407),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1454),
.B(n_1313),
.Y(n_1539)
);

AO21x2_ASAP7_75t_L g1540 ( 
.A1(n_1450),
.A2(n_1355),
.B(n_1405),
.Y(n_1540)
);

INVxp67_ASAP7_75t_L g1541 ( 
.A(n_1457),
.Y(n_1541)
);

NOR2xp33_ASAP7_75t_L g1542 ( 
.A(n_1473),
.B(n_1405),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1454),
.B(n_1329),
.Y(n_1543)
);

OAI21xp5_ASAP7_75t_L g1544 ( 
.A1(n_1464),
.A2(n_1480),
.B(n_1468),
.Y(n_1544)
);

AO32x2_ASAP7_75t_L g1545 ( 
.A1(n_1449),
.A2(n_1505),
.A3(n_1507),
.B1(n_1428),
.B2(n_1482),
.Y(n_1545)
);

AND2x4_ASAP7_75t_L g1546 ( 
.A(n_1433),
.B(n_1434),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1458),
.B(n_1462),
.Y(n_1547)
);

OAI21xp5_ASAP7_75t_L g1548 ( 
.A1(n_1464),
.A2(n_1480),
.B(n_1436),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1458),
.B(n_1462),
.Y(n_1549)
);

AOI22xp5_ASAP7_75t_L g1550 ( 
.A1(n_1476),
.A2(n_1501),
.B1(n_1499),
.B2(n_1498),
.Y(n_1550)
);

OAI211xp5_ASAP7_75t_L g1551 ( 
.A1(n_1436),
.A2(n_1457),
.B(n_1492),
.C(n_1446),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1509),
.B(n_1490),
.Y(n_1552)
);

BUFx12f_ASAP7_75t_L g1553 ( 
.A(n_1444),
.Y(n_1553)
);

A2O1A1Ixp33_ASAP7_75t_L g1554 ( 
.A1(n_1498),
.A2(n_1492),
.B(n_1501),
.C(n_1483),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1451),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1508),
.B(n_1486),
.Y(n_1556)
);

OAI22xp5_ASAP7_75t_L g1557 ( 
.A1(n_1428),
.A2(n_1482),
.B1(n_1499),
.B2(n_1481),
.Y(n_1557)
);

AOI22xp5_ASAP7_75t_L g1558 ( 
.A1(n_1499),
.A2(n_1497),
.B1(n_1495),
.B2(n_1450),
.Y(n_1558)
);

AND2x4_ASAP7_75t_L g1559 ( 
.A(n_1434),
.B(n_1461),
.Y(n_1559)
);

O2A1O1Ixp33_ASAP7_75t_SL g1560 ( 
.A1(n_1470),
.A2(n_1491),
.B(n_1441),
.C(n_1475),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1465),
.B(n_1467),
.Y(n_1561)
);

AOI22x1_ASAP7_75t_SL g1562 ( 
.A1(n_1443),
.A2(n_1506),
.B1(n_1482),
.B2(n_1444),
.Y(n_1562)
);

AND2x4_ASAP7_75t_L g1563 ( 
.A(n_1434),
.B(n_1461),
.Y(n_1563)
);

OAI21xp5_ASAP7_75t_L g1564 ( 
.A1(n_1487),
.A2(n_1477),
.B(n_1475),
.Y(n_1564)
);

NOR2xp33_ASAP7_75t_L g1565 ( 
.A(n_1510),
.B(n_1470),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1439),
.B(n_1442),
.Y(n_1566)
);

OA21x2_ASAP7_75t_L g1567 ( 
.A1(n_1477),
.A2(n_1487),
.B(n_1481),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1510),
.B(n_1470),
.Y(n_1568)
);

O2A1O1Ixp33_ASAP7_75t_L g1569 ( 
.A1(n_1474),
.A2(n_1495),
.B(n_1497),
.C(n_1502),
.Y(n_1569)
);

AO32x2_ASAP7_75t_L g1570 ( 
.A1(n_1449),
.A2(n_1507),
.A3(n_1505),
.B1(n_1437),
.B2(n_1456),
.Y(n_1570)
);

OA21x2_ASAP7_75t_L g1571 ( 
.A1(n_1452),
.A2(n_1453),
.B(n_1489),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1556),
.B(n_1446),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1517),
.Y(n_1573)
);

BUFx2_ASAP7_75t_L g1574 ( 
.A(n_1545),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1555),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1570),
.B(n_1446),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1541),
.B(n_1469),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1541),
.B(n_1469),
.Y(n_1578)
);

INVxp67_ASAP7_75t_SL g1579 ( 
.A(n_1571),
.Y(n_1579)
);

HB1xp67_ASAP7_75t_L g1580 ( 
.A(n_1571),
.Y(n_1580)
);

AND2x4_ASAP7_75t_L g1581 ( 
.A(n_1559),
.B(n_1459),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1551),
.B(n_1471),
.Y(n_1582)
);

NAND3xp33_ASAP7_75t_L g1583 ( 
.A(n_1548),
.B(n_1516),
.C(n_1544),
.Y(n_1583)
);

OAI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1554),
.A2(n_1499),
.B1(n_1446),
.B2(n_1438),
.Y(n_1584)
);

INVxp67_ASAP7_75t_SL g1585 ( 
.A(n_1571),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1565),
.B(n_1568),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1565),
.B(n_1472),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1566),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1559),
.B(n_1459),
.Y(n_1589)
);

BUFx2_ASAP7_75t_L g1590 ( 
.A(n_1545),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1542),
.B(n_1440),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1547),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1550),
.A2(n_1500),
.B1(n_1456),
.B2(n_1463),
.Y(n_1593)
);

AOI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1554),
.A2(n_1438),
.B1(n_1460),
.B2(n_1448),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1549),
.B(n_1437),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1561),
.Y(n_1596)
);

INVx1_ASAP7_75t_SL g1597 ( 
.A(n_1514),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1542),
.B(n_1447),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1568),
.B(n_1472),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1552),
.B(n_1445),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1570),
.Y(n_1601)
);

AOI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1558),
.A2(n_1438),
.B1(n_1460),
.B2(n_1448),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1570),
.Y(n_1603)
);

AND2x4_ASAP7_75t_L g1604 ( 
.A(n_1563),
.B(n_1463),
.Y(n_1604)
);

BUFx3_ASAP7_75t_L g1605 ( 
.A(n_1526),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1576),
.Y(n_1606)
);

OR2x2_ASAP7_75t_L g1607 ( 
.A(n_1574),
.B(n_1567),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1574),
.B(n_1570),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1573),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1590),
.B(n_1545),
.Y(n_1610)
);

INVx3_ASAP7_75t_L g1611 ( 
.A(n_1581),
.Y(n_1611)
);

INVx2_ASAP7_75t_L g1612 ( 
.A(n_1576),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1576),
.Y(n_1613)
);

INVxp67_ASAP7_75t_SL g1614 ( 
.A(n_1580),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1590),
.B(n_1545),
.Y(n_1615)
);

OR2x6_ASAP7_75t_L g1616 ( 
.A(n_1584),
.B(n_1429),
.Y(n_1616)
);

NOR3xp33_ASAP7_75t_L g1617 ( 
.A(n_1583),
.B(n_1516),
.C(n_1519),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1580),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1573),
.Y(n_1619)
);

INVx4_ASAP7_75t_L g1620 ( 
.A(n_1605),
.Y(n_1620)
);

HB1xp67_ASAP7_75t_L g1621 ( 
.A(n_1601),
.Y(n_1621)
);

HB1xp67_ASAP7_75t_L g1622 ( 
.A(n_1601),
.Y(n_1622)
);

OAI221xp5_ASAP7_75t_L g1623 ( 
.A1(n_1583),
.A2(n_1521),
.B1(n_1569),
.B2(n_1529),
.C(n_1557),
.Y(n_1623)
);

NAND3xp33_ASAP7_75t_L g1624 ( 
.A(n_1582),
.B(n_1529),
.C(n_1564),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1575),
.Y(n_1625)
);

OAI21xp5_ASAP7_75t_SL g1626 ( 
.A1(n_1594),
.A2(n_1533),
.B(n_1521),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1577),
.B(n_1567),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1575),
.Y(n_1628)
);

HB1xp67_ASAP7_75t_L g1629 ( 
.A(n_1603),
.Y(n_1629)
);

AOI21xp5_ASAP7_75t_L g1630 ( 
.A1(n_1584),
.A2(n_1560),
.B(n_1579),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1577),
.B(n_1523),
.Y(n_1631)
);

HB1xp67_ASAP7_75t_L g1632 ( 
.A(n_1603),
.Y(n_1632)
);

AOI222xp33_ASAP7_75t_SL g1633 ( 
.A1(n_1597),
.A2(n_1447),
.B1(n_1562),
.B2(n_1553),
.C1(n_1531),
.C2(n_1537),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1588),
.B(n_1528),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1572),
.B(n_1523),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1572),
.B(n_1523),
.Y(n_1636)
);

AND2x4_ASAP7_75t_L g1637 ( 
.A(n_1581),
.B(n_1546),
.Y(n_1637)
);

HB1xp67_ASAP7_75t_L g1638 ( 
.A(n_1587),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1578),
.B(n_1534),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1638),
.B(n_1592),
.Y(n_1640)
);

NAND2x1_ASAP7_75t_L g1641 ( 
.A(n_1611),
.B(n_1604),
.Y(n_1641)
);

HB1xp67_ASAP7_75t_L g1642 ( 
.A(n_1634),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1638),
.B(n_1587),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1610),
.B(n_1597),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1639),
.B(n_1599),
.Y(n_1645)
);

NOR2x1_ASAP7_75t_L g1646 ( 
.A(n_1626),
.B(n_1513),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1610),
.B(n_1586),
.Y(n_1647)
);

INVx2_ASAP7_75t_SL g1648 ( 
.A(n_1634),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1606),
.B(n_1588),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1627),
.B(n_1592),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1610),
.B(n_1586),
.Y(n_1651)
);

INVx2_ASAP7_75t_SL g1652 ( 
.A(n_1634),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1615),
.B(n_1604),
.Y(n_1653)
);

INVxp67_ASAP7_75t_SL g1654 ( 
.A(n_1617),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1609),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1609),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1609),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1627),
.B(n_1596),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1615),
.B(n_1604),
.Y(n_1659)
);

INVx4_ASAP7_75t_L g1660 ( 
.A(n_1620),
.Y(n_1660)
);

NOR2xp67_ASAP7_75t_L g1661 ( 
.A(n_1630),
.B(n_1553),
.Y(n_1661)
);

AND2x4_ASAP7_75t_L g1662 ( 
.A(n_1611),
.B(n_1581),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1639),
.B(n_1599),
.Y(n_1663)
);

INVx2_ASAP7_75t_L g1664 ( 
.A(n_1618),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1606),
.B(n_1595),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1606),
.B(n_1595),
.Y(n_1666)
);

AND2x4_ASAP7_75t_L g1667 ( 
.A(n_1611),
.B(n_1604),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1619),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1619),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1618),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1615),
.B(n_1589),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1619),
.Y(n_1672)
);

NOR2x1_ASAP7_75t_L g1673 ( 
.A(n_1626),
.B(n_1513),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1625),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1618),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1606),
.B(n_1600),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1637),
.B(n_1589),
.Y(n_1677)
);

HB1xp67_ASAP7_75t_L g1678 ( 
.A(n_1625),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1654),
.B(n_1617),
.Y(n_1679)
);

AOI32xp33_ASAP7_75t_L g1680 ( 
.A1(n_1646),
.A2(n_1608),
.A3(n_1636),
.B1(n_1635),
.B2(n_1623),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1678),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1661),
.B(n_1608),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1661),
.B(n_1677),
.Y(n_1683)
);

INVxp67_ASAP7_75t_L g1684 ( 
.A(n_1646),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1655),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1677),
.B(n_1608),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1647),
.B(n_1608),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1655),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_L g1689 ( 
.A(n_1660),
.B(n_1531),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1647),
.B(n_1611),
.Y(n_1690)
);

HB1xp67_ASAP7_75t_L g1691 ( 
.A(n_1642),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1651),
.B(n_1624),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1651),
.B(n_1624),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1656),
.Y(n_1694)
);

NOR2x1_ASAP7_75t_L g1695 ( 
.A(n_1660),
.B(n_1620),
.Y(n_1695)
);

NAND2x1p5_ASAP7_75t_L g1696 ( 
.A(n_1673),
.B(n_1526),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1664),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1656),
.Y(n_1698)
);

AND2x4_ASAP7_75t_L g1699 ( 
.A(n_1660),
.B(n_1611),
.Y(n_1699)
);

AND2x4_ASAP7_75t_L g1700 ( 
.A(n_1660),
.B(n_1611),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1645),
.B(n_1607),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1657),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1657),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1664),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1648),
.B(n_1624),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_SL g1706 ( 
.A(n_1673),
.B(n_1526),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1668),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1664),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1653),
.B(n_1659),
.Y(n_1709)
);

NAND2xp67_ASAP7_75t_SL g1710 ( 
.A(n_1644),
.B(n_1520),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1648),
.B(n_1631),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1668),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1669),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1670),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1653),
.B(n_1659),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_R g1716 ( 
.A(n_1652),
.B(n_1536),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1669),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1672),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1672),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1670),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1674),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1690),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1679),
.B(n_1652),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1692),
.B(n_1663),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1709),
.B(n_1662),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_SL g1726 ( 
.A(n_1680),
.B(n_1630),
.Y(n_1726)
);

INVxp67_ASAP7_75t_L g1727 ( 
.A(n_1691),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1685),
.Y(n_1728)
);

AOI22xp5_ASAP7_75t_L g1729 ( 
.A1(n_1693),
.A2(n_1623),
.B1(n_1616),
.B2(n_1594),
.Y(n_1729)
);

NOR2x1_ASAP7_75t_L g1730 ( 
.A(n_1710),
.B(n_1641),
.Y(n_1730)
);

NOR2x1p5_ASAP7_75t_SL g1731 ( 
.A(n_1697),
.B(n_1670),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1687),
.B(n_1643),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1705),
.B(n_1644),
.Y(n_1733)
);

NAND4xp25_ASAP7_75t_L g1734 ( 
.A(n_1689),
.B(n_1522),
.C(n_1620),
.D(n_1535),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1709),
.B(n_1671),
.Y(n_1735)
);

NAND4xp75_ASAP7_75t_L g1736 ( 
.A(n_1682),
.B(n_1635),
.C(n_1636),
.D(n_1602),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1685),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1715),
.B(n_1671),
.Y(n_1738)
);

AND2x4_ASAP7_75t_L g1739 ( 
.A(n_1715),
.B(n_1683),
.Y(n_1739)
);

NOR2x1_ASAP7_75t_SL g1740 ( 
.A(n_1683),
.B(n_1506),
.Y(n_1740)
);

AO22x1_ASAP7_75t_L g1741 ( 
.A1(n_1684),
.A2(n_1614),
.B1(n_1598),
.B2(n_1526),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1681),
.B(n_1640),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1688),
.Y(n_1743)
);

NOR2xp67_ASAP7_75t_SL g1744 ( 
.A(n_1682),
.B(n_1532),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1681),
.B(n_1640),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1688),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1686),
.B(n_1662),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1694),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_L g1749 ( 
.A(n_1701),
.B(n_1591),
.Y(n_1749)
);

NAND2x1p5_ASAP7_75t_L g1750 ( 
.A(n_1695),
.B(n_1532),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1694),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_L g1752 ( 
.A(n_1701),
.B(n_1525),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1686),
.B(n_1631),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1711),
.B(n_1650),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1698),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1690),
.B(n_1650),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1698),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1702),
.B(n_1658),
.Y(n_1758)
);

INVx1_ASAP7_75t_SL g1759 ( 
.A(n_1723),
.Y(n_1759)
);

OAI22xp33_ASAP7_75t_SL g1760 ( 
.A1(n_1726),
.A2(n_1710),
.B1(n_1706),
.B2(n_1607),
.Y(n_1760)
);

NAND2xp5_ASAP7_75t_L g1761 ( 
.A(n_1749),
.B(n_1612),
.Y(n_1761)
);

NAND3xp33_ASAP7_75t_L g1762 ( 
.A(n_1726),
.B(n_1729),
.C(n_1727),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1749),
.B(n_1703),
.Y(n_1763)
);

OAI322xp33_ASAP7_75t_L g1764 ( 
.A1(n_1727),
.A2(n_1607),
.A3(n_1614),
.B1(n_1696),
.B2(n_1721),
.C1(n_1717),
.C2(n_1718),
.Y(n_1764)
);

AOI22xp33_ASAP7_75t_L g1765 ( 
.A1(n_1733),
.A2(n_1616),
.B1(n_1636),
.B2(n_1635),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1728),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1737),
.Y(n_1767)
);

OAI221xp5_ASAP7_75t_L g1768 ( 
.A1(n_1730),
.A2(n_1696),
.B1(n_1616),
.B2(n_1585),
.C(n_1582),
.Y(n_1768)
);

OAI21xp33_ASAP7_75t_SL g1769 ( 
.A1(n_1736),
.A2(n_1712),
.B(n_1707),
.Y(n_1769)
);

AND2x4_ASAP7_75t_L g1770 ( 
.A(n_1739),
.B(n_1699),
.Y(n_1770)
);

A2O1A1Ixp33_ASAP7_75t_L g1771 ( 
.A1(n_1731),
.A2(n_1613),
.B(n_1612),
.C(n_1585),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1743),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1746),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1724),
.B(n_1707),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1748),
.Y(n_1775)
);

NAND4xp25_ASAP7_75t_L g1776 ( 
.A(n_1739),
.B(n_1699),
.C(n_1700),
.D(n_1719),
.Y(n_1776)
);

NAND2xp5_ASAP7_75t_SL g1777 ( 
.A(n_1739),
.B(n_1696),
.Y(n_1777)
);

AOI222xp33_ASAP7_75t_L g1778 ( 
.A1(n_1752),
.A2(n_1593),
.B1(n_1629),
.B2(n_1622),
.C1(n_1621),
.C2(n_1632),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1751),
.Y(n_1779)
);

AOI322xp5_ASAP7_75t_L g1780 ( 
.A1(n_1752),
.A2(n_1613),
.A3(n_1612),
.B1(n_1632),
.B2(n_1629),
.C1(n_1622),
.C2(n_1621),
.Y(n_1780)
);

OAI222xp33_ASAP7_75t_L g1781 ( 
.A1(n_1753),
.A2(n_1616),
.B1(n_1602),
.B2(n_1612),
.C1(n_1613),
.C2(n_1704),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1747),
.Y(n_1782)
);

OAI21xp33_ASAP7_75t_L g1783 ( 
.A1(n_1754),
.A2(n_1716),
.B(n_1713),
.Y(n_1783)
);

OAI21xp33_ASAP7_75t_L g1784 ( 
.A1(n_1756),
.A2(n_1716),
.B(n_1713),
.Y(n_1784)
);

INVxp67_ASAP7_75t_SL g1785 ( 
.A(n_1760),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1766),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1770),
.Y(n_1787)
);

OAI211xp5_ASAP7_75t_L g1788 ( 
.A1(n_1769),
.A2(n_1722),
.B(n_1745),
.C(n_1742),
.Y(n_1788)
);

NAND3xp33_ASAP7_75t_L g1789 ( 
.A(n_1762),
.B(n_1757),
.C(n_1755),
.Y(n_1789)
);

A2O1A1Ixp33_ASAP7_75t_SL g1790 ( 
.A1(n_1768),
.A2(n_1773),
.B(n_1775),
.C(n_1767),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1763),
.B(n_1732),
.Y(n_1791)
);

AOI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1778),
.A2(n_1616),
.B1(n_1633),
.B2(n_1538),
.Y(n_1792)
);

A2O1A1Ixp33_ASAP7_75t_L g1793 ( 
.A1(n_1783),
.A2(n_1758),
.B(n_1613),
.C(n_1744),
.Y(n_1793)
);

INVxp67_ASAP7_75t_SL g1794 ( 
.A(n_1763),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1759),
.B(n_1722),
.Y(n_1795)
);

HB1xp67_ASAP7_75t_L g1796 ( 
.A(n_1782),
.Y(n_1796)
);

NOR4xp25_ASAP7_75t_SL g1797 ( 
.A(n_1777),
.B(n_1741),
.C(n_1740),
.D(n_1712),
.Y(n_1797)
);

INVxp67_ASAP7_75t_SL g1798 ( 
.A(n_1774),
.Y(n_1798)
);

OR2x2_ASAP7_75t_L g1799 ( 
.A(n_1774),
.B(n_1735),
.Y(n_1799)
);

NOR2xp33_ASAP7_75t_L g1800 ( 
.A(n_1776),
.B(n_1734),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1772),
.B(n_1738),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1770),
.B(n_1725),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1779),
.B(n_1747),
.Y(n_1803)
);

INVxp67_ASAP7_75t_L g1804 ( 
.A(n_1761),
.Y(n_1804)
);

AO22x2_ASAP7_75t_L g1805 ( 
.A1(n_1785),
.A2(n_1794),
.B1(n_1798),
.B2(n_1789),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1796),
.Y(n_1806)
);

OAI21xp5_ASAP7_75t_L g1807 ( 
.A1(n_1785),
.A2(n_1780),
.B(n_1784),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1795),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1798),
.B(n_1725),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1799),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1791),
.Y(n_1811)
);

OAI322xp33_ASAP7_75t_L g1812 ( 
.A1(n_1800),
.A2(n_1804),
.A3(n_1786),
.B1(n_1792),
.B2(n_1801),
.C1(n_1803),
.C2(n_1787),
.Y(n_1812)
);

OAI221xp5_ASAP7_75t_SL g1813 ( 
.A1(n_1788),
.A2(n_1765),
.B1(n_1771),
.B2(n_1764),
.C(n_1616),
.Y(n_1813)
);

INVx2_ASAP7_75t_L g1814 ( 
.A(n_1802),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1804),
.B(n_1658),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1793),
.Y(n_1816)
);

AOI221xp5_ASAP7_75t_L g1817 ( 
.A1(n_1805),
.A2(n_1790),
.B1(n_1781),
.B2(n_1714),
.C(n_1697),
.Y(n_1817)
);

NAND4xp25_ASAP7_75t_L g1818 ( 
.A(n_1807),
.B(n_1797),
.C(n_1699),
.D(n_1700),
.Y(n_1818)
);

NOR2xp33_ASAP7_75t_L g1819 ( 
.A(n_1809),
.B(n_1700),
.Y(n_1819)
);

NOR3xp33_ASAP7_75t_L g1820 ( 
.A(n_1812),
.B(n_1708),
.C(n_1704),
.Y(n_1820)
);

OAI211xp5_ASAP7_75t_L g1821 ( 
.A1(n_1816),
.A2(n_1641),
.B(n_1620),
.C(n_1718),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1805),
.Y(n_1822)
);

NOR2x1_ASAP7_75t_L g1823 ( 
.A(n_1806),
.B(n_1717),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1808),
.Y(n_1824)
);

OAI211xp5_ASAP7_75t_L g1825 ( 
.A1(n_1811),
.A2(n_1620),
.B(n_1721),
.C(n_1719),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1814),
.B(n_1667),
.Y(n_1826)
);

NOR2x1_ASAP7_75t_L g1827 ( 
.A(n_1810),
.B(n_1675),
.Y(n_1827)
);

O2A1O1Ixp5_ASAP7_75t_SL g1828 ( 
.A1(n_1822),
.A2(n_1815),
.B(n_1812),
.C(n_1813),
.Y(n_1828)
);

AOI221x1_ASAP7_75t_L g1829 ( 
.A1(n_1820),
.A2(n_1720),
.B1(n_1714),
.B2(n_1708),
.C(n_1675),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1824),
.B(n_1720),
.Y(n_1830)
);

O2A1O1Ixp33_ASAP7_75t_L g1831 ( 
.A1(n_1817),
.A2(n_1675),
.B(n_1618),
.C(n_1616),
.Y(n_1831)
);

OAI22xp5_ASAP7_75t_L g1832 ( 
.A1(n_1819),
.A2(n_1750),
.B1(n_1649),
.B2(n_1674),
.Y(n_1832)
);

NAND2x1p5_ASAP7_75t_L g1833 ( 
.A(n_1826),
.B(n_1488),
.Y(n_1833)
);

OAI22xp33_ASAP7_75t_R g1834 ( 
.A1(n_1828),
.A2(n_1818),
.B1(n_1823),
.B2(n_1821),
.Y(n_1834)
);

BUFx8_ASAP7_75t_SL g1835 ( 
.A(n_1830),
.Y(n_1835)
);

AOI21xp5_ASAP7_75t_L g1836 ( 
.A1(n_1831),
.A2(n_1827),
.B(n_1825),
.Y(n_1836)
);

O2A1O1Ixp33_ASAP7_75t_L g1837 ( 
.A1(n_1833),
.A2(n_1750),
.B(n_1616),
.C(n_1543),
.Y(n_1837)
);

NAND3xp33_ASAP7_75t_SL g1838 ( 
.A(n_1832),
.B(n_1633),
.C(n_1539),
.Y(n_1838)
);

OAI211xp5_ASAP7_75t_L g1839 ( 
.A1(n_1829),
.A2(n_1493),
.B(n_1620),
.C(n_1532),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1835),
.Y(n_1840)
);

NAND4xp75_ASAP7_75t_L g1841 ( 
.A(n_1836),
.B(n_1524),
.C(n_1527),
.D(n_1530),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1839),
.B(n_1837),
.Y(n_1842)
);

XNOR2xp5_ASAP7_75t_L g1843 ( 
.A(n_1838),
.B(n_1488),
.Y(n_1843)
);

NOR2x1_ASAP7_75t_L g1844 ( 
.A(n_1834),
.B(n_1667),
.Y(n_1844)
);

OR3x1_ASAP7_75t_L g1845 ( 
.A(n_1840),
.B(n_1628),
.C(n_1625),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1844),
.Y(n_1846)
);

OR2x2_ASAP7_75t_L g1847 ( 
.A(n_1841),
.B(n_1649),
.Y(n_1847)
);

OA22x2_ASAP7_75t_L g1848 ( 
.A1(n_1846),
.A2(n_1843),
.B1(n_1842),
.B2(n_1845),
.Y(n_1848)
);

BUFx6f_ASAP7_75t_L g1849 ( 
.A(n_1848),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1849),
.Y(n_1850)
);

AO22x1_ASAP7_75t_L g1851 ( 
.A1(n_1849),
.A2(n_1847),
.B1(n_1532),
.B2(n_1667),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1850),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1851),
.Y(n_1853)
);

AOI22xp33_ASAP7_75t_L g1854 ( 
.A1(n_1853),
.A2(n_1849),
.B1(n_1493),
.B2(n_1540),
.Y(n_1854)
);

OAI21xp5_ASAP7_75t_SL g1855 ( 
.A1(n_1852),
.A2(n_1512),
.B(n_1518),
.Y(n_1855)
);

AOI21xp5_ASAP7_75t_L g1856 ( 
.A1(n_1854),
.A2(n_1855),
.B(n_1493),
.Y(n_1856)
);

AO21x2_ASAP7_75t_L g1857 ( 
.A1(n_1856),
.A2(n_1666),
.B(n_1665),
.Y(n_1857)
);

INVx2_ASAP7_75t_L g1858 ( 
.A(n_1857),
.Y(n_1858)
);

OAI221xp5_ASAP7_75t_R g1859 ( 
.A1(n_1858),
.A2(n_1493),
.B1(n_1667),
.B2(n_1662),
.C(n_1676),
.Y(n_1859)
);

AOI211xp5_ASAP7_75t_L g1860 ( 
.A1(n_1859),
.A2(n_1493),
.B(n_1560),
.C(n_1515),
.Y(n_1860)
);


endmodule