module fake_aes_9371_n_647 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_647);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_647;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_446;
wire n_420;
wire n_423;
wire n_342;
wire n_165;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_570;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g78 ( .A(n_9), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_25), .Y(n_79) );
CKINVDCx16_ASAP7_75t_R g80 ( .A(n_23), .Y(n_80) );
CKINVDCx20_ASAP7_75t_R g81 ( .A(n_27), .Y(n_81) );
NOR2xp67_ASAP7_75t_L g82 ( .A(n_53), .B(n_2), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_8), .Y(n_83) );
INVxp67_ASAP7_75t_SL g84 ( .A(n_65), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_6), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_74), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_48), .Y(n_87) );
BUFx3_ASAP7_75t_L g88 ( .A(n_64), .Y(n_88) );
CKINVDCx14_ASAP7_75t_R g89 ( .A(n_59), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_46), .Y(n_90) );
INVxp33_ASAP7_75t_L g91 ( .A(n_10), .Y(n_91) );
CKINVDCx14_ASAP7_75t_R g92 ( .A(n_8), .Y(n_92) );
INVxp33_ASAP7_75t_SL g93 ( .A(n_33), .Y(n_93) );
INVx2_ASAP7_75t_SL g94 ( .A(n_60), .Y(n_94) );
BUFx6f_ASAP7_75t_L g95 ( .A(n_28), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_24), .Y(n_96) );
INVxp67_ASAP7_75t_L g97 ( .A(n_52), .Y(n_97) );
CKINVDCx16_ASAP7_75t_R g98 ( .A(n_72), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_35), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_55), .Y(n_100) );
BUFx6f_ASAP7_75t_L g101 ( .A(n_67), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_68), .Y(n_102) );
HB1xp67_ASAP7_75t_L g103 ( .A(n_6), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_47), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_20), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_29), .Y(n_106) );
CKINVDCx14_ASAP7_75t_R g107 ( .A(n_45), .Y(n_107) );
BUFx5_ASAP7_75t_L g108 ( .A(n_73), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_18), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_62), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_38), .Y(n_111) );
INVxp33_ASAP7_75t_SL g112 ( .A(n_77), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_63), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_2), .Y(n_114) );
INVxp33_ASAP7_75t_SL g115 ( .A(n_40), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_17), .Y(n_116) );
AND2x4_ASAP7_75t_L g117 ( .A(n_94), .B(n_0), .Y(n_117) );
INVx3_ASAP7_75t_L g118 ( .A(n_99), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_108), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_79), .Y(n_120) );
INVx2_ASAP7_75t_SL g121 ( .A(n_88), .Y(n_121) );
INVx3_ASAP7_75t_L g122 ( .A(n_99), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_87), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_91), .B(n_0), .Y(n_124) );
HB1xp67_ASAP7_75t_L g125 ( .A(n_92), .Y(n_125) );
OA21x2_ASAP7_75t_L g126 ( .A1(n_96), .A2(n_34), .B(n_75), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_100), .Y(n_127) );
AND2x4_ASAP7_75t_L g128 ( .A(n_88), .B(n_116), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_102), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_104), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_108), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_95), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_80), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_95), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_106), .Y(n_135) );
AND2x2_ASAP7_75t_L g136 ( .A(n_91), .B(n_1), .Y(n_136) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_95), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_110), .Y(n_138) );
AND2x4_ASAP7_75t_L g139 ( .A(n_78), .B(n_1), .Y(n_139) );
NOR2xp33_ASAP7_75t_L g140 ( .A(n_113), .B(n_3), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_83), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_95), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_85), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_114), .Y(n_144) );
AND2x2_ASAP7_75t_L g145 ( .A(n_92), .B(n_3), .Y(n_145) );
AND2x2_ASAP7_75t_L g146 ( .A(n_89), .B(n_107), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_84), .Y(n_147) );
HB1xp67_ASAP7_75t_L g148 ( .A(n_103), .Y(n_148) );
HB1xp67_ASAP7_75t_L g149 ( .A(n_98), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_128), .B(n_108), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_132), .Y(n_151) );
HB1xp67_ASAP7_75t_L g152 ( .A(n_125), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_132), .Y(n_153) );
INVx4_ASAP7_75t_L g154 ( .A(n_117), .Y(n_154) );
AND2x6_ASAP7_75t_L g155 ( .A(n_145), .B(n_101), .Y(n_155) );
AND2x2_ASAP7_75t_SL g156 ( .A(n_139), .B(n_101), .Y(n_156) );
AND2x4_ASAP7_75t_L g157 ( .A(n_128), .B(n_82), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_132), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_128), .B(n_108), .Y(n_159) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_125), .B(n_97), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_119), .Y(n_161) );
INVx6_ASAP7_75t_L g162 ( .A(n_128), .Y(n_162) );
INVx2_ASAP7_75t_SL g163 ( .A(n_121), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_132), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_132), .Y(n_165) );
INVx3_ASAP7_75t_L g166 ( .A(n_139), .Y(n_166) );
INVx1_ASAP7_75t_SL g167 ( .A(n_149), .Y(n_167) );
INVx2_ASAP7_75t_SL g168 ( .A(n_121), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_132), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g170 ( .A(n_146), .B(n_93), .Y(n_170) );
BUFx3_ASAP7_75t_L g171 ( .A(n_117), .Y(n_171) );
AND2x2_ASAP7_75t_SL g172 ( .A(n_139), .B(n_101), .Y(n_172) );
INVxp67_ASAP7_75t_SL g173 ( .A(n_148), .Y(n_173) );
INVxp67_ASAP7_75t_L g174 ( .A(n_148), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_132), .Y(n_175) );
AO22x2_ASAP7_75t_L g176 ( .A1(n_139), .A2(n_93), .B1(n_81), .B2(n_111), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_119), .Y(n_177) );
BUFx3_ASAP7_75t_L g178 ( .A(n_117), .Y(n_178) );
BUFx3_ASAP7_75t_L g179 ( .A(n_117), .Y(n_179) );
INVx3_ASAP7_75t_L g180 ( .A(n_118), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_119), .Y(n_181) );
AO22x2_ASAP7_75t_L g182 ( .A1(n_145), .A2(n_81), .B1(n_105), .B2(n_111), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_131), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_131), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_131), .Y(n_185) );
AND2x4_ASAP7_75t_L g186 ( .A(n_147), .B(n_101), .Y(n_186) );
INVx4_ASAP7_75t_L g187 ( .A(n_126), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_134), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_156), .B(n_146), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_170), .B(n_147), .Y(n_190) );
INVx3_ASAP7_75t_L g191 ( .A(n_162), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_174), .B(n_149), .Y(n_192) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_171), .Y(n_193) );
AND2x4_ASAP7_75t_L g194 ( .A(n_173), .B(n_136), .Y(n_194) );
NAND2x1p5_ASAP7_75t_L g195 ( .A(n_167), .B(n_145), .Y(n_195) );
NAND3xp33_ASAP7_75t_SL g196 ( .A(n_167), .B(n_133), .C(n_105), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g197 ( .A(n_156), .B(n_136), .Y(n_197) );
NOR2xp33_ASAP7_75t_SL g198 ( .A(n_174), .B(n_136), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_173), .B(n_124), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_162), .Y(n_200) );
HB1xp67_ASAP7_75t_L g201 ( .A(n_152), .Y(n_201) );
INVx1_ASAP7_75t_SL g202 ( .A(n_155), .Y(n_202) );
AND2x6_ASAP7_75t_L g203 ( .A(n_171), .B(n_178), .Y(n_203) );
NOR2xp33_ASAP7_75t_R g204 ( .A(n_156), .B(n_172), .Y(n_204) );
INVx2_ASAP7_75t_SL g205 ( .A(n_155), .Y(n_205) );
AO21x2_ASAP7_75t_L g206 ( .A1(n_150), .A2(n_124), .B(n_120), .Y(n_206) );
OAI21xp5_ASAP7_75t_L g207 ( .A1(n_187), .A2(n_126), .B(n_120), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_160), .B(n_123), .Y(n_208) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_172), .B(n_112), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_162), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_163), .Y(n_211) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_162), .B(n_123), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_157), .B(n_127), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_157), .B(n_127), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_162), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_157), .B(n_130), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_172), .B(n_138), .Y(n_217) );
AOI22xp5_ASAP7_75t_L g218 ( .A1(n_176), .A2(n_140), .B1(n_129), .B2(n_130), .Y(n_218) );
AOI22xp33_ASAP7_75t_SL g219 ( .A1(n_182), .A2(n_176), .B1(n_155), .B2(n_154), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_157), .B(n_138), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_163), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g222 ( .A(n_154), .B(n_129), .Y(n_222) );
OAI22xp5_ASAP7_75t_SL g223 ( .A1(n_182), .A2(n_144), .B1(n_143), .B2(n_141), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_154), .B(n_135), .Y(n_224) );
INVx2_ASAP7_75t_SL g225 ( .A(n_155), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_186), .Y(n_226) );
HB1xp67_ASAP7_75t_L g227 ( .A(n_155), .Y(n_227) );
NAND3xp33_ASAP7_75t_L g228 ( .A(n_187), .B(n_135), .C(n_126), .Y(n_228) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_171), .Y(n_229) );
CKINVDCx5p33_ASAP7_75t_R g230 ( .A(n_155), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_154), .B(n_144), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_186), .Y(n_232) );
AOI22xp33_ASAP7_75t_L g233 ( .A1(n_166), .A2(n_143), .B1(n_141), .B2(n_118), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_186), .Y(n_234) );
BUFx2_ASAP7_75t_L g235 ( .A(n_176), .Y(n_235) );
AND2x4_ASAP7_75t_L g236 ( .A(n_178), .B(n_121), .Y(n_236) );
NOR2x1p5_ASAP7_75t_L g237 ( .A(n_182), .B(n_122), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_166), .B(n_115), .Y(n_238) );
INVx2_ASAP7_75t_SL g239 ( .A(n_201), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_222), .A2(n_166), .B(n_187), .Y(n_240) );
INVx3_ASAP7_75t_L g241 ( .A(n_193), .Y(n_241) );
INVx3_ASAP7_75t_L g242 ( .A(n_193), .Y(n_242) );
A2O1A1Ixp33_ASAP7_75t_SL g243 ( .A1(n_238), .A2(n_166), .B(n_107), .C(n_89), .Y(n_243) );
INVx5_ASAP7_75t_L g244 ( .A(n_203), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_231), .Y(n_245) );
BUFx3_ASAP7_75t_L g246 ( .A(n_203), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_222), .A2(n_187), .B(n_178), .Y(n_247) );
AOI22xp5_ASAP7_75t_L g248 ( .A1(n_198), .A2(n_176), .B1(n_182), .B2(n_155), .Y(n_248) );
O2A1O1Ixp33_ASAP7_75t_SL g249 ( .A1(n_207), .A2(n_168), .B(n_163), .C(n_150), .Y(n_249) );
NOR2xp33_ASAP7_75t_SL g250 ( .A(n_201), .B(n_155), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_192), .B(n_179), .Y(n_251) );
INVx4_ASAP7_75t_L g252 ( .A(n_203), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_224), .Y(n_253) );
INVx3_ASAP7_75t_L g254 ( .A(n_193), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_226), .Y(n_255) );
INVx3_ASAP7_75t_L g256 ( .A(n_193), .Y(n_256) );
BUFx2_ASAP7_75t_L g257 ( .A(n_195), .Y(n_257) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_229), .Y(n_258) );
AND2x4_ASAP7_75t_L g259 ( .A(n_194), .B(n_186), .Y(n_259) );
BUFx3_ASAP7_75t_L g260 ( .A(n_203), .Y(n_260) );
BUFx3_ASAP7_75t_L g261 ( .A(n_203), .Y(n_261) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_195), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_199), .B(n_179), .Y(n_263) );
OR2x6_ASAP7_75t_L g264 ( .A(n_237), .B(n_182), .Y(n_264) );
AND2x4_ASAP7_75t_L g265 ( .A(n_194), .B(n_179), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_228), .A2(n_159), .B(n_168), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_238), .A2(n_159), .B(n_168), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_232), .Y(n_268) );
NAND2xp5_ASAP7_75t_SL g269 ( .A(n_229), .B(n_161), .Y(n_269) );
AO22x1_ASAP7_75t_L g270 ( .A1(n_235), .A2(n_176), .B1(n_90), .B2(n_109), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_229), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_229), .Y(n_272) );
OAI221xp5_ASAP7_75t_L g273 ( .A1(n_218), .A2(n_180), .B1(n_185), .B2(n_184), .C(n_183), .Y(n_273) );
INVxp67_ASAP7_75t_L g274 ( .A(n_196), .Y(n_274) );
BUFx2_ASAP7_75t_L g275 ( .A(n_204), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_234), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_200), .Y(n_277) );
OAI22xp5_ASAP7_75t_L g278 ( .A1(n_197), .A2(n_219), .B1(n_217), .B2(n_208), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_210), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_215), .Y(n_280) );
INVx2_ASAP7_75t_SL g281 ( .A(n_213), .Y(n_281) );
BUFx2_ASAP7_75t_L g282 ( .A(n_204), .Y(n_282) );
CKINVDCx14_ASAP7_75t_R g283 ( .A(n_223), .Y(n_283) );
A2O1A1Ixp33_ASAP7_75t_L g284 ( .A1(n_190), .A2(n_180), .B(n_122), .C(n_118), .Y(n_284) );
NAND2xp5_ASAP7_75t_SL g285 ( .A(n_211), .B(n_161), .Y(n_285) );
NAND2x1_ASAP7_75t_L g286 ( .A(n_252), .B(n_205), .Y(n_286) );
OAI21x1_ASAP7_75t_L g287 ( .A1(n_266), .A2(n_267), .B(n_240), .Y(n_287) );
OAI21x1_ASAP7_75t_L g288 ( .A1(n_247), .A2(n_126), .B(n_221), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_245), .B(n_206), .Y(n_289) );
NAND2x1p5_ASAP7_75t_L g290 ( .A(n_252), .B(n_225), .Y(n_290) );
AOI21xp5_ASAP7_75t_L g291 ( .A1(n_249), .A2(n_217), .B(n_214), .Y(n_291) );
AO32x2_ASAP7_75t_L g292 ( .A1(n_278), .A2(n_206), .A3(n_126), .B1(n_118), .B2(n_122), .Y(n_292) );
NOR2xp33_ASAP7_75t_L g293 ( .A(n_239), .B(n_190), .Y(n_293) );
OR2x2_ASAP7_75t_L g294 ( .A(n_257), .B(n_216), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_281), .B(n_220), .Y(n_295) );
AOI22xp5_ASAP7_75t_L g296 ( .A1(n_248), .A2(n_197), .B1(n_189), .B2(n_209), .Y(n_296) );
AOI22xp33_ASAP7_75t_L g297 ( .A1(n_264), .A2(n_189), .B1(n_191), .B2(n_236), .Y(n_297) );
OAI21x1_ASAP7_75t_L g298 ( .A1(n_241), .A2(n_233), .B(n_122), .Y(n_298) );
AOI22xp33_ASAP7_75t_L g299 ( .A1(n_264), .A2(n_191), .B1(n_236), .B2(n_212), .Y(n_299) );
OAI21x1_ASAP7_75t_L g300 ( .A1(n_241), .A2(n_233), .B(n_180), .Y(n_300) );
OAI22x1_ASAP7_75t_L g301 ( .A1(n_274), .A2(n_230), .B1(n_227), .B2(n_180), .Y(n_301) );
INVx3_ASAP7_75t_L g302 ( .A(n_252), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_258), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_265), .B(n_212), .Y(n_304) );
BUFx2_ASAP7_75t_L g305 ( .A(n_246), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_265), .B(n_227), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_259), .Y(n_307) );
OAI21x1_ASAP7_75t_L g308 ( .A1(n_241), .A2(n_177), .B(n_181), .Y(n_308) );
AOI21xp33_ASAP7_75t_L g309 ( .A1(n_251), .A2(n_202), .B(n_185), .Y(n_309) );
AO21x2_ASAP7_75t_L g310 ( .A1(n_249), .A2(n_177), .B(n_184), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_258), .Y(n_311) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_262), .Y(n_312) );
AOI21xp33_ASAP7_75t_SL g313 ( .A1(n_264), .A2(n_4), .B(n_5), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g314 ( .A1(n_285), .A2(n_181), .B(n_183), .Y(n_314) );
OAI221xp5_ASAP7_75t_L g315 ( .A1(n_264), .A2(n_263), .B1(n_253), .B2(n_284), .C(n_273), .Y(n_315) );
OAI21x1_ASAP7_75t_L g316 ( .A1(n_242), .A2(n_188), .B(n_175), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_265), .B(n_86), .Y(n_317) );
OAI21x1_ASAP7_75t_L g318 ( .A1(n_242), .A2(n_188), .B(n_175), .Y(n_318) );
OAI21x1_ASAP7_75t_SL g319 ( .A1(n_271), .A2(n_108), .B(n_5), .Y(n_319) );
AOI21xp5_ASAP7_75t_L g320 ( .A1(n_310), .A2(n_243), .B(n_269), .Y(n_320) );
BUFx4f_ASAP7_75t_SL g321 ( .A(n_294), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_293), .B(n_259), .Y(n_322) );
INVx3_ASAP7_75t_L g323 ( .A(n_302), .Y(n_323) );
A2O1A1Ixp33_ASAP7_75t_L g324 ( .A1(n_289), .A2(n_284), .B(n_283), .C(n_255), .Y(n_324) );
AOI21xp33_ASAP7_75t_L g325 ( .A1(n_315), .A2(n_243), .B(n_250), .Y(n_325) );
BUFx2_ASAP7_75t_L g326 ( .A(n_312), .Y(n_326) );
AOI22xp33_ASAP7_75t_SL g327 ( .A1(n_319), .A2(n_283), .B1(n_275), .B2(n_282), .Y(n_327) );
INVx4_ASAP7_75t_L g328 ( .A(n_305), .Y(n_328) );
BUFx8_ASAP7_75t_L g329 ( .A(n_307), .Y(n_329) );
AO221x2_ASAP7_75t_L g330 ( .A1(n_301), .A2(n_270), .B1(n_7), .B2(n_9), .C(n_10), .Y(n_330) );
OAI21x1_ASAP7_75t_L g331 ( .A1(n_287), .A2(n_256), .B(n_254), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_308), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_295), .Y(n_333) );
AOI22xp5_ASAP7_75t_L g334 ( .A1(n_299), .A2(n_259), .B1(n_268), .B2(n_276), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_308), .Y(n_335) );
NOR2x1_ASAP7_75t_SL g336 ( .A(n_289), .B(n_244), .Y(n_336) );
OAI21xp33_ASAP7_75t_L g337 ( .A1(n_313), .A2(n_280), .B(n_279), .Y(n_337) );
OAI221xp5_ASAP7_75t_L g338 ( .A1(n_297), .A2(n_277), .B1(n_279), .B2(n_246), .C(n_260), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_294), .B(n_260), .Y(n_339) );
AOI22xp33_ASAP7_75t_L g340 ( .A1(n_296), .A2(n_277), .B1(n_261), .B2(n_244), .Y(n_340) );
OAI22xp5_ASAP7_75t_L g341 ( .A1(n_304), .A2(n_244), .B1(n_261), .B2(n_258), .Y(n_341) );
OR2x6_ASAP7_75t_L g342 ( .A(n_305), .B(n_258), .Y(n_342) );
INVx3_ASAP7_75t_L g343 ( .A(n_302), .Y(n_343) );
OAI22xp5_ASAP7_75t_L g344 ( .A1(n_306), .A2(n_244), .B1(n_256), .B2(n_242), .Y(n_344) );
OAI211xp5_ASAP7_75t_SL g345 ( .A1(n_317), .A2(n_269), .B(n_285), .C(n_256), .Y(n_345) );
AOI22xp33_ASAP7_75t_SL g346 ( .A1(n_319), .A2(n_244), .B1(n_254), .B2(n_108), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_300), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_332), .Y(n_348) );
OAI211xp5_ASAP7_75t_L g349 ( .A1(n_327), .A2(n_291), .B(n_309), .C(n_314), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_332), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_335), .Y(n_351) );
AOI31xp33_ASAP7_75t_L g352 ( .A1(n_333), .A2(n_290), .A3(n_303), .B(n_311), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_335), .Y(n_353) );
AND2x4_ASAP7_75t_L g354 ( .A(n_336), .B(n_303), .Y(n_354) );
INVx3_ASAP7_75t_L g355 ( .A(n_342), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_330), .B(n_292), .Y(n_356) );
OR2x2_ASAP7_75t_L g357 ( .A(n_326), .B(n_310), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_347), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_347), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_331), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_330), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_330), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_342), .Y(n_363) );
BUFx2_ASAP7_75t_L g364 ( .A(n_328), .Y(n_364) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_321), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_321), .B(n_301), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_342), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_323), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_323), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_324), .B(n_292), .Y(n_370) );
INVxp67_ASAP7_75t_L g371 ( .A(n_339), .Y(n_371) );
INVxp67_ASAP7_75t_L g372 ( .A(n_339), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_343), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_343), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_324), .B(n_292), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_328), .Y(n_376) );
BUFx3_ASAP7_75t_L g377 ( .A(n_329), .Y(n_377) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_364), .Y(n_378) );
AOI21xp5_ASAP7_75t_L g379 ( .A1(n_352), .A2(n_320), .B(n_325), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_356), .B(n_292), .Y(n_380) );
OAI31xp33_ASAP7_75t_L g381 ( .A1(n_361), .A2(n_337), .A3(n_322), .B(n_345), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_348), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_356), .B(n_292), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_348), .Y(n_384) );
NAND2xp5_ASAP7_75t_SL g385 ( .A(n_364), .B(n_346), .Y(n_385) );
INVx2_ASAP7_75t_SL g386 ( .A(n_377), .Y(n_386) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_376), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_348), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_371), .B(n_334), .Y(n_389) );
OR2x2_ASAP7_75t_L g390 ( .A(n_357), .B(n_310), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_350), .Y(n_391) );
AOI31xp33_ASAP7_75t_L g392 ( .A1(n_361), .A2(n_340), .A3(n_341), .B(n_344), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_370), .B(n_300), .Y(n_393) );
OAI31xp33_ASAP7_75t_L g394 ( .A1(n_362), .A2(n_338), .A3(n_340), .B(n_302), .Y(n_394) );
AO21x2_ASAP7_75t_L g395 ( .A1(n_360), .A2(n_288), .B(n_298), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_372), .B(n_329), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_370), .B(n_108), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_362), .B(n_298), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_375), .B(n_311), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_377), .A2(n_329), .B1(n_287), .B2(n_254), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_350), .Y(n_401) );
AND2x6_ASAP7_75t_SL g402 ( .A(n_366), .B(n_4), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_365), .B(n_7), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_351), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_351), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_353), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_353), .Y(n_407) );
AND2x2_ASAP7_75t_SL g408 ( .A(n_375), .B(n_271), .Y(n_408) );
OR2x2_ASAP7_75t_L g409 ( .A(n_357), .B(n_11), .Y(n_409) );
OAI22xp5_ASAP7_75t_L g410 ( .A1(n_377), .A2(n_272), .B1(n_290), .B2(n_286), .Y(n_410) );
OAI31xp33_ASAP7_75t_L g411 ( .A1(n_349), .A2(n_290), .A3(n_272), .B(n_13), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_358), .Y(n_412) );
INVxp67_ASAP7_75t_SL g413 ( .A(n_376), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_358), .Y(n_414) );
HB1xp67_ASAP7_75t_L g415 ( .A(n_354), .Y(n_415) );
OR2x2_ASAP7_75t_L g416 ( .A(n_363), .B(n_11), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_359), .Y(n_417) );
AOI33xp33_ASAP7_75t_L g418 ( .A1(n_368), .A2(n_12), .A3(n_13), .B1(n_14), .B2(n_15), .B3(n_16), .Y(n_418) );
INVx5_ASAP7_75t_L g419 ( .A(n_354), .Y(n_419) );
NAND3xp33_ASAP7_75t_L g420 ( .A(n_368), .B(n_134), .C(n_137), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_409), .B(n_355), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_380), .B(n_359), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_391), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_382), .Y(n_424) );
OR2x2_ASAP7_75t_L g425 ( .A(n_390), .B(n_409), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_390), .B(n_363), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_380), .B(n_360), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_391), .Y(n_428) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_378), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_383), .B(n_367), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_397), .B(n_355), .Y(n_431) );
CKINVDCx16_ASAP7_75t_R g432 ( .A(n_386), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_383), .B(n_367), .Y(n_433) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_387), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_413), .Y(n_435) );
INVx5_ASAP7_75t_SL g436 ( .A(n_408), .Y(n_436) );
OR2x6_ASAP7_75t_L g437 ( .A(n_415), .B(n_363), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_393), .B(n_367), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_397), .B(n_355), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_389), .B(n_355), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_401), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_401), .Y(n_442) );
NAND4xp25_ASAP7_75t_L g443 ( .A(n_411), .B(n_374), .C(n_373), .D(n_369), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_382), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_404), .B(n_374), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_393), .B(n_374), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_386), .B(n_373), .Y(n_447) );
OAI21xp33_ASAP7_75t_SL g448 ( .A1(n_411), .A2(n_373), .B(n_369), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_399), .B(n_369), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_405), .Y(n_450) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_404), .Y(n_451) );
AND2x4_ASAP7_75t_L g452 ( .A(n_419), .B(n_354), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_399), .B(n_354), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_404), .B(n_134), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_405), .B(n_12), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_406), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_382), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_406), .Y(n_458) );
INVx3_ASAP7_75t_L g459 ( .A(n_419), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_412), .Y(n_460) );
INVx1_ASAP7_75t_SL g461 ( .A(n_419), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_412), .B(n_14), .Y(n_462) );
NAND2x1p5_ASAP7_75t_L g463 ( .A(n_419), .B(n_318), .Y(n_463) );
INVx1_ASAP7_75t_SL g464 ( .A(n_419), .Y(n_464) );
INVx3_ASAP7_75t_L g465 ( .A(n_419), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_414), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_407), .B(n_142), .Y(n_467) );
INVx1_ASAP7_75t_SL g468 ( .A(n_396), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_407), .B(n_142), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_414), .B(n_15), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_384), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_407), .B(n_142), .Y(n_472) );
INVx2_ASAP7_75t_SL g473 ( .A(n_417), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_416), .B(n_16), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_417), .B(n_142), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_416), .B(n_17), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_417), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_434), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_429), .B(n_432), .Y(n_479) );
INVx4_ASAP7_75t_L g480 ( .A(n_459), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_423), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_427), .B(n_398), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_438), .B(n_388), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_423), .Y(n_484) );
HB1xp67_ASAP7_75t_L g485 ( .A(n_435), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_438), .B(n_388), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_430), .B(n_388), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_430), .B(n_384), .Y(n_488) );
INVxp67_ASAP7_75t_L g489 ( .A(n_468), .Y(n_489) );
NOR3xp33_ASAP7_75t_SL g490 ( .A(n_448), .B(n_403), .C(n_385), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_433), .B(n_384), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_428), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_433), .B(n_408), .Y(n_493) );
INVxp67_ASAP7_75t_SL g494 ( .A(n_451), .Y(n_494) );
OR2x2_ASAP7_75t_L g495 ( .A(n_425), .B(n_398), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_427), .B(n_408), .Y(n_496) );
INVx3_ASAP7_75t_SL g497 ( .A(n_452), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_425), .B(n_418), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_422), .B(n_402), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_422), .B(n_402), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_446), .B(n_395), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_446), .B(n_395), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_428), .B(n_441), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_441), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_442), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_442), .B(n_400), .Y(n_506) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_440), .B(n_392), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_466), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_449), .B(n_395), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_466), .B(n_381), .Y(n_510) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_473), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_426), .B(n_395), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_450), .B(n_381), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_449), .B(n_379), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_456), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_453), .B(n_394), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_458), .B(n_394), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_473), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_453), .B(n_142), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_460), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_439), .B(n_142), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_477), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_439), .B(n_142), .Y(n_523) );
INVx2_ASAP7_75t_SL g524 ( .A(n_459), .Y(n_524) );
OR2x2_ASAP7_75t_L g525 ( .A(n_426), .B(n_431), .Y(n_525) );
NOR3xp33_ASAP7_75t_SL g526 ( .A(n_443), .B(n_410), .C(n_420), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_421), .B(n_392), .Y(n_527) );
CKINVDCx16_ASAP7_75t_R g528 ( .A(n_452), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_445), .Y(n_529) );
AND2x4_ASAP7_75t_L g530 ( .A(n_459), .B(n_420), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_455), .B(n_410), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_462), .B(n_137), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_445), .Y(n_533) );
AOI22xp5_ASAP7_75t_L g534 ( .A1(n_474), .A2(n_288), .B1(n_134), .B2(n_137), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_470), .B(n_137), .Y(n_535) );
AOI221x1_ASAP7_75t_L g536 ( .A1(n_499), .A2(n_476), .B1(n_465), .B2(n_447), .C(n_472), .Y(n_536) );
NAND2x1p5_ASAP7_75t_L g537 ( .A(n_480), .B(n_465), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_485), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_510), .B(n_424), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_478), .Y(n_540) );
AOI22xp5_ASAP7_75t_L g541 ( .A1(n_507), .A2(n_437), .B1(n_436), .B2(n_452), .Y(n_541) );
AOI31xp33_ASAP7_75t_L g542 ( .A1(n_479), .A2(n_461), .A3(n_464), .B(n_463), .Y(n_542) );
OAI222xp33_ASAP7_75t_L g543 ( .A1(n_480), .A2(n_437), .B1(n_465), .B2(n_463), .C1(n_436), .C2(n_444), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_503), .Y(n_544) );
OAI211xp5_ASAP7_75t_L g545 ( .A1(n_490), .A2(n_475), .B(n_472), .C(n_454), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_513), .B(n_424), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_528), .B(n_437), .Y(n_547) );
O2A1O1Ixp5_ASAP7_75t_L g548 ( .A1(n_480), .A2(n_457), .B(n_471), .C(n_444), .Y(n_548) );
AOI21xp33_ASAP7_75t_L g549 ( .A1(n_498), .A2(n_437), .B(n_475), .Y(n_549) );
OAI22xp5_ASAP7_75t_L g550 ( .A1(n_497), .A2(n_436), .B1(n_463), .B2(n_457), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_525), .B(n_471), .Y(n_551) );
OAI22xp33_ASAP7_75t_L g552 ( .A1(n_497), .A2(n_436), .B1(n_467), .B2(n_454), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_514), .B(n_467), .Y(n_553) );
O2A1O1Ixp33_ASAP7_75t_SL g554 ( .A1(n_489), .A2(n_469), .B(n_21), .C(n_22), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_514), .B(n_469), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_530), .A2(n_318), .B(n_316), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_515), .Y(n_557) );
OAI21xp33_ASAP7_75t_L g558 ( .A1(n_507), .A2(n_134), .B(n_137), .Y(n_558) );
AND2x4_ASAP7_75t_L g559 ( .A(n_524), .B(n_137), .Y(n_559) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_530), .A2(n_316), .B(n_134), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_511), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_516), .A2(n_134), .B1(n_137), .B2(n_169), .Y(n_562) );
AOI221xp5_ASAP7_75t_L g563 ( .A1(n_527), .A2(n_188), .B1(n_175), .B2(n_169), .C(n_165), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_520), .Y(n_564) );
OAI221xp5_ASAP7_75t_L g565 ( .A1(n_500), .A2(n_169), .B1(n_165), .B2(n_164), .C(n_158), .Y(n_565) );
INVxp67_ASAP7_75t_L g566 ( .A(n_519), .Y(n_566) );
OAI21xp33_ASAP7_75t_SL g567 ( .A1(n_524), .A2(n_19), .B(n_26), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_481), .Y(n_568) );
AOI21xp33_ASAP7_75t_L g569 ( .A1(n_531), .A2(n_30), .B(n_31), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_484), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_509), .B(n_32), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_492), .Y(n_572) );
INVx1_ASAP7_75t_SL g573 ( .A(n_519), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_504), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_483), .B(n_36), .Y(n_575) );
OAI21xp5_ASAP7_75t_L g576 ( .A1(n_526), .A2(n_165), .B(n_164), .Y(n_576) );
AOI211xp5_ASAP7_75t_L g577 ( .A1(n_516), .A2(n_164), .B(n_158), .C(n_153), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_495), .B(n_37), .Y(n_578) );
OAI21xp5_ASAP7_75t_L g579 ( .A1(n_530), .A2(n_158), .B(n_153), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_538), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_546), .Y(n_581) );
XOR2xp5_ASAP7_75t_L g582 ( .A(n_541), .B(n_495), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_557), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_564), .Y(n_584) );
AOI221xp5_ASAP7_75t_L g585 ( .A1(n_540), .A2(n_517), .B1(n_533), .B2(n_529), .C(n_506), .Y(n_585) );
XOR2x2_ASAP7_75t_L g586 ( .A(n_537), .B(n_496), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_539), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_548), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_544), .B(n_509), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_568), .Y(n_590) );
AOI222xp33_ASAP7_75t_L g591 ( .A1(n_566), .A2(n_501), .B1(n_502), .B2(n_521), .C1(n_523), .C2(n_496), .Y(n_591) );
XNOR2xp5_ASAP7_75t_L g592 ( .A(n_547), .B(n_493), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_570), .Y(n_593) );
OA21x2_ASAP7_75t_SL g594 ( .A1(n_573), .A2(n_482), .B(n_535), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_572), .B(n_502), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_574), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_551), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_573), .B(n_501), .Y(n_598) );
AND2x2_ASAP7_75t_L g599 ( .A(n_555), .B(n_483), .Y(n_599) );
INVxp67_ASAP7_75t_L g600 ( .A(n_561), .Y(n_600) );
AND2x2_ASAP7_75t_L g601 ( .A(n_553), .B(n_486), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_537), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_536), .B(n_494), .Y(n_603) );
NAND3xp33_ASAP7_75t_L g604 ( .A(n_577), .B(n_523), .C(n_521), .Y(n_604) );
OAI21xp5_ASAP7_75t_SL g605 ( .A1(n_542), .A2(n_493), .B(n_486), .Y(n_605) );
OAI22xp5_ASAP7_75t_L g606 ( .A1(n_542), .A2(n_518), .B1(n_512), .B2(n_522), .Y(n_606) );
AOI21x1_ASAP7_75t_L g607 ( .A1(n_606), .A2(n_559), .B(n_560), .Y(n_607) );
AOI221xp5_ASAP7_75t_L g608 ( .A1(n_585), .A2(n_549), .B1(n_543), .B2(n_565), .C(n_545), .Y(n_608) );
OAI211xp5_ASAP7_75t_L g609 ( .A1(n_605), .A2(n_567), .B(n_558), .C(n_562), .Y(n_609) );
OA211x2_ASAP7_75t_L g610 ( .A1(n_585), .A2(n_571), .B(n_579), .C(n_563), .Y(n_610) );
INVx1_ASAP7_75t_SL g611 ( .A(n_586), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_581), .Y(n_612) );
NAND3xp33_ASAP7_75t_SL g613 ( .A(n_603), .B(n_550), .C(n_578), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_587), .Y(n_614) );
O2A1O1Ixp33_ASAP7_75t_SL g615 ( .A1(n_606), .A2(n_552), .B(n_569), .C(n_579), .Y(n_615) );
AOI21xp33_ASAP7_75t_L g616 ( .A1(n_588), .A2(n_559), .B(n_532), .Y(n_616) );
INVxp67_ASAP7_75t_L g617 ( .A(n_580), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_592), .A2(n_575), .B1(n_518), .B2(n_512), .Y(n_618) );
AND2x4_ASAP7_75t_L g619 ( .A(n_602), .B(n_508), .Y(n_619) );
OAI31xp33_ASAP7_75t_L g620 ( .A1(n_582), .A2(n_554), .A3(n_505), .B(n_491), .Y(n_620) );
OAI22xp33_ASAP7_75t_L g621 ( .A1(n_603), .A2(n_488), .B1(n_491), .B2(n_487), .Y(n_621) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_604), .A2(n_488), .B1(n_487), .B2(n_534), .Y(n_622) );
OAI311xp33_ASAP7_75t_L g623 ( .A1(n_608), .A2(n_591), .A3(n_594), .B1(n_600), .C1(n_589), .Y(n_623) );
OAI211xp5_ASAP7_75t_SL g624 ( .A1(n_620), .A2(n_589), .B(n_584), .C(n_583), .Y(n_624) );
OAI22xp33_ASAP7_75t_SL g625 ( .A1(n_611), .A2(n_593), .B1(n_590), .B2(n_596), .Y(n_625) );
NAND3xp33_ASAP7_75t_L g626 ( .A(n_615), .B(n_576), .C(n_595), .Y(n_626) );
AOI221xp5_ASAP7_75t_L g627 ( .A1(n_621), .A2(n_613), .B1(n_616), .B2(n_622), .C(n_617), .Y(n_627) );
OAI322xp33_ASAP7_75t_L g628 ( .A1(n_618), .A2(n_595), .A3(n_597), .B1(n_598), .B2(n_601), .C1(n_599), .C2(n_556), .Y(n_628) );
NOR4xp25_ASAP7_75t_L g629 ( .A(n_609), .B(n_153), .C(n_151), .D(n_42), .Y(n_629) );
OAI22xp5_ASAP7_75t_L g630 ( .A1(n_607), .A2(n_151), .B1(n_41), .B2(n_43), .Y(n_630) );
AOI221xp5_ASAP7_75t_L g631 ( .A1(n_612), .A2(n_151), .B1(n_44), .B2(n_49), .C(n_50), .Y(n_631) );
OAI211xp5_ASAP7_75t_L g632 ( .A1(n_627), .A2(n_610), .B(n_614), .C(n_619), .Y(n_632) );
OAI21xp33_ASAP7_75t_L g633 ( .A1(n_624), .A2(n_619), .B(n_51), .Y(n_633) );
AND2x4_ASAP7_75t_L g634 ( .A(n_626), .B(n_39), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_625), .B(n_54), .Y(n_635) );
NAND3xp33_ASAP7_75t_SL g636 ( .A(n_629), .B(n_56), .C(n_57), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_634), .B(n_630), .Y(n_637) );
NAND3xp33_ASAP7_75t_SL g638 ( .A(n_632), .B(n_623), .C(n_631), .Y(n_638) );
OAI22x1_ASAP7_75t_L g639 ( .A1(n_635), .A2(n_628), .B1(n_61), .B2(n_66), .Y(n_639) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_637), .Y(n_640) );
INVxp67_ASAP7_75t_SL g641 ( .A(n_639), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_640), .Y(n_642) );
AOI21xp33_ASAP7_75t_SL g643 ( .A1(n_641), .A2(n_633), .B(n_638), .Y(n_643) );
BUFx6f_ASAP7_75t_L g644 ( .A(n_642), .Y(n_644) );
AOI22xp33_ASAP7_75t_R g645 ( .A1(n_644), .A2(n_643), .B1(n_636), .B2(n_70), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_645), .A2(n_644), .B1(n_69), .B2(n_71), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g647 ( .A1(n_646), .A2(n_644), .B1(n_58), .B2(n_76), .Y(n_647) );
endmodule