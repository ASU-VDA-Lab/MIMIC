module fake_netlist_5_1250_n_757 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_757);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_757;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_684;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_667;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_452;
wire n_397;
wire n_525;
wire n_493;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_155;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_378;
wire n_551;
wire n_688;
wire n_581;
wire n_382;
wire n_554;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_372;
wire n_293;
wire n_443;
wire n_244;
wire n_677;
wire n_173;
wire n_198;
wire n_714;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_373;
wire n_307;
wire n_633;
wire n_439;
wire n_150;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_576;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_563;
wire n_171;
wire n_153;
wire n_756;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_752;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_325;
wire n_449;
wire n_724;
wire n_546;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_152;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_654;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_379;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_156;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_219;
wire n_442;
wire n_157;
wire n_192;
wire n_636;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_158;
wire n_655;
wire n_704;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_183;
wire n_243;
wire n_185;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_696;
wire n_215;
wire n_350;
wire n_196;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_473;
wire n_422;
wire n_475;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_670;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_521;
wire n_614;
wire n_663;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_553;
wire n_727;
wire n_311;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_749;
wire n_691;
wire n_717;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_517;
wire n_482;
wire n_588;
wire n_361;
wire n_464;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_149;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_693;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_151;
wire n_306;
wire n_575;
wire n_722;
wire n_458;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_474;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_736;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_745;
wire n_627;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_729;
wire n_730;
wire n_176;
wire n_557;
wire n_182;
wire n_354;
wire n_607;
wire n_647;
wire n_480;
wire n_679;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_707;
wire n_710;
wire n_695;
wire n_180;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_720;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_565;
wire n_426;
wire n_520;
wire n_566;
wire n_409;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_154;
wire n_148;
wire n_300;
wire n_651;
wire n_435;
wire n_159;
wire n_334;
wire n_599;
wire n_541;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_538;
wire n_666;
wire n_262;
wire n_238;
wire n_639;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_200;
wire n_162;
wire n_222;
wire n_438;
wire n_713;
wire n_324;
wire n_634;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;

INVx2_ASAP7_75t_SL g148 ( 
.A(n_103),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_65),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g150 ( 
.A(n_131),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_54),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_93),
.Y(n_152)
);

BUFx10_ASAP7_75t_L g153 ( 
.A(n_35),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_117),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_91),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

BUFx10_ASAP7_75t_L g157 ( 
.A(n_37),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_120),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_7),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_82),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_61),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_90),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_80),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_135),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_42),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_77),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_134),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_63),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_122),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_14),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_92),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_84),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_79),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_41),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_76),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_75),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_64),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_44),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_32),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_115),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_19),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_21),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_23),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_100),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_114),
.Y(n_186)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_16),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_142),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_145),
.Y(n_189)
);

BUFx10_ASAP7_75t_L g190 ( 
.A(n_133),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_81),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_144),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_46),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_40),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_104),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_89),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_119),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_138),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_129),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_121),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_25),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_159),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_170),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_152),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g205 ( 
.A(n_182),
.Y(n_205)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_156),
.Y(n_206)
);

OAI22x1_ASAP7_75t_R g207 ( 
.A1(n_172),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_0),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_1),
.Y(n_209)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_148),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_187),
.Y(n_211)
);

OAI21x1_ASAP7_75t_L g212 ( 
.A1(n_160),
.A2(n_2),
.B(n_3),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_152),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_155),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_156),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_199),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_160),
.B(n_3),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_155),
.Y(n_218)
);

AND2x6_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_22),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_156),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g221 ( 
.A(n_157),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_193),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_4),
.Y(n_223)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_157),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_193),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_164),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_156),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_172),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_156),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_149),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_171),
.B(n_5),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_178),
.Y(n_232)
);

OA21x2_ASAP7_75t_L g233 ( 
.A1(n_151),
.A2(n_6),
.B(n_7),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_158),
.Y(n_234)
);

OA21x2_ASAP7_75t_L g235 ( 
.A1(n_163),
.A2(n_8),
.B(n_9),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_156),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_166),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_168),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_169),
.Y(n_239)
);

INVxp33_ASAP7_75t_SL g240 ( 
.A(n_150),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_175),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_240),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_240),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_232),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_232),
.Y(n_245)
);

BUFx10_ASAP7_75t_L g246 ( 
.A(n_208),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_228),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_228),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_221),
.B(n_176),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_204),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_224),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_202),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_211),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_211),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_204),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_205),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_205),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_221),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_216),
.Y(n_259)
);

AND2x6_ASAP7_75t_L g260 ( 
.A(n_206),
.B(n_179),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_222),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_R g262 ( 
.A(n_213),
.B(n_154),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_237),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_209),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_204),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_204),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_204),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_214),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_214),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_225),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_214),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_214),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_210),
.B(n_180),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_214),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_218),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_218),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_238),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_218),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_218),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_218),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_234),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_239),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_234),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_239),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_239),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_239),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_230),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_239),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_271),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_256),
.B(n_231),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_288),
.B(n_210),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_251),
.B(n_153),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_257),
.B(n_210),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_265),
.B(n_210),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_258),
.B(n_153),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_287),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_284),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_261),
.B(n_210),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_268),
.Y(n_299)
);

NAND3xp33_ASAP7_75t_L g300 ( 
.A(n_270),
.B(n_223),
.C(n_217),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_272),
.B(n_241),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_281),
.B(n_241),
.Y(n_302)
);

INVxp67_ASAP7_75t_SL g303 ( 
.A(n_266),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_283),
.B(n_241),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_275),
.B(n_241),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_276),
.B(n_241),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_278),
.B(n_161),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_263),
.B(n_153),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_250),
.B(n_162),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_255),
.B(n_165),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_267),
.B(n_167),
.Y(n_311)
);

XOR2x2_ASAP7_75t_L g312 ( 
.A(n_252),
.B(n_226),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_269),
.Y(n_313)
);

INVx1_ASAP7_75t_SL g314 ( 
.A(n_248),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_262),
.Y(n_315)
);

NAND3xp33_ASAP7_75t_L g316 ( 
.A(n_249),
.B(n_203),
.C(n_174),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_266),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_266),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_253),
.B(n_190),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_286),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_274),
.B(n_173),
.Y(n_321)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_282),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_254),
.B(n_246),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_279),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_266),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_280),
.B(n_177),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_285),
.Y(n_327)
);

OAI21xp33_ASAP7_75t_L g328 ( 
.A1(n_259),
.A2(n_188),
.B(n_196),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_242),
.B(n_181),
.Y(n_329)
);

INVx2_ASAP7_75t_SL g330 ( 
.A(n_246),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_285),
.B(n_183),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_243),
.B(n_184),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_273),
.B(n_185),
.Y(n_333)
);

NAND2xp33_ASAP7_75t_L g334 ( 
.A(n_260),
.B(n_219),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_264),
.B(n_244),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_260),
.B(n_186),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_245),
.B(n_189),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_247),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_282),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_260),
.B(n_191),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_260),
.B(n_192),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_282),
.B(n_194),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_277),
.B(n_190),
.Y(n_343)
);

AND2x4_ASAP7_75t_L g344 ( 
.A(n_260),
.B(n_212),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_282),
.A2(n_197),
.B1(n_198),
.B2(n_200),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_288),
.B(n_219),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_256),
.B(n_190),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_288),
.B(n_219),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_256),
.B(n_206),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_287),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_271),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_288),
.B(n_219),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_297),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_349),
.B(n_219),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_349),
.A2(n_219),
.B1(n_235),
.B2(n_233),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_344),
.B(n_233),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_344),
.B(n_233),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_302),
.B(n_235),
.Y(n_358)
);

INVx1_ASAP7_75t_SL g359 ( 
.A(n_314),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_299),
.B(n_236),
.Y(n_360)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_299),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_296),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_302),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_335),
.A2(n_207),
.B1(n_235),
.B2(n_10),
.Y(n_364)
);

INVx5_ASAP7_75t_L g365 ( 
.A(n_322),
.Y(n_365)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_297),
.Y(n_366)
);

OR2x2_ASAP7_75t_L g367 ( 
.A(n_290),
.B(n_212),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_329),
.B(n_332),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_350),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_320),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_320),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_304),
.Y(n_372)
);

O2A1O1Ixp33_ASAP7_75t_L g373 ( 
.A1(n_328),
.A2(n_334),
.B(n_352),
.C(n_348),
.Y(n_373)
);

AND2x4_ASAP7_75t_L g374 ( 
.A(n_300),
.B(n_24),
.Y(n_374)
);

OAI221xp5_ASAP7_75t_L g375 ( 
.A1(n_345),
.A2(n_236),
.B1(n_229),
.B2(n_227),
.C(n_220),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_289),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_304),
.B(n_215),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_289),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_301),
.B(n_215),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_305),
.B(n_220),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_337),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_329),
.B(n_8),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_325),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_351),
.Y(n_384)
);

NOR2x2_ASAP7_75t_L g385 ( 
.A(n_312),
.B(n_9),
.Y(n_385)
);

AND2x6_ASAP7_75t_SL g386 ( 
.A(n_335),
.B(n_10),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_351),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_306),
.B(n_227),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_313),
.B(n_229),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_337),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g391 ( 
.A(n_338),
.Y(n_391)
);

INVx3_ASAP7_75t_L g392 ( 
.A(n_325),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_327),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_332),
.B(n_11),
.Y(n_394)
);

INVx5_ASAP7_75t_L g395 ( 
.A(n_322),
.Y(n_395)
);

AND2x4_ASAP7_75t_L g396 ( 
.A(n_315),
.B(n_26),
.Y(n_396)
);

BUFx3_ASAP7_75t_L g397 ( 
.A(n_330),
.Y(n_397)
);

A2O1A1Ixp33_ASAP7_75t_SL g398 ( 
.A1(n_342),
.A2(n_78),
.B(n_147),
.C(n_146),
.Y(n_398)
);

AOI22xp33_ASAP7_75t_L g399 ( 
.A1(n_324),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_339),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_317),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_292),
.B(n_12),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_333),
.B(n_27),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_318),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_293),
.B(n_13),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_347),
.B(n_14),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_323),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_293),
.B(n_15),
.Y(n_408)
);

AND2x4_ASAP7_75t_L g409 ( 
.A(n_316),
.B(n_28),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_295),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_308),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_342),
.A2(n_85),
.B1(n_143),
.B2(n_140),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_303),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_319),
.B(n_15),
.Y(n_414)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_346),
.Y(n_415)
);

OR2x6_ASAP7_75t_L g416 ( 
.A(n_343),
.B(n_16),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_298),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_307),
.A2(n_86),
.B1(n_139),
.B2(n_137),
.Y(n_418)
);

OR2x2_ASAP7_75t_SL g419 ( 
.A(n_331),
.B(n_17),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_309),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_298),
.B(n_17),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_356),
.A2(n_321),
.B(n_310),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_368),
.A2(n_326),
.B1(n_311),
.B2(n_336),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_390),
.B(n_294),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_362),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_353),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_370),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_356),
.A2(n_341),
.B(n_340),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_383),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_372),
.B(n_291),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_381),
.B(n_18),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_363),
.B(n_18),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_357),
.A2(n_83),
.B1(n_136),
.B2(n_29),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_420),
.B(n_19),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_377),
.B(n_20),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_357),
.A2(n_87),
.B1(n_30),
.B2(n_31),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_361),
.B(n_20),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_376),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_361),
.B(n_33),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_383),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_378),
.Y(n_441)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_379),
.A2(n_34),
.B(n_36),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_359),
.Y(n_443)
);

OAI21xp33_ASAP7_75t_L g444 ( 
.A1(n_382),
.A2(n_38),
.B(n_39),
.Y(n_444)
);

AO21x1_ASAP7_75t_L g445 ( 
.A1(n_394),
.A2(n_403),
.B(n_355),
.Y(n_445)
);

AOI21xp5_ASAP7_75t_L g446 ( 
.A1(n_379),
.A2(n_43),
.B(n_45),
.Y(n_446)
);

OAI21x1_ASAP7_75t_L g447 ( 
.A1(n_415),
.A2(n_47),
.B(n_48),
.Y(n_447)
);

A2O1A1Ixp33_ASAP7_75t_L g448 ( 
.A1(n_367),
.A2(n_49),
.B(n_50),
.C(n_51),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_396),
.B(n_52),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_410),
.B(n_53),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_380),
.A2(n_55),
.B(n_56),
.Y(n_451)
);

OR2x6_ASAP7_75t_L g452 ( 
.A(n_391),
.B(n_57),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_377),
.B(n_358),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_373),
.A2(n_58),
.B(n_59),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_374),
.A2(n_409),
.B1(n_360),
.B2(n_369),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_371),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_380),
.B(n_60),
.Y(n_457)
);

INVx6_ASAP7_75t_SL g458 ( 
.A(n_416),
.Y(n_458)
);

O2A1O1Ixp33_ASAP7_75t_L g459 ( 
.A1(n_405),
.A2(n_408),
.B(n_421),
.C(n_406),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_415),
.B(n_62),
.Y(n_460)
);

BUFx2_ASAP7_75t_L g461 ( 
.A(n_359),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_387),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_384),
.Y(n_463)
);

A2O1A1Ixp33_ASAP7_75t_L g464 ( 
.A1(n_414),
.A2(n_66),
.B(n_67),
.C(n_68),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_388),
.A2(n_354),
.B(n_413),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_417),
.B(n_69),
.Y(n_466)
);

OR2x6_ASAP7_75t_L g467 ( 
.A(n_416),
.B(n_70),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_374),
.B(n_71),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_403),
.A2(n_72),
.B(n_73),
.Y(n_469)
);

O2A1O1Ixp33_ASAP7_75t_L g470 ( 
.A1(n_402),
.A2(n_74),
.B(n_88),
.C(n_94),
.Y(n_470)
);

OR2x6_ASAP7_75t_L g471 ( 
.A(n_416),
.B(n_95),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_396),
.B(n_96),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_383),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_409),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_474)
);

A2O1A1Ixp33_ASAP7_75t_L g475 ( 
.A1(n_393),
.A2(n_101),
.B(n_102),
.C(n_105),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_389),
.B(n_106),
.Y(n_476)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_397),
.B(n_107),
.Y(n_477)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_461),
.Y(n_478)
);

CKINVDCx11_ASAP7_75t_R g479 ( 
.A(n_452),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g480 ( 
.A(n_430),
.B(n_407),
.Y(n_480)
);

INVxp67_ASAP7_75t_SL g481 ( 
.A(n_429),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_L g482 ( 
.A1(n_453),
.A2(n_389),
.B(n_366),
.Y(n_482)
);

AO21x2_ASAP7_75t_L g483 ( 
.A1(n_445),
.A2(n_398),
.B(n_400),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_455),
.B(n_401),
.Y(n_484)
);

AO21x2_ASAP7_75t_L g485 ( 
.A1(n_454),
.A2(n_412),
.B(n_418),
.Y(n_485)
);

BUFx2_ASAP7_75t_SL g486 ( 
.A(n_429),
.Y(n_486)
);

INVx2_ASAP7_75t_SL g487 ( 
.A(n_443),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_456),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_425),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_426),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_465),
.A2(n_365),
.B(n_395),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_429),
.Y(n_492)
);

OAI21x1_ASAP7_75t_SL g493 ( 
.A1(n_468),
.A2(n_399),
.B(n_419),
.Y(n_493)
);

INVx2_ASAP7_75t_SL g494 ( 
.A(n_473),
.Y(n_494)
);

INVx5_ASAP7_75t_L g495 ( 
.A(n_473),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_463),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_427),
.Y(n_497)
);

INVx4_ASAP7_75t_L g498 ( 
.A(n_473),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_438),
.Y(n_499)
);

INVx2_ASAP7_75t_SL g500 ( 
.A(n_440),
.Y(n_500)
);

NAND2x1p5_ASAP7_75t_L g501 ( 
.A(n_447),
.B(n_392),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_441),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_462),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_452),
.Y(n_504)
);

CKINVDCx11_ASAP7_75t_R g505 ( 
.A(n_467),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_477),
.Y(n_506)
);

OAI21x1_ASAP7_75t_L g507 ( 
.A1(n_428),
.A2(n_392),
.B(n_404),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_435),
.Y(n_508)
);

AOI21x1_ASAP7_75t_L g509 ( 
.A1(n_457),
.A2(n_366),
.B(n_404),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_440),
.Y(n_510)
);

AOI22x1_ASAP7_75t_L g511 ( 
.A1(n_422),
.A2(n_411),
.B1(n_375),
.B2(n_364),
.Y(n_511)
);

OAI21x1_ASAP7_75t_L g512 ( 
.A1(n_460),
.A2(n_395),
.B(n_365),
.Y(n_512)
);

NAND2x1p5_ASAP7_75t_L g513 ( 
.A(n_439),
.B(n_472),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_L g514 ( 
.A1(n_449),
.A2(n_395),
.B1(n_365),
.B2(n_385),
.Y(n_514)
);

AND2x4_ASAP7_75t_L g515 ( 
.A(n_467),
.B(n_395),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_476),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_434),
.Y(n_517)
);

HB1xp67_ASAP7_75t_L g518 ( 
.A(n_471),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_433),
.Y(n_519)
);

BUFx4_ASAP7_75t_SL g520 ( 
.A(n_471),
.Y(n_520)
);

OA21x2_ASAP7_75t_L g521 ( 
.A1(n_448),
.A2(n_365),
.B(n_109),
.Y(n_521)
);

OR2x6_ASAP7_75t_L g522 ( 
.A(n_459),
.B(n_108),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_480),
.A2(n_506),
.B1(n_478),
.B2(n_431),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_L g524 ( 
.A1(n_511),
.A2(n_432),
.B1(n_474),
.B2(n_444),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_508),
.B(n_424),
.Y(n_525)
);

NAND2x1p5_ASAP7_75t_L g526 ( 
.A(n_495),
.B(n_498),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_488),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_495),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_488),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_496),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_496),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_489),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_487),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_503),
.Y(n_534)
);

OR2x6_ASAP7_75t_L g535 ( 
.A(n_486),
.B(n_470),
.Y(n_535)
);

CKINVDCx6p67_ASAP7_75t_R g536 ( 
.A(n_504),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_503),
.Y(n_537)
);

OAI21x1_ASAP7_75t_L g538 ( 
.A1(n_512),
.A2(n_469),
.B(n_446),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_490),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_490),
.Y(n_540)
);

AOI21x1_ASAP7_75t_L g541 ( 
.A1(n_509),
.A2(n_442),
.B(n_451),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_495),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_L g543 ( 
.A1(n_511),
.A2(n_437),
.B1(n_450),
.B2(n_466),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_508),
.B(n_423),
.Y(n_544)
);

INVx1_ASAP7_75t_SL g545 ( 
.A(n_487),
.Y(n_545)
);

INVx4_ASAP7_75t_L g546 ( 
.A(n_495),
.Y(n_546)
);

AOI22xp5_ASAP7_75t_L g547 ( 
.A1(n_480),
.A2(n_436),
.B1(n_464),
.B2(n_475),
.Y(n_547)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_518),
.A2(n_458),
.B1(n_386),
.B2(n_112),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_497),
.Y(n_549)
);

INVx3_ASAP7_75t_SL g550 ( 
.A(n_504),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_495),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_497),
.Y(n_552)
);

OA21x2_ASAP7_75t_L g553 ( 
.A1(n_507),
.A2(n_458),
.B(n_111),
.Y(n_553)
);

CKINVDCx11_ASAP7_75t_R g554 ( 
.A(n_479),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_517),
.A2(n_110),
.B1(n_113),
.B2(n_116),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_499),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_517),
.B(n_118),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_499),
.Y(n_558)
);

BUFx2_ASAP7_75t_L g559 ( 
.A(n_481),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_520),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_502),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_525),
.B(n_514),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_527),
.Y(n_563)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_533),
.Y(n_564)
);

HB1xp67_ASAP7_75t_L g565 ( 
.A(n_533),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_523),
.B(n_502),
.Y(n_566)
);

OR2x6_ASAP7_75t_L g567 ( 
.A(n_535),
.B(n_522),
.Y(n_567)
);

AO32x1_ASAP7_75t_L g568 ( 
.A1(n_530),
.A2(n_519),
.A3(n_516),
.B1(n_500),
.B2(n_510),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_544),
.B(n_493),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_557),
.B(n_515),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_527),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_R g572 ( 
.A(n_560),
.B(n_505),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_529),
.Y(n_573)
);

INVx5_ASAP7_75t_L g574 ( 
.A(n_528),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_R g575 ( 
.A(n_554),
.B(n_495),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_529),
.Y(n_576)
);

OR2x6_ASAP7_75t_L g577 ( 
.A(n_535),
.B(n_522),
.Y(n_577)
);

NAND2xp33_ASAP7_75t_R g578 ( 
.A(n_535),
.B(n_521),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_SL g579 ( 
.A(n_550),
.B(n_515),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_554),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_R g581 ( 
.A(n_550),
.B(n_492),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_536),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_531),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_L g584 ( 
.A1(n_543),
.A2(n_493),
.B1(n_522),
.B2(n_485),
.Y(n_584)
);

AOI21xp5_ASAP7_75t_L g585 ( 
.A1(n_543),
.A2(n_485),
.B(n_516),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_532),
.B(n_515),
.Y(n_586)
);

INVx4_ASAP7_75t_L g587 ( 
.A(n_528),
.Y(n_587)
);

INVxp67_ASAP7_75t_L g588 ( 
.A(n_545),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_534),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_537),
.B(n_515),
.Y(n_590)
);

OAI21x1_ASAP7_75t_L g591 ( 
.A1(n_538),
.A2(n_512),
.B(n_509),
.Y(n_591)
);

A2O1A1Ixp33_ASAP7_75t_L g592 ( 
.A1(n_524),
.A2(n_519),
.B(n_482),
.C(n_484),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_548),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_539),
.Y(n_594)
);

CKINVDCx16_ASAP7_75t_R g595 ( 
.A(n_559),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_L g596 ( 
.A1(n_524),
.A2(n_522),
.B1(n_513),
.B2(n_484),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_552),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_L g598 ( 
.A1(n_547),
.A2(n_522),
.B1(n_485),
.B2(n_513),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_556),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_540),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_540),
.Y(n_601)
);

AOI22xp33_ASAP7_75t_L g602 ( 
.A1(n_555),
.A2(n_484),
.B1(n_513),
.B2(n_521),
.Y(n_602)
);

NOR3xp33_ASAP7_75t_SL g603 ( 
.A(n_558),
.B(n_510),
.C(n_491),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_561),
.B(n_492),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_549),
.B(n_492),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_549),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_551),
.B(n_484),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_583),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_573),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_563),
.B(n_553),
.Y(n_610)
);

AND2x2_ASAP7_75t_L g611 ( 
.A(n_571),
.B(n_553),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_576),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_589),
.B(n_553),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_564),
.Y(n_614)
);

NAND3xp33_ASAP7_75t_L g615 ( 
.A(n_593),
.B(n_521),
.C(n_500),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_600),
.Y(n_616)
);

OR2x2_ASAP7_75t_L g617 ( 
.A(n_569),
.B(n_483),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_568),
.Y(n_618)
);

BUFx3_ASAP7_75t_L g619 ( 
.A(n_586),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_606),
.Y(n_620)
);

AOI22xp33_ASAP7_75t_SL g621 ( 
.A1(n_596),
.A2(n_521),
.B1(n_551),
.B2(n_542),
.Y(n_621)
);

BUFx2_ASAP7_75t_L g622 ( 
.A(n_564),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_594),
.B(n_483),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_568),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_607),
.B(n_546),
.Y(n_625)
);

AND2x4_ASAP7_75t_L g626 ( 
.A(n_567),
.B(n_546),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_565),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_562),
.B(n_494),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_601),
.Y(n_629)
);

HB1xp67_ASAP7_75t_L g630 ( 
.A(n_565),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_SL g631 ( 
.A1(n_595),
.A2(n_542),
.B1(n_528),
.B2(n_486),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_597),
.B(n_599),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_568),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_591),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_566),
.B(n_605),
.Y(n_635)
);

OR2x2_ASAP7_75t_L g636 ( 
.A(n_567),
.B(n_483),
.Y(n_636)
);

OAI221xp5_ASAP7_75t_L g637 ( 
.A1(n_598),
.A2(n_501),
.B1(n_541),
.B2(n_494),
.C(n_526),
.Y(n_637)
);

AOI22xp5_ASAP7_75t_L g638 ( 
.A1(n_570),
.A2(n_498),
.B1(n_528),
.B2(n_542),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_588),
.B(n_498),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_603),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_604),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_603),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_592),
.Y(n_643)
);

INVx4_ASAP7_75t_L g644 ( 
.A(n_626),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_623),
.B(n_577),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_609),
.Y(n_646)
);

NOR2xp67_ASAP7_75t_L g647 ( 
.A(n_614),
.B(n_588),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_609),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_630),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_623),
.B(n_577),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_635),
.B(n_636),
.Y(n_651)
);

OR2x2_ASAP7_75t_L g652 ( 
.A(n_636),
.B(n_567),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_635),
.B(n_585),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_622),
.Y(n_654)
);

OR2x2_ASAP7_75t_L g655 ( 
.A(n_617),
.B(n_577),
.Y(n_655)
);

NAND2xp33_ASAP7_75t_R g656 ( 
.A(n_639),
.B(n_572),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_608),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_622),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_617),
.B(n_584),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_628),
.B(n_584),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_627),
.Y(n_661)
);

OAI22xp5_ASAP7_75t_L g662 ( 
.A1(n_631),
.A2(n_602),
.B1(n_592),
.B2(n_582),
.Y(n_662)
);

NAND2xp67_ASAP7_75t_L g663 ( 
.A(n_632),
.B(n_590),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_613),
.B(n_602),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_632),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_613),
.B(n_507),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_641),
.B(n_587),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_641),
.B(n_587),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_620),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_SL g670 ( 
.A(n_626),
.B(n_580),
.Y(n_670)
);

AND2x2_ASAP7_75t_SL g671 ( 
.A(n_644),
.B(n_626),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_646),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_651),
.B(n_643),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_657),
.Y(n_674)
);

OR2x2_ASAP7_75t_L g675 ( 
.A(n_651),
.B(n_642),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_646),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_660),
.B(n_649),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_648),
.Y(n_678)
);

OR2x2_ASAP7_75t_L g679 ( 
.A(n_655),
.B(n_642),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_645),
.B(n_618),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_657),
.Y(n_681)
);

INVx4_ASAP7_75t_L g682 ( 
.A(n_644),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_669),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_645),
.B(n_618),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_653),
.B(n_643),
.Y(n_685)
);

OR2x2_ASAP7_75t_L g686 ( 
.A(n_655),
.B(n_640),
.Y(n_686)
);

OAI22xp5_ASAP7_75t_L g687 ( 
.A1(n_677),
.A2(n_662),
.B1(n_640),
.B2(n_652),
.Y(n_687)
);

AND2x4_ASAP7_75t_L g688 ( 
.A(n_682),
.B(n_644),
.Y(n_688)
);

OAI22xp5_ASAP7_75t_L g689 ( 
.A1(n_685),
.A2(n_652),
.B1(n_638),
.B2(n_621),
.Y(n_689)
);

OAI32xp33_ASAP7_75t_L g690 ( 
.A1(n_675),
.A2(n_656),
.A3(n_578),
.B1(n_615),
.B2(n_658),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_672),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_680),
.B(n_650),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_672),
.Y(n_693)
);

XNOR2xp5_ASAP7_75t_L g694 ( 
.A(n_671),
.B(n_663),
.Y(n_694)
);

AND2x4_ASAP7_75t_L g695 ( 
.A(n_682),
.B(n_665),
.Y(n_695)
);

OAI22xp5_ASAP7_75t_L g696 ( 
.A1(n_671),
.A2(n_647),
.B1(n_619),
.B2(n_637),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_674),
.Y(n_697)
);

AOI22xp5_ASAP7_75t_L g698 ( 
.A1(n_687),
.A2(n_670),
.B1(n_659),
.B2(n_650),
.Y(n_698)
);

AOI21xp33_ASAP7_75t_SL g699 ( 
.A1(n_694),
.A2(n_686),
.B(n_679),
.Y(n_699)
);

NAND3xp33_ASAP7_75t_L g700 ( 
.A(n_696),
.B(n_654),
.C(n_683),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_697),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_688),
.B(n_673),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_701),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_699),
.B(n_692),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_702),
.Y(n_705)
);

AO22x2_ASAP7_75t_L g706 ( 
.A1(n_700),
.A2(n_688),
.B1(n_682),
.B2(n_695),
.Y(n_706)
);

AOI21xp33_ASAP7_75t_L g707 ( 
.A1(n_698),
.A2(n_690),
.B(n_689),
.Y(n_707)
);

INVx3_ASAP7_75t_SL g708 ( 
.A(n_706),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_705),
.B(n_695),
.Y(n_709)
);

NOR3xp33_ASAP7_75t_L g710 ( 
.A(n_707),
.B(n_704),
.C(n_703),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_705),
.B(n_680),
.Y(n_711)
);

OAI22xp5_ASAP7_75t_L g712 ( 
.A1(n_708),
.A2(n_684),
.B1(n_681),
.B2(n_664),
.Y(n_712)
);

AOI21xp33_ASAP7_75t_L g713 ( 
.A1(n_709),
.A2(n_690),
.B(n_661),
.Y(n_713)
);

AOI21xp5_ASAP7_75t_L g714 ( 
.A1(n_710),
.A2(n_579),
.B(n_691),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_711),
.B(n_663),
.Y(n_715)
);

AOI221xp5_ASAP7_75t_L g716 ( 
.A1(n_713),
.A2(n_572),
.B1(n_693),
.B2(n_664),
.C(n_684),
.Y(n_716)
);

OAI221xp5_ASAP7_75t_L g717 ( 
.A1(n_712),
.A2(n_578),
.B1(n_676),
.B2(n_678),
.C(n_619),
.Y(n_717)
);

AOI221xp5_ASAP7_75t_L g718 ( 
.A1(n_714),
.A2(n_659),
.B1(n_676),
.B2(n_678),
.C(n_667),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_715),
.Y(n_719)
);

NOR2x1_ASAP7_75t_L g720 ( 
.A(n_719),
.B(n_575),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_717),
.Y(n_721)
);

INVx1_ASAP7_75t_SL g722 ( 
.A(n_716),
.Y(n_722)
);

NOR2x1_ASAP7_75t_L g723 ( 
.A(n_718),
.B(n_575),
.Y(n_723)
);

NOR2x1_ASAP7_75t_L g724 ( 
.A(n_719),
.B(n_581),
.Y(n_724)
);

AND2x2_ASAP7_75t_SL g725 ( 
.A(n_719),
.B(n_581),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_725),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_720),
.B(n_668),
.Y(n_727)
);

AOI21xp5_ASAP7_75t_L g728 ( 
.A1(n_724),
.A2(n_612),
.B(n_668),
.Y(n_728)
);

OR2x2_ASAP7_75t_L g729 ( 
.A(n_722),
.B(n_667),
.Y(n_729)
);

OAI21xp5_ASAP7_75t_L g730 ( 
.A1(n_721),
.A2(n_625),
.B(n_612),
.Y(n_730)
);

NAND4xp25_ASAP7_75t_L g731 ( 
.A(n_723),
.B(n_625),
.C(n_648),
.D(n_620),
.Y(n_731)
);

XNOR2x1_ASAP7_75t_L g732 ( 
.A(n_726),
.B(n_123),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_729),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_R g734 ( 
.A(n_727),
.B(n_124),
.Y(n_734)
);

INVx1_ASAP7_75t_SL g735 ( 
.A(n_730),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_728),
.B(n_624),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_731),
.Y(n_737)
);

INVx1_ASAP7_75t_SL g738 ( 
.A(n_729),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_726),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_733),
.Y(n_740)
);

AOI22xp5_ASAP7_75t_L g741 ( 
.A1(n_739),
.A2(n_625),
.B1(n_629),
.B2(n_634),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_738),
.B(n_126),
.Y(n_742)
);

HB1xp67_ASAP7_75t_L g743 ( 
.A(n_734),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_737),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_732),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_735),
.A2(n_629),
.B1(n_634),
.B2(n_624),
.Y(n_746)
);

AOI22xp5_ASAP7_75t_L g747 ( 
.A1(n_744),
.A2(n_736),
.B1(n_574),
.B2(n_633),
.Y(n_747)
);

INVx4_ASAP7_75t_L g748 ( 
.A(n_740),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_743),
.B(n_666),
.Y(n_749)
);

OAI22xp5_ASAP7_75t_L g750 ( 
.A1(n_745),
.A2(n_742),
.B1(n_741),
.B2(n_746),
.Y(n_750)
);

AOI22xp5_ASAP7_75t_L g751 ( 
.A1(n_750),
.A2(n_574),
.B1(n_542),
.B2(n_666),
.Y(n_751)
);

OAI22x1_ASAP7_75t_L g752 ( 
.A1(n_748),
.A2(n_747),
.B1(n_749),
.B2(n_574),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_751),
.A2(n_574),
.B1(n_526),
.B2(n_616),
.Y(n_753)
);

OAI21xp5_ASAP7_75t_L g754 ( 
.A1(n_753),
.A2(n_752),
.B(n_538),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_754),
.A2(n_611),
.B1(n_610),
.B2(n_616),
.Y(n_755)
);

OR2x6_ASAP7_75t_L g756 ( 
.A(n_755),
.B(n_127),
.Y(n_756)
);

AOI211xp5_ASAP7_75t_L g757 ( 
.A1(n_756),
.A2(n_128),
.B(n_130),
.C(n_132),
.Y(n_757)
);


endmodule