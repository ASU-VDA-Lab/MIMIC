module real_jpeg_30019_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_249;
wire n_78;
wire n_83;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_173;
wire n_105;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_268;
wire n_42;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_258;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_191;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_167;
wire n_213;
wire n_128;
wire n_179;
wire n_202;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_256;
wire n_101;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_0),
.A2(n_61),
.B1(n_62),
.B2(n_68),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_0),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_0),
.A2(n_58),
.B1(n_59),
.B2(n_68),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_0),
.A2(n_38),
.B1(n_39),
.B2(n_68),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_0),
.A2(n_25),
.B1(n_30),
.B2(n_68),
.Y(n_218)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_1),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_2),
.A2(n_38),
.B1(n_39),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_2),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_2),
.A2(n_25),
.B1(n_30),
.B2(n_48),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_2),
.A2(n_48),
.B1(n_58),
.B2(n_59),
.Y(n_111)
);

O2A1O1Ixp33_ASAP7_75t_SL g139 ( 
.A1(n_3),
.A2(n_57),
.B(n_62),
.C(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_3),
.Y(n_141)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_3),
.A2(n_61),
.B1(n_62),
.B2(n_141),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_3),
.B(n_55),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_3),
.B(n_38),
.Y(n_203)
);

A2O1A1O1Ixp25_ASAP7_75t_L g205 ( 
.A1(n_3),
.A2(n_38),
.B(n_42),
.C(n_203),
.D(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_3),
.B(n_72),
.Y(n_210)
);

OAI21xp33_ASAP7_75t_L g234 ( 
.A1(n_3),
.A2(n_24),
.B(n_216),
.Y(n_234)
);

A2O1A1O1Ixp25_ASAP7_75t_L g246 ( 
.A1(n_3),
.A2(n_59),
.B(n_71),
.C(n_152),
.D(n_247),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_3),
.B(n_59),
.Y(n_247)
);

BUFx12_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_5),
.A2(n_25),
.B1(n_30),
.B2(n_35),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_5),
.A2(n_35),
.B1(n_38),
.B2(n_39),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_8),
.A2(n_58),
.B1(n_59),
.B2(n_77),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_8),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_8),
.A2(n_38),
.B1(n_39),
.B2(n_77),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_8),
.A2(n_61),
.B1(n_62),
.B2(n_77),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g190 ( 
.A1(n_8),
.A2(n_25),
.B1(n_30),
.B2(n_77),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_9),
.A2(n_61),
.B1(n_62),
.B2(n_97),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_9),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_9),
.A2(n_58),
.B1(n_59),
.B2(n_97),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_9),
.A2(n_38),
.B1(n_39),
.B2(n_97),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_9),
.A2(n_25),
.B1(n_30),
.B2(n_97),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_10),
.A2(n_61),
.B1(n_62),
.B2(n_65),
.Y(n_64)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_10),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_10),
.A2(n_58),
.B1(n_59),
.B2(n_65),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_10),
.A2(n_25),
.B1(n_30),
.B2(n_65),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_10),
.A2(n_38),
.B1(n_39),
.B2(n_65),
.Y(n_250)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_11),
.B(n_38),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_11),
.A2(n_25),
.B1(n_30),
.B2(n_44),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_11),
.B(n_25),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_12),
.A2(n_25),
.B1(n_30),
.B2(n_31),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_12),
.A2(n_31),
.B1(n_38),
.B2(n_39),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_13),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_13),
.A2(n_40),
.B1(n_58),
.B2(n_59),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_13),
.A2(n_25),
.B1(n_30),
.B2(n_40),
.Y(n_146)
);

BUFx24_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_15),
.A2(n_58),
.B1(n_59),
.B2(n_73),
.Y(n_75)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_16),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_126),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_124),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_103),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_20),
.B(n_103),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_81),
.C(n_88),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_21),
.B(n_81),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_50),
.B1(n_51),
.B2(n_80),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_22),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_36),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_23),
.B(n_36),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_29),
.B1(n_32),
.B2(n_34),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_24),
.A2(n_32),
.B(n_34),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_24),
.A2(n_29),
.B1(n_32),
.B2(n_91),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_24),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_24),
.A2(n_146),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_24),
.A2(n_215),
.B(n_216),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_24),
.B(n_218),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_28),
.Y(n_24)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_28),
.A2(n_223),
.B(n_231),
.Y(n_230)
);

AOI32xp33_ASAP7_75t_L g202 ( 
.A1(n_30),
.A2(n_39),
.A3(n_44),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_30),
.B(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_32),
.Y(n_225)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_33),
.A2(n_92),
.B1(n_144),
.B2(n_145),
.Y(n_143)
);

INVx5_ASAP7_75t_SL g191 ( 
.A(n_33),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_33),
.B(n_217),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_33),
.A2(n_232),
.B(n_253),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.B1(n_47),
.B2(n_49),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_37),
.A2(n_41),
.B1(n_49),
.B2(n_94),
.Y(n_93)
);

O2A1O1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_43),
.B(n_45),
.C(n_46),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_38),
.A2(n_39),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

AOI32xp33_ASAP7_75t_L g254 ( 
.A1(n_38),
.A2(n_58),
.A3(n_247),
.B1(n_255),
.B2(n_256),
.Y(n_254)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp33_ASAP7_75t_SL g256 ( 
.A(n_39),
.B(n_74),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_41),
.A2(n_267),
.B(n_268),
.Y(n_266)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_42),
.A2(n_46),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_42),
.A2(n_46),
.B1(n_85),
.B2(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_42),
.B(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_42),
.A2(n_46),
.B1(n_249),
.B2(n_250),
.Y(n_248)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_47),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_49),
.A2(n_94),
.B(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_49),
.B(n_168),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_49),
.A2(n_166),
.B(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_49),
.B(n_141),
.Y(n_229)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_SL g51 ( 
.A(n_52),
.B(n_69),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_52),
.B(n_69),
.C(n_80),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_63),
.B(n_66),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_54),
.A2(n_55),
.B1(n_64),
.B2(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_54),
.B(n_67),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_54),
.A2(n_170),
.B(n_171),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_60),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_55),
.B(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_56),
.A2(n_57),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

OAI21xp33_ASAP7_75t_L g140 ( 
.A1(n_56),
.A2(n_59),
.B(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_61),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_66),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_76),
.B1(n_78),
.B2(n_79),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_70),
.A2(n_149),
.B(n_151),
.Y(n_148)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_71),
.B(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_71),
.A2(n_72),
.B1(n_110),
.B2(n_111),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_71),
.A2(n_72),
.B1(n_150),
.B2(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

INVx6_ASAP7_75t_L g255 ( 
.A(n_74),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_76),
.A2(n_78),
.B(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_78),
.B(n_102),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_78),
.A2(n_100),
.B(n_174),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_79),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_86),
.B2(n_87),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_87),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_86),
.A2(n_87),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_88),
.B(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_95),
.C(n_98),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_89),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_93),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_90),
.B(n_93),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_95),
.A2(n_98),
.B1(n_99),
.B2(n_131),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_95),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_96),
.Y(n_137)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_123),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_113),
.B1(n_114),
.B2(n_122),
.Y(n_104)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

OAI21xp33_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_109),
.B(n_112),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_109),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_121),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_119),
.B(n_120),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_118),
.A2(n_120),
.B(n_137),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_155),
.B(n_277),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_153),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_128),
.B(n_153),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_132),
.C(n_133),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_129),
.B(n_132),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_133),
.A2(n_134),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_138),
.C(n_147),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_135),
.A2(n_136),
.B1(n_147),
.B2(n_148),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_142),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_139),
.A2(n_142),
.B1(n_143),
.B2(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_139),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_141),
.B(n_237),
.Y(n_236)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_144),
.A2(n_222),
.B1(n_224),
.B2(n_225),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_195),
.Y(n_155)
);

INVxp33_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_178),
.B(n_194),
.Y(n_157)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_158),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_175),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_159),
.B(n_175),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_162),
.C(n_163),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_163),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_169),
.C(n_172),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_164),
.A2(n_165),
.B1(n_172),
.B2(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_169),
.B(n_183),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_172),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_176),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_179),
.B(n_181),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_185),
.C(n_187),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_182),
.B(n_273),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_185),
.B(n_187),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.C(n_192),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_188),
.B(n_262),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_189),
.A2(n_192),
.B1(n_193),
.B2(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_189),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_190),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

NOR3xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_275),
.C(n_276),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_270),
.B(n_274),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_258),
.B(n_269),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_242),
.B(n_257),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_200),
.A2(n_219),
.B(n_241),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_207),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_201),
.B(n_207),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_205),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_205),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_206),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_214),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_211),
.B2(n_212),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_209),
.B(n_212),
.C(n_214),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_213),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_215),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_227),
.B(n_240),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_226),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_221),
.B(n_226),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_233),
.B(n_239),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_229),
.B(n_230),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_243),
.B(n_244),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_251),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_248),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_248),
.C(n_251),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_250),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_254),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_254),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_259),
.B(n_260),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_264),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_265),
.C(n_266),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_271),
.B(n_272),
.Y(n_274)
);


endmodule