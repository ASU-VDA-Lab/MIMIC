module real_aes_3710_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_977;
wire n_943;
wire n_287;
wire n_635;
wire n_357;
wire n_503;
wire n_386;
wire n_905;
wire n_673;
wire n_518;
wire n_254;
wire n_792;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_979;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_974;
wire n_132;
wire n_857;
wire n_919;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_952;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_963;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_955;
wire n_889;
wire n_975;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_958;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_961;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_953;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_121;
wire n_352;
wire n_935;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_951;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_931;
wire n_780;
wire n_174;
wire n_904;
wire n_570;
wire n_675;
wire n_840;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_962;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_656;
wire n_153;
wire n_316;
wire n_532;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_119;
wire n_725;
wire n_455;
wire n_504;
wire n_960;
wire n_164;
wire n_671;
wire n_973;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_950;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_142;
wire n_970;
wire n_947;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_964;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_917;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_957;
wire n_296;
wire n_702;
wire n_954;
wire n_969;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_945;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_133;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_965;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_972;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_978;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_899;
wire n_243;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_926;
wire n_922;
wire n_149;
wire n_942;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_959;
wire n_715;
wire n_134;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_639;
wire n_587;
wire n_546;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_888;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_967;
wire n_566;
wire n_719;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_175;
wire n_168;
wire n_241;
wire n_687;
wire n_844;
wire n_968;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_554;
wire n_475;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_668;
wire n_237;
wire n_797;
wire n_862;
INVx1_ASAP7_75t_L g702 ( .A(n_0), .Y(n_702) );
OAI22x1_ASAP7_75t_SL g114 ( .A1(n_1), .A2(n_54), .B1(n_115), .B2(n_116), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_1), .Y(n_116) );
AOI22xp5_ASAP7_75t_L g127 ( .A1(n_2), .A2(n_21), .B1(n_128), .B2(n_131), .Y(n_127) );
INVx1_ASAP7_75t_L g272 ( .A(n_3), .Y(n_272) );
AOI22xp33_ASAP7_75t_L g105 ( .A1(n_4), .A2(n_106), .B1(n_970), .B2(n_979), .Y(n_105) );
INVx2_ASAP7_75t_L g298 ( .A(n_5), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_6), .B(n_601), .Y(n_658) );
INVx1_ASAP7_75t_SL g248 ( .A(n_7), .Y(n_248) );
INVxp67_ASAP7_75t_L g551 ( .A(n_8), .Y(n_551) );
INVx1_ASAP7_75t_L g582 ( .A(n_8), .Y(n_582) );
BUFx2_ASAP7_75t_L g586 ( .A(n_8), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g659 ( .A(n_9), .B(n_205), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_10), .A2(n_44), .B1(n_600), .B2(n_645), .Y(n_644) );
AOI22xp5_ASAP7_75t_L g725 ( .A1(n_11), .A2(n_50), .B1(n_192), .B2(n_619), .Y(n_725) );
XOR2xp5_ASAP7_75t_R g571 ( .A(n_12), .B(n_572), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g686 ( .A1(n_13), .A2(n_71), .B1(n_680), .B2(n_681), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_14), .B(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_15), .B(n_209), .Y(n_208) );
INVx1_ASAP7_75t_L g697 ( .A(n_16), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_17), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g536 ( .A(n_17), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g203 ( .A1(n_18), .A2(n_59), .B1(n_204), .B2(n_205), .Y(n_203) );
INVx1_ASAP7_75t_L g700 ( .A(n_19), .Y(n_700) );
OA21x2_ASAP7_75t_L g143 ( .A1(n_20), .A2(n_76), .B(n_144), .Y(n_143) );
OA21x2_ASAP7_75t_L g150 ( .A1(n_20), .A2(n_76), .B(n_144), .Y(n_150) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_22), .A2(n_74), .B1(n_680), .B2(n_681), .Y(n_679) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_23), .B(n_129), .Y(n_159) );
AOI22xp5_ASAP7_75t_L g292 ( .A1(n_24), .A2(n_86), .B1(n_293), .B2(n_294), .Y(n_292) );
INVx2_ASAP7_75t_L g197 ( .A(n_25), .Y(n_197) );
CKINVDCx5p33_ASAP7_75t_R g583 ( .A(n_26), .Y(n_583) );
OAI22xp5_ASAP7_75t_R g570 ( .A1(n_27), .A2(n_571), .B1(n_575), .B2(n_576), .Y(n_570) );
CKINVDCx5p33_ASAP7_75t_R g575 ( .A(n_27), .Y(n_575) );
INVx1_ASAP7_75t_L g694 ( .A(n_28), .Y(n_694) );
AOI22xp5_ASAP7_75t_L g134 ( .A1(n_29), .A2(n_33), .B1(n_135), .B2(n_137), .Y(n_134) );
BUFx3_ASAP7_75t_L g109 ( .A(n_30), .Y(n_109) );
O2A1O1Ixp5_ASAP7_75t_L g191 ( .A1(n_31), .A2(n_132), .B(n_192), .C(n_194), .Y(n_191) );
AOI22xp33_ASAP7_75t_L g296 ( .A1(n_32), .A2(n_68), .B1(n_157), .B2(n_193), .Y(n_296) );
CKINVDCx5p33_ASAP7_75t_R g234 ( .A(n_34), .Y(n_234) );
AO22x1_ASAP7_75t_L g655 ( .A1(n_35), .A2(n_84), .B1(n_252), .B2(n_656), .Y(n_655) );
CKINVDCx5p33_ASAP7_75t_R g604 ( .A(n_36), .Y(n_604) );
AND2x2_ASAP7_75t_L g618 ( .A(n_37), .B(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_38), .B(n_252), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g211 ( .A1(n_39), .A2(n_87), .B1(n_212), .B2(n_215), .Y(n_211) );
INVx1_ASAP7_75t_L g556 ( .A(n_40), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g975 ( .A(n_40), .B(n_85), .Y(n_975) );
INVx1_ASAP7_75t_L g185 ( .A(n_41), .Y(n_185) );
AOI22x1_ASAP7_75t_L g727 ( .A1(n_42), .A2(n_101), .B1(n_641), .B2(n_680), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_43), .B(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g977 ( .A(n_45), .B(n_978), .Y(n_977) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_46), .B(n_181), .Y(n_267) );
INVx2_ASAP7_75t_L g195 ( .A(n_47), .Y(n_195) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_48), .Y(n_236) );
NAND2xp5_ASAP7_75t_SL g627 ( .A(n_49), .B(n_628), .Y(n_627) );
INVx2_ASAP7_75t_L g158 ( .A(n_51), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_52), .B(n_265), .Y(n_264) );
INVx1_ASAP7_75t_SL g251 ( .A(n_53), .Y(n_251) );
INVx1_ASAP7_75t_L g115 ( .A(n_54), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_55), .B(n_137), .Y(n_670) );
INVx1_ASAP7_75t_L g229 ( .A(n_56), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_57), .B(n_187), .Y(n_607) );
INVx1_ASAP7_75t_L g144 ( .A(n_58), .Y(n_144) );
AND2x4_ASAP7_75t_L g146 ( .A(n_60), .B(n_147), .Y(n_146) );
AND2x4_ASAP7_75t_L g189 ( .A(n_60), .B(n_147), .Y(n_189) );
INVx1_ASAP7_75t_L g255 ( .A(n_61), .Y(n_255) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_62), .Y(n_133) );
INVx2_ASAP7_75t_L g683 ( .A(n_63), .Y(n_683) );
AOI22xp5_ASAP7_75t_L g572 ( .A1(n_64), .A2(n_102), .B1(n_573), .B2(n_574), .Y(n_572) );
INVx1_ASAP7_75t_L g574 ( .A(n_64), .Y(n_574) );
AOI22xp33_ASAP7_75t_L g640 ( .A1(n_65), .A2(n_79), .B1(n_600), .B2(n_641), .Y(n_640) );
CKINVDCx14_ASAP7_75t_R g661 ( .A(n_66), .Y(n_661) );
AND2x2_ASAP7_75t_L g625 ( .A(n_67), .B(n_252), .Y(n_625) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_69), .B(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_70), .B(n_265), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_72), .B(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_73), .B(n_259), .Y(n_664) );
NAND2x1p5_ASAP7_75t_L g629 ( .A(n_75), .B(n_613), .Y(n_629) );
CKINVDCx14_ASAP7_75t_R g543 ( .A(n_77), .Y(n_543) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_78), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g183 ( .A(n_80), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_81), .B(n_601), .Y(n_668) );
OR2x6_ASAP7_75t_L g553 ( .A(n_82), .B(n_554), .Y(n_553) );
NAND3xp33_ASAP7_75t_L g976 ( .A(n_82), .B(n_551), .C(n_977), .Y(n_976) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_83), .B(n_138), .Y(n_253) );
INVx1_ASAP7_75t_L g555 ( .A(n_85), .Y(n_555) );
INVx1_ASAP7_75t_L g978 ( .A(n_88), .Y(n_978) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_89), .Y(n_130) );
BUFx5_ASAP7_75t_L g136 ( .A(n_89), .Y(n_136) );
INVx1_ASAP7_75t_L g165 ( .A(n_89), .Y(n_165) );
INVx2_ASAP7_75t_L g704 ( .A(n_90), .Y(n_704) );
NOR2xp33_ASAP7_75t_L g249 ( .A(n_91), .B(n_167), .Y(n_249) );
OAI22xp5_ASAP7_75t_L g542 ( .A1(n_92), .A2(n_543), .B1(n_544), .B2(n_545), .Y(n_542) );
INVx1_ASAP7_75t_L g544 ( .A(n_92), .Y(n_544) );
INVx2_ASAP7_75t_L g162 ( .A(n_93), .Y(n_162) );
INVx1_ASAP7_75t_L g172 ( .A(n_94), .Y(n_172) );
NAND2xp33_ASAP7_75t_L g621 ( .A(n_95), .B(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g238 ( .A(n_96), .Y(n_238) );
INVx2_ASAP7_75t_SL g147 ( .A(n_97), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_98), .B(n_227), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_99), .B(n_628), .Y(n_667) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_100), .B(n_259), .Y(n_258) );
CKINVDCx5p33_ASAP7_75t_R g573 ( .A(n_102), .Y(n_573) );
AO32x2_ASAP7_75t_L g125 ( .A1(n_103), .A2(n_126), .A3(n_141), .B1(n_145), .B2(n_148), .Y(n_125) );
AO22x2_ASAP7_75t_L g309 ( .A1(n_103), .A2(n_126), .B1(n_310), .B2(n_312), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_104), .B(n_611), .Y(n_610) );
OA21x2_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_110), .B(n_565), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
HB1xp67_ASAP7_75t_L g567 ( .A(n_109), .Y(n_567) );
OAI21xp5_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_540), .B(n_557), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVxp67_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AOI21xp33_ASAP7_75t_SL g557 ( .A1(n_113), .A2(n_558), .B(n_561), .Y(n_557) );
XNOR2x1_ASAP7_75t_L g113 ( .A(n_114), .B(n_117), .Y(n_113) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_117), .A2(n_585), .B1(n_587), .B2(n_966), .Y(n_584) );
OR2x2_ASAP7_75t_L g117 ( .A(n_118), .B(n_533), .Y(n_117) );
NOR3xp33_ASAP7_75t_L g118 ( .A(n_119), .B(n_407), .C(n_465), .Y(n_118) );
OAI21xp5_ASAP7_75t_L g534 ( .A1(n_119), .A2(n_535), .B(n_536), .Y(n_534) );
NAND4xp75_ASAP7_75t_L g119 ( .A(n_120), .B(n_324), .C(n_355), .D(n_388), .Y(n_119) );
AND2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_299), .Y(n_120) );
AOI22xp5_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_198), .B1(n_274), .B2(n_280), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OR2x2_ASAP7_75t_L g123 ( .A(n_124), .B(n_151), .Y(n_123) );
BUFx3_ASAP7_75t_L g338 ( .A(n_124), .Y(n_338) );
AND2x4_ASAP7_75t_L g348 ( .A(n_124), .B(n_349), .Y(n_348) );
AND2x2_ASAP7_75t_L g371 ( .A(n_124), .B(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_SL g385 ( .A(n_124), .B(n_152), .Y(n_385) );
AND2x2_ASAP7_75t_L g454 ( .A(n_124), .B(n_426), .Y(n_454) );
AND2x2_ASAP7_75t_L g493 ( .A(n_124), .B(n_401), .Y(n_493) );
BUFx8_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx2_ASAP7_75t_L g282 ( .A(n_125), .Y(n_282) );
AND2x2_ASAP7_75t_L g483 ( .A(n_125), .B(n_484), .Y(n_483) );
OAI22xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_132), .B1(n_134), .B2(n_139), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_128), .B(n_195), .Y(n_194) );
INVx2_ASAP7_75t_SL g128 ( .A(n_129), .Y(n_128) );
INVx1_ASAP7_75t_L g157 ( .A(n_129), .Y(n_157) );
INVx2_ASAP7_75t_L g179 ( .A(n_129), .Y(n_179) );
INVx2_ASAP7_75t_L g235 ( .A(n_129), .Y(n_235) );
INVx1_ASAP7_75t_L g622 ( .A(n_129), .Y(n_622) );
INVx1_ASAP7_75t_L g628 ( .A(n_129), .Y(n_628) );
INVx6_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g131 ( .A(n_130), .Y(n_131) );
INVx3_ASAP7_75t_L g138 ( .A(n_130), .Y(n_138) );
INVx2_ASAP7_75t_L g214 ( .A(n_130), .Y(n_214) );
INVx2_ASAP7_75t_L g187 ( .A(n_131), .Y(n_187) );
INVxp67_ASAP7_75t_SL g215 ( .A(n_131), .Y(n_215) );
INVx4_ASAP7_75t_L g232 ( .A(n_132), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_132), .A2(n_262), .B(n_264), .Y(n_261) );
OAI22xp5_ASAP7_75t_L g599 ( .A1(n_132), .A2(n_600), .B1(n_602), .B2(n_605), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_132), .B(n_639), .Y(n_638) );
AOI21xp5_ASAP7_75t_L g666 ( .A1(n_132), .A2(n_667), .B(n_668), .Y(n_666) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_133), .Y(n_140) );
INVx3_ASAP7_75t_L g160 ( .A(n_133), .Y(n_160) );
INVx4_ASAP7_75t_L g182 ( .A(n_133), .Y(n_182) );
INVx1_ASAP7_75t_L g217 ( .A(n_133), .Y(n_217) );
INVxp67_ASAP7_75t_L g623 ( .A(n_133), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_133), .B(n_694), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_133), .B(n_697), .Y(n_696) );
OAI22xp33_ASAP7_75t_L g233 ( .A1(n_135), .A2(n_234), .B1(n_235), .B2(n_236), .Y(n_233) );
INVx2_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx2_ASAP7_75t_L g204 ( .A(n_136), .Y(n_204) );
INVx2_ASAP7_75t_L g252 ( .A(n_136), .Y(n_252) );
INVx2_ASAP7_75t_L g265 ( .A(n_136), .Y(n_265) );
INVx1_ASAP7_75t_L g269 ( .A(n_136), .Y(n_269) );
INVx2_ASAP7_75t_L g601 ( .A(n_136), .Y(n_601) );
INVx1_ASAP7_75t_L g247 ( .A(n_137), .Y(n_247) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx1_ASAP7_75t_L g205 ( .A(n_138), .Y(n_205) );
INVx1_ASAP7_75t_L g263 ( .A(n_138), .Y(n_263) );
INVx2_ASAP7_75t_L g294 ( .A(n_138), .Y(n_294) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
A2O1A1Ixp33_ASAP7_75t_L g161 ( .A1(n_140), .A2(n_162), .B(n_163), .C(n_166), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_140), .B(n_207), .Y(n_206) );
A2O1A1Ixp33_ASAP7_75t_L g246 ( .A1(n_140), .A2(n_247), .B(n_248), .C(n_249), .Y(n_246) );
INVx1_ASAP7_75t_L g295 ( .A(n_140), .Y(n_295) );
INVxp67_ASAP7_75t_L g609 ( .A(n_140), .Y(n_609) );
INVx2_ASAP7_75t_SL g631 ( .A(n_140), .Y(n_631) );
INVx1_ASAP7_75t_L g672 ( .A(n_140), .Y(n_672) );
AO31x2_ASAP7_75t_L g175 ( .A1(n_141), .A2(n_176), .A3(n_190), .B(n_196), .Y(n_175) );
INVx2_ASAP7_75t_L g312 ( .A(n_141), .Y(n_312) );
BUFx3_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
NOR2xp33_ASAP7_75t_L g196 ( .A(n_142), .B(n_197), .Y(n_196) );
INVx3_ASAP7_75t_L g259 ( .A(n_142), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_142), .B(n_298), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_142), .B(n_704), .Y(n_703) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx4_ASAP7_75t_L g245 ( .A(n_143), .Y(n_245) );
BUFx3_ASAP7_75t_L g305 ( .A(n_143), .Y(n_305) );
OAI21x1_ASAP7_75t_L g598 ( .A1(n_145), .A2(n_599), .B(n_606), .Y(n_598) );
AO31x2_ASAP7_75t_L g723 ( .A1(n_145), .A2(n_724), .A3(n_728), .B(n_729), .Y(n_723) );
AO31x2_ASAP7_75t_L g742 ( .A1(n_145), .A2(n_724), .A3(n_728), .B(n_729), .Y(n_742) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx3_ASAP7_75t_L g170 ( .A(n_146), .Y(n_170) );
AND2x2_ASAP7_75t_L g289 ( .A(n_146), .B(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g310 ( .A(n_146), .B(n_311), .Y(n_310) );
INVx3_ASAP7_75t_L g634 ( .A(n_146), .Y(n_634) );
INVx1_ASAP7_75t_L g653 ( .A(n_146), .Y(n_653) );
INVxp67_ASAP7_75t_L g219 ( .A(n_148), .Y(n_219) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_149), .B(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g169 ( .A(n_150), .B(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g173 ( .A(n_150), .Y(n_173) );
NOR2xp67_ASAP7_75t_L g207 ( .A(n_150), .B(n_170), .Y(n_207) );
BUFx3_ASAP7_75t_L g209 ( .A(n_150), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g273 ( .A(n_150), .B(n_170), .Y(n_273) );
INVx1_ASAP7_75t_L g311 ( .A(n_150), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_150), .B(n_170), .Y(n_639) );
INVx2_ASAP7_75t_L g678 ( .A(n_150), .Y(n_678) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g485 ( .A(n_152), .Y(n_485) );
AND2x2_ASAP7_75t_L g515 ( .A(n_152), .B(n_315), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_152), .B(n_435), .Y(n_522) );
AND2x4_ASAP7_75t_L g152 ( .A(n_153), .B(n_174), .Y(n_152) );
AND2x4_ASAP7_75t_L g281 ( .A(n_153), .B(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g307 ( .A(n_153), .B(n_175), .Y(n_307) );
INVx2_ASAP7_75t_L g319 ( .A(n_153), .Y(n_319) );
INVx1_ASAP7_75t_L g361 ( .A(n_153), .Y(n_361) );
BUFx3_ASAP7_75t_L g396 ( .A(n_153), .Y(n_396) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AO31x2_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_161), .A3(n_169), .B(n_171), .Y(n_154) );
A2O1A1Ixp33_ASAP7_75t_L g155 ( .A1(n_156), .A2(n_158), .B(n_159), .C(n_160), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx3_ASAP7_75t_L g225 ( .A(n_160), .Y(n_225) );
A2O1A1Ixp33_ASAP7_75t_L g250 ( .A1(n_160), .A2(n_251), .B(n_252), .C(n_253), .Y(n_250) );
NOR2xp67_ASAP7_75t_L g222 ( .A(n_163), .B(n_223), .Y(n_222) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g293 ( .A(n_164), .Y(n_293) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g168 ( .A(n_165), .Y(n_168) );
INVx1_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g193 ( .A(n_168), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_170), .B(n_244), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_172), .B(n_173), .Y(n_171) );
NOR2xp33_ASAP7_75t_SL g254 ( .A(n_173), .B(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g647 ( .A(n_173), .Y(n_647) );
INVx1_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_175), .B(n_332), .Y(n_331) );
INVx2_ASAP7_75t_L g350 ( .A(n_175), .Y(n_350) );
OR2x2_ASAP7_75t_L g364 ( .A(n_175), .B(n_332), .Y(n_364) );
AND2x2_ASAP7_75t_L g426 ( .A(n_175), .B(n_319), .Y(n_426) );
AOI221x1_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_180), .B1(n_184), .B2(n_186), .C(n_188), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AND2x2_ASAP7_75t_L g180 ( .A(n_181), .B(n_183), .Y(n_180) );
AND2x2_ASAP7_75t_L g184 ( .A(n_181), .B(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_182), .B(n_272), .Y(n_271) );
NAND3xp33_ASAP7_75t_SL g677 ( .A(n_182), .B(n_633), .C(n_678), .Y(n_677) );
NOR2xp33_ASAP7_75t_SL g699 ( .A(n_182), .B(n_700), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g701 ( .A(n_182), .B(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_187), .B(n_696), .Y(n_695) );
AOI22xp5_ASAP7_75t_L g698 ( .A1(n_187), .A2(n_252), .B1(n_699), .B2(n_701), .Y(n_698) );
NOR2xp33_ASAP7_75t_L g224 ( .A(n_188), .B(n_225), .Y(n_224) );
NOR3xp33_ASAP7_75t_L g228 ( .A(n_188), .B(n_225), .C(n_229), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_188), .B(n_232), .Y(n_231) );
INVx4_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx1_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx3_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
AND2x4_ASAP7_75t_L g198 ( .A(n_199), .B(n_239), .Y(n_198) );
AND2x2_ASAP7_75t_L g448 ( .A(n_199), .B(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g512 ( .A(n_199), .B(n_392), .Y(n_512) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_218), .Y(n_199) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_200), .Y(n_342) );
AND2x2_ASAP7_75t_L g437 ( .A(n_200), .B(n_438), .Y(n_437) );
BUFx2_ASAP7_75t_L g457 ( .A(n_200), .Y(n_457) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g279 ( .A(n_201), .Y(n_279) );
AND2x2_ASAP7_75t_L g301 ( .A(n_201), .B(n_257), .Y(n_301) );
INVx1_ASAP7_75t_L g368 ( .A(n_201), .Y(n_368) );
AND2x2_ASAP7_75t_L g375 ( .A(n_201), .B(n_345), .Y(n_375) );
NAND2x1p5_ASAP7_75t_L g201 ( .A(n_202), .B(n_210), .Y(n_201) );
AND2x2_ASAP7_75t_SL g422 ( .A(n_202), .B(n_210), .Y(n_422) );
OA21x2_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_206), .B(n_208), .Y(n_202) );
INVx2_ASAP7_75t_L g680 ( .A(n_204), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_207), .B(n_217), .Y(n_216) );
OR2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_216), .Y(n_210) );
INVx1_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g227 ( .A(n_214), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_217), .B(n_639), .Y(n_643) );
INVx1_ASAP7_75t_L g726 ( .A(n_217), .Y(n_726) );
AND2x2_ASAP7_75t_L g322 ( .A(n_218), .B(n_323), .Y(n_322) );
OR2x2_ASAP7_75t_L g344 ( .A(n_218), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g369 ( .A(n_218), .B(n_242), .Y(n_369) );
AND2x2_ASAP7_75t_L g514 ( .A(n_218), .B(n_421), .Y(n_514) );
AO21x2_ASAP7_75t_L g218 ( .A1(n_219), .A2(n_220), .B(n_237), .Y(n_218) );
AO21x2_ASAP7_75t_L g303 ( .A1(n_220), .A2(n_237), .B(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_221), .B(n_230), .Y(n_220) );
AOI22xp5_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_224), .B1(n_226), .B2(n_228), .Y(n_221) );
OAI22xp5_ASAP7_75t_L g291 ( .A1(n_225), .A2(n_292), .B1(n_295), .B2(n_296), .Y(n_291) );
NAND3xp33_ASAP7_75t_L g685 ( .A(n_225), .B(n_633), .C(n_678), .Y(n_685) );
INVx1_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_231), .B(n_233), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_232), .B(n_603), .Y(n_602) );
OAI22x1_ASAP7_75t_L g724 ( .A1(n_232), .A2(n_725), .B1(n_726), .B2(n_727), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_235), .B(n_271), .Y(n_270) );
INVx2_ASAP7_75t_L g619 ( .A(n_235), .Y(n_619) );
AND2x2_ASAP7_75t_L g239 ( .A(n_240), .B(n_256), .Y(n_239) );
AND2x2_ASAP7_75t_L g321 ( .A(n_240), .B(n_279), .Y(n_321) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_240), .Y(n_327) );
INVx2_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx2_ASAP7_75t_L g285 ( .A(n_242), .Y(n_285) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_242), .Y(n_347) );
OR2x2_ASAP7_75t_L g381 ( .A(n_242), .B(n_303), .Y(n_381) );
INVx2_ASAP7_75t_L g393 ( .A(n_242), .Y(n_393) );
INVx1_ASAP7_75t_L g450 ( .A(n_242), .Y(n_450) );
AO31x2_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_246), .A3(n_250), .B(n_254), .Y(n_242) );
INVx2_ASAP7_75t_L g290 ( .A(n_244), .Y(n_290) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx3_ASAP7_75t_L g613 ( .A(n_245), .Y(n_613) );
INVx1_ASAP7_75t_L g463 ( .A(n_256), .Y(n_463) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
INVx1_ASAP7_75t_L g277 ( .A(n_257), .Y(n_277) );
INVx1_ASAP7_75t_L g323 ( .A(n_257), .Y(n_323) );
INVx2_ASAP7_75t_L g345 ( .A(n_257), .Y(n_345) );
AND2x2_ASAP7_75t_L g392 ( .A(n_257), .B(n_393), .Y(n_392) );
AND2x4_ASAP7_75t_L g257 ( .A(n_258), .B(n_260), .Y(n_257) );
NOR2x1_ASAP7_75t_L g673 ( .A(n_259), .B(n_634), .Y(n_673) );
OAI21xp5_ASAP7_75t_L g260 ( .A1(n_261), .A2(n_266), .B(n_273), .Y(n_260) );
OAI21xp5_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_268), .B(n_270), .Y(n_266) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVxp67_ASAP7_75t_SL g274 ( .A(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_276), .B(n_278), .Y(n_275) );
INVx2_ASAP7_75t_L g328 ( .A(n_276), .Y(n_328) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g497 ( .A(n_277), .B(n_422), .Y(n_497) );
INVx1_ASAP7_75t_L g507 ( .A(n_278), .Y(n_507) );
BUFx3_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g280 ( .A(n_281), .B(n_283), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_281), .B(n_316), .Y(n_474) );
INVx2_ASAP7_75t_L g490 ( .A(n_281), .Y(n_490) );
AND2x2_ASAP7_75t_L g510 ( .A(n_281), .B(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g400 ( .A(n_282), .B(n_401), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_282), .B(n_350), .Y(n_461) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
AND2x2_ASAP7_75t_L g336 ( .A(n_285), .B(n_303), .Y(n_336) );
INVxp67_ASAP7_75t_SL g477 ( .A(n_285), .Y(n_477) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_285), .Y(n_525) );
AND2x2_ASAP7_75t_L g373 ( .A(n_286), .B(n_360), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_286), .B(n_401), .Y(n_429) );
BUFx3_ASAP7_75t_L g446 ( .A(n_286), .Y(n_446) );
AND2x2_ASAP7_75t_L g464 ( .A(n_286), .B(n_426), .Y(n_464) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
HB1xp67_ASAP7_75t_L g335 ( .A(n_287), .Y(n_335) );
AND2x2_ASAP7_75t_L g349 ( .A(n_287), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g492 ( .A(n_287), .B(n_319), .Y(n_492) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g317 ( .A(n_288), .Y(n_317) );
INVx1_ASAP7_75t_L g332 ( .A(n_288), .Y(n_332) );
AOI21x1_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_291), .B(n_297), .Y(n_288) );
AOI21xp33_ASAP7_75t_SL g632 ( .A1(n_290), .A2(n_633), .B(n_635), .Y(n_632) );
INVx2_ASAP7_75t_L g656 ( .A(n_293), .Y(n_656) );
INVx1_ASAP7_75t_L g645 ( .A(n_294), .Y(n_645) );
INVx1_ASAP7_75t_L g681 ( .A(n_294), .Y(n_681) );
AOI21x1_ASAP7_75t_L g654 ( .A1(n_295), .A2(n_655), .B(n_657), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g299 ( .A1(n_300), .A2(n_306), .B1(n_313), .B2(n_320), .Y(n_299) );
NAND2x1p5_ASAP7_75t_L g352 ( .A(n_300), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
INVx1_ASAP7_75t_L g339 ( .A(n_301), .Y(n_339) );
AND2x2_ASAP7_75t_L g346 ( .A(n_301), .B(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g427 ( .A(n_301), .B(n_369), .Y(n_427) );
AND2x2_ASAP7_75t_L g518 ( .A(n_301), .B(n_336), .Y(n_518) );
INVx2_ASAP7_75t_L g417 ( .A(n_302), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_302), .B(n_375), .Y(n_469) );
BUFx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx2_ASAP7_75t_L g438 ( .A(n_303), .Y(n_438) );
OR2x2_ASAP7_75t_L g660 ( .A(n_304), .B(n_661), .Y(n_660) );
NOR2xp67_ASAP7_75t_SL g729 ( .A(n_304), .B(n_543), .Y(n_729) );
INVx3_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
OA21x2_ASAP7_75t_L g597 ( .A1(n_305), .A2(n_598), .B(n_610), .Y(n_597) );
OA21x2_ASAP7_75t_L g713 ( .A1(n_305), .A2(n_598), .B(n_610), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_306), .B(n_480), .Y(n_479) );
AND2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
NAND2x1p5_ASAP7_75t_L g354 ( .A(n_307), .B(n_315), .Y(n_354) );
INVx2_ASAP7_75t_L g403 ( .A(n_307), .Y(n_403) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x4_ASAP7_75t_L g318 ( .A(n_309), .B(n_319), .Y(n_318) );
INVx1_ASAP7_75t_L g362 ( .A(n_309), .Y(n_362) );
AND2x4_ASAP7_75t_L g395 ( .A(n_309), .B(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g435 ( .A(n_309), .B(n_332), .Y(n_435) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_318), .Y(n_314) );
AND2x4_ASAP7_75t_L g399 ( .A(n_315), .B(n_400), .Y(n_399) );
INVx4_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g425 ( .A(n_316), .B(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g511 ( .A(n_316), .Y(n_511) );
BUFx3_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g484 ( .A(n_317), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_318), .B(n_330), .Y(n_329) );
INVx4_ASAP7_75t_L g423 ( .A(n_318), .Y(n_423) );
AND2x4_ASAP7_75t_L g471 ( .A(n_318), .B(n_472), .Y(n_471) );
AND2x4_ASAP7_75t_L g503 ( .A(n_318), .B(n_363), .Y(n_503) );
AOI22xp5_ASAP7_75t_L g424 ( .A1(n_320), .A2(n_425), .B1(n_427), .B2(n_428), .Y(n_424) );
AND2x4_ASAP7_75t_L g320 ( .A(n_321), .B(n_322), .Y(n_320) );
AND2x2_ASAP7_75t_L g413 ( .A(n_321), .B(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g449 ( .A(n_323), .B(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g506 ( .A(n_323), .Y(n_506) );
NOR3x1_ASAP7_75t_L g324 ( .A(n_325), .B(n_340), .C(n_351), .Y(n_324) );
OAI21xp5_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_329), .B(n_333), .Y(n_325) );
NOR3xp33_ASAP7_75t_L g415 ( .A(n_326), .B(n_416), .C(n_420), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
AND2x2_ASAP7_75t_L g440 ( .A(n_330), .B(n_423), .Y(n_440) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g372 ( .A(n_331), .Y(n_372) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_332), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_334), .B(n_337), .Y(n_333) );
AND2x4_ASAP7_75t_L g334 ( .A(n_335), .B(n_336), .Y(n_334) );
NAND2x1p5_ASAP7_75t_L g442 ( .A(n_336), .B(n_443), .Y(n_442) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_338), .B(n_339), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g523 ( .A(n_339), .B(n_524), .Y(n_523) );
OA21x2_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_346), .B(n_348), .Y(n_340) );
AND2x4_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
INVxp67_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g414 ( .A(n_344), .Y(n_414) );
OR2x6_ASAP7_75t_L g476 ( .A(n_344), .B(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g453 ( .A(n_349), .B(n_360), .Y(n_453) );
INVx2_ASAP7_75t_SL g401 ( .A(n_350), .Y(n_401) );
INVx1_ASAP7_75t_L g419 ( .A(n_350), .Y(n_419) );
BUFx3_ASAP7_75t_L g472 ( .A(n_350), .Y(n_472) );
INVxp67_ASAP7_75t_SL g351 ( .A(n_352), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_353), .A2(n_505), .B1(n_528), .B2(n_530), .Y(n_527) );
INVx3_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
NOR2x1_ASAP7_75t_L g355 ( .A(n_356), .B(n_376), .Y(n_355) );
OAI21xp5_ASAP7_75t_SL g356 ( .A1(n_357), .A2(n_365), .B(n_370), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_360), .B(n_363), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g434 ( .A(n_360), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g447 ( .A(n_360), .Y(n_447) );
AND2x4_ASAP7_75t_SL g360 ( .A(n_361), .B(n_362), .Y(n_360) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
OAI22xp5_ASAP7_75t_L g473 ( .A1(n_364), .A2(n_474), .B1(n_475), .B2(n_476), .Y(n_473) );
OAI21xp5_ASAP7_75t_SL g489 ( .A1(n_364), .A2(n_490), .B(n_491), .Y(n_489) );
INVx2_ASAP7_75t_L g532 ( .A(n_364), .Y(n_532) );
INVx1_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_367), .B(n_369), .Y(n_366) );
OR2x2_ASAP7_75t_L g387 ( .A(n_367), .B(n_381), .Y(n_387) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g391 ( .A(n_368), .B(n_392), .Y(n_391) );
AND2x2_ASAP7_75t_L g374 ( .A(n_369), .B(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g456 ( .A(n_369), .B(n_457), .Y(n_456) );
OAI21xp33_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_373), .B(n_374), .Y(n_370) );
INVxp67_ASAP7_75t_SL g377 ( .A(n_373), .Y(n_377) );
BUFx3_ASAP7_75t_L g383 ( .A(n_375), .Y(n_383) );
NAND2xp67_ASAP7_75t_L g405 ( .A(n_375), .B(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_375), .B(n_417), .Y(n_475) );
OAI21xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_378), .B(n_384), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_379), .B(n_382), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx2_ASAP7_75t_L g406 ( .A(n_381), .Y(n_406) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
OA21x2_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_394), .B(n_398), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AOI22xp5_ASAP7_75t_L g458 ( .A1(n_390), .A2(n_459), .B1(n_462), .B2(n_464), .Y(n_458) );
BUFx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g470 ( .A(n_391), .Y(n_470) );
AND2x2_ASAP7_75t_L g436 ( .A(n_392), .B(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g496 ( .A(n_393), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_395), .B(n_397), .Y(n_394) );
INVx2_ASAP7_75t_L g433 ( .A(n_395), .Y(n_433) );
OAI21xp33_ASAP7_75t_L g445 ( .A1(n_395), .A2(n_446), .B(n_447), .Y(n_445) );
NAND3xp33_ASAP7_75t_L g504 ( .A(n_395), .B(n_505), .C(n_507), .Y(n_504) );
AND2x2_ASAP7_75t_L g526 ( .A(n_395), .B(n_511), .Y(n_526) );
INVx2_ASAP7_75t_SL g531 ( .A(n_396), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_397), .B(n_421), .Y(n_420) );
OR2x2_ASAP7_75t_L g460 ( .A(n_397), .B(n_461), .Y(n_460) );
OAI21xp33_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_402), .B(n_404), .Y(n_398) );
INVx1_ASAP7_75t_L g412 ( .A(n_401), .Y(n_412) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g538 ( .A(n_408), .Y(n_538) );
NOR3x1_ASAP7_75t_L g408 ( .A(n_409), .B(n_430), .C(n_451), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_410), .B(n_424), .Y(n_409) );
A2O1A1Ixp33_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_413), .B(n_415), .C(n_423), .Y(n_410) );
INVxp67_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g529 ( .A(n_414), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g443 ( .A(n_422), .Y(n_443) );
OAI21xp5_ASAP7_75t_L g516 ( .A1(n_428), .A2(n_517), .B(n_518), .Y(n_516) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
NAND3xp33_ASAP7_75t_L g430 ( .A(n_431), .B(n_439), .C(n_444), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_432), .B(n_436), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .Y(n_432) );
AND2x4_ASAP7_75t_L g462 ( .A(n_437), .B(n_463), .Y(n_462) );
AND2x4_ASAP7_75t_L g495 ( .A(n_438), .B(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_440), .B(n_441), .Y(n_439) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_443), .B(n_495), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_445), .B(n_448), .Y(n_444) );
INVx1_ASAP7_75t_L g480 ( .A(n_446), .Y(n_480) );
INVx1_ASAP7_75t_L g486 ( .A(n_449), .Y(n_486) );
AND2x4_ASAP7_75t_L g513 ( .A(n_449), .B(n_514), .Y(n_513) );
OAI21xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_455), .B(n_458), .Y(n_451) );
NOR2x1_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
AOI22xp5_ASAP7_75t_L g500 ( .A1(n_454), .A2(n_462), .B1(n_501), .B2(n_503), .Y(n_500) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AOI22xp5_ASAP7_75t_L g520 ( .A1(n_456), .A2(n_521), .B1(n_523), .B2(n_526), .Y(n_520) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
NAND2xp33_ASAP7_75t_L g465 ( .A(n_466), .B(n_498), .Y(n_465) );
NOR3xp33_ASAP7_75t_L g466 ( .A(n_467), .B(n_478), .C(n_487), .Y(n_466) );
OR3x1_ASAP7_75t_L g535 ( .A(n_467), .B(n_478), .C(n_487), .Y(n_535) );
AO21x1_ASAP7_75t_L g467 ( .A1(n_468), .A2(n_471), .B(n_473), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_472), .B(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g517 ( .A(n_472), .B(n_492), .Y(n_517) );
AOI21xp33_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_481), .B(n_486), .Y(n_478) );
OR2x2_ASAP7_75t_L g481 ( .A(n_482), .B(n_485), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
OAI21xp33_ASAP7_75t_L g488 ( .A1(n_489), .A2(n_493), .B(n_494), .Y(n_488) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_497), .Y(n_494) );
AND2x4_ASAP7_75t_L g505 ( .A(n_495), .B(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g539 ( .A(n_498), .Y(n_539) );
NOR3xp33_ASAP7_75t_SL g498 ( .A(n_499), .B(n_508), .C(n_519), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_500), .B(n_504), .Y(n_499) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g508 ( .A(n_509), .B(n_516), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_512), .B1(n_513), .B2(n_515), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_520), .B(n_527), .Y(n_519) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_532), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_534), .B(n_537), .Y(n_533) );
OAI21xp5_ASAP7_75t_L g537 ( .A1(n_536), .A2(n_538), .B(n_539), .Y(n_537) );
CKINVDCx5p33_ASAP7_75t_R g540 ( .A(n_541), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g541 ( .A(n_542), .B(n_546), .Y(n_541) );
CKINVDCx5p33_ASAP7_75t_R g559 ( .A(n_542), .Y(n_559) );
CKINVDCx5p33_ASAP7_75t_R g545 ( .A(n_543), .Y(n_545) );
BUFx3_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
BUFx3_ASAP7_75t_L g560 ( .A(n_547), .Y(n_560) );
INVx3_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
BUFx12f_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
BUFx8_ASAP7_75t_SL g564 ( .A(n_549), .Y(n_564) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
INVx8_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
OR2x6_ASAP7_75t_L g581 ( .A(n_553), .B(n_582), .Y(n_581) );
INVxp67_ASAP7_75t_L g968 ( .A(n_553), .Y(n_968) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_555), .B(n_556), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g566 ( .A(n_562), .B(n_567), .Y(n_566) );
CKINVDCx5p33_ASAP7_75t_R g563 ( .A(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_566), .B(n_568), .Y(n_565) );
OAI21xp5_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_584), .B(n_967), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_570), .B(n_577), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g969 ( .A(n_570), .B(n_578), .Y(n_969) );
INVxp67_ASAP7_75t_R g576 ( .A(n_571), .Y(n_576) );
AOI22xp5_ASAP7_75t_L g967 ( .A1(n_577), .A2(n_584), .B1(n_968), .B2(n_969), .Y(n_967) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
NOR2xp33_ASAP7_75t_SL g578 ( .A(n_579), .B(n_583), .Y(n_578) );
CKINVDCx5p33_ASAP7_75t_R g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
CKINVDCx5p33_ASAP7_75t_R g585 ( .A(n_586), .Y(n_585) );
BUFx8_ASAP7_75t_L g966 ( .A(n_586), .Y(n_966) );
INVx2_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
NAND3x1_ASAP7_75t_L g589 ( .A(n_590), .B(n_829), .C(n_905), .Y(n_589) );
NOR2x1_ASAP7_75t_L g590 ( .A(n_591), .B(n_758), .Y(n_590) );
NAND3xp33_ASAP7_75t_L g591 ( .A(n_592), .B(n_714), .C(n_738), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
OAI22xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_648), .B1(n_705), .B2(n_709), .Y(n_593) );
OR2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_614), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_595), .B(n_777), .Y(n_927) );
AND3x2_ASAP7_75t_L g933 ( .A(n_595), .B(n_711), .C(n_813), .Y(n_933) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g766 ( .A(n_596), .B(n_723), .Y(n_766) );
AND2x2_ASAP7_75t_L g803 ( .A(n_596), .B(n_636), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g881 ( .A(n_596), .B(n_846), .Y(n_881) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g753 ( .A(n_597), .Y(n_753) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
AOI21xp5_ASAP7_75t_L g606 ( .A1(n_607), .A2(n_608), .B(n_609), .Y(n_606) );
OR2x2_ASAP7_75t_L g652 ( .A(n_611), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
OR2x2_ASAP7_75t_L g682 ( .A(n_612), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_615), .B(n_636), .Y(n_614) );
INVx1_ASAP7_75t_L g964 ( .A(n_615), .Y(n_964) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVxp67_ASAP7_75t_L g711 ( .A(n_616), .Y(n_711) );
AND2x2_ASAP7_75t_L g721 ( .A(n_616), .B(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g765 ( .A(n_616), .Y(n_765) );
AO21x2_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_624), .B(n_632), .Y(n_616) );
AO21x2_ASAP7_75t_L g745 ( .A1(n_617), .A2(n_624), .B(n_632), .Y(n_745) );
OAI21x1_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_620), .B(n_623), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_619), .B(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVx2_ASAP7_75t_L g641 ( .A(n_622), .Y(n_641) );
OAI21x1_ASAP7_75t_SL g624 ( .A1(n_625), .A2(n_626), .B(n_630), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_627), .B(n_629), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_629), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g635 ( .A(n_629), .Y(n_635) );
AOI21x1_ASAP7_75t_L g657 ( .A1(n_631), .A2(n_658), .B(n_659), .Y(n_657) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g712 ( .A(n_636), .B(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g750 ( .A(n_636), .Y(n_750) );
INVx1_ASAP7_75t_L g790 ( .A(n_636), .Y(n_790) );
INVx2_ASAP7_75t_L g846 ( .A(n_636), .Y(n_846) );
NAND2x1p5_ASAP7_75t_L g636 ( .A(n_637), .B(n_642), .Y(n_636) );
AND2x2_ASAP7_75t_L g719 ( .A(n_637), .B(n_642), .Y(n_719) );
OR2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_640), .Y(n_637) );
OA21x2_ASAP7_75t_L g642 ( .A1(n_643), .A2(n_644), .B(n_646), .Y(n_642) );
INVx1_ASAP7_75t_L g728 ( .A(n_647), .Y(n_728) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AND2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_674), .Y(n_649) );
INVx2_ASAP7_75t_L g773 ( .A(n_650), .Y(n_773) );
AND2x4_ASAP7_75t_L g809 ( .A(n_650), .B(n_810), .Y(n_809) );
AND2x2_ASAP7_75t_L g895 ( .A(n_650), .B(n_794), .Y(n_895) );
AND2x2_ASAP7_75t_L g650 ( .A(n_651), .B(n_662), .Y(n_650) );
AND2x2_ASAP7_75t_L g707 ( .A(n_651), .B(n_663), .Y(n_707) );
INVx2_ASAP7_75t_SL g737 ( .A(n_651), .Y(n_737) );
OAI21x1_ASAP7_75t_L g651 ( .A1(n_652), .A2(n_654), .B(n_660), .Y(n_651) );
OAI21xp5_ASAP7_75t_L g852 ( .A1(n_652), .A2(n_654), .B(n_660), .Y(n_852) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_653), .B(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g782 ( .A(n_662), .Y(n_782) );
AND2x2_ASAP7_75t_L g904 ( .A(n_662), .B(n_675), .Y(n_904) );
INVx3_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx2_ASAP7_75t_L g733 ( .A(n_663), .Y(n_733) );
AND2x2_ASAP7_75t_L g825 ( .A(n_663), .B(n_737), .Y(n_825) );
AND2x4_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
OAI21x1_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_669), .B(n_673), .Y(n_665) );
AOI21xp5_ASAP7_75t_L g669 ( .A1(n_670), .A2(n_671), .B(n_672), .Y(n_669) );
INVx2_ASAP7_75t_L g708 ( .A(n_674), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_674), .B(n_816), .Y(n_815) );
HB1xp67_ASAP7_75t_L g860 ( .A(n_674), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g958 ( .A(n_674), .B(n_959), .Y(n_958) );
AND2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_687), .Y(n_674) );
INVx1_ASAP7_75t_L g734 ( .A(n_675), .Y(n_734) );
INVx1_ASAP7_75t_L g772 ( .A(n_675), .Y(n_772) );
INVx1_ASAP7_75t_L g780 ( .A(n_675), .Y(n_780) );
INVx2_ASAP7_75t_L g795 ( .A(n_675), .Y(n_795) );
NOR2x1_ASAP7_75t_L g810 ( .A(n_675), .B(n_811), .Y(n_810) );
AND2x2_ASAP7_75t_L g821 ( .A(n_675), .B(n_688), .Y(n_821) );
OR2x6_ASAP7_75t_L g675 ( .A(n_676), .B(n_684), .Y(n_675) );
OAI21x1_ASAP7_75t_L g676 ( .A1(n_677), .A2(n_679), .B(n_682), .Y(n_676) );
INVx1_ASAP7_75t_L g690 ( .A(n_678), .Y(n_690) );
NOR2xp67_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
AND2x2_ASAP7_75t_L g794 ( .A(n_687), .B(n_795), .Y(n_794) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
AND2x2_ASAP7_75t_L g736 ( .A(n_688), .B(n_737), .Y(n_736) );
INVxp67_ASAP7_75t_L g757 ( .A(n_688), .Y(n_757) );
INVx1_ASAP7_75t_L g806 ( .A(n_688), .Y(n_806) );
INVx1_ASAP7_75t_L g811 ( .A(n_688), .Y(n_811) );
OR2x2_ASAP7_75t_L g851 ( .A(n_688), .B(n_852), .Y(n_851) );
AO21x2_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_691), .B(n_703), .Y(n_688) );
NAND3xp33_ASAP7_75t_SL g691 ( .A(n_692), .B(n_695), .C(n_698), .Y(n_691) );
NAND2xp33_ASAP7_75t_SL g876 ( .A(n_705), .B(n_877), .Y(n_876) );
OR2x2_ASAP7_75t_L g705 ( .A(n_706), .B(n_708), .Y(n_705) );
INVx2_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_L g828 ( .A(n_707), .B(n_821), .Y(n_828) );
AND2x2_ASAP7_75t_L g843 ( .A(n_707), .B(n_771), .Y(n_843) );
AND2x2_ASAP7_75t_L g856 ( .A(n_707), .B(n_857), .Y(n_856) );
HB1xp67_ASAP7_75t_L g951 ( .A(n_708), .Y(n_951) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_709), .B(n_716), .Y(n_715) );
INVx2_ASAP7_75t_SL g709 ( .A(n_710), .Y(n_709) );
AND2x2_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_712), .B(n_768), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g900 ( .A(n_712), .B(n_901), .Y(n_900) );
AND2x2_ASAP7_75t_L g960 ( .A(n_712), .B(n_961), .Y(n_960) );
AND2x2_ASAP7_75t_L g718 ( .A(n_713), .B(n_719), .Y(n_718) );
AND2x2_ASAP7_75t_L g744 ( .A(n_713), .B(n_745), .Y(n_744) );
NAND2x1_ASAP7_75t_L g787 ( .A(n_713), .B(n_722), .Y(n_787) );
NAND2xp5_ASAP7_75t_SL g714 ( .A(n_715), .B(n_730), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_717), .B(n_720), .Y(n_716) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
AND2x4_ASAP7_75t_L g776 ( .A(n_718), .B(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g869 ( .A(n_718), .Y(n_869) );
AND2x2_ASAP7_75t_L g889 ( .A(n_718), .B(n_768), .Y(n_889) );
INVx2_ASAP7_75t_SL g747 ( .A(n_719), .Y(n_747) );
BUFx3_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_721), .B(n_863), .Y(n_862) );
AND2x2_ASAP7_75t_L g919 ( .A(n_721), .B(n_813), .Y(n_919) );
AOI32xp33_ASAP7_75t_L g929 ( .A1(n_721), .A2(n_850), .A3(n_930), .B1(n_931), .B2(n_933), .Y(n_929) );
INVx2_ASAP7_75t_L g755 ( .A(n_722), .Y(n_755) );
INVx1_ASAP7_75t_L g961 ( .A(n_722), .Y(n_961) );
INVx3_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
OAI321xp33_ASAP7_75t_L g948 ( .A1(n_731), .A2(n_949), .A3(n_951), .B1(n_952), .B2(n_954), .C(n_955), .Y(n_948) );
NAND2x2_ASAP7_75t_L g731 ( .A(n_732), .B(n_735), .Y(n_731) );
AND2x2_ASAP7_75t_L g912 ( .A(n_732), .B(n_850), .Y(n_912) );
AND2x2_ASAP7_75t_L g732 ( .A(n_733), .B(n_734), .Y(n_732) );
NOR2xp33_ASAP7_75t_L g756 ( .A(n_733), .B(n_757), .Y(n_756) );
INVx2_ASAP7_75t_L g793 ( .A(n_733), .Y(n_793) );
HB1xp67_ASAP7_75t_L g849 ( .A(n_733), .Y(n_849) );
OR2x2_ASAP7_75t_L g868 ( .A(n_733), .B(n_851), .Y(n_868) );
OR2x2_ASAP7_75t_L g891 ( .A(n_734), .B(n_773), .Y(n_891) );
AND2x2_ASAP7_75t_L g939 ( .A(n_734), .B(n_825), .Y(n_939) );
BUFx3_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_736), .B(n_780), .Y(n_799) );
AND2x4_ASAP7_75t_L g903 ( .A(n_736), .B(n_904), .Y(n_903) );
INVx1_ASAP7_75t_L g783 ( .A(n_737), .Y(n_783) );
INVx1_ASAP7_75t_L g816 ( .A(n_737), .Y(n_816) );
OAI21xp5_ASAP7_75t_L g738 ( .A1(n_739), .A2(n_748), .B(n_756), .Y(n_738) );
AND2x2_ASAP7_75t_L g739 ( .A(n_740), .B(n_743), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_741), .B(n_753), .Y(n_884) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
OR2x2_ASAP7_75t_L g769 ( .A(n_742), .B(n_745), .Y(n_769) );
AND2x4_ASAP7_75t_L g777 ( .A(n_742), .B(n_765), .Y(n_777) );
AND2x2_ASAP7_75t_L g791 ( .A(n_742), .B(n_745), .Y(n_791) );
INVx2_ASAP7_75t_L g826 ( .A(n_743), .Y(n_826) );
AND2x2_ASAP7_75t_L g743 ( .A(n_744), .B(n_746), .Y(n_743) );
INVx2_ASAP7_75t_L g874 ( .A(n_744), .Y(n_874) );
AND2x2_ASAP7_75t_L g892 ( .A(n_744), .B(n_754), .Y(n_892) );
AND2x4_ASAP7_75t_L g752 ( .A(n_745), .B(n_753), .Y(n_752) );
INVx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
OR2x2_ASAP7_75t_L g786 ( .A(n_747), .B(n_787), .Y(n_786) );
INVx2_ASAP7_75t_L g813 ( .A(n_747), .Y(n_813) );
AND2x2_ASAP7_75t_L g875 ( .A(n_747), .B(n_755), .Y(n_875) );
AND2x2_ASAP7_75t_L g748 ( .A(n_749), .B(n_751), .Y(n_748) );
AND2x2_ASAP7_75t_L g930 ( .A(n_749), .B(n_804), .Y(n_930) );
INVx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
AOI221xp5_ASAP7_75t_L g808 ( .A1(n_751), .A2(n_809), .B1(n_812), .B2(n_814), .C(n_817), .Y(n_808) );
AND2x2_ASAP7_75t_L g751 ( .A(n_752), .B(n_754), .Y(n_751) );
AND2x2_ASAP7_75t_L g845 ( .A(n_752), .B(n_846), .Y(n_845) );
BUFx3_ASAP7_75t_L g886 ( .A(n_752), .Y(n_886) );
INVxp67_ASAP7_75t_SL g909 ( .A(n_753), .Y(n_909) );
INVx1_ASAP7_75t_L g941 ( .A(n_754), .Y(n_941) );
INVx2_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g834 ( .A(n_755), .Y(n_834) );
AND2x2_ASAP7_75t_L g937 ( .A(n_756), .B(n_916), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_759), .B(n_808), .Y(n_758) );
NOR3xp33_ASAP7_75t_L g759 ( .A(n_760), .B(n_774), .C(n_796), .Y(n_759) );
NOR2xp33_ASAP7_75t_L g760 ( .A(n_761), .B(n_770), .Y(n_760) );
AND2x2_ASAP7_75t_L g761 ( .A(n_762), .B(n_767), .Y(n_761) );
OAI21xp33_ASAP7_75t_L g796 ( .A1(n_762), .A2(n_797), .B(n_800), .Y(n_796) );
NAND2x1p5_ASAP7_75t_L g762 ( .A(n_763), .B(n_766), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g954 ( .A(n_766), .Y(n_954) );
INVx2_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
INVx2_ASAP7_75t_L g819 ( .A(n_769), .Y(n_819) );
INVx1_ASAP7_75t_L g871 ( .A(n_770), .Y(n_871) );
OR2x2_ASAP7_75t_SL g770 ( .A(n_771), .B(n_773), .Y(n_770) );
INVx2_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
AND2x2_ASAP7_75t_L g956 ( .A(n_772), .B(n_947), .Y(n_956) );
OR2x2_ASAP7_75t_L g837 ( .A(n_773), .B(n_838), .Y(n_837) );
OAI21xp33_ASAP7_75t_L g774 ( .A1(n_775), .A2(n_778), .B(n_784), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
BUFx3_ASAP7_75t_L g807 ( .A(n_777), .Y(n_807) );
AND2x2_ASAP7_75t_L g812 ( .A(n_777), .B(n_813), .Y(n_812) );
NOR2xp67_ASAP7_75t_L g841 ( .A(n_777), .B(n_802), .Y(n_841) );
INVx3_ASAP7_75t_L g901 ( .A(n_777), .Y(n_901) );
OR2x2_ASAP7_75t_L g778 ( .A(n_779), .B(n_781), .Y(n_778) );
HB1xp67_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
AND2x2_ASAP7_75t_L g916 ( .A(n_780), .B(n_917), .Y(n_916) );
OR2x2_ASAP7_75t_L g781 ( .A(n_782), .B(n_783), .Y(n_781) );
INVx1_ASAP7_75t_L g804 ( .A(n_782), .Y(n_804) );
INVxp67_ASAP7_75t_SL g866 ( .A(n_783), .Y(n_866) );
OAI21xp33_ASAP7_75t_L g784 ( .A1(n_785), .A2(n_788), .B(n_792), .Y(n_784) );
INVx2_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
AND2x2_ASAP7_75t_L g788 ( .A(n_789), .B(n_791), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g857 ( .A(n_790), .Y(n_857) );
INVx1_ASAP7_75t_L g935 ( .A(n_790), .Y(n_935) );
NOR3xp33_ASAP7_75t_L g897 ( .A(n_791), .B(n_819), .C(n_875), .Y(n_897) );
INVx2_ASAP7_75t_L g936 ( .A(n_791), .Y(n_936) );
AOI22xp5_ASAP7_75t_L g938 ( .A1(n_791), .A2(n_939), .B1(n_940), .B2(n_943), .Y(n_938) );
AND2x2_ASAP7_75t_L g953 ( .A(n_791), .B(n_813), .Y(n_953) );
INVx2_ASAP7_75t_L g922 ( .A(n_792), .Y(n_922) );
AND2x2_ASAP7_75t_L g792 ( .A(n_793), .B(n_794), .Y(n_792) );
AND2x2_ASAP7_75t_L g915 ( .A(n_793), .B(n_806), .Y(n_915) );
INVx1_ASAP7_75t_L g959 ( .A(n_793), .Y(n_959) );
AND2x2_ASAP7_75t_L g899 ( .A(n_794), .B(n_825), .Y(n_899) );
INVx1_ASAP7_75t_L g932 ( .A(n_794), .Y(n_932) );
OAI21xp33_ASAP7_75t_L g962 ( .A1(n_797), .A2(n_963), .B(n_965), .Y(n_962) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
NAND4xp25_ASAP7_75t_L g800 ( .A(n_801), .B(n_804), .C(n_805), .D(n_807), .Y(n_800) );
INVx2_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVx2_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g835 ( .A(n_803), .Y(n_835) );
INVx1_ASAP7_75t_L g950 ( .A(n_804), .Y(n_950) );
INVx2_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx2_ASAP7_75t_L g877 ( .A(n_809), .Y(n_877) );
NAND2x1_ASAP7_75t_L g818 ( .A(n_813), .B(n_819), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g965 ( .A(n_814), .B(n_845), .Y(n_965) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
OAI32xp33_ASAP7_75t_L g817 ( .A1(n_818), .A2(n_820), .A3(n_822), .B1(n_826), .B2(n_827), .Y(n_817) );
INVx1_ASAP7_75t_L g831 ( .A(n_818), .Y(n_831) );
A2O1A1Ixp33_ASAP7_75t_L g934 ( .A1(n_819), .A2(n_935), .B(n_936), .C(n_937), .Y(n_934) );
HB1xp67_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx1_ASAP7_75t_L g838 ( .A(n_821), .Y(n_838) );
AND2x2_ASAP7_75t_L g865 ( .A(n_821), .B(n_866), .Y(n_865) );
NAND2x1_ASAP7_75t_SL g887 ( .A(n_821), .B(n_825), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g923 ( .A(n_821), .B(n_924), .Y(n_923) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx2_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx2_ASAP7_75t_L g827 ( .A(n_828), .Y(n_827) );
AND4x1_ASAP7_75t_L g829 ( .A(n_830), .B(n_853), .C(n_870), .D(n_888), .Y(n_829) );
O2A1O1Ixp5_ASAP7_75t_L g830 ( .A1(n_831), .A2(n_832), .B(n_836), .C(n_839), .Y(n_830) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
OR2x2_ASAP7_75t_L g833 ( .A(n_834), .B(n_835), .Y(n_833) );
NAND2xp5_ASAP7_75t_SL g855 ( .A(n_834), .B(n_856), .Y(n_855) );
INVx2_ASAP7_75t_SL g836 ( .A(n_837), .Y(n_836) );
OAI22xp5_ASAP7_75t_L g839 ( .A1(n_840), .A2(n_842), .B1(n_844), .B2(n_847), .Y(n_839) );
INVx1_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
INVx2_ASAP7_75t_L g844 ( .A(n_845), .Y(n_844) );
INVx1_ASAP7_75t_L g863 ( .A(n_846), .Y(n_863) );
INVx1_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
AND2x2_ASAP7_75t_L g848 ( .A(n_849), .B(n_850), .Y(n_848) );
INVx1_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx2_ASAP7_75t_L g947 ( .A(n_851), .Y(n_947) );
BUFx2_ASAP7_75t_L g917 ( .A(n_852), .Y(n_917) );
AOI21xp5_ASAP7_75t_L g853 ( .A1(n_854), .A2(n_858), .B(n_861), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
OR2x2_ASAP7_75t_L g883 ( .A(n_857), .B(n_884), .Y(n_883) );
INVx1_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVx1_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
OAI22xp5_ASAP7_75t_SL g861 ( .A1(n_862), .A2(n_864), .B1(n_867), .B2(n_869), .Y(n_861) );
INVx1_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
HB1xp67_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
AOI221xp5_ASAP7_75t_L g870 ( .A1(n_871), .A2(n_872), .B1(n_876), .B2(n_878), .C(n_882), .Y(n_870) );
AND2x4_ASAP7_75t_L g872 ( .A(n_873), .B(n_875), .Y(n_872) );
INVx1_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
INVx1_ASAP7_75t_L g942 ( .A(n_874), .Y(n_942) );
INVx1_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
INVx1_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
OR2x2_ASAP7_75t_L g963 ( .A(n_881), .B(n_964), .Y(n_963) );
AOI21xp33_ASAP7_75t_SL g882 ( .A1(n_883), .A2(n_885), .B(n_887), .Y(n_882) );
INVx2_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
AOI221xp5_ASAP7_75t_L g888 ( .A1(n_889), .A2(n_890), .B1(n_892), .B2(n_893), .C(n_896), .Y(n_888) );
INVx1_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
INVx1_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
INVx2_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
OAI22xp33_ASAP7_75t_L g896 ( .A1(n_897), .A2(n_898), .B1(n_900), .B2(n_902), .Y(n_896) );
INVx2_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
INVx1_ASAP7_75t_L g910 ( .A(n_901), .Y(n_910) );
INVx2_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
INVx2_ASAP7_75t_L g945 ( .A(n_904), .Y(n_945) );
NOR4xp25_ASAP7_75t_L g905 ( .A(n_906), .B(n_928), .C(n_948), .D(n_962), .Y(n_905) );
OAI322xp33_ASAP7_75t_L g906 ( .A1(n_907), .A2(n_910), .A3(n_911), .B1(n_913), .B2(n_918), .C1(n_920), .C2(n_926), .Y(n_906) );
INVx1_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
INVx1_ASAP7_75t_L g908 ( .A(n_909), .Y(n_908) );
INVx1_ASAP7_75t_L g911 ( .A(n_912), .Y(n_911) );
INVx1_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
AND2x2_ASAP7_75t_L g914 ( .A(n_915), .B(n_916), .Y(n_914) );
INVx1_ASAP7_75t_L g925 ( .A(n_917), .Y(n_925) );
INVx1_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
INVx1_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_922), .B(n_923), .Y(n_921) );
INVxp67_ASAP7_75t_L g924 ( .A(n_925), .Y(n_924) );
HB1xp67_ASAP7_75t_L g926 ( .A(n_927), .Y(n_926) );
NAND3xp33_ASAP7_75t_SL g928 ( .A(n_929), .B(n_934), .C(n_938), .Y(n_928) );
INVx1_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
AND2x2_ASAP7_75t_L g940 ( .A(n_941), .B(n_942), .Y(n_940) );
INVx1_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
OR2x2_ASAP7_75t_L g944 ( .A(n_945), .B(n_946), .Y(n_944) );
INVx1_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
INVx1_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
INVx1_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
OAI21xp5_ASAP7_75t_L g955 ( .A1(n_956), .A2(n_957), .B(n_960), .Y(n_955) );
INVx1_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
INVx4_ASAP7_75t_SL g970 ( .A(n_971), .Y(n_970) );
INVx2_ASAP7_75t_SL g971 ( .A(n_972), .Y(n_971) );
INVx1_ASAP7_75t_L g972 ( .A(n_973), .Y(n_972) );
BUFx2_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
BUFx3_ASAP7_75t_L g979 ( .A(n_974), .Y(n_979) );
OR2x2_ASAP7_75t_SL g974 ( .A(n_975), .B(n_976), .Y(n_974) );
endmodule