module fake_netlist_5_1825_n_1273 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1273);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1273;

wire n_924;
wire n_1263;
wire n_977;
wire n_611;
wire n_1126;
wire n_1166;
wire n_469;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_667;
wire n_790;
wire n_1055;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1198;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_688;
wire n_800;
wire n_671;
wire n_819;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_292;
wire n_625;
wire n_854;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_373;
wire n_307;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_191;
wire n_1104;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_709;
wire n_317;
wire n_1236;
wire n_569;
wire n_227;
wire n_920;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_308;
wire n_297;
wire n_1078;
wire n_775;
wire n_219;
wire n_600;
wire n_223;
wire n_264;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_436;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_958;
wire n_1034;
wire n_670;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_214;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_197;
wire n_1069;
wire n_1075;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_907;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1002;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_596;
wire n_558;
wire n_702;
wire n_822;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_409;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_759;
wire n_806;
wire n_324;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_649;
wire n_547;
wire n_1191;
wire n_284;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_254;
wire n_1233;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1121;
wire n_314;
wire n_368;
wire n_604;
wire n_433;
wire n_949;
wire n_1008;
wire n_946;
wire n_1001;
wire n_498;
wire n_689;
wire n_738;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1054;
wire n_1269;
wire n_1095;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_374;
wire n_185;
wire n_396;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_473;
wire n_1043;
wire n_355;
wire n_486;
wire n_614;
wire n_337;
wire n_1177;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1132;
wire n_388;
wire n_1127;
wire n_761;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_582;
wire n_309;
wire n_512;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_987;
wire n_261;
wire n_767;
wire n_993;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_513;
wire n_1094;
wire n_560;
wire n_340;
wire n_1205;
wire n_1044;
wire n_346;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1037;
wire n_1080;
wire n_426;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_960;
wire n_222;
wire n_1123;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_256;
wire n_950;
wire n_380;
wire n_419;
wire n_444;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_376;
wire n_967;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_280;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_690;
wire n_583;
wire n_302;
wire n_1203;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_385;
wire n_212;
wire n_507;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1214;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1077;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1096;
wire n_234;
wire n_833;
wire n_225;
wire n_988;
wire n_814;
wire n_192;
wire n_1201;
wire n_1114;
wire n_655;
wire n_669;
wire n_472;
wire n_1176;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_577;
wire n_338;
wire n_693;
wire n_836;
wire n_990;
wire n_975;
wire n_1256;
wire n_567;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1102;
wire n_711;
wire n_1187;
wire n_1164;
wire n_489;
wire n_1174;
wire n_617;
wire n_876;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1212;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1059;
wire n_1133;
wire n_557;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_393;
wire n_487;
wire n_665;
wire n_421;
wire n_910;
wire n_768;
wire n_205;
wire n_1136;
wire n_754;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_202;
wire n_427;
wire n_791;
wire n_732;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1155;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_194;
wire n_855;
wire n_1178;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_605;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_780;
wire n_998;
wire n_467;
wire n_1227;
wire n_840;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_997;
wire n_932;
wire n_612;
wire n_788;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_737;
wire n_986;
wire n_509;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_733;
wire n_941;
wire n_981;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1108;
wire n_782;
wire n_1100;
wire n_862;
wire n_760;
wire n_381;
wire n_220;
wire n_390;
wire n_481;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_570;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_522;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_221;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_432;
wire n_839;
wire n_1210;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_772;
wire n_499;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_236;
wire n_1012;
wire n_903;
wire n_740;
wire n_203;
wire n_384;
wire n_277;
wire n_1061;
wire n_333;
wire n_462;
wire n_1193;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_632;
wire n_699;
wire n_979;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_312;
wire n_1076;
wire n_1091;
wire n_494;
wire n_641;
wire n_730;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1220;
wire n_229;
wire n_437;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_863;
wire n_805;
wire n_712;
wire n_246;
wire n_1042;
wire n_269;
wire n_285;
wire n_412;
wire n_657;
wire n_644;
wire n_1160;
wire n_491;
wire n_1258;
wire n_1074;
wire n_251;
wire n_566;
wire n_565;
wire n_597;
wire n_1181;
wire n_1196;
wire n_651;
wire n_334;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_20),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_76),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_6),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_51),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_147),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_90),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_45),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_113),
.Y(n_186)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_14),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_69),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_170),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_54),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_151),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_29),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_96),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_173),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_26),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_94),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_81),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_59),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_141),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_106),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_10),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_41),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_130),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_85),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_82),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_128),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_40),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_92),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_137),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_9),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_46),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_57),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_8),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_102),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_153),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_103),
.Y(n_216)
);

BUFx5_ASAP7_75t_L g217 ( 
.A(n_3),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_35),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_149),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_166),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_116),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_58),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_150),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_55),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g225 ( 
.A(n_145),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_49),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_24),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_13),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_118),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_138),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_43),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_78),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_87),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_36),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_169),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_167),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_179),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_201),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_225),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_227),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_228),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_181),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_217),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_217),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_182),
.Y(n_245)
);

BUFx5_ASAP7_75t_L g246 ( 
.A(n_180),
.Y(n_246)
);

BUFx10_ASAP7_75t_L g247 ( 
.A(n_191),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_183),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_217),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_217),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_225),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_184),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_185),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_217),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_217),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_217),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_192),
.Y(n_257)
);

BUFx10_ASAP7_75t_L g258 ( 
.A(n_195),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g259 ( 
.A(n_181),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_187),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_187),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_187),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_195),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_189),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_195),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_190),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_242),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_258),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_245),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_248),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_259),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_258),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_252),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_263),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_265),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_262),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_262),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_260),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_255),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_261),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_258),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_253),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_257),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_243),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_244),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_249),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_264),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_264),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_250),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_266),
.Y(n_290)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_255),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_254),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_256),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_237),
.Y(n_294)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_237),
.Y(n_295)
);

BUFx2_ASAP7_75t_SL g296 ( 
.A(n_247),
.Y(n_296)
);

INVx2_ASAP7_75t_SL g297 ( 
.A(n_247),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_246),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_246),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_246),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_246),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_246),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_238),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_246),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_246),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_266),
.Y(n_306)
);

INVx2_ASAP7_75t_SL g307 ( 
.A(n_247),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_238),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_240),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_240),
.Y(n_310)
);

INVxp67_ASAP7_75t_SL g311 ( 
.A(n_239),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_251),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_241),
.Y(n_313)
);

BUFx10_ASAP7_75t_L g314 ( 
.A(n_241),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_263),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_245),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_263),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_263),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_279),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_271),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_283),
.Y(n_321)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_283),
.Y(n_322)
);

INVxp67_ASAP7_75t_SL g323 ( 
.A(n_302),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_271),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_279),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_284),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_296),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_285),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_291),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_272),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_272),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_267),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_312),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_286),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_289),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_294),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_291),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_292),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_294),
.Y(n_339)
);

INVxp67_ASAP7_75t_SL g340 ( 
.A(n_302),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_293),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_312),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_297),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_291),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_303),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_272),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_303),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_278),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_280),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_318),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_274),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_267),
.Y(n_352)
);

INVxp67_ASAP7_75t_SL g353 ( 
.A(n_272),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g354 ( 
.A(n_268),
.Y(n_354)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_308),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_269),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_275),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_308),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_315),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_309),
.Y(n_360)
);

INVx4_ASAP7_75t_R g361 ( 
.A(n_297),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_268),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_317),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g364 ( 
.A(n_295),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_276),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_307),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_309),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_277),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_307),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_319),
.B(n_298),
.Y(n_370)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_330),
.Y(n_371)
);

BUFx3_ASAP7_75t_L g372 ( 
.A(n_330),
.Y(n_372)
);

INVx3_ASAP7_75t_L g373 ( 
.A(n_329),
.Y(n_373)
);

AND2x4_ASAP7_75t_L g374 ( 
.A(n_348),
.B(n_233),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_319),
.B(n_325),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_325),
.Y(n_376)
);

NOR2x1_ASAP7_75t_L g377 ( 
.A(n_326),
.B(n_310),
.Y(n_377)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_364),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_326),
.B(n_313),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_323),
.B(n_299),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_344),
.Y(n_381)
);

AND2x4_ASAP7_75t_L g382 ( 
.A(n_348),
.B(n_233),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_340),
.B(n_300),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_337),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_343),
.B(n_288),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_328),
.B(n_314),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_337),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_338),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_328),
.B(n_301),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_334),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_365),
.B(n_314),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g392 ( 
.A(n_334),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_366),
.B(n_288),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_344),
.Y(n_394)
);

BUFx2_ASAP7_75t_L g395 ( 
.A(n_324),
.Y(n_395)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_335),
.Y(n_396)
);

INVx5_ASAP7_75t_L g397 ( 
.A(n_346),
.Y(n_397)
);

BUFx8_ASAP7_75t_SL g398 ( 
.A(n_336),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_365),
.B(n_314),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_368),
.Y(n_400)
);

INVx5_ASAP7_75t_L g401 ( 
.A(n_353),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_368),
.Y(n_402)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_335),
.Y(n_403)
);

AND2x4_ASAP7_75t_L g404 ( 
.A(n_349),
.B(n_186),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_369),
.B(n_306),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_341),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_341),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_349),
.B(n_311),
.Y(n_408)
);

INVx5_ASAP7_75t_L g409 ( 
.A(n_331),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_350),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_350),
.B(n_304),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_351),
.B(n_270),
.Y(n_412)
);

AND2x6_ASAP7_75t_L g413 ( 
.A(n_351),
.B(n_204),
.Y(n_413)
);

BUFx3_ASAP7_75t_L g414 ( 
.A(n_359),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_359),
.Y(n_415)
);

OAI22x1_ASAP7_75t_SL g416 ( 
.A1(n_398),
.A2(n_321),
.B1(n_345),
.B2(n_339),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_402),
.Y(n_417)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_379),
.B(n_327),
.Y(n_418)
);

BUFx2_ASAP7_75t_L g419 ( 
.A(n_395),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_402),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_381),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_381),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_402),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_371),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_379),
.B(n_322),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_394),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_379),
.B(n_354),
.Y(n_427)
);

INVx2_ASAP7_75t_SL g428 ( 
.A(n_390),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_390),
.Y(n_429)
);

BUFx8_ASAP7_75t_L g430 ( 
.A(n_395),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_394),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_403),
.B(n_357),
.Y(n_432)
);

AND2x2_ASAP7_75t_SL g433 ( 
.A(n_403),
.B(n_204),
.Y(n_433)
);

OAI22x1_ASAP7_75t_SL g434 ( 
.A1(n_400),
.A2(n_321),
.B1(n_358),
.B2(n_347),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_376),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_392),
.B(n_414),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_376),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_403),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_387),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_371),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_387),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_390),
.B(n_356),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_371),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_392),
.B(n_363),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_385),
.B(n_282),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_387),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_393),
.B(n_316),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_405),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_378),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_378),
.A2(n_367),
.B1(n_332),
.B2(n_352),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_408),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_400),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_373),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_412),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_392),
.B(n_270),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_375),
.Y(n_456)
);

NAND2xp33_ASAP7_75t_SL g457 ( 
.A(n_390),
.B(n_356),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_373),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_386),
.B(n_362),
.Y(n_459)
);

OA21x2_ASAP7_75t_L g460 ( 
.A1(n_370),
.A2(n_305),
.B(n_218),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_377),
.A2(n_306),
.B1(n_287),
.B2(n_290),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_373),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_414),
.B(n_273),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_373),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_372),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_375),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_415),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g468 ( 
.A(n_408),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_390),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_415),
.Y(n_470)
);

INVx4_ASAP7_75t_L g471 ( 
.A(n_390),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_396),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_414),
.B(n_194),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_377),
.A2(n_273),
.B1(n_212),
.B2(n_197),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_372),
.Y(n_475)
);

INVx5_ASAP7_75t_L g476 ( 
.A(n_413),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_396),
.Y(n_477)
);

INVx5_ASAP7_75t_L g478 ( 
.A(n_413),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_372),
.Y(n_479)
);

AND2x4_ASAP7_75t_L g480 ( 
.A(n_415),
.B(n_200),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_408),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_396),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_396),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_396),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_396),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_388),
.B(n_205),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_412),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_406),
.Y(n_488)
);

AOI22x1_ASAP7_75t_SL g489 ( 
.A1(n_386),
.A2(n_342),
.B1(n_333),
.B2(n_360),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_406),
.B(n_207),
.Y(n_490)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_386),
.Y(n_491)
);

BUFx3_ASAP7_75t_L g492 ( 
.A(n_406),
.Y(n_492)
);

NOR2x1_ASAP7_75t_L g493 ( 
.A(n_391),
.B(n_399),
.Y(n_493)
);

BUFx3_ASAP7_75t_L g494 ( 
.A(n_406),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_406),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_406),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_407),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_407),
.Y(n_498)
);

INVx3_ASAP7_75t_L g499 ( 
.A(n_407),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g500 ( 
.A(n_407),
.Y(n_500)
);

AND2x4_ASAP7_75t_L g501 ( 
.A(n_388),
.B(n_208),
.Y(n_501)
);

HB1xp67_ASAP7_75t_L g502 ( 
.A(n_391),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_407),
.B(n_214),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_407),
.Y(n_504)
);

AND2x4_ASAP7_75t_L g505 ( 
.A(n_388),
.B(n_222),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_410),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_410),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_410),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_410),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_410),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_436),
.B(n_410),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_436),
.B(n_404),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_421),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_422),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_426),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_417),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_419),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_431),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_435),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_437),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_495),
.Y(n_521)
);

AND2x4_ASAP7_75t_L g522 ( 
.A(n_436),
.B(n_404),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_416),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_417),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_420),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_495),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_456),
.B(n_399),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_420),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_423),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_423),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_438),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_438),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_495),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_471),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_439),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_430),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_430),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_430),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_495),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_R g540 ( 
.A(n_448),
.B(n_333),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_466),
.B(n_451),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_489),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_452),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_R g544 ( 
.A(n_448),
.B(n_342),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_439),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_419),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_468),
.B(n_481),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_418),
.B(n_404),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_441),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_434),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_441),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_450),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_446),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_445),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_445),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_454),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_446),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_432),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_453),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_453),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_487),
.B(n_388),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_449),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_425),
.B(n_427),
.Y(n_563)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_425),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_458),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_471),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_458),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_462),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_418),
.B(n_447),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_R g570 ( 
.A(n_457),
.B(n_355),
.Y(n_570)
);

AND2x4_ASAP7_75t_L g571 ( 
.A(n_493),
.B(n_404),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_471),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_500),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_474),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_462),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_464),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_464),
.Y(n_577)
);

NAND2xp33_ASAP7_75t_L g578 ( 
.A(n_554),
.B(n_424),
.Y(n_578)
);

BUFx2_ASAP7_75t_L g579 ( 
.A(n_517),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_516),
.Y(n_580)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_516),
.Y(n_581)
);

AOI21x1_ASAP7_75t_L g582 ( 
.A1(n_511),
.A2(n_503),
.B(n_490),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_535),
.Y(n_583)
);

BUFx2_ASAP7_75t_L g584 ( 
.A(n_546),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_528),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_528),
.Y(n_586)
);

NAND2xp33_ASAP7_75t_L g587 ( 
.A(n_555),
.B(n_424),
.Y(n_587)
);

OA22x2_ASAP7_75t_L g588 ( 
.A1(n_569),
.A2(n_491),
.B1(n_502),
.B2(n_461),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_535),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_562),
.B(n_447),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_545),
.Y(n_591)
);

BUFx6f_ASAP7_75t_SL g592 ( 
.A(n_512),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_545),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_562),
.B(n_455),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_534),
.Y(n_595)
);

OAI22xp33_ASAP7_75t_L g596 ( 
.A1(n_574),
.A2(n_463),
.B1(n_320),
.B2(n_444),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_568),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_568),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_524),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_563),
.B(n_427),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_525),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_529),
.Y(n_602)
);

AO21x2_ASAP7_75t_L g603 ( 
.A1(n_511),
.A2(n_442),
.B(n_486),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_530),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_549),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_531),
.Y(n_606)
);

NAND3xp33_ASAP7_75t_L g607 ( 
.A(n_527),
.B(n_459),
.C(n_457),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_556),
.B(n_540),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_551),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_558),
.B(n_459),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_553),
.Y(n_611)
);

BUFx2_ASAP7_75t_L g612 ( 
.A(n_556),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_574),
.B(n_442),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_541),
.B(n_473),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_564),
.B(n_473),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_557),
.Y(n_616)
);

INVx8_ASAP7_75t_L g617 ( 
.A(n_512),
.Y(n_617)
);

NAND2xp33_ASAP7_75t_L g618 ( 
.A(n_614),
.B(n_540),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_597),
.Y(n_619)
);

OAI22x1_ASAP7_75t_L g620 ( 
.A1(n_613),
.A2(n_552),
.B1(n_550),
.B2(n_523),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_596),
.B(n_548),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_600),
.B(n_547),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_597),
.Y(n_623)
);

BUFx10_ASAP7_75t_L g624 ( 
.A(n_592),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_609),
.Y(n_625)
);

BUFx3_ASAP7_75t_L g626 ( 
.A(n_579),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_609),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_599),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_607),
.B(n_571),
.Y(n_629)
);

NAND2xp33_ASAP7_75t_L g630 ( 
.A(n_610),
.B(n_544),
.Y(n_630)
);

XNOR2x2_ASAP7_75t_SL g631 ( 
.A(n_607),
.B(n_210),
.Y(n_631)
);

BUFx2_ASAP7_75t_L g632 ( 
.A(n_612),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_600),
.B(n_561),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_597),
.Y(n_634)
);

AND2x6_ASAP7_75t_L g635 ( 
.A(n_595),
.B(n_571),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_612),
.Y(n_636)
);

CKINVDCx6p67_ASAP7_75t_R g637 ( 
.A(n_608),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_590),
.A2(n_570),
.B1(n_571),
.B2(n_473),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_598),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_610),
.A2(n_588),
.B1(n_594),
.B2(n_615),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_598),
.Y(n_641)
);

BUFx4f_ASAP7_75t_L g642 ( 
.A(n_617),
.Y(n_642)
);

INVx5_ASAP7_75t_L g643 ( 
.A(n_595),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_579),
.B(n_570),
.Y(n_644)
);

BUFx3_ASAP7_75t_L g645 ( 
.A(n_584),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_599),
.Y(n_646)
);

BUFx4f_ASAP7_75t_L g647 ( 
.A(n_617),
.Y(n_647)
);

AOI22xp33_ASAP7_75t_L g648 ( 
.A1(n_588),
.A2(n_480),
.B1(n_561),
.B2(n_514),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_588),
.B(n_388),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_SL g650 ( 
.A(n_592),
.B(n_536),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_584),
.B(n_513),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_581),
.Y(n_652)
);

BUFx2_ASAP7_75t_L g653 ( 
.A(n_617),
.Y(n_653)
);

BUFx6f_ASAP7_75t_SL g654 ( 
.A(n_580),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_601),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_601),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_617),
.B(n_515),
.Y(n_657)
);

AND2x2_ASAP7_75t_L g658 ( 
.A(n_602),
.B(n_512),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_581),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_SL g660 ( 
.A1(n_578),
.A2(n_544),
.B1(n_538),
.B2(n_537),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_602),
.B(n_388),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_617),
.B(n_518),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_604),
.B(n_500),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_604),
.B(n_519),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_595),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_606),
.B(n_520),
.Y(n_666)
);

OAI22xp33_ASAP7_75t_SL g667 ( 
.A1(n_606),
.A2(n_543),
.B1(n_213),
.B2(n_480),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_605),
.B(n_500),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_605),
.B(n_522),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_585),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_585),
.Y(n_671)
);

INVxp67_ASAP7_75t_SL g672 ( 
.A(n_605),
.Y(n_672)
);

OAI22xp33_ASAP7_75t_L g673 ( 
.A1(n_616),
.A2(n_467),
.B1(n_470),
.B2(n_542),
.Y(n_673)
);

INVx4_ASAP7_75t_L g674 ( 
.A(n_592),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_583),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_611),
.Y(n_676)
);

AOI22x1_ASAP7_75t_L g677 ( 
.A1(n_616),
.A2(n_480),
.B1(n_501),
.B2(n_486),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_592),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_583),
.Y(n_679)
);

AOI22xp33_ASAP7_75t_L g680 ( 
.A1(n_611),
.A2(n_213),
.B1(n_382),
.B2(n_374),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_611),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_616),
.B(n_500),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_583),
.Y(n_683)
);

OR2x6_ASAP7_75t_L g684 ( 
.A(n_595),
.B(n_534),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_580),
.B(n_522),
.Y(n_685)
);

INVx2_ASAP7_75t_SL g686 ( 
.A(n_586),
.Y(n_686)
);

AOI22xp33_ASAP7_75t_SL g687 ( 
.A1(n_587),
.A2(n_199),
.B1(n_234),
.B2(n_188),
.Y(n_687)
);

INVx6_ASAP7_75t_L g688 ( 
.A(n_586),
.Y(n_688)
);

AND3x1_ASAP7_75t_L g689 ( 
.A(n_589),
.B(n_281),
.C(n_361),
.Y(n_689)
);

INVx3_ASAP7_75t_L g690 ( 
.A(n_591),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_589),
.Y(n_691)
);

NAND3xp33_ASAP7_75t_L g692 ( 
.A(n_593),
.B(n_522),
.C(n_382),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_591),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_593),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_591),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_603),
.Y(n_696)
);

HB1xp67_ASAP7_75t_L g697 ( 
.A(n_603),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_603),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g699 ( 
.A(n_582),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_582),
.B(n_424),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_609),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_613),
.B(n_424),
.Y(n_702)
);

BUFx3_ASAP7_75t_L g703 ( 
.A(n_579),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_688),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_625),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_627),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_701),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_672),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_622),
.B(n_198),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_688),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_618),
.B(n_215),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_702),
.B(n_224),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_672),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_676),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_681),
.Y(n_715)
);

CKINVDCx20_ASAP7_75t_R g716 ( 
.A(n_637),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_640),
.B(n_532),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_691),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_694),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_SL g720 ( 
.A(n_674),
.B(n_440),
.Y(n_720)
);

XOR2xp5_ASAP7_75t_L g721 ( 
.A(n_620),
.B(n_486),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_628),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_646),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_655),
.Y(n_724)
);

NAND2x1p5_ASAP7_75t_L g725 ( 
.A(n_631),
.B(n_534),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_702),
.B(n_501),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_658),
.B(n_501),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_656),
.Y(n_728)
);

OR2x6_ASAP7_75t_L g729 ( 
.A(n_629),
.B(n_440),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_695),
.Y(n_730)
);

OAI21xp5_ASAP7_75t_L g731 ( 
.A1(n_621),
.A2(n_433),
.B(n_505),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_633),
.B(n_505),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_687),
.B(n_374),
.Y(n_733)
);

AOI21xp5_ASAP7_75t_L g734 ( 
.A1(n_677),
.A2(n_433),
.B(n_566),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_SL g735 ( 
.A(n_674),
.B(n_440),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_640),
.B(n_559),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_619),
.Y(n_737)
);

INVx4_ASAP7_75t_L g738 ( 
.A(n_642),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_621),
.B(n_440),
.Y(n_739)
);

XNOR2xp5_ASAP7_75t_L g740 ( 
.A(n_687),
.B(n_374),
.Y(n_740)
);

AND2x4_ASAP7_75t_L g741 ( 
.A(n_678),
.B(n_573),
.Y(n_741)
);

INVx4_ASAP7_75t_L g742 ( 
.A(n_642),
.Y(n_742)
);

BUFx6f_ASAP7_75t_L g743 ( 
.A(n_626),
.Y(n_743)
);

AND2x2_ASAP7_75t_L g744 ( 
.A(n_636),
.B(n_505),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_623),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_634),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_675),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_679),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_632),
.B(n_374),
.Y(n_749)
);

INVxp67_ASAP7_75t_L g750 ( 
.A(n_645),
.Y(n_750)
);

CKINVDCx11_ASAP7_75t_R g751 ( 
.A(n_703),
.Y(n_751)
);

AOI21xp5_ASAP7_75t_L g752 ( 
.A1(n_631),
.A2(n_629),
.B(n_661),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_683),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_693),
.Y(n_754)
);

BUFx3_ASAP7_75t_L g755 ( 
.A(n_651),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_688),
.Y(n_756)
);

XOR2xp5_ASAP7_75t_L g757 ( 
.A(n_660),
.B(n_382),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_664),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_666),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_686),
.Y(n_760)
);

XNOR2xp5_ASAP7_75t_L g761 ( 
.A(n_660),
.B(n_382),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_639),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_641),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_624),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_644),
.B(n_196),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_652),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_659),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_670),
.Y(n_768)
);

OAI21xp5_ASAP7_75t_L g769 ( 
.A1(n_692),
.A2(n_648),
.B(n_700),
.Y(n_769)
);

INVxp67_ASAP7_75t_SL g770 ( 
.A(n_690),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_624),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_671),
.Y(n_772)
);

NAND2x1p5_ASAP7_75t_L g773 ( 
.A(n_643),
.B(n_566),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_630),
.B(n_202),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_690),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_650),
.B(n_203),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_L g777 ( 
.A(n_657),
.B(n_206),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_657),
.B(n_211),
.Y(n_778)
);

INVx2_ASAP7_75t_SL g779 ( 
.A(n_647),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_696),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_669),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_662),
.B(n_216),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_698),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_697),
.Y(n_784)
);

AND2x6_ASAP7_75t_L g785 ( 
.A(n_678),
.B(n_566),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_662),
.B(n_219),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_697),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_668),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_665),
.Y(n_789)
);

AO21x1_ASAP7_75t_L g790 ( 
.A1(n_673),
.A2(n_218),
.B(n_209),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_647),
.Y(n_791)
);

AO21x2_ASAP7_75t_L g792 ( 
.A1(n_769),
.A2(n_649),
.B(n_700),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_711),
.B(n_673),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_755),
.B(n_648),
.Y(n_794)
);

OR2x2_ASAP7_75t_L g795 ( 
.A(n_708),
.B(n_713),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_760),
.Y(n_796)
);

BUFx10_ASAP7_75t_L g797 ( 
.A(n_776),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_781),
.B(n_649),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_758),
.B(n_759),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_705),
.Y(n_800)
);

INVxp67_ASAP7_75t_L g801 ( 
.A(n_743),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_733),
.A2(n_638),
.B1(n_654),
.B2(n_667),
.Y(n_802)
);

NAND3xp33_ASAP7_75t_L g803 ( 
.A(n_712),
.B(n_689),
.C(n_638),
.Y(n_803)
);

AOI22xp5_ASAP7_75t_L g804 ( 
.A1(n_721),
.A2(n_654),
.B1(n_635),
.B2(n_653),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_706),
.Y(n_805)
);

INVxp67_ASAP7_75t_L g806 ( 
.A(n_743),
.Y(n_806)
);

INVx2_ASAP7_75t_SL g807 ( 
.A(n_743),
.Y(n_807)
);

AO221x1_ASAP7_75t_L g808 ( 
.A1(n_784),
.A2(n_699),
.B1(n_665),
.B2(n_195),
.C(n_526),
.Y(n_808)
);

INVxp67_ASAP7_75t_SL g809 ( 
.A(n_770),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_707),
.Y(n_810)
);

INVxp67_ASAP7_75t_L g811 ( 
.A(n_704),
.Y(n_811)
);

NAND3xp33_ASAP7_75t_L g812 ( 
.A(n_709),
.B(n_685),
.C(n_230),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_757),
.A2(n_635),
.B1(n_680),
.B2(n_229),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_722),
.B(n_665),
.Y(n_814)
);

OAI22xp5_ASAP7_75t_L g815 ( 
.A1(n_740),
.A2(n_680),
.B1(n_684),
.B2(n_643),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_750),
.B(n_221),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_723),
.B(n_665),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_718),
.Y(n_818)
);

NOR3xp33_ASAP7_75t_L g819 ( 
.A(n_774),
.B(n_663),
.C(n_668),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_777),
.B(n_643),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_761),
.A2(n_635),
.B1(n_226),
.B2(n_231),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_SL g822 ( 
.A(n_738),
.B(n_635),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_719),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_778),
.B(n_782),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_786),
.B(n_643),
.Y(n_825)
);

BUFx2_ASAP7_75t_L g826 ( 
.A(n_764),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_724),
.B(n_699),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_728),
.B(n_699),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_732),
.B(n_699),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_751),
.B(n_223),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_762),
.Y(n_831)
);

OAI22xp33_ASAP7_75t_L g832 ( 
.A1(n_752),
.A2(n_684),
.B1(n_465),
.B2(n_475),
.Y(n_832)
);

AOI22xp5_ASAP7_75t_L g833 ( 
.A1(n_765),
.A2(n_635),
.B1(n_235),
.B2(n_236),
.Y(n_833)
);

CKINVDCx20_ASAP7_75t_R g834 ( 
.A(n_716),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_763),
.B(n_682),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_749),
.B(n_232),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_766),
.B(n_682),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_710),
.B(n_209),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_771),
.B(n_738),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_734),
.A2(n_661),
.B(n_684),
.Y(n_840)
);

INVx2_ASAP7_75t_SL g841 ( 
.A(n_756),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_771),
.B(n_663),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_742),
.B(n_443),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_742),
.B(n_443),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_752),
.B(n_720),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_720),
.B(n_443),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_726),
.B(n_0),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_789),
.B(n_573),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_731),
.A2(n_572),
.B(n_478),
.Y(n_849)
);

INVx8_ASAP7_75t_L g850 ( 
.A(n_785),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_780),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_767),
.B(n_560),
.Y(n_852)
);

O2A1O1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_790),
.A2(n_411),
.B(n_389),
.C(n_575),
.Y(n_853)
);

BUFx2_ASAP7_75t_L g854 ( 
.A(n_785),
.Y(n_854)
);

OAI22xp5_ASAP7_75t_L g855 ( 
.A1(n_725),
.A2(n_572),
.B1(n_482),
.B2(n_507),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_768),
.B(n_565),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_772),
.B(n_567),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_791),
.B(n_0),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_783),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_714),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_739),
.B(n_576),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_715),
.B(n_577),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_741),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_737),
.B(n_1),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_745),
.B(n_1),
.Y(n_865)
);

NOR2xp33_ASAP7_75t_L g866 ( 
.A(n_779),
.B(n_2),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_796),
.B(n_799),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_824),
.B(n_744),
.Y(n_868)
);

NAND3xp33_ASAP7_75t_L g869 ( 
.A(n_793),
.B(n_769),
.C(n_731),
.Y(n_869)
);

AOI21xp5_ASAP7_75t_L g870 ( 
.A1(n_849),
.A2(n_735),
.B(n_729),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_831),
.B(n_788),
.Y(n_871)
);

OAI21xp5_ASAP7_75t_L g872 ( 
.A1(n_812),
.A2(n_803),
.B(n_845),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_797),
.B(n_741),
.Y(n_873)
);

AOI22xp5_ASAP7_75t_L g874 ( 
.A1(n_815),
.A2(n_727),
.B1(n_735),
.B2(n_729),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_797),
.B(n_826),
.Y(n_875)
);

AOI22xp5_ASAP7_75t_L g876 ( 
.A1(n_815),
.A2(n_729),
.B1(n_736),
.B2(n_717),
.Y(n_876)
);

NOR2x1p5_ASAP7_75t_L g877 ( 
.A(n_794),
.B(n_736),
.Y(n_877)
);

O2A1O1Ixp5_ASAP7_75t_L g878 ( 
.A1(n_820),
.A2(n_717),
.B(n_787),
.C(n_730),
.Y(n_878)
);

NAND2xp33_ASAP7_75t_L g879 ( 
.A(n_819),
.B(n_785),
.Y(n_879)
);

NAND2x1_ASAP7_75t_L g880 ( 
.A(n_808),
.B(n_785),
.Y(n_880)
);

OAI22xp5_ASAP7_75t_L g881 ( 
.A1(n_813),
.A2(n_725),
.B1(n_773),
.B2(n_775),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_830),
.B(n_746),
.Y(n_882)
);

OAI22xp5_ASAP7_75t_L g883 ( 
.A1(n_821),
.A2(n_773),
.B1(n_754),
.B2(n_753),
.Y(n_883)
);

AOI22xp5_ASAP7_75t_L g884 ( 
.A1(n_802),
.A2(n_748),
.B1(n_747),
.B2(n_389),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_834),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_804),
.B(n_443),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_801),
.B(n_2),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_L g888 ( 
.A(n_806),
.B(n_3),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_811),
.B(n_193),
.Y(n_889)
);

AOI22xp33_ASAP7_75t_L g890 ( 
.A1(n_825),
.A2(n_193),
.B1(n_220),
.B2(n_475),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_800),
.Y(n_891)
);

INVx8_ASAP7_75t_L g892 ( 
.A(n_850),
.Y(n_892)
);

AND2x4_ASAP7_75t_SL g893 ( 
.A(n_863),
.B(n_465),
.Y(n_893)
);

INVxp67_ASAP7_75t_L g894 ( 
.A(n_841),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_809),
.B(n_4),
.Y(n_895)
);

AOI22xp33_ASAP7_75t_L g896 ( 
.A1(n_847),
.A2(n_193),
.B1(n_220),
.B2(n_475),
.Y(n_896)
);

OAI21xp5_ASAP7_75t_L g897 ( 
.A1(n_833),
.A2(n_411),
.B(n_483),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_805),
.Y(n_898)
);

INVx2_ASAP7_75t_SL g899 ( 
.A(n_807),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_810),
.B(n_4),
.Y(n_900)
);

AOI22xp5_ASAP7_75t_SL g901 ( 
.A1(n_854),
.A2(n_858),
.B1(n_866),
.B2(n_863),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_822),
.A2(n_572),
.B(n_428),
.Y(n_902)
);

AOI22xp5_ASAP7_75t_L g903 ( 
.A1(n_822),
.A2(n_465),
.B1(n_479),
.B2(n_475),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_863),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_818),
.B(n_5),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_851),
.B(n_573),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_823),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_816),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_836),
.B(n_838),
.Y(n_909)
);

OAI22xp5_ASAP7_75t_L g910 ( 
.A1(n_832),
.A2(n_479),
.B1(n_465),
.B2(n_484),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_839),
.B(n_479),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_860),
.B(n_5),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_829),
.B(n_6),
.Y(n_913)
);

AOI22xp33_ASAP7_75t_L g914 ( 
.A1(n_792),
.A2(n_193),
.B1(n_220),
.B2(n_479),
.Y(n_914)
);

AOI22xp33_ASAP7_75t_SL g915 ( 
.A1(n_850),
.A2(n_220),
.B1(n_533),
.B2(n_526),
.Y(n_915)
);

OAI22xp5_ASAP7_75t_L g916 ( 
.A1(n_798),
.A2(n_508),
.B1(n_498),
.B2(n_496),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_859),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_814),
.B(n_7),
.Y(n_918)
);

AOI22xp5_ASAP7_75t_L g919 ( 
.A1(n_855),
.A2(n_413),
.B1(n_488),
.B2(n_472),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_795),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_817),
.B(n_7),
.Y(n_921)
);

CKINVDCx20_ASAP7_75t_R g922 ( 
.A(n_850),
.Y(n_922)
);

AOI22xp5_ASAP7_75t_L g923 ( 
.A1(n_792),
.A2(n_413),
.B1(n_497),
.B2(n_472),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_842),
.B(n_521),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_835),
.B(n_8),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_864),
.B(n_9),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_843),
.A2(n_413),
.B1(n_497),
.B2(n_477),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_837),
.B(n_10),
.Y(n_928)
);

OAI22xp5_ASAP7_75t_L g929 ( 
.A1(n_865),
.A2(n_533),
.B1(n_526),
.B2(n_521),
.Y(n_929)
);

AOI22xp5_ASAP7_75t_L g930 ( 
.A1(n_844),
.A2(n_413),
.B1(n_510),
.B2(n_477),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_827),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_846),
.A2(n_428),
.B(n_476),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_840),
.B(n_521),
.Y(n_933)
);

HB1xp67_ASAP7_75t_L g934 ( 
.A(n_828),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_862),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_848),
.Y(n_936)
);

OAI22xp5_ASAP7_75t_L g937 ( 
.A1(n_861),
.A2(n_533),
.B1(n_526),
.B2(n_521),
.Y(n_937)
);

AOI22xp33_ASAP7_75t_L g938 ( 
.A1(n_852),
.A2(n_413),
.B1(n_409),
.B2(n_492),
.Y(n_938)
);

AND2x4_ASAP7_75t_L g939 ( 
.A(n_856),
.B(n_533),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_857),
.B(n_11),
.Y(n_940)
);

AND2x2_ASAP7_75t_L g941 ( 
.A(n_853),
.B(n_11),
.Y(n_941)
);

AOI22xp5_ASAP7_75t_L g942 ( 
.A1(n_824),
.A2(n_510),
.B1(n_469),
.B2(n_429),
.Y(n_942)
);

AOI22xp33_ASAP7_75t_L g943 ( 
.A1(n_824),
.A2(n_409),
.B1(n_504),
.B2(n_494),
.Y(n_943)
);

AOI22xp33_ASAP7_75t_L g944 ( 
.A1(n_824),
.A2(n_409),
.B1(n_504),
.B2(n_494),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_824),
.B(n_12),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_891),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_892),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_934),
.B(n_12),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_872),
.B(n_13),
.Y(n_949)
);

AOI22xp5_ASAP7_75t_L g950 ( 
.A1(n_869),
.A2(n_539),
.B1(n_460),
.B2(n_429),
.Y(n_950)
);

AND2x6_ASAP7_75t_L g951 ( 
.A(n_941),
.B(n_539),
.Y(n_951)
);

NAND2x1p5_ASAP7_75t_L g952 ( 
.A(n_933),
.B(n_539),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_877),
.B(n_14),
.Y(n_953)
);

NOR3xp33_ASAP7_75t_SL g954 ( 
.A(n_945),
.B(n_15),
.C(n_16),
.Y(n_954)
);

INVx3_ASAP7_75t_L g955 ( 
.A(n_936),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_878),
.B(n_539),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_L g957 ( 
.A1(n_879),
.A2(n_460),
.B1(n_429),
.B2(n_499),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_885),
.Y(n_958)
);

INVxp67_ASAP7_75t_L g959 ( 
.A(n_898),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_907),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_870),
.B(n_506),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_917),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_935),
.B(n_15),
.Y(n_963)
);

NOR2x1p5_ASAP7_75t_L g964 ( 
.A(n_913),
.B(n_469),
.Y(n_964)
);

INVx3_ASAP7_75t_L g965 ( 
.A(n_936),
.Y(n_965)
);

AOI22xp33_ASAP7_75t_L g966 ( 
.A1(n_926),
.A2(n_485),
.B1(n_499),
.B2(n_469),
.Y(n_966)
);

OR2x6_ASAP7_75t_L g967 ( 
.A(n_892),
.B(n_506),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_931),
.B(n_16),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_920),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_936),
.B(n_17),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_871),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_867),
.Y(n_972)
);

AND2x6_ASAP7_75t_L g973 ( 
.A(n_874),
.B(n_506),
.Y(n_973)
);

INVxp67_ASAP7_75t_L g974 ( 
.A(n_889),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_900),
.Y(n_975)
);

HB1xp67_ASAP7_75t_L g976 ( 
.A(n_894),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_876),
.B(n_17),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_899),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_906),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_892),
.Y(n_980)
);

HB1xp67_ASAP7_75t_L g981 ( 
.A(n_905),
.Y(n_981)
);

INVx4_ASAP7_75t_L g982 ( 
.A(n_904),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_875),
.B(n_901),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_906),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_882),
.B(n_18),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_868),
.B(n_18),
.Y(n_986)
);

INVx2_ASAP7_75t_L g987 ( 
.A(n_939),
.Y(n_987)
);

AOI22xp33_ASAP7_75t_L g988 ( 
.A1(n_909),
.A2(n_485),
.B1(n_499),
.B2(n_492),
.Y(n_988)
);

AOI22xp33_ASAP7_75t_L g989 ( 
.A1(n_896),
.A2(n_485),
.B1(n_460),
.B2(n_384),
.Y(n_989)
);

BUFx3_ASAP7_75t_L g990 ( 
.A(n_922),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_912),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_939),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_895),
.B(n_19),
.Y(n_993)
);

OAI22xp5_ASAP7_75t_L g994 ( 
.A1(n_915),
.A2(n_509),
.B1(n_506),
.B2(n_409),
.Y(n_994)
);

INVxp33_ASAP7_75t_L g995 ( 
.A(n_873),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_925),
.B(n_19),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_928),
.B(n_20),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_918),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_924),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_880),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_921),
.B(n_940),
.Y(n_1001)
);

INVx3_ASAP7_75t_L g1002 ( 
.A(n_893),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_937),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_881),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_959),
.Y(n_1005)
);

AND2x4_ASAP7_75t_L g1006 ( 
.A(n_974),
.B(n_911),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_959),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_946),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_987),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_947),
.Y(n_1010)
);

HB1xp67_ASAP7_75t_L g1011 ( 
.A(n_976),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_962),
.Y(n_1012)
);

BUFx2_ASAP7_75t_L g1013 ( 
.A(n_976),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_981),
.B(n_929),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_981),
.B(n_923),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_972),
.B(n_998),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_955),
.B(n_886),
.Y(n_1017)
);

INVx3_ASAP7_75t_L g1018 ( 
.A(n_982),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_971),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_992),
.Y(n_1020)
);

INVx2_ASAP7_75t_SL g1021 ( 
.A(n_982),
.Y(n_1021)
);

AOI21xp33_ASAP7_75t_L g1022 ( 
.A1(n_949),
.A2(n_888),
.B(n_887),
.Y(n_1022)
);

INVxp67_ASAP7_75t_L g1023 ( 
.A(n_953),
.Y(n_1023)
);

INVx2_ASAP7_75t_SL g1024 ( 
.A(n_990),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_975),
.B(n_884),
.Y(n_1025)
);

INVx4_ASAP7_75t_L g1026 ( 
.A(n_947),
.Y(n_1026)
);

OR2x6_ASAP7_75t_L g1027 ( 
.A(n_961),
.B(n_902),
.Y(n_1027)
);

A2O1A1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_949),
.A2(n_908),
.B(n_883),
.C(n_914),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_979),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_969),
.Y(n_1030)
);

AND2x4_ASAP7_75t_L g1031 ( 
.A(n_974),
.B(n_903),
.Y(n_1031)
);

AOI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_954),
.A2(n_890),
.B1(n_942),
.B2(n_910),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_960),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_991),
.B(n_916),
.Y(n_1034)
);

BUFx3_ASAP7_75t_L g1035 ( 
.A(n_958),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_SL g1036 ( 
.A(n_947),
.B(n_919),
.Y(n_1036)
);

INVx3_ASAP7_75t_L g1037 ( 
.A(n_947),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_1004),
.B(n_932),
.Y(n_1038)
);

BUFx4f_ASAP7_75t_L g1039 ( 
.A(n_980),
.Y(n_1039)
);

BUFx2_ASAP7_75t_L g1040 ( 
.A(n_951),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_999),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_1001),
.B(n_943),
.Y(n_1042)
);

AOI22xp33_ASAP7_75t_L g1043 ( 
.A1(n_973),
.A2(n_897),
.B1(n_944),
.B2(n_938),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_984),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_955),
.Y(n_1045)
);

INVx3_ASAP7_75t_L g1046 ( 
.A(n_980),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_1003),
.B(n_927),
.Y(n_1047)
);

CKINVDCx5p33_ASAP7_75t_R g1048 ( 
.A(n_980),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_980),
.Y(n_1049)
);

AND2x4_ASAP7_75t_L g1050 ( 
.A(n_978),
.B(n_930),
.Y(n_1050)
);

NOR3xp33_ASAP7_75t_SL g1051 ( 
.A(n_983),
.B(n_961),
.C(n_977),
.Y(n_1051)
);

BUFx3_ASAP7_75t_L g1052 ( 
.A(n_970),
.Y(n_1052)
);

OR2x6_ASAP7_75t_L g1053 ( 
.A(n_956),
.B(n_509),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_1000),
.Y(n_1054)
);

INVx3_ASAP7_75t_L g1055 ( 
.A(n_965),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_1001),
.B(n_951),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_948),
.Y(n_1057)
);

NAND3xp33_ASAP7_75t_SL g1058 ( 
.A(n_983),
.B(n_21),
.C(n_22),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_968),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_965),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_951),
.B(n_995),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_956),
.B(n_21),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_967),
.B(n_22),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_SL g1064 ( 
.A(n_1000),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_963),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_952),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_952),
.Y(n_1067)
);

NOR2xp67_ASAP7_75t_L g1068 ( 
.A(n_1000),
.B(n_23),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_951),
.B(n_23),
.Y(n_1069)
);

INVx4_ASAP7_75t_L g1070 ( 
.A(n_1000),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_1058),
.A2(n_985),
.B(n_993),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_1055),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_1023),
.B(n_996),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_1028),
.A2(n_1022),
.B(n_1056),
.Y(n_1074)
);

INVxp67_ASAP7_75t_SL g1075 ( 
.A(n_1011),
.Y(n_1075)
);

NOR3xp33_ASAP7_75t_L g1076 ( 
.A(n_1022),
.B(n_997),
.C(n_986),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_1018),
.B(n_951),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_1010),
.Y(n_1078)
);

BUFx3_ASAP7_75t_L g1079 ( 
.A(n_1035),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_1027),
.A2(n_966),
.B(n_994),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_1018),
.B(n_966),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_1051),
.B(n_954),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_SL g1083 ( 
.A(n_1054),
.B(n_1038),
.Y(n_1083)
);

OAI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_1068),
.A2(n_973),
.B(n_957),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_1065),
.B(n_1002),
.Y(n_1085)
);

O2A1O1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_1062),
.A2(n_1069),
.B(n_1042),
.C(n_1025),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_1057),
.B(n_1002),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1059),
.B(n_973),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_L g1089 ( 
.A1(n_1072),
.A2(n_1061),
.B(n_1055),
.Y(n_1089)
);

INVx3_ASAP7_75t_L g1090 ( 
.A(n_1078),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_1082),
.A2(n_1068),
.B(n_1062),
.Y(n_1091)
);

INVx3_ASAP7_75t_L g1092 ( 
.A(n_1078),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_1086),
.B(n_1074),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1075),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_1079),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_1071),
.A2(n_1038),
.B(n_1027),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_1083),
.A2(n_1014),
.B(n_1007),
.Y(n_1097)
);

OAI21x1_ASAP7_75t_L g1098 ( 
.A1(n_1088),
.A2(n_1005),
.B(n_1045),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_1073),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1076),
.B(n_1019),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_1080),
.A2(n_1013),
.B(n_1039),
.C(n_1032),
.Y(n_1101)
);

A2O1A1Ixp33_ASAP7_75t_L g1102 ( 
.A1(n_1084),
.A2(n_1039),
.B(n_1032),
.C(n_1040),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_1085),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_SL g1104 ( 
.A1(n_1077),
.A2(n_1064),
.B(n_1063),
.Y(n_1104)
);

AOI21x1_ASAP7_75t_SL g1105 ( 
.A1(n_1081),
.A2(n_1015),
.B(n_1034),
.Y(n_1105)
);

NOR2x1_ASAP7_75t_L g1106 ( 
.A(n_1087),
.B(n_1070),
.Y(n_1106)
);

AOI21x1_ASAP7_75t_L g1107 ( 
.A1(n_1082),
.A2(n_1021),
.B(n_1060),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1086),
.B(n_1016),
.Y(n_1108)
);

AOI21x1_ASAP7_75t_L g1109 ( 
.A1(n_1082),
.A2(n_1063),
.B(n_1041),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_1082),
.A2(n_1027),
.B(n_1043),
.Y(n_1110)
);

OAI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_1082),
.A2(n_1053),
.B1(n_1047),
.B2(n_1064),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_1082),
.A2(n_1036),
.B(n_1047),
.Y(n_1112)
);

AO31x2_ASAP7_75t_L g1113 ( 
.A1(n_1074),
.A2(n_1070),
.A3(n_1026),
.B(n_1008),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1094),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_1095),
.B(n_1037),
.Y(n_1115)
);

OR2x2_ASAP7_75t_L g1116 ( 
.A(n_1100),
.B(n_1037),
.Y(n_1116)
);

INVx4_ASAP7_75t_L g1117 ( 
.A(n_1090),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1090),
.Y(n_1118)
);

INVxp67_ASAP7_75t_SL g1119 ( 
.A(n_1093),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_SL g1120 ( 
.A(n_1101),
.B(n_1054),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1120),
.A2(n_1108),
.B(n_1102),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_SL g1122 ( 
.A1(n_1119),
.A2(n_1110),
.B(n_1111),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_1121),
.A2(n_1107),
.B(n_1109),
.Y(n_1123)
);

A2O1A1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_1122),
.A2(n_1110),
.B(n_1096),
.C(n_1120),
.Y(n_1124)
);

BUFx3_ASAP7_75t_L g1125 ( 
.A(n_1123),
.Y(n_1125)
);

AOI22xp33_ASAP7_75t_L g1126 ( 
.A1(n_1124),
.A2(n_1119),
.B1(n_1117),
.B2(n_1118),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1123),
.Y(n_1127)
);

INVx1_ASAP7_75t_SL g1128 ( 
.A(n_1125),
.Y(n_1128)
);

HB1xp67_ASAP7_75t_L g1129 ( 
.A(n_1125),
.Y(n_1129)
);

AND2x4_ASAP7_75t_L g1130 ( 
.A(n_1127),
.B(n_1117),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1129),
.Y(n_1131)
);

NOR2x1_ASAP7_75t_SL g1132 ( 
.A(n_1130),
.B(n_1127),
.Y(n_1132)
);

INVx3_ASAP7_75t_L g1133 ( 
.A(n_1131),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_1132),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_1134),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1133),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1136),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1135),
.B(n_1130),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1138),
.Y(n_1139)
);

INVxp67_ASAP7_75t_L g1140 ( 
.A(n_1137),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_1139),
.Y(n_1141)
);

HB1xp67_ASAP7_75t_L g1142 ( 
.A(n_1140),
.Y(n_1142)
);

AND2x4_ASAP7_75t_L g1143 ( 
.A(n_1141),
.B(n_1133),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1142),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_1141),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1143),
.Y(n_1146)
);

NAND4xp25_ASAP7_75t_L g1147 ( 
.A(n_1144),
.B(n_1128),
.C(n_1126),
.D(n_1132),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_1145),
.B(n_1114),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_1148),
.B(n_1115),
.Y(n_1149)
);

AND2x2_ASAP7_75t_SL g1150 ( 
.A(n_1146),
.B(n_1116),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1150),
.B(n_1147),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_1149),
.B(n_1103),
.Y(n_1152)
);

HB1xp67_ASAP7_75t_L g1153 ( 
.A(n_1151),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_1152),
.Y(n_1154)
);

NAND2x1_ASAP7_75t_L g1155 ( 
.A(n_1154),
.B(n_1153),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1154),
.Y(n_1156)
);

AO221x2_ASAP7_75t_L g1157 ( 
.A1(n_1156),
.A2(n_1111),
.B1(n_1108),
.B2(n_1100),
.C(n_1104),
.Y(n_1157)
);

AOI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_1155),
.A2(n_1099),
.B1(n_1092),
.B2(n_1106),
.Y(n_1158)
);

NAND2xp33_ASAP7_75t_L g1159 ( 
.A(n_1158),
.B(n_1092),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_1157),
.Y(n_1160)
);

OR2x2_ASAP7_75t_L g1161 ( 
.A(n_1160),
.B(n_1113),
.Y(n_1161)
);

INVxp67_ASAP7_75t_SL g1162 ( 
.A(n_1159),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1160),
.Y(n_1163)
);

NOR2xp67_ASAP7_75t_L g1164 ( 
.A(n_1163),
.B(n_24),
.Y(n_1164)
);

OR2x2_ASAP7_75t_L g1165 ( 
.A(n_1161),
.B(n_1113),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1162),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_L g1167 ( 
.A(n_1166),
.B(n_25),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1164),
.B(n_1091),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1168),
.Y(n_1169)
);

AOI322xp5_ASAP7_75t_L g1170 ( 
.A1(n_1167),
.A2(n_1165),
.A3(n_1046),
.B1(n_1048),
.B2(n_1024),
.C1(n_1049),
.C2(n_1010),
.Y(n_1170)
);

OAI211xp5_ASAP7_75t_SL g1171 ( 
.A1(n_1169),
.A2(n_25),
.B(n_26),
.C(n_27),
.Y(n_1171)
);

INVxp67_ASAP7_75t_L g1172 ( 
.A(n_1170),
.Y(n_1172)
);

OR2x2_ASAP7_75t_L g1173 ( 
.A(n_1172),
.B(n_27),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1171),
.Y(n_1174)
);

NAND2x1p5_ASAP7_75t_L g1175 ( 
.A(n_1174),
.B(n_1097),
.Y(n_1175)
);

OAI322xp33_ASAP7_75t_L g1176 ( 
.A1(n_1173),
.A2(n_1112),
.A3(n_29),
.B1(n_30),
.B2(n_31),
.C1(n_32),
.C2(n_33),
.Y(n_1176)
);

INVx1_ASAP7_75t_SL g1177 ( 
.A(n_1176),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1175),
.Y(n_1178)
);

INVxp67_ASAP7_75t_L g1179 ( 
.A(n_1178),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1177),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1178),
.Y(n_1181)
);

OAI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1179),
.A2(n_1098),
.B(n_1089),
.Y(n_1182)
);

OAI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1181),
.A2(n_28),
.B(n_30),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1180),
.B(n_1113),
.Y(n_1184)
);

NOR3xp33_ASAP7_75t_L g1185 ( 
.A(n_1184),
.B(n_305),
.C(n_28),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1183),
.Y(n_1186)
);

AOI22xp33_ASAP7_75t_L g1187 ( 
.A1(n_1186),
.A2(n_1182),
.B1(n_1049),
.B2(n_1010),
.Y(n_1187)
);

O2A1O1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_1185),
.A2(n_31),
.B(n_32),
.C(n_33),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_SL g1189 ( 
.A1(n_1187),
.A2(n_1049),
.B1(n_1026),
.B2(n_34),
.Y(n_1189)
);

O2A1O1Ixp33_ASAP7_75t_L g1190 ( 
.A1(n_1188),
.A2(n_34),
.B(n_1046),
.C(n_370),
.Y(n_1190)
);

OAI31xp33_ASAP7_75t_L g1191 ( 
.A1(n_1190),
.A2(n_1105),
.A3(n_1052),
.B(n_39),
.Y(n_1191)
);

AOI211xp5_ASAP7_75t_SL g1192 ( 
.A1(n_1189),
.A2(n_37),
.B(n_38),
.C(n_42),
.Y(n_1192)
);

NOR5xp2_ASAP7_75t_L g1193 ( 
.A(n_1192),
.B(n_44),
.C(n_47),
.D(n_48),
.E(n_50),
.Y(n_1193)
);

OAI221xp5_ASAP7_75t_L g1194 ( 
.A1(n_1191),
.A2(n_52),
.B1(n_53),
.B2(n_56),
.C(n_60),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1194),
.A2(n_409),
.B(n_62),
.Y(n_1195)
);

HB1xp67_ASAP7_75t_L g1196 ( 
.A(n_1193),
.Y(n_1196)
);

NOR2x1_ASAP7_75t_L g1197 ( 
.A(n_1196),
.B(n_1054),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1195),
.Y(n_1198)
);

AND3x4_ASAP7_75t_L g1199 ( 
.A(n_1196),
.B(n_61),
.C(n_63),
.Y(n_1199)
);

NOR3xp33_ASAP7_75t_SL g1200 ( 
.A(n_1198),
.B(n_64),
.C(n_65),
.Y(n_1200)
);

OR2x2_ASAP7_75t_L g1201 ( 
.A(n_1197),
.B(n_66),
.Y(n_1201)
);

NOR3xp33_ASAP7_75t_SL g1202 ( 
.A(n_1199),
.B(n_67),
.C(n_68),
.Y(n_1202)
);

NOR3xp33_ASAP7_75t_L g1203 ( 
.A(n_1201),
.B(n_70),
.C(n_71),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1202),
.Y(n_1204)
);

XNOR2xp5_ASAP7_75t_L g1205 ( 
.A(n_1204),
.B(n_1200),
.Y(n_1205)
);

O2A1O1Ixp33_ASAP7_75t_SL g1206 ( 
.A1(n_1203),
.A2(n_72),
.B(n_73),
.C(n_74),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1205),
.Y(n_1207)
);

NAND4xp75_ASAP7_75t_L g1208 ( 
.A(n_1206),
.B(n_75),
.C(n_77),
.D(n_79),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1207),
.Y(n_1209)
);

AND2x4_ASAP7_75t_L g1210 ( 
.A(n_1208),
.B(n_80),
.Y(n_1210)
);

AOI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1209),
.A2(n_409),
.B1(n_84),
.B2(n_86),
.Y(n_1211)
);

AOI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1210),
.A2(n_409),
.B1(n_88),
.B2(n_89),
.Y(n_1212)
);

NAND2x1_ASAP7_75t_L g1213 ( 
.A(n_1212),
.B(n_83),
.Y(n_1213)
);

AOI211xp5_ASAP7_75t_L g1214 ( 
.A1(n_1211),
.A2(n_91),
.B(n_93),
.C(n_95),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1213),
.Y(n_1215)
);

OAI31xp33_ASAP7_75t_L g1216 ( 
.A1(n_1214),
.A2(n_97),
.A3(n_98),
.B(n_99),
.Y(n_1216)
);

OAI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1213),
.A2(n_100),
.B(n_101),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1215),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1216),
.B(n_104),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1217),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1218),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_1220),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1221),
.Y(n_1223)
);

OAI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_1222),
.A2(n_1219),
.B1(n_967),
.B2(n_108),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1223),
.Y(n_1225)
);

HB1xp67_ASAP7_75t_L g1226 ( 
.A(n_1224),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_SL g1227 ( 
.A1(n_1225),
.A2(n_967),
.B1(n_107),
.B2(n_109),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1226),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1228),
.A2(n_105),
.B(n_110),
.Y(n_1229)
);

AOI221xp5_ASAP7_75t_L g1230 ( 
.A1(n_1227),
.A2(n_111),
.B1(n_112),
.B2(n_114),
.C(n_115),
.Y(n_1230)
);

AOI21xp33_ASAP7_75t_L g1231 ( 
.A1(n_1228),
.A2(n_117),
.B(n_119),
.Y(n_1231)
);

XNOR2xp5_ASAP7_75t_L g1232 ( 
.A(n_1230),
.B(n_120),
.Y(n_1232)
);

NOR2xp67_ASAP7_75t_L g1233 ( 
.A(n_1229),
.B(n_121),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1231),
.B(n_122),
.Y(n_1234)
);

AOI22x1_ASAP7_75t_L g1235 ( 
.A1(n_1232),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_1235)
);

AOI22xp5_ASAP7_75t_L g1236 ( 
.A1(n_1233),
.A2(n_126),
.B1(n_127),
.B2(n_129),
.Y(n_1236)
);

AOI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1234),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_1237)
);

AOI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1232),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1235),
.A2(n_139),
.B(n_140),
.Y(n_1239)
);

AOI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1238),
.A2(n_142),
.B(n_143),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1237),
.Y(n_1241)
);

AOI22xp5_ASAP7_75t_L g1242 ( 
.A1(n_1236),
.A2(n_144),
.B1(n_146),
.B2(n_148),
.Y(n_1242)
);

NAND3xp33_ASAP7_75t_L g1243 ( 
.A(n_1235),
.B(n_152),
.C(n_154),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1235),
.A2(n_155),
.B(n_156),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1235),
.Y(n_1245)
);

AOI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1238),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_1246)
);

OAI22x1_ASAP7_75t_L g1247 ( 
.A1(n_1235),
.A2(n_160),
.B1(n_161),
.B2(n_162),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1235),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1235),
.A2(n_168),
.B(n_171),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1235),
.B(n_172),
.Y(n_1250)
);

NAND3xp33_ASAP7_75t_L g1251 ( 
.A(n_1241),
.B(n_174),
.C(n_175),
.Y(n_1251)
);

NAND3xp33_ASAP7_75t_L g1252 ( 
.A(n_1245),
.B(n_176),
.C(n_177),
.Y(n_1252)
);

AND2x2_ASAP7_75t_L g1253 ( 
.A(n_1250),
.B(n_1240),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1239),
.B(n_178),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1244),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_SL g1256 ( 
.A(n_1249),
.B(n_401),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1243),
.A2(n_380),
.B(n_383),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1247),
.B(n_384),
.Y(n_1258)
);

AOI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1255),
.A2(n_1248),
.B1(n_1242),
.B2(n_1246),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1253),
.A2(n_384),
.B1(n_397),
.B2(n_401),
.Y(n_1260)
);

AOI322xp5_ASAP7_75t_L g1261 ( 
.A1(n_1258),
.A2(n_380),
.A3(n_383),
.B1(n_1006),
.B2(n_1031),
.C1(n_988),
.C2(n_1067),
.Y(n_1261)
);

AOI22x1_ASAP7_75t_L g1262 ( 
.A1(n_1257),
.A2(n_964),
.B1(n_1006),
.B2(n_509),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1256),
.Y(n_1263)
);

AOI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1254),
.A2(n_1031),
.B1(n_1017),
.B2(n_509),
.Y(n_1264)
);

OAI21xp5_ASAP7_75t_SL g1265 ( 
.A1(n_1259),
.A2(n_1252),
.B(n_1251),
.Y(n_1265)
);

OAI211xp5_ASAP7_75t_SL g1266 ( 
.A1(n_1263),
.A2(n_1066),
.B(n_988),
.C(n_1033),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_L g1267 ( 
.A1(n_1264),
.A2(n_1053),
.B(n_1012),
.Y(n_1267)
);

OR2x6_ASAP7_75t_L g1268 ( 
.A(n_1262),
.B(n_1053),
.Y(n_1268)
);

AOI221xp5_ASAP7_75t_L g1269 ( 
.A1(n_1265),
.A2(n_1261),
.B1(n_1260),
.B2(n_1050),
.C(n_1030),
.Y(n_1269)
);

AOI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1269),
.A2(n_1268),
.B1(n_1267),
.B2(n_1266),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_L g1271 ( 
.A1(n_1270),
.A2(n_973),
.B1(n_1050),
.B2(n_1020),
.Y(n_1271)
);

AOI211xp5_ASAP7_75t_L g1272 ( 
.A1(n_1271),
.A2(n_1009),
.B(n_1029),
.C(n_1044),
.Y(n_1272)
);

AOI211xp5_ASAP7_75t_L g1273 ( 
.A1(n_1272),
.A2(n_973),
.B(n_950),
.C(n_989),
.Y(n_1273)
);


endmodule