module fake_jpeg_14388_n_188 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_188);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_188;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_23),
.B(n_8),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_37),
.B(n_48),
.Y(n_58)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_31),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_39),
.A2(n_43),
.B1(n_19),
.B2(n_27),
.Y(n_66)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

OA22x2_ASAP7_75t_L g43 ( 
.A1(n_22),
.A2(n_17),
.B1(n_26),
.B2(n_30),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

NAND2xp33_ASAP7_75t_SL g47 ( 
.A(n_20),
.B(n_1),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_33),
.C(n_32),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_28),
.B(n_2),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_68),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_26),
.B1(n_30),
.B2(n_16),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_55),
.A2(n_38),
.B1(n_42),
.B2(n_44),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_23),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_56),
.B(n_64),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_25),
.B1(n_33),
.B2(n_32),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_60),
.A2(n_38),
.B1(n_36),
.B2(n_35),
.Y(n_94)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_61),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_63),
.B(n_18),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_48),
.B(n_25),
.Y(n_64)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_43),
.B(n_19),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_65),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_66),
.A2(n_69),
.B(n_34),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_16),
.Y(n_68)
);

CKINVDCx6p67_ASAP7_75t_R g69 ( 
.A(n_35),
.Y(n_69)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_72),
.Y(n_82)
);

AOI21xp33_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_43),
.B(n_24),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_73),
.B(n_62),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_50),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_79),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_55),
.B(n_41),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_67),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_78),
.A2(n_58),
.B1(n_62),
.B2(n_52),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_69),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g98 ( 
.A1(n_80),
.A2(n_95),
.B(n_77),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_91),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_54),
.B(n_44),
.C(n_42),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_90),
.Y(n_102)
);

OAI21xp33_ASAP7_75t_SL g87 ( 
.A1(n_66),
.A2(n_29),
.B(n_24),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_94),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_29),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_50),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_74),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_51),
.A2(n_36),
.B1(n_18),
.B2(n_4),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_96),
.A2(n_34),
.B1(n_3),
.B2(n_4),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_100),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_98),
.A2(n_99),
.B(n_76),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_80),
.A2(n_71),
.B(n_61),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_57),
.Y(n_100)
);

AOI21xp33_ASAP7_75t_L g119 ( 
.A1(n_101),
.A2(n_114),
.B(n_111),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_67),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_116),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_106),
.Y(n_117)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_107),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_109),
.A2(n_89),
.B1(n_52),
.B2(n_62),
.Y(n_133)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

MAJx2_ASAP7_75t_L g112 ( 
.A(n_83),
.B(n_61),
.C(n_13),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_79),
.C(n_91),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_86),
.B(n_85),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_113),
.B(n_114),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_73),
.B(n_12),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_84),
.B(n_2),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_118),
.B(n_132),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_119),
.A2(n_123),
.B(n_126),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_108),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_133),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_101),
.A2(n_93),
.B1(n_82),
.B2(n_74),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_100),
.C(n_112),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_128),
.B(n_134),
.C(n_104),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_102),
.B(n_92),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_129),
.B(n_131),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_99),
.A2(n_89),
.B(n_82),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_130),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_116),
.B(n_11),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_11),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_98),
.B(n_88),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_107),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_140),
.C(n_118),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_97),
.Y(n_138)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_138),
.Y(n_152)
);

A2O1A1O1Ixp25_ASAP7_75t_L g142 ( 
.A1(n_127),
.A2(n_104),
.B(n_105),
.C(n_75),
.D(n_88),
.Y(n_142)
);

NOR3xp33_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_130),
.C(n_120),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_117),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_143),
.B(n_147),
.Y(n_151)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_125),
.Y(n_144)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_122),
.Y(n_145)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_145),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_124),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_110),
.Y(n_148)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_149),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_140),
.C(n_137),
.Y(n_163)
);

NOR3xp33_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_160),
.C(n_142),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_148),
.A2(n_121),
.B1(n_126),
.B2(n_134),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_155),
.A2(n_139),
.B1(n_138),
.B2(n_136),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_144),
.Y(n_157)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_157),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_139),
.A2(n_121),
.B(n_110),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_151),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_162),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_153),
.B(n_145),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_163),
.B(n_164),
.C(n_169),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_146),
.C(n_136),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_160),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_165),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_166),
.A2(n_153),
.B(n_152),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_168),
.B(n_155),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_159),
.A2(n_141),
.B1(n_135),
.B2(n_103),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_164),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_173),
.Y(n_178)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_169),
.A2(n_156),
.B(n_158),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_175),
.B(n_171),
.C(n_170),
.Y(n_180)
);

A2O1A1Ixp33_ASAP7_75t_SL g176 ( 
.A1(n_174),
.A2(n_168),
.B(n_152),
.C(n_167),
.Y(n_176)
);

A2O1A1Ixp33_ASAP7_75t_SL g183 ( 
.A1(n_176),
.A2(n_115),
.B(n_14),
.C(n_15),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_177),
.B(n_180),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_170),
.A2(n_157),
.B1(n_163),
.B2(n_103),
.Y(n_179)
);

AOI322xp5_ASAP7_75t_L g181 ( 
.A1(n_179),
.A2(n_75),
.A3(n_52),
.B1(n_115),
.B2(n_5),
.C1(n_3),
.C2(n_15),
.Y(n_181)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_181),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_183),
.B(n_184),
.C(n_176),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_178),
.B(n_176),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_186),
.B(n_182),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_185),
.Y(n_188)
);


endmodule