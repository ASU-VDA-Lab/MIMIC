module fake_jpeg_5042_n_102 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_102);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_102;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_32),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_14),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_13),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_25),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_5),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_3),
.Y(n_59)
);

INVx4_ASAP7_75t_SL g60 ( 
.A(n_58),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_61),
.Y(n_71)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_46),
.B(n_1),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_66),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_1),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_63),
.B(n_41),
.Y(n_72)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_65),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_49),
.Y(n_66)
);

AO22x1_ASAP7_75t_SL g67 ( 
.A1(n_62),
.A2(n_51),
.B1(n_41),
.B2(n_56),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_67),
.A2(n_73),
.B1(n_53),
.B2(n_50),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_47),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_63),
.A2(n_56),
.B1(n_57),
.B2(n_59),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_71),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_74),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_69),
.B(n_54),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_75),
.B(n_78),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_76),
.A2(n_77),
.B1(n_2),
.B2(n_4),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_69),
.A2(n_44),
.B1(n_40),
.B2(n_48),
.Y(n_77)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_76),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_80),
.B(n_82),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_76),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_43),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_76),
.A2(n_70),
.B1(n_68),
.B2(n_7),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_84),
.A2(n_85),
.B1(n_9),
.B2(n_10),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_12),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_87),
.A2(n_89),
.B(n_81),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_91),
.B(n_84),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g93 ( 
.A(n_92),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_93),
.A2(n_88),
.B1(n_79),
.B2(n_90),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_94),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_19),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_20),
.Y(n_97)
);

A2O1A1O1Ixp25_ASAP7_75t_L g98 ( 
.A1(n_97),
.A2(n_22),
.B(n_24),
.C(n_29),
.D(n_30),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_31),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_33),
.B(n_35),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_36),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_37),
.Y(n_102)
);


endmodule