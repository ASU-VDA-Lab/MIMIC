module fake_jpeg_1047_n_194 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_194);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_194;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

INVx13_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx4f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

HB1xp67_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_31),
.Y(n_73)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_19),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_38),
.B(n_22),
.Y(n_64)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_44),
.Y(n_54)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_41),
.Y(n_70)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_42),
.Y(n_53)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_45),
.Y(n_46)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_31),
.A2(n_18),
.B1(n_28),
.B2(n_25),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_49),
.A2(n_51),
.B1(n_29),
.B2(n_4),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_38),
.A2(n_18),
.B1(n_17),
.B2(n_25),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_50),
.A2(n_52),
.B1(n_62),
.B2(n_65),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_43),
.A2(n_28),
.B1(n_17),
.B2(n_22),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_36),
.A2(n_18),
.B1(n_24),
.B2(n_23),
.Y(n_52)
);

CKINVDCx12_ASAP7_75t_R g55 ( 
.A(n_29),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_39),
.B(n_27),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_64),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_32),
.B(n_13),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_61),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_13),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_34),
.A2(n_41),
.B1(n_40),
.B2(n_37),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_33),
.A2(n_27),
.B1(n_24),
.B2(n_23),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_42),
.A2(n_21),
.B1(n_20),
.B2(n_14),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_68),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_34),
.B(n_21),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_69),
.B(n_6),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_45),
.A2(n_41),
.B1(n_20),
.B2(n_35),
.Y(n_71)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_71),
.A2(n_29),
.B1(n_2),
.B2(n_3),
.Y(n_80)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_75),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_54),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_82),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_56),
.B(n_0),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_81),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_80),
.A2(n_87),
.B1(n_95),
.B2(n_89),
.Y(n_126)
);

AND2x2_ASAP7_75t_SL g81 ( 
.A(n_56),
.B(n_47),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_70),
.Y(n_82)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_11),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_92),
.Y(n_113)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

INVx6_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_1),
.B1(n_4),
.B2(n_6),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_88),
.A2(n_90),
.B1(n_79),
.B2(n_97),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_73),
.A2(n_1),
.B1(n_4),
.B2(n_6),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_98),
.Y(n_123)
);

NAND2x1_ASAP7_75t_L g96 ( 
.A(n_60),
.B(n_7),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_96),
.A2(n_76),
.B(n_89),
.Y(n_115)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_99),
.Y(n_127)
);

AOI21xp33_ASAP7_75t_L g100 ( 
.A1(n_60),
.A2(n_65),
.B(n_52),
.Y(n_100)
);

FAx1_ASAP7_75t_SL g119 ( 
.A(n_100),
.B(n_96),
.CI(n_81),
.CON(n_119),
.SN(n_119)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_101),
.Y(n_120)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_102),
.B(n_72),
.Y(n_109)
);

OR2x2_ASAP7_75t_SL g104 ( 
.A(n_50),
.B(n_60),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_104),
.A2(n_72),
.B(n_9),
.C(n_7),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_103),
.B(n_94),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_76),
.A2(n_10),
.B(n_11),
.C(n_59),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_107),
.A2(n_106),
.B(n_108),
.C(n_115),
.Y(n_143)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_109),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_114),
.A2(n_78),
.B1(n_102),
.B2(n_86),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_115),
.A2(n_119),
.B(n_104),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_81),
.B(n_76),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_124),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_83),
.B(n_74),
.Y(n_124)
);

NOR2x1_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_103),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_117),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_128),
.B(n_136),
.Y(n_151)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_123),
.Y(n_130)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_108),
.Y(n_148)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_134),
.A2(n_137),
.B1(n_143),
.B2(n_107),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_122),
.B(n_124),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_109),
.C(n_127),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_117),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_105),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_138),
.B(n_139),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_103),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_141),
.Y(n_153)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_142),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_147),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_148),
.B(n_150),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_112),
.C(n_119),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_152),
.B(n_154),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_119),
.C(n_118),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_141),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_156),
.B(n_121),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_140),
.Y(n_158)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_158),
.Y(n_171)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_153),
.Y(n_159)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_159),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_160),
.B(n_162),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_146),
.A2(n_132),
.B(n_137),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_161),
.A2(n_147),
.B(n_154),
.Y(n_169)
);

OAI322xp33_ASAP7_75t_L g162 ( 
.A1(n_155),
.A2(n_143),
.A3(n_140),
.B1(n_113),
.B2(n_135),
.C1(n_130),
.C2(n_129),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_133),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_163),
.B(n_165),
.Y(n_173)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_151),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_121),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_167),
.A2(n_127),
.B1(n_118),
.B2(n_120),
.Y(n_172)
);

XNOR2x1_ASAP7_75t_L g168 ( 
.A(n_166),
.B(n_148),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_166),
.C(n_157),
.Y(n_178)
);

OAI21xp33_ASAP7_75t_L g180 ( 
.A1(n_169),
.A2(n_114),
.B(n_145),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_175),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_164),
.A2(n_134),
.B1(n_126),
.B2(n_152),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_169),
.A2(n_161),
.B(n_158),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_176),
.A2(n_179),
.B(n_171),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_178),
.B(n_180),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_170),
.A2(n_163),
.B(n_159),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_177),
.A2(n_171),
.B1(n_173),
.B2(n_175),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_181),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_182),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_180),
.A2(n_174),
.B1(n_168),
.B2(n_145),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_183),
.B(n_125),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_186),
.B(n_181),
.Y(n_189)
);

OR2x6_ASAP7_75t_SL g188 ( 
.A(n_187),
.B(n_184),
.Y(n_188)
);

OAI21x1_ASAP7_75t_L g190 ( 
.A1(n_188),
.A2(n_189),
.B(n_185),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_190),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_188),
.A2(n_183),
.B1(n_125),
.B2(n_111),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_191),
.C(n_110),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_110),
.Y(n_194)
);


endmodule