module fake_jpeg_11970_n_648 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_648);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_648;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_442;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_587;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_538;
wire n_47;
wire n_312;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVx6_ASAP7_75t_SL g26 ( 
.A(n_11),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

CKINVDCx11_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_12),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_15),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_1),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g211 ( 
.A(n_63),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_64),
.Y(n_141)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_65),
.Y(n_196)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_66),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_67),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_68),
.Y(n_168)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx11_ASAP7_75t_L g145 ( 
.A(n_69),
.Y(n_145)
);

INVx13_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g207 ( 
.A(n_70),
.Y(n_207)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_71),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_33),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_72),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_73),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_74),
.Y(n_192)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_75),
.Y(n_133)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_76),
.Y(n_135)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_77),
.Y(n_144)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_78),
.Y(n_157)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_79),
.Y(n_136)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_80),
.Y(n_143)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_22),
.Y(n_81)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_81),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_82),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_83),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_84),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_18),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_85),
.B(n_95),
.Y(n_161)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_86),
.Y(n_149)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_20),
.Y(n_87)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_87),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_88),
.Y(n_156)
);

INVx6_ASAP7_75t_SL g89 ( 
.A(n_22),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g162 ( 
.A(n_89),
.Y(n_162)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_21),
.Y(n_90)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_90),
.Y(n_165)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_91),
.Y(n_173)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_24),
.Y(n_92)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_92),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_93),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_59),
.B(n_18),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_94),
.B(n_112),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_48),
.B(n_17),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_96),
.Y(n_213)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_97),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

INVx8_ASAP7_75t_L g185 ( 
.A(n_98),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_99),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_53),
.Y(n_100)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_100),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_40),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_102),
.Y(n_154)
);

BUFx12_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_103),
.Y(n_202)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_56),
.Y(n_104)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_104),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_39),
.Y(n_105)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_23),
.Y(n_106)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_106),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_39),
.Y(n_107)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_107),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_56),
.B(n_0),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_108),
.B(n_3),
.Y(n_170)
);

INVx4_ASAP7_75t_SL g109 ( 
.A(n_51),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_109),
.B(n_113),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_37),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_110),
.B(n_120),
.Y(n_147)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_30),
.Y(n_111)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_111),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_51),
.B(n_0),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_30),
.B(n_1),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_49),
.Y(n_114)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_114),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_44),
.B(n_1),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_115),
.B(n_125),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_52),
.Y(n_116)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_116),
.Y(n_194)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_44),
.Y(n_117)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_117),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_52),
.Y(n_118)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_118),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_25),
.Y(n_119)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_119),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g120 ( 
.A(n_37),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_46),
.Y(n_121)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_121),
.Y(n_176)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_46),
.Y(n_122)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_122),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_25),
.Y(n_123)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_123),
.Y(n_188)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_61),
.Y(n_124)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_124),
.Y(n_193)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_49),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_29),
.B(n_3),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_128),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_49),
.Y(n_127)
);

NAND2xp33_ASAP7_75t_SL g146 ( 
.A(n_127),
.B(n_130),
.Y(n_146)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_61),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_57),
.B(n_3),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_129),
.B(n_8),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_54),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_71),
.A2(n_27),
.B1(n_32),
.B2(n_55),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_138),
.A2(n_148),
.B1(n_153),
.B2(n_160),
.Y(n_223)
);

OA22x2_ASAP7_75t_L g139 ( 
.A1(n_97),
.A2(n_58),
.B1(n_27),
.B2(n_29),
.Y(n_139)
);

OA22x2_ASAP7_75t_L g282 ( 
.A1(n_139),
.A2(n_103),
.B1(n_14),
.B2(n_16),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_64),
.A2(n_32),
.B1(n_55),
.B2(n_58),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_105),
.A2(n_54),
.B1(n_45),
.B2(n_43),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_152),
.A2(n_167),
.B1(n_187),
.B2(n_201),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_86),
.A2(n_45),
.B1(n_57),
.B2(n_60),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_67),
.A2(n_43),
.B1(n_31),
.B2(n_60),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_86),
.A2(n_60),
.B1(n_57),
.B2(n_31),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_166),
.A2(n_172),
.B1(n_190),
.B2(n_205),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_68),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_170),
.B(n_13),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_72),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_113),
.B(n_5),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_174),
.B(n_179),
.Y(n_277)
);

AND2x2_ASAP7_75t_SL g177 ( 
.A(n_89),
.B(n_5),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_177),
.B(n_109),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_115),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_178),
.B(n_197),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_78),
.B(n_6),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_107),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_189),
.B(n_127),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_96),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_114),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_81),
.B(n_16),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_199),
.B(n_208),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_73),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_63),
.B(n_69),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_203),
.B(n_204),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_84),
.B(n_88),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_96),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_87),
.B(n_13),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_82),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_214),
.A2(n_101),
.B1(n_99),
.B2(n_118),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_215),
.B(n_250),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_177),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_216),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_184),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_217),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_135),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g296 ( 
.A(n_218),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_219),
.B(n_228),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_152),
.A2(n_106),
.B1(n_75),
.B2(n_123),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_220),
.Y(n_308)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_184),
.Y(n_221)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_221),
.Y(n_292)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_136),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g342 ( 
.A(n_224),
.Y(n_342)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_141),
.Y(n_225)
);

INVx6_ASAP7_75t_L g315 ( 
.A(n_225),
.Y(n_315)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_135),
.Y(n_227)
);

INVx4_ASAP7_75t_L g343 ( 
.A(n_227),
.Y(n_343)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_161),
.B(n_76),
.Y(n_228)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_143),
.Y(n_229)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_229),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_155),
.B(n_66),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_230),
.B(n_247),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g231 ( 
.A(n_211),
.Y(n_231)
);

INVx5_ASAP7_75t_L g347 ( 
.A(n_231),
.Y(n_347)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_151),
.Y(n_232)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_232),
.Y(n_294)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_141),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_233),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_177),
.A2(n_80),
.B(n_125),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_234),
.B(n_245),
.C(n_246),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_187),
.A2(n_119),
.B1(n_65),
.B2(n_74),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g349 ( 
.A1(n_235),
.A2(n_268),
.B1(n_270),
.B2(n_274),
.Y(n_349)
);

OAI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_197),
.A2(n_100),
.B1(n_98),
.B2(n_93),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_236),
.A2(n_269),
.B1(n_198),
.B2(n_185),
.Y(n_313)
);

INVx8_ASAP7_75t_L g237 ( 
.A(n_133),
.Y(n_237)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_237),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_143),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g327 ( 
.A(n_238),
.Y(n_327)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_180),
.Y(n_239)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_239),
.Y(n_300)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_173),
.Y(n_241)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_241),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_150),
.Y(n_242)
);

INVx8_ASAP7_75t_L g312 ( 
.A(n_242),
.Y(n_312)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_173),
.Y(n_243)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_243),
.Y(n_299)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_157),
.Y(n_244)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_244),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_158),
.B(n_91),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_158),
.B(n_120),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_164),
.B(n_70),
.Y(n_247)
);

INVx6_ASAP7_75t_L g248 ( 
.A(n_150),
.Y(n_248)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_248),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_145),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_249),
.B(n_252),
.Y(n_331)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_137),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_176),
.Y(n_251)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_251),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_202),
.B(n_120),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_140),
.Y(n_253)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_253),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_168),
.Y(n_254)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_254),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_196),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_255),
.Y(n_329)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_168),
.Y(n_256)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_256),
.Y(n_321)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_140),
.Y(n_257)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_257),
.Y(n_324)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_182),
.Y(n_258)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_258),
.Y(n_334)
);

INVx6_ASAP7_75t_L g259 ( 
.A(n_210),
.Y(n_259)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_259),
.Y(n_344)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_145),
.Y(n_260)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_260),
.Y(n_350)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_182),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_262),
.B(n_263),
.Y(n_330)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_194),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_193),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g352 ( 
.A(n_264),
.B(n_266),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_169),
.A2(n_130),
.B1(n_110),
.B2(n_83),
.Y(n_265)
);

OA21x2_ASAP7_75t_L g340 ( 
.A1(n_265),
.A2(n_283),
.B(n_285),
.Y(n_340)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_149),
.Y(n_266)
);

BUFx5_ASAP7_75t_L g267 ( 
.A(n_133),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_267),
.Y(n_318)
);

INVx6_ASAP7_75t_L g268 ( 
.A(n_210),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_185),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_271),
.B(n_273),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_169),
.B(n_116),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_272),
.B(n_278),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_139),
.B(n_110),
.Y(n_273)
);

INVx6_ASAP7_75t_L g274 ( 
.A(n_132),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_157),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_275),
.Y(n_339)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_175),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_276),
.Y(n_335)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_175),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_139),
.B(n_13),
.Y(n_279)
);

NAND2x1p5_ASAP7_75t_L g310 ( 
.A(n_279),
.B(n_282),
.Y(n_310)
);

INVx5_ASAP7_75t_L g280 ( 
.A(n_149),
.Y(n_280)
);

AND2x2_ASAP7_75t_SL g291 ( 
.A(n_280),
.B(n_289),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_146),
.A2(n_103),
.B1(n_102),
.B2(n_16),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_281),
.A2(n_290),
.B1(n_205),
.B2(n_190),
.Y(n_302)
);

INVx13_ASAP7_75t_L g283 ( 
.A(n_162),
.Y(n_283)
);

OAI21xp33_ASAP7_75t_L g285 ( 
.A1(n_178),
.A2(n_14),
.B(n_146),
.Y(n_285)
);

INVx6_ASAP7_75t_L g286 ( 
.A(n_132),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g333 ( 
.A1(n_286),
.A2(n_287),
.B1(n_288),
.B2(n_162),
.Y(n_333)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_159),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_147),
.Y(n_288)
);

INVx5_ASAP7_75t_L g289 ( 
.A(n_213),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_188),
.A2(n_183),
.B1(n_192),
.B2(n_213),
.Y(n_290)
);

AO22x2_ASAP7_75t_L g295 ( 
.A1(n_234),
.A2(n_142),
.B1(n_206),
.B2(n_198),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_295),
.B(n_336),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_222),
.A2(n_153),
.B1(n_212),
.B2(n_194),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_301),
.A2(n_306),
.B1(n_311),
.B2(n_319),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_302),
.A2(n_325),
.B1(n_328),
.B2(n_215),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_222),
.A2(n_166),
.B1(n_131),
.B2(n_195),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_216),
.A2(n_131),
.B1(n_195),
.B2(n_206),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_313),
.A2(n_317),
.B1(n_346),
.B2(n_250),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_269),
.A2(n_163),
.B1(n_200),
.B2(n_209),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_228),
.A2(n_191),
.B1(n_165),
.B2(n_144),
.Y(n_319)
);

OAI22xp33_ASAP7_75t_SL g325 ( 
.A1(n_282),
.A2(n_154),
.B1(n_183),
.B2(n_142),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_284),
.A2(n_163),
.B1(n_200),
.B2(n_209),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_326),
.A2(n_351),
.B1(n_301),
.B2(n_340),
.Y(n_385)
);

OAI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_282),
.A2(n_154),
.B1(n_134),
.B2(n_156),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_333),
.Y(n_356)
);

A2O1A1Ixp33_ASAP7_75t_L g336 ( 
.A1(n_215),
.A2(n_207),
.B(n_186),
.C(n_171),
.Y(n_336)
);

O2A1O1Ixp33_ASAP7_75t_SL g338 ( 
.A1(n_279),
.A2(n_181),
.B(n_207),
.C(n_192),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_338),
.B(n_241),
.Y(n_383)
);

MAJx2_ASAP7_75t_L g341 ( 
.A(n_277),
.B(n_134),
.C(n_156),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_341),
.B(n_283),
.C(n_280),
.Y(n_388)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_273),
.A2(n_211),
.B1(n_279),
.B2(n_223),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_265),
.A2(n_240),
.B1(n_282),
.B2(n_273),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_345),
.B(n_341),
.C(n_322),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_353),
.B(n_363),
.C(n_386),
.Y(n_412)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_291),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_354),
.B(n_364),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_330),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_355),
.B(n_367),
.Y(n_411)
);

AOI22xp33_ASAP7_75t_SL g358 ( 
.A1(n_308),
.A2(n_288),
.B1(n_237),
.B2(n_261),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_358),
.A2(n_359),
.B1(n_361),
.B2(n_382),
.Y(n_405)
);

AOI22xp33_ASAP7_75t_SL g361 ( 
.A1(n_308),
.A2(n_231),
.B1(n_260),
.B2(n_227),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_293),
.Y(n_362)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_362),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_298),
.B(n_345),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_304),
.B(n_226),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_365),
.A2(n_366),
.B1(n_372),
.B2(n_374),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_313),
.A2(n_285),
.B1(n_226),
.B2(n_274),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_330),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_332),
.B(n_245),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_368),
.B(n_369),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_332),
.B(n_245),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g370 ( 
.A(n_323),
.B(n_246),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_370),
.B(n_388),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_310),
.B(n_246),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_371),
.B(n_376),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_317),
.A2(n_286),
.B1(n_225),
.B2(n_248),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_350),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_373),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_310),
.A2(n_259),
.B1(n_256),
.B2(n_233),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_342),
.Y(n_375)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_375),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_330),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_310),
.A2(n_268),
.B1(n_254),
.B2(n_242),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_377),
.A2(n_387),
.B1(n_390),
.B2(n_365),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_329),
.B(n_278),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_378),
.B(n_379),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_352),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_342),
.Y(n_380)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_380),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_298),
.B(n_276),
.Y(n_381)
);

CKINVDCx14_ASAP7_75t_R g437 ( 
.A(n_381),
.Y(n_437)
);

AOI22xp33_ASAP7_75t_SL g382 ( 
.A1(n_306),
.A2(n_229),
.B1(n_243),
.B2(n_244),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_383),
.A2(n_389),
.B(n_327),
.Y(n_424)
);

INVx2_ASAP7_75t_SL g384 ( 
.A(n_350),
.Y(n_384)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_384),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_385),
.A2(n_397),
.B1(n_359),
.B2(n_360),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_323),
.B(n_218),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_351),
.A2(n_270),
.B1(n_238),
.B2(n_266),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_309),
.B(n_289),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_349),
.A2(n_267),
.B1(n_338),
.B2(n_322),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_342),
.Y(n_391)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_391),
.Y(n_416)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_300),
.Y(n_392)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_392),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_319),
.B(n_323),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_393),
.B(n_396),
.Y(n_432)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_300),
.Y(n_394)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_394),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_331),
.B(n_338),
.Y(n_395)
);

NOR2x1_ASAP7_75t_L g422 ( 
.A(n_395),
.B(n_352),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_295),
.B(n_311),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_340),
.A2(n_295),
.B1(n_336),
.B2(n_307),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_307),
.Y(n_398)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_398),
.Y(n_440)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_324),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g428 ( 
.A(n_399),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_295),
.B(n_335),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_400),
.B(n_334),
.Y(n_439)
);

AOI22xp33_ASAP7_75t_L g401 ( 
.A1(n_396),
.A2(n_340),
.B1(n_295),
.B2(n_337),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_401),
.A2(n_414),
.B1(n_395),
.B2(n_368),
.Y(n_449)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_362),
.Y(n_402)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_402),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_385),
.A2(n_321),
.B1(n_344),
.B2(n_337),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_403),
.A2(n_417),
.B1(n_436),
.B2(n_408),
.Y(n_467)
);

INVx2_ASAP7_75t_SL g413 ( 
.A(n_399),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_413),
.B(n_439),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_415),
.A2(n_386),
.B1(n_384),
.B2(n_375),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_400),
.A2(n_321),
.B1(n_344),
.B2(n_320),
.Y(n_417)
);

INVx4_ASAP7_75t_L g418 ( 
.A(n_373),
.Y(n_418)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_418),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_363),
.B(n_339),
.C(n_334),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_421),
.B(n_353),
.C(n_388),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_SL g454 ( 
.A(n_422),
.B(n_434),
.C(n_369),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_357),
.B(n_291),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_423),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_424),
.B(n_422),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_378),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_425),
.B(n_426),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_383),
.A2(n_296),
.B(n_347),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_430),
.A2(n_354),
.B(n_397),
.Y(n_443)
);

BUFx2_ASAP7_75t_L g433 ( 
.A(n_372),
.Y(n_433)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_433),
.Y(n_458)
);

NOR2x1_ASAP7_75t_L g434 ( 
.A(n_371),
.B(n_352),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_360),
.A2(n_320),
.B1(n_314),
.B2(n_315),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_366),
.A2(n_291),
.B1(n_293),
.B2(n_315),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_438),
.A2(n_382),
.B1(n_409),
.B2(n_414),
.Y(n_445)
);

OAI21xp33_ASAP7_75t_SL g441 ( 
.A1(n_357),
.A2(n_347),
.B(n_305),
.Y(n_441)
);

OAI21xp33_ASAP7_75t_SL g457 ( 
.A1(n_441),
.A2(n_411),
.B(n_408),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_443),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_445),
.A2(n_449),
.B1(n_452),
.B2(n_456),
.Y(n_481)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_446),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_447),
.B(n_464),
.C(n_471),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_SL g506 ( 
.A1(n_448),
.A2(n_455),
.B(n_318),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_425),
.B(n_367),
.Y(n_450)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_450),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_409),
.A2(n_353),
.B1(n_393),
.B2(n_358),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g453 ( 
.A1(n_430),
.A2(n_361),
.B(n_355),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g486 ( 
.A1(n_453),
.A2(n_468),
.B(n_423),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_454),
.B(n_403),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_405),
.A2(n_390),
.B1(n_387),
.B2(n_374),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_433),
.A2(n_376),
.B1(n_379),
.B2(n_377),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_457),
.A2(n_460),
.B1(n_461),
.B2(n_474),
.Y(n_492)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_419),
.Y(n_459)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_459),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_433),
.A2(n_381),
.B1(n_356),
.B2(n_389),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_438),
.A2(n_384),
.B1(n_364),
.B2(n_380),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_437),
.B(n_398),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_462),
.B(n_463),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_411),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_412),
.B(n_406),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_465),
.A2(n_467),
.B1(n_428),
.B2(n_407),
.Y(n_499)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_419),
.Y(n_466)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_466),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_424),
.A2(n_384),
.B(n_391),
.Y(n_468)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_435),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_470),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_412),
.B(n_386),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_417),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_472),
.Y(n_503)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_435),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_473),
.B(n_475),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_427),
.A2(n_394),
.B1(n_392),
.B2(n_370),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_440),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_410),
.B(n_370),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_476),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_SL g477 ( 
.A(n_427),
.B(n_343),
.Y(n_477)
);

AOI21xp33_ASAP7_75t_L g508 ( 
.A1(n_477),
.A2(n_418),
.B(n_429),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_410),
.B(n_303),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_SL g509 ( 
.A(n_478),
.B(n_343),
.Y(n_509)
);

OAI211xp5_ASAP7_75t_SL g483 ( 
.A1(n_454),
.A2(n_431),
.B(n_432),
.C(n_439),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_483),
.B(n_510),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_464),
.B(n_406),
.C(n_421),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_484),
.B(n_491),
.C(n_497),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_SL g534 ( 
.A1(n_486),
.A2(n_453),
.B(n_455),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_SL g487 ( 
.A(n_471),
.B(n_420),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_SL g515 ( 
.A(n_487),
.B(n_494),
.Y(n_515)
);

O2A1O1Ixp33_ASAP7_75t_L g489 ( 
.A1(n_469),
.A2(n_423),
.B(n_431),
.C(n_432),
.Y(n_489)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_489),
.Y(n_522)
);

XOR2x2_ASAP7_75t_L g490 ( 
.A(n_452),
.B(n_434),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_490),
.A2(n_502),
.B(n_506),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_464),
.B(n_404),
.C(n_407),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_SL g495 ( 
.A(n_471),
.B(n_440),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_SL g517 ( 
.A(n_495),
.B(n_500),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_L g496 ( 
.A1(n_472),
.A2(n_413),
.B1(n_436),
.B2(n_428),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_496),
.A2(n_499),
.B1(n_445),
.B2(n_458),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_447),
.B(n_416),
.C(n_404),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_447),
.B(n_416),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_498),
.B(n_444),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_SL g500 ( 
.A(n_448),
.B(n_413),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_443),
.A2(n_429),
.B(n_402),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_508),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_509),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_446),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_476),
.B(n_444),
.C(n_474),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_511),
.B(n_460),
.C(n_456),
.Y(n_530)
);

CKINVDCx16_ASAP7_75t_R g512 ( 
.A(n_468),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_512),
.B(n_468),
.Y(n_516)
);

XNOR2x1_ASAP7_75t_L g513 ( 
.A(n_494),
.B(n_449),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_513),
.B(n_518),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_491),
.B(n_465),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_514),
.B(n_521),
.Y(n_548)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_516),
.Y(n_545)
);

XOR2xp5_ASAP7_75t_L g520 ( 
.A(n_482),
.B(n_457),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g567 ( 
.A(n_520),
.B(n_527),
.Y(n_567)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_498),
.B(n_461),
.Y(n_521)
);

NOR3xp33_ASAP7_75t_SL g523 ( 
.A(n_479),
.B(n_450),
.C(n_463),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_SL g552 ( 
.A(n_523),
.B(n_485),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_481),
.A2(n_455),
.B1(n_467),
.B2(n_453),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_524),
.A2(n_538),
.B1(n_496),
.B2(n_502),
.Y(n_553)
);

INVxp33_ASAP7_75t_SL g526 ( 
.A(n_480),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_526),
.B(n_534),
.Y(n_565)
);

XOR2xp5_ASAP7_75t_L g527 ( 
.A(n_482),
.B(n_462),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_510),
.B(n_478),
.Y(n_528)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_528),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_530),
.B(n_543),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_L g549 ( 
.A1(n_533),
.A2(n_492),
.B1(n_505),
.B2(n_485),
.Y(n_549)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_480),
.Y(n_535)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_535),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_497),
.B(n_451),
.C(n_467),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_536),
.B(n_537),
.C(n_539),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_484),
.B(n_477),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_SL g538 ( 
.A1(n_481),
.A2(n_458),
.B1(n_475),
.B2(n_470),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_495),
.B(n_473),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_504),
.Y(n_540)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_540),
.Y(n_556)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_504),
.Y(n_541)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_541),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_487),
.B(n_451),
.C(n_459),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_542),
.B(n_500),
.C(n_490),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_504),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_519),
.B(n_479),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_SL g589 ( 
.A(n_546),
.B(n_550),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_549),
.A2(n_528),
.B1(n_520),
.B2(n_523),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_519),
.B(n_492),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_L g580 ( 
.A(n_551),
.B(n_515),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_L g571 ( 
.A1(n_552),
.A2(n_555),
.B1(n_558),
.B2(n_563),
.Y(n_571)
);

OAI22xp5_ASAP7_75t_SL g575 ( 
.A1(n_553),
.A2(n_564),
.B1(n_568),
.B2(n_525),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g555 ( 
.A1(n_524),
.A2(n_490),
.B1(n_503),
.B2(n_501),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_538),
.A2(n_503),
.B1(n_531),
.B2(n_522),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_529),
.B(n_511),
.C(n_501),
.Y(n_559)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_559),
.B(n_561),
.C(n_562),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_529),
.B(n_486),
.C(n_505),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_527),
.B(n_536),
.C(n_537),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_522),
.A2(n_489),
.B1(n_507),
.B2(n_506),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_530),
.A2(n_507),
.B1(n_483),
.B2(n_488),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g568 ( 
.A1(n_532),
.A2(n_493),
.B1(n_488),
.B2(n_466),
.Y(n_568)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_569),
.Y(n_601)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_557),
.Y(n_570)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_570),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_554),
.B(n_542),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_SL g606 ( 
.A(n_572),
.B(n_573),
.Y(n_606)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_556),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g599 ( 
.A1(n_575),
.A2(n_577),
.B1(n_578),
.B2(n_587),
.Y(n_599)
);

OAI21xp5_ASAP7_75t_L g576 ( 
.A1(n_565),
.A2(n_525),
.B(n_534),
.Y(n_576)
);

XNOR2xp5_ASAP7_75t_L g607 ( 
.A(n_576),
.B(n_580),
.Y(n_607)
);

OAI22xp5_ASAP7_75t_SL g577 ( 
.A1(n_553),
.A2(n_533),
.B1(n_513),
.B2(n_493),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_L g578 ( 
.A1(n_558),
.A2(n_521),
.B1(n_517),
.B2(n_514),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_562),
.B(n_518),
.C(n_539),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_579),
.B(n_583),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g581 ( 
.A1(n_545),
.A2(n_509),
.B1(n_517),
.B2(n_515),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_L g596 ( 
.A1(n_581),
.A2(n_585),
.B1(n_560),
.B2(n_565),
.Y(n_596)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_556),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_582),
.B(n_568),
.Y(n_602)
);

XNOR2xp5_ASAP7_75t_L g583 ( 
.A(n_548),
.B(n_442),
.Y(n_583)
);

XOR2xp5_ASAP7_75t_L g584 ( 
.A(n_548),
.B(n_442),
.Y(n_584)
);

XOR2xp5_ASAP7_75t_L g594 ( 
.A(n_584),
.B(n_566),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_545),
.A2(n_312),
.B1(n_297),
.B2(n_314),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_564),
.B(n_297),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_586),
.B(n_588),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_L g587 ( 
.A1(n_555),
.A2(n_312),
.B1(n_303),
.B2(n_299),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_544),
.B(n_299),
.C(n_324),
.Y(n_588)
);

MAJx2_ASAP7_75t_L g590 ( 
.A(n_580),
.B(n_561),
.C(n_551),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_L g613 ( 
.A(n_590),
.B(n_596),
.Y(n_613)
);

OAI22xp5_ASAP7_75t_L g591 ( 
.A1(n_569),
.A2(n_589),
.B1(n_570),
.B2(n_547),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_591),
.B(n_592),
.Y(n_611)
);

OAI22xp5_ASAP7_75t_L g592 ( 
.A1(n_589),
.A2(n_547),
.B1(n_563),
.B2(n_560),
.Y(n_592)
);

XOR2xp5_ASAP7_75t_L g612 ( 
.A(n_594),
.B(n_567),
.Y(n_612)
);

CKINVDCx20_ASAP7_75t_R g597 ( 
.A(n_571),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_597),
.B(n_600),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_574),
.B(n_559),
.C(n_544),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_602),
.B(n_573),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g603 ( 
.A(n_574),
.B(n_567),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_SL g610 ( 
.A(n_603),
.B(n_605),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_579),
.B(n_584),
.C(n_583),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_604),
.B(n_578),
.C(n_581),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g605 ( 
.A(n_588),
.B(n_566),
.Y(n_605)
);

OAI21xp5_ASAP7_75t_L g608 ( 
.A1(n_601),
.A2(n_576),
.B(n_575),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_L g631 ( 
.A1(n_608),
.A2(n_609),
.B(n_596),
.Y(n_631)
);

OAI21xp5_ASAP7_75t_L g609 ( 
.A1(n_601),
.A2(n_577),
.B(n_582),
.Y(n_609)
);

XOR2xp5_ASAP7_75t_L g630 ( 
.A(n_612),
.B(n_620),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_614),
.B(n_616),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_615),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_606),
.B(n_585),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_606),
.B(n_587),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_617),
.B(n_621),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_SL g619 ( 
.A(n_600),
.B(n_305),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_SL g626 ( 
.A(n_619),
.B(n_593),
.Y(n_626)
);

XOR2xp5_ASAP7_75t_L g620 ( 
.A(n_607),
.B(n_348),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g621 ( 
.A(n_604),
.B(n_348),
.C(n_316),
.Y(n_621)
);

OAI21xp5_ASAP7_75t_SL g624 ( 
.A1(n_618),
.A2(n_614),
.B(n_610),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g634 ( 
.A1(n_624),
.A2(n_627),
.B(n_629),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g625 ( 
.A(n_613),
.B(n_595),
.C(n_590),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_625),
.B(n_626),
.Y(n_632)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_613),
.B(n_597),
.C(n_599),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_611),
.B(n_598),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_SL g636 ( 
.A1(n_631),
.A2(n_620),
.B(n_599),
.Y(n_636)
);

MAJIxp5_ASAP7_75t_L g633 ( 
.A(n_622),
.B(n_608),
.C(n_621),
.Y(n_633)
);

INVxp33_ASAP7_75t_L g642 ( 
.A(n_633),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_625),
.A2(n_607),
.B(n_609),
.Y(n_635)
);

OAI21xp5_ASAP7_75t_L g640 ( 
.A1(n_635),
.A2(n_636),
.B(n_638),
.Y(n_640)
);

MAJIxp5_ASAP7_75t_L g637 ( 
.A(n_623),
.B(n_612),
.C(n_593),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_637),
.B(n_628),
.Y(n_641)
);

OAI21xp5_ASAP7_75t_L g638 ( 
.A1(n_631),
.A2(n_594),
.B(n_292),
.Y(n_638)
);

NOR2xp67_ASAP7_75t_L g639 ( 
.A(n_634),
.B(n_627),
.Y(n_639)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_639),
.Y(n_643)
);

AOI321xp33_ASAP7_75t_L g644 ( 
.A1(n_641),
.A2(n_632),
.A3(n_630),
.B1(n_292),
.B2(n_316),
.C(n_294),
.Y(n_644)
);

OAI21xp5_ASAP7_75t_L g645 ( 
.A1(n_644),
.A2(n_640),
.B(n_642),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_645),
.B(n_643),
.Y(n_646)
);

XNOR2xp5_ASAP7_75t_L g647 ( 
.A(n_646),
.B(n_630),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_SL g648 ( 
.A(n_647),
.B(n_294),
.Y(n_648)
);


endmodule