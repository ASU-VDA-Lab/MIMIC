module real_jpeg_32579_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_666, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_666;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_657;
wire n_656;
wire n_643;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_640;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_620;
wire n_456;
wire n_578;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_393;
wire n_221;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_631;
wire n_175;
wire n_653;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_411;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_579;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_638;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_307;
wire n_316;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_586;
wire n_412;
wire n_405;
wire n_572;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_537;
wire n_318;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_662;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_545;
wire n_201;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_660;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_625;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_0),
.Y(n_205)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_0),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_0),
.Y(n_351)
);

BUFx12f_ASAP7_75t_L g491 ( 
.A(n_0),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_1),
.A2(n_66),
.B1(n_72),
.B2(n_73),
.Y(n_65)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_1),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_1),
.A2(n_72),
.B1(n_178),
.B2(n_182),
.Y(n_177)
);

OAI22x1_ASAP7_75t_L g293 ( 
.A1(n_1),
.A2(n_72),
.B1(n_294),
.B2(n_299),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g353 ( 
.A1(n_1),
.A2(n_72),
.B1(n_354),
.B2(n_358),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_3),
.A2(n_114),
.B1(n_118),
.B2(n_119),
.Y(n_113)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_3),
.Y(n_118)
);

AO22x1_ASAP7_75t_SL g212 ( 
.A1(n_3),
.A2(n_118),
.B1(n_213),
.B2(n_215),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_3),
.A2(n_118),
.B1(n_251),
.B2(n_256),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_4),
.A2(n_323),
.B1(n_325),
.B2(n_326),
.Y(n_322)
);

INVx1_ASAP7_75t_SL g325 ( 
.A(n_4),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_4),
.A2(n_325),
.B1(n_384),
.B2(n_385),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_SL g520 ( 
.A1(n_4),
.A2(n_325),
.B1(n_521),
.B2(n_523),
.Y(n_520)
);

AOI22xp33_ASAP7_75t_L g541 ( 
.A1(n_4),
.A2(n_325),
.B1(n_542),
.B2(n_545),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_5),
.B(n_75),
.Y(n_286)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_5),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_5),
.B(n_79),
.Y(n_424)
);

OAI32xp33_ASAP7_75t_L g502 ( 
.A1(n_5),
.A2(n_503),
.A3(n_505),
.B1(n_510),
.B2(n_514),
.Y(n_502)
);

OAI21xp33_ASAP7_75t_L g578 ( 
.A1(n_5),
.A2(n_348),
.B(n_579),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g628 ( 
.A1(n_5),
.A2(n_403),
.B1(n_629),
.B2(n_633),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_6),
.A2(n_56),
.B1(n_60),
.B2(n_61),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_6),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_6),
.A2(n_60),
.B1(n_224),
.B2(n_363),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_6),
.A2(n_60),
.B1(n_376),
.B2(n_379),
.Y(n_375)
);

AO22x1_ASAP7_75t_L g427 ( 
.A1(n_6),
.A2(n_60),
.B1(n_428),
.B2(n_431),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_7),
.A2(n_314),
.B1(n_315),
.B2(n_317),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_7),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_7),
.A2(n_314),
.B1(n_407),
.B2(n_410),
.Y(n_406)
);

AOI22xp33_ASAP7_75t_SL g534 ( 
.A1(n_7),
.A2(n_314),
.B1(n_535),
.B2(n_537),
.Y(n_534)
);

AOI22xp33_ASAP7_75t_SL g606 ( 
.A1(n_7),
.A2(n_314),
.B1(n_607),
.B2(n_610),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_8),
.Y(n_196)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_9),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_9),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_10),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_10),
.Y(n_94)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_10),
.Y(n_211)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_10),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_11),
.A2(n_156),
.B1(n_159),
.B2(n_160),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_11),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_11),
.A2(n_159),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g341 ( 
.A1(n_11),
.A2(n_159),
.B1(n_342),
.B2(n_345),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_12),
.A2(n_193),
.B1(n_197),
.B2(n_198),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_12),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_12),
.A2(n_197),
.B1(n_333),
.B2(n_334),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_12),
.A2(n_197),
.B1(n_393),
.B2(n_395),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g494 ( 
.A1(n_12),
.A2(n_197),
.B1(n_495),
.B2(n_500),
.Y(n_494)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_13),
.Y(n_90)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_13),
.Y(n_106)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_13),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_14),
.A2(n_149),
.B1(n_151),
.B2(n_152),
.Y(n_148)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_14),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_14),
.A2(n_151),
.B1(n_221),
.B2(n_224),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_14),
.A2(n_151),
.B1(n_239),
.B2(n_242),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_14),
.A2(n_151),
.B1(n_307),
.B2(n_309),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_15),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_15),
.Y(n_662)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_16),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_16),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_16),
.Y(n_117)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_16),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g659 ( 
.A(n_17),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_18),
.Y(n_140)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_18),
.Y(n_154)
);

OAI311xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_265),
.A3(n_656),
.B1(n_660),
.C1(n_663),
.Y(n_19)
);

INVxp67_ASAP7_75t_SL g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_21),
.B(n_656),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_264),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_227),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_24),
.B(n_227),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_167),
.C(n_186),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g653 ( 
.A(n_26),
.B(n_167),
.Y(n_653)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_80),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_27),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_55),
.B1(n_65),
.B2(n_78),
.Y(n_27)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_28),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2x1_ASAP7_75t_L g191 ( 
.A(n_29),
.B(n_192),
.Y(n_191)
);

AO22x1_ASAP7_75t_L g382 ( 
.A1(n_29),
.A2(n_79),
.B1(n_313),
.B2(n_383),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_29),
.B(n_401),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_29),
.B(n_383),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_45),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_34),
.B1(n_37),
.B2(n_41),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_33),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_33),
.Y(n_285)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_35),
.Y(n_281)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g244 ( 
.A(n_38),
.Y(n_244)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_38),
.Y(n_384)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_42),
.Y(n_41)
);

INVx4_ASAP7_75t_SL g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_44),
.Y(n_291)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

AOI22x1_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_48),
.Y(n_150)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx5_ASAP7_75t_L g288 ( 
.A(n_53),
.Y(n_288)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_54),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_54),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_55),
.B(n_79),
.Y(n_190)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_65),
.Y(n_236)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_71),
.Y(n_386)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_78),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_79),
.B(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_79),
.B(n_192),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_124),
.B2(n_166),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_81),
.A2(n_82),
.B1(n_247),
.B2(n_260),
.Y(n_246)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp33_ASAP7_75t_R g229 ( 
.A(n_82),
.B(n_166),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_82),
.B(n_166),
.Y(n_232)
);

OA21x2_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_97),
.B(n_113),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_83),
.A2(n_97),
.B1(n_113),
.B2(n_170),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_83),
.A2(n_97),
.B1(n_392),
.B2(n_397),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_83),
.B(n_392),
.Y(n_524)
);

INVx1_ASAP7_75t_SL g593 ( 
.A(n_83),
.Y(n_593)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_84),
.Y(n_219)
);

OAI22x1_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_88),
.B1(n_91),
.B2(n_95),
.Y(n_84)
);

INVx4_ASAP7_75t_L g544 ( 
.A(n_85),
.Y(n_544)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_87),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_87),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g536 ( 
.A(n_87),
.Y(n_536)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_90),
.Y(n_96)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_93),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g308 ( 
.A(n_93),
.Y(n_308)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_94),
.Y(n_566)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_97),
.B(n_571),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_97),
.B(n_392),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g623 ( 
.A1(n_97),
.A2(n_624),
.B1(n_625),
.B2(n_626),
.Y(n_623)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_98),
.A2(n_171),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_98),
.A2(n_219),
.B1(n_220),
.B2(n_353),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_98),
.A2(n_219),
.B1(n_353),
.B2(n_362),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g519 ( 
.A1(n_98),
.A2(n_520),
.B(n_524),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_103),
.B1(n_107),
.B2(n_110),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_102),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_102),
.Y(n_357)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_102),
.Y(n_366)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx6_ASAP7_75t_L g561 ( 
.A(n_105),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_112),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_112),
.Y(n_609)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_116),
.Y(n_172)
);

BUFx2_ASAP7_75t_L g358 ( 
.A(n_116),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g394 ( 
.A(n_116),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_117),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_117),
.Y(n_225)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_122),
.Y(n_133)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_122),
.Y(n_522)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_124),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_148),
.B1(n_155),
.B2(n_163),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_125),
.A2(n_148),
.B1(n_163),
.B2(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_125),
.Y(n_249)
);

AOI22x1_ASAP7_75t_L g405 ( 
.A1(n_125),
.A2(n_163),
.B1(n_406),
.B2(n_411),
.Y(n_405)
);

NAND2xp33_ASAP7_75t_SL g423 ( 
.A(n_125),
.B(n_332),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_125),
.A2(n_165),
.B1(n_177),
.B2(n_375),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_137),
.Y(n_125)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_126),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_130),
.B1(n_133),
.B2(n_134),
.Y(n_126)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_128),
.Y(n_517)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g575 ( 
.A(n_129),
.Y(n_575)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_132),
.Y(n_146)
);

INVx5_ASAP7_75t_SL g134 ( 
.A(n_135),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_136),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_141),
.B1(n_144),
.B2(n_147),
.Y(n_137)
);

INVx2_ASAP7_75t_SL g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_139),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_139),
.Y(n_409)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_139),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_140),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_140),
.Y(n_279)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_140),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_140),
.Y(n_632)
);

INVx2_ASAP7_75t_SL g141 ( 
.A(n_142),
.Y(n_141)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_143),
.Y(n_513)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_153),
.Y(n_185)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_153),
.Y(n_324)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_153),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_154),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_154),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_155),
.A2(n_163),
.B1(n_248),
.B2(n_250),
.Y(n_247)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g373 ( 
.A(n_164),
.B(n_374),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_164),
.A2(n_422),
.B(n_423),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g604 ( 
.A(n_164),
.B(n_403),
.Y(n_604)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_165),
.B(n_332),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

NAND2x1_ASAP7_75t_L g442 ( 
.A(n_168),
.B(n_443),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_176),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g443 ( 
.A(n_169),
.B(n_176),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g568 ( 
.A(n_174),
.Y(n_568)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_175),
.Y(n_396)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g652 ( 
.A(n_187),
.B(n_653),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_200),
.B1(n_226),
.B2(n_666),
.Y(n_187)
);

HB1xp67_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g445 ( 
.A(n_189),
.B(n_226),
.Y(n_445)
);

NAND2x1_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_191),
.B(n_312),
.Y(n_311)
);

INVx3_ASAP7_75t_SL g193 ( 
.A(n_194),
.Y(n_193)
);

INVx4_ASAP7_75t_SL g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_196),
.Y(n_241)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_196),
.Y(n_319)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_198),
.Y(n_402)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XNOR2x1_ASAP7_75t_L g444 ( 
.A(n_200),
.B(n_445),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_218),
.Y(n_200)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_201),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_201),
.A2(n_218),
.B1(n_226),
.B2(n_459),
.Y(n_458)
);

OA21x2_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_206),
.B(n_212),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_205),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_205),
.Y(n_584)
);

HB1xp67_ASAP7_75t_L g596 ( 
.A(n_205),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_205),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_206),
.A2(n_293),
.B1(n_302),
.B2(n_306),
.Y(n_292)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_206),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_206),
.B(n_494),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g532 ( 
.A1(n_206),
.A2(n_433),
.B1(n_533),
.B2(n_540),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_207),
.A2(n_341),
.B1(n_348),
.B2(n_368),
.Y(n_367)
);

INVx3_ASAP7_75t_SL g433 ( 
.A(n_207),
.Y(n_433)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_211),
.Y(n_217)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_211),
.Y(n_298)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_211),
.Y(n_344)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_211),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g556 ( 
.A(n_211),
.Y(n_556)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_212),
.Y(n_349)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_215),
.Y(n_309)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g539 ( 
.A(n_217),
.Y(n_539)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_218),
.Y(n_459)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_219),
.Y(n_625)
);

INVx1_ASAP7_75t_SL g610 ( 
.A(n_221),
.Y(n_610)
);

INVx4_ASAP7_75t_SL g221 ( 
.A(n_222),
.Y(n_221)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_233),
.B1(n_234),
.B2(n_261),
.Y(n_227)
);

OAI21xp33_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_230),
.B(n_231),
.Y(n_228)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_229),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_230),
.B(n_232),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_230),
.A2(n_232),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_230),
.Y(n_262)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_246),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_238),
.B2(n_245),
.Y(n_235)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_247),
.Y(n_260)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_249),
.A2(n_322),
.B(n_331),
.Y(n_321)
);

OAI21x1_ASAP7_75t_L g371 ( 
.A1(n_249),
.A2(n_372),
.B(n_373),
.Y(n_371)
);

OA21x2_ASAP7_75t_L g627 ( 
.A1(n_249),
.A2(n_331),
.B(n_628),
.Y(n_627)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_253),
.B(n_511),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_255),
.Y(n_504)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_258),
.Y(n_333)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_265),
.B(n_664),
.Y(n_663)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_648),
.B(n_654),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_267),
.Y(n_266)
);

NAND2x1_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_475),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_269),
.A2(n_437),
.B(n_471),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_387),
.C(n_414),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g477 ( 
.A1(n_271),
.A2(n_478),
.B(n_479),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_337),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_273),
.B(n_339),
.C(n_470),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_310),
.C(n_320),
.Y(n_273)
);

XNOR2x1_ASAP7_75t_L g388 ( 
.A(n_274),
.B(n_389),
.Y(n_388)
);

OR2x2_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_292),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_275),
.B(n_292),
.Y(n_418)
);

AOI32xp33_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_280),
.A3(n_282),
.B1(n_286),
.B2(n_287),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx11_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

BUFx12f_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx3_ASAP7_75t_SL g316 ( 
.A(n_285),
.Y(n_316)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_286),
.Y(n_404)
);

NAND2xp33_ASAP7_75t_R g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_293),
.B(n_433),
.Y(n_432)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_SL g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_305),
.Y(n_590)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_306),
.Y(n_368)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_310),
.A2(n_311),
.B1(n_320),
.B2(n_321),
.Y(n_389)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_322),
.Y(n_411)
);

INVx1_ASAP7_75t_SL g323 ( 
.A(n_324),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVxp67_ASAP7_75t_SL g372 ( 
.A(n_332),
.Y(n_372)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_359),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_352),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g447 ( 
.A(n_340),
.B(n_352),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_341),
.A2(n_348),
.B1(n_349),
.B2(n_350),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g585 ( 
.A(n_342),
.B(n_586),
.Y(n_585)
);

INVx5_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g345 ( 
.A(n_346),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx4_ASAP7_75t_L g430 ( 
.A(n_347),
.Y(n_430)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_348),
.A2(n_427),
.B(n_432),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g602 ( 
.A1(n_348),
.A2(n_541),
.B(n_579),
.Y(n_602)
);

INVx5_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx5_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_357),
.Y(n_523)
);

INVxp67_ASAP7_75t_SL g470 ( 
.A(n_359),
.Y(n_470)
);

XNOR2x1_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_369),
.Y(n_359)
);

MAJx2_ASAP7_75t_L g456 ( 
.A(n_360),
.B(n_382),
.C(n_457),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_367),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_SL g413 ( 
.A(n_361),
.B(n_367),
.Y(n_413)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_362),
.Y(n_397)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

BUFx4f_ASAP7_75t_SL g364 ( 
.A(n_365),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

AOI22x1_ASAP7_75t_L g369 ( 
.A1(n_370),
.A2(n_371),
.B1(n_381),
.B2(n_382),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g457 ( 
.A(n_371),
.Y(n_457)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx8_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_387),
.Y(n_478)
);

MAJx2_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_390),
.C(n_412),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_388),
.B(n_435),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_390),
.A2(n_412),
.B1(n_413),
.B2(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_390),
.Y(n_436)
);

MAJx2_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_398),
.C(n_405),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_391),
.B(n_405),
.Y(n_417)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx2_ASAP7_75t_SL g395 ( 
.A(n_396),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_398),
.B(n_417),
.Y(n_416)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_400),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_399),
.B(n_450),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_402),
.A2(n_403),
.B(n_404),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_403),
.B(n_515),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_403),
.B(n_508),
.Y(n_553)
);

OAI21xp33_ASAP7_75t_L g571 ( 
.A1(n_403),
.A2(n_553),
.B(n_572),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g586 ( 
.A(n_403),
.B(n_587),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_SL g592 ( 
.A(n_403),
.B(n_593),
.Y(n_592)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_406),
.Y(n_422)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx4_ASAP7_75t_L g410 ( 
.A(n_409),
.Y(n_410)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

OR2x2_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_434),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_415),
.B(n_434),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_418),
.C(n_419),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_416),
.B(n_483),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_418),
.A2(n_419),
.B1(n_420),
.B2(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_418),
.Y(n_484)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_424),
.C(n_425),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_421),
.B(n_527),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_424),
.B(n_426),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_R g488 ( 
.A(n_427),
.B(n_489),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g619 ( 
.A1(n_427),
.A2(n_493),
.B(n_620),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g428 ( 
.A(n_429),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_430),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_438),
.B(n_477),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_439),
.A2(n_454),
.B(n_465),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_439),
.B(n_454),
.Y(n_474)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_440),
.B(n_455),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_446),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_444),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g650 ( 
.A(n_442),
.B(n_444),
.C(n_651),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_446),
.Y(n_651)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_448),
.C(n_451),
.Y(n_446)
);

XNOR2x1_ASAP7_75t_L g462 ( 
.A(n_447),
.B(n_463),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_449),
.A2(n_452),
.B1(n_453),
.B2(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_449),
.Y(n_464)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_458),
.C(n_460),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_456),
.B(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_458),
.Y(n_468)
);

INVxp67_ASAP7_75t_SL g460 ( 
.A(n_461),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_462),
.B(n_468),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_469),
.Y(n_465)
);

OR2x2_ASAP7_75t_L g472 ( 
.A(n_466),
.B(n_469),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_L g471 ( 
.A1(n_472),
.A2(n_473),
.B(n_474),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_480),
.Y(n_475)
);

OAI21x1_ASAP7_75t_L g480 ( 
.A1(n_481),
.A2(n_528),
.B(n_646),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_485),
.Y(n_481)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_482),
.Y(n_647)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_486),
.B(n_647),
.Y(n_646)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_518),
.C(n_525),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g640 ( 
.A1(n_487),
.A2(n_518),
.B1(n_519),
.B2(n_641),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_487),
.Y(n_641)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_488),
.A2(n_492),
.B(n_502),
.Y(n_487)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx8_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVxp67_ASAP7_75t_SL g492 ( 
.A(n_493),
.Y(n_492)
);

OAI21xp33_ASAP7_75t_SL g594 ( 
.A1(n_493),
.A2(n_534),
.B(n_595),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_494),
.B(n_580),
.Y(n_579)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

BUFx3_ASAP7_75t_L g496 ( 
.A(n_497),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_499),
.Y(n_549)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g618 ( 
.A(n_502),
.B(n_619),
.Y(n_618)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_504),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

INVx4_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_520),
.Y(n_626)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_524),
.B(n_570),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g639 ( 
.A(n_526),
.B(n_640),
.Y(n_639)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_529),
.A2(n_637),
.B(n_645),
.Y(n_528)
);

O2A1O1Ixp5_ASAP7_75t_L g529 ( 
.A1(n_530),
.A2(n_599),
.B(n_612),
.C(n_613),
.Y(n_529)
);

AOI21x1_ASAP7_75t_L g530 ( 
.A1(n_531),
.A2(n_576),
.B(n_598),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_532),
.B(n_550),
.Y(n_531)
);

NOR2xp67_ASAP7_75t_L g598 ( 
.A(n_532),
.B(n_550),
.Y(n_598)
);

INVxp67_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g535 ( 
.A(n_536),
.Y(n_535)
);

INVx1_ASAP7_75t_SL g537 ( 
.A(n_538),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

INVxp33_ASAP7_75t_SL g540 ( 
.A(n_541),
.Y(n_540)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_551),
.B(n_569),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_551),
.B(n_569),
.Y(n_600)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_552),
.A2(n_554),
.B1(n_562),
.B2(n_567),
.Y(n_551)
);

INVxp67_ASAP7_75t_SL g552 ( 
.A(n_553),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_555),
.B(n_557),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_556),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_557),
.B(n_568),
.Y(n_567)
);

BUFx2_ASAP7_75t_L g557 ( 
.A(n_558),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_559),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

INVx1_ASAP7_75t_SL g562 ( 
.A(n_563),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_564),
.Y(n_563)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_565),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_566),
.Y(n_565)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_573),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_574),
.Y(n_573)
);

INVx4_ASAP7_75t_L g574 ( 
.A(n_575),
.Y(n_574)
);

OAI21xp33_ASAP7_75t_L g576 ( 
.A1(n_577),
.A2(n_591),
.B(n_597),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_578),
.B(n_585),
.Y(n_577)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_581),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_582),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_583),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g583 ( 
.A(n_584),
.Y(n_583)
);

INVx4_ASAP7_75t_L g587 ( 
.A(n_588),
.Y(n_587)
);

INVx4_ASAP7_75t_L g588 ( 
.A(n_589),
.Y(n_588)
);

INVx2_ASAP7_75t_SL g589 ( 
.A(n_590),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_592),
.B(n_594),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_592),
.B(n_594),
.Y(n_597)
);

OAI21xp5_ASAP7_75t_L g605 ( 
.A1(n_593),
.A2(n_606),
.B(n_611),
.Y(n_605)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_596),
.Y(n_595)
);

NOR2xp67_ASAP7_75t_L g599 ( 
.A(n_600),
.B(n_601),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_600),
.B(n_601),
.Y(n_612)
);

XNOR2xp5_ASAP7_75t_SL g601 ( 
.A(n_602),
.B(n_603),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_602),
.B(n_615),
.C(n_616),
.Y(n_614)
);

XNOR2xp5_ASAP7_75t_L g603 ( 
.A(n_604),
.B(n_605),
.Y(n_603)
);

HB1xp67_ASAP7_75t_L g616 ( 
.A(n_604),
.Y(n_616)
);

HB1xp67_ASAP7_75t_L g615 ( 
.A(n_605),
.Y(n_615)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_606),
.Y(n_624)
);

INVx1_ASAP7_75t_SL g607 ( 
.A(n_608),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_609),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_614),
.B(n_617),
.Y(n_613)
);

OR2x2_ASAP7_75t_L g644 ( 
.A(n_614),
.B(n_617),
.Y(n_644)
);

XOR2xp5_ASAP7_75t_L g617 ( 
.A(n_618),
.B(n_622),
.Y(n_617)
);

INVxp67_ASAP7_75t_L g643 ( 
.A(n_618),
.Y(n_643)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_621),
.Y(n_620)
);

XNOR2xp5_ASAP7_75t_L g622 ( 
.A(n_623),
.B(n_627),
.Y(n_622)
);

MAJIxp5_ASAP7_75t_L g642 ( 
.A(n_623),
.B(n_627),
.C(n_643),
.Y(n_642)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_630),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_631),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_632),
.Y(n_631)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_634),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_635),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_636),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_638),
.B(n_644),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_639),
.B(n_642),
.Y(n_638)
);

OR2x2_ASAP7_75t_L g645 ( 
.A(n_639),
.B(n_642),
.Y(n_645)
);

INVxp33_ASAP7_75t_L g648 ( 
.A(n_649),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_650),
.B(n_652),
.Y(n_649)
);

NOR2xp67_ASAP7_75t_L g655 ( 
.A(n_650),
.B(n_652),
.Y(n_655)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_655),
.Y(n_654)
);

INVxp67_ASAP7_75t_L g661 ( 
.A(n_656),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_657),
.B(n_659),
.Y(n_656)
);

INVx6_ASAP7_75t_L g657 ( 
.A(n_658),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_661),
.B(n_662),
.Y(n_660)
);


endmodule