module fake_jpeg_28767_n_37 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_37);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_37;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_36;
wire n_25;
wire n_17;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_15;

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_8),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx3_ASAP7_75t_SL g15 ( 
.A(n_3),
.Y(n_15)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx24_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_1),
.B(n_6),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_22),
.A2(n_9),
.B1(n_2),
.B2(n_5),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_25),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_31)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_28),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_15),
.A2(n_5),
.B1(n_12),
.B2(n_21),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g28 ( 
.A1(n_23),
.A2(n_14),
.B(n_18),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_13),
.B(n_24),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_19),
.A2(n_17),
.B1(n_18),
.B2(n_16),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_25),
.C(n_12),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_34),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_31),
.B(n_27),
.C(n_20),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_31),
.Y(n_36)
);

NOR2x1_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_20),
.Y(n_37)
);


endmodule