module real_jpeg_22746_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_346, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_346;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_1),
.A2(n_86),
.B(n_87),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_1),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_1),
.B(n_79),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_L g167 ( 
.A1(n_1),
.A2(n_35),
.B1(n_36),
.B2(n_89),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_1),
.B(n_30),
.C(n_31),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_1),
.B(n_69),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_1),
.A2(n_45),
.B1(n_188),
.B2(n_195),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx8_ASAP7_75t_SL g80 ( 
.A(n_4),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_5),
.A2(n_66),
.B1(n_68),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_5),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_5),
.A2(n_71),
.B1(n_92),
.B2(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_5),
.A2(n_35),
.B1(n_36),
.B2(n_71),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_71),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_51),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_6),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_6),
.A2(n_35),
.B1(n_36),
.B2(n_51),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_6),
.A2(n_51),
.B1(n_66),
.B2(n_68),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_6),
.A2(n_51),
.B1(n_86),
.B2(n_234),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_7),
.A2(n_35),
.B1(n_36),
.B2(n_58),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_7),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_7),
.A2(n_58),
.B1(n_66),
.B2(n_68),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_58),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_7),
.A2(n_58),
.B1(n_86),
.B2(n_92),
.Y(n_259)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_8),
.Y(n_65)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_9),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_10),
.A2(n_83),
.B1(n_92),
.B2(n_93),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_10),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_10),
.A2(n_66),
.B1(n_68),
.B2(n_93),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_10),
.A2(n_35),
.B1(n_36),
.B2(n_93),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_93),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_11),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_37),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_11),
.A2(n_37),
.B1(n_66),
.B2(n_68),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_L g297 ( 
.A1(n_11),
.A2(n_37),
.B1(n_101),
.B2(n_298),
.Y(n_297)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_13),
.A2(n_66),
.B1(n_68),
.B2(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_13),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_13),
.A2(n_35),
.B1(n_36),
.B2(n_73),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g178 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_73),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_13),
.A2(n_73),
.B1(n_101),
.B2(n_234),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_14),
.A2(n_35),
.B1(n_36),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_43),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_14),
.A2(n_43),
.B1(n_66),
.B2(n_68),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_14),
.A2(n_43),
.B1(n_83),
.B2(n_92),
.Y(n_284)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_15),
.Y(n_115)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_15),
.Y(n_189)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_15),
.Y(n_202)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_339),
.C(n_343),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_337),
.B(n_342),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_327),
.B(n_336),
.Y(n_18)
);

OAI321xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_292),
.A3(n_322),
.B1(n_325),
.B2(n_326),
.C(n_346),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_268),
.B(n_291),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_244),
.B(n_267),
.Y(n_21)
);

O2A1O1Ixp33_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_131),
.B(n_217),
.C(n_243),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_116),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_24),
.B(n_116),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_96),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_54),
.B1(n_94),
.B2(n_95),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_26),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_26),
.B(n_95),
.C(n_96),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_44),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_27),
.B(n_44),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_34),
.B(n_38),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_40),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_28),
.B(n_42),
.Y(n_59)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_28),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_28),
.B(n_160),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_28),
.B(n_89),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_28),
.A2(n_160),
.B(n_309),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_29),
.B(n_47),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_29),
.B(n_201),
.Y(n_200)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_L g40 ( 
.A1(n_31),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_40)
);

BUFx24_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_34),
.Y(n_226)
);

AO22x1_ASAP7_75t_L g69 ( 
.A1(n_35),
.A2(n_36),
.B1(n_64),
.B2(n_65),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_35),
.B(n_64),
.Y(n_140)
);

INVx2_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

OAI32xp33_ASAP7_75t_L g138 ( 
.A1(n_36),
.A2(n_65),
.A3(n_68),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_36),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_38),
.B(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_41),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_57),
.B(n_59),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_39),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_39),
.A2(n_148),
.B(n_159),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_39),
.A2(n_147),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_39),
.A2(n_146),
.B1(n_147),
.B2(n_168),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_39),
.A2(n_147),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_39),
.A2(n_59),
.B(n_227),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_39),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g44 ( 
.A1(n_45),
.A2(n_49),
.B(n_52),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_45),
.A2(n_52),
.B(n_142),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_45),
.A2(n_178),
.B(n_179),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_45),
.A2(n_185),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_45),
.A2(n_142),
.B(n_196),
.Y(n_252)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_46),
.A2(n_50),
.B1(n_112),
.B2(n_114),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_46),
.B(n_53),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_46),
.A2(n_184),
.B1(n_186),
.B2(n_187),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_47),
.B(n_53),
.Y(n_52)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g180 ( 
.A(n_48),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_60),
.C(n_75),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_55),
.A2(n_56),
.B1(n_60),
.B2(n_119),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_57),
.Y(n_160)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_70),
.B1(n_72),
.B2(n_74),
.Y(n_60)
);

OAI21xp33_ASAP7_75t_L g104 ( 
.A1(n_61),
.A2(n_72),
.B(n_105),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_61),
.A2(n_70),
.B1(n_74),
.B2(n_129),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_61),
.A2(n_237),
.B(n_238),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_61),
.A2(n_74),
.B1(n_262),
.B2(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_62),
.A2(n_69),
.B1(n_130),
.B2(n_139),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_62),
.B(n_239),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_62),
.A2(n_305),
.B(n_306),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g334 ( 
.A1(n_62),
.A2(n_69),
.B(n_106),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_69),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_65),
.B1(n_66),
.B2(n_68),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_66),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_66),
.A2(n_68),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g108 ( 
.A1(n_66),
.A2(n_81),
.B(n_88),
.C(n_109),
.Y(n_108)
);

HAxp5_ASAP7_75t_SL g139 ( 
.A(n_66),
.B(n_89),
.CON(n_139),
.SN(n_139)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

NAND3xp33_ASAP7_75t_L g109 ( 
.A(n_68),
.B(n_80),
.C(n_102),
.Y(n_109)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_69),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_69),
.B(n_239),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_74),
.A2(n_262),
.B(n_263),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_75),
.B(n_118),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_76),
.A2(n_78),
.B1(n_85),
.B2(n_90),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_77),
.A2(n_79),
.B1(n_91),
.B2(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_77),
.A2(n_79),
.B1(n_100),
.B2(n_233),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_77),
.A2(n_233),
.B(n_258),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_77),
.A2(n_282),
.B(n_283),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_77),
.B(n_300),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_77),
.A2(n_79),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_77),
.A2(n_283),
.B(n_316),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_77),
.A2(n_79),
.B(n_282),
.Y(n_343)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_82),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_78),
.B(n_259),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_78),
.B(n_284),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_78),
.A2(n_297),
.B(n_299),
.Y(n_296)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_L g82 ( 
.A1(n_80),
.A2(n_81),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

INVx8_ASAP7_75t_L g298 ( 
.A(n_83),
.Y(n_298)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_84),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_84),
.B(n_89),
.Y(n_88)
);

INVx8_ASAP7_75t_L g234 ( 
.A(n_86),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_89),
.B(n_202),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_107),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_103),
.B2(n_104),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_99),
.B(n_103),
.C(n_107),
.Y(n_241)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_105),
.B(n_263),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_106),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_110),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_108),
.A2(n_110),
.B1(n_111),
.B2(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g123 ( 
.A1(n_113),
.A2(n_124),
.B(n_125),
.Y(n_123)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_114),
.Y(n_124)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_115),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_120),
.C(n_122),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_117),
.B(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_120),
.B(n_122),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_126),
.C(n_128),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_123),
.A2(n_126),
.B1(n_127),
.B2(n_153),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_123),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_125),
.B(n_179),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_212),
.B(n_216),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_162),
.B(n_211),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_149),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_136),
.B(n_149),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_144),
.C(n_145),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_137),
.B(n_209),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_141),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_141),
.Y(n_156)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_143),
.B(n_180),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_144),
.B(n_145),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_151),
.B1(n_154),
.B2(n_155),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_150),
.B(n_157),
.C(n_161),
.Y(n_213)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_158),
.B2(n_161),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_156),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_159),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_206),
.B(n_210),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_181),
.B(n_205),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_171),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_165),
.B(n_171),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_169),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_177),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_173),
.B(n_176),
.C(n_177),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_175),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_178),
.Y(n_186)
);

AOI21xp33_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_191),
.B(n_204),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_190),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_190),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_192),
.A2(n_198),
.B(n_203),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_193),
.B(n_194),
.Y(n_203)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_207),
.B(n_208),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_213),
.B(n_214),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_219),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_241),
.B2(n_242),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_229),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_229),
.C(n_242),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_225),
.B2(n_228),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_223),
.B(n_228),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_225),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_240),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_232),
.B1(n_235),
.B2(n_236),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_232),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_232),
.B(n_235),
.C(n_240),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_238),
.Y(n_306)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_241),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_245),
.B(n_246),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_266),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_253),
.B1(n_264),
.B2(n_265),
.Y(n_247)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_248),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_265),
.C(n_266),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_251),
.B2(n_252),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_250),
.B(n_251),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_251),
.A2(n_252),
.B1(n_281),
.B2(n_285),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_251),
.A2(n_285),
.B(n_286),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_253),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_254),
.B(n_257),
.C(n_260),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_257),
.B1(n_260),
.B2(n_261),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g340 ( 
.A(n_258),
.Y(n_340)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_259),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_269),
.B(n_270),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_289),
.B2(n_290),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_279),
.B1(n_287),
.B2(n_288),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_273),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_273),
.B(n_288),
.C(n_290),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_276),
.B(n_278),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_276),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_277),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_294),
.C(n_310),
.Y(n_293)
);

FAx1_ASAP7_75t_SL g324 ( 
.A(n_278),
.B(n_294),
.CI(n_310),
.CON(n_324),
.SN(n_324)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_279),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_286),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_281),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_284),
.Y(n_300)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_289),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_311),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_293),
.B(n_311),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_301),
.B2(n_302),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_295),
.A2(n_296),
.B1(n_313),
.B2(n_320),
.Y(n_312)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_296),
.B(n_304),
.C(n_307),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_296),
.B(n_320),
.C(n_321),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_297),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_299),
.B(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_304),
.B1(n_307),
.B2(n_308),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_304),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_307),
.A2(n_308),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_308),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_308),
.B(n_314),
.C(n_318),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_321),
.Y(n_311)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_313),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_314),
.B(n_317),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_319),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_323),
.B(n_324),
.Y(n_325)
);

BUFx24_ASAP7_75t_SL g345 ( 
.A(n_324),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_328),
.B(n_329),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_335),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_331),
.A2(n_332),
.B1(n_333),
.B2(n_334),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_331),
.B(n_334),
.C(n_335),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_332),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_334),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_338),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_341),
.Y(n_338)
);

OR2x2_ASAP7_75t_L g342 ( 
.A(n_339),
.B(n_341),
.Y(n_342)
);


endmodule