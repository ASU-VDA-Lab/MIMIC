module fake_ariane_1487_n_1253 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1253);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1253;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_423;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_690;
wire n_416;
wire n_1109;
wire n_525;
wire n_187;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_232;
wire n_568;
wire n_1088;
wire n_766;
wire n_377;
wire n_520;
wire n_870;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1018;
wire n_259;
wire n_953;
wire n_1224;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_200;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_868;
wire n_884;
wire n_1034;
wire n_1085;
wire n_277;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_611;
wire n_365;
wire n_238;
wire n_1013;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_440;
wire n_273;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_491;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_461;
wire n_1121;
wire n_209;
wire n_490;
wire n_225;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_555;
wire n_804;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_513;
wire n_288;
wire n_1178;
wire n_1026;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_746;
wire n_292;
wire n_1079;
wire n_615;
wire n_1139;
wire n_517;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1101;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_299;
wire n_836;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_776;
wire n_424;
wire n_466;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_327;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_855;
wire n_808;
wire n_553;
wire n_814;
wire n_578;
wire n_405;
wire n_320;
wire n_1134;
wire n_647;
wire n_481;
wire n_600;
wire n_1053;
wire n_529;
wire n_502;
wire n_218;
wire n_247;
wire n_1105;
wire n_547;
wire n_604;
wire n_439;
wire n_677;
wire n_478;
wire n_703;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_545;
wire n_1015;
wire n_1162;
wire n_536;
wire n_325;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_233;
wire n_957;
wire n_388;
wire n_1242;
wire n_1218;
wire n_321;
wire n_221;
wire n_861;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_845;
wire n_888;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_769;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_999;
wire n_456;
wire n_852;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1243;
wire n_342;
wire n_358;
wire n_608;
wire n_1037;
wire n_317;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_687;
wire n_797;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_602;
wire n_592;
wire n_854;
wire n_393;
wire n_474;
wire n_805;
wire n_295;
wire n_190;
wire n_1072;
wire n_695;
wire n_180;
wire n_730;
wire n_386;
wire n_516;
wire n_1137;
wire n_640;
wire n_197;
wire n_463;
wire n_1118;
wire n_943;
wire n_678;
wire n_651;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_752;
wire n_985;
wire n_421;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_649;
wire n_374;
wire n_643;
wire n_226;
wire n_682;
wire n_819;
wire n_586;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_818;
wire n_779;
wire n_594;
wire n_1052;
wire n_272;
wire n_833;
wire n_879;
wire n_1117;
wire n_422;
wire n_597;
wire n_1047;
wire n_1050;
wire n_566;
wire n_1201;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_224;
wire n_894;
wire n_420;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1128;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1065;
wire n_453;
wire n_810;
wire n_181;
wire n_617;
wire n_543;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_743;
wire n_1194;
wire n_907;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_571;
wire n_414;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_613;
wire n_1022;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_820;
wire n_872;
wire n_254;
wire n_1157;
wire n_234;
wire n_848;
wire n_280;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_213;
wire n_1014;
wire n_724;
wire n_493;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1124;
wire n_932;
wire n_1183;
wire n_981;
wire n_1110;
wire n_243;
wire n_185;
wire n_1204;
wire n_994;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_353;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_828;
wire n_322;
wire n_558;
wire n_653;
wire n_783;
wire n_556;
wire n_1127;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1167;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_318;
wire n_244;
wire n_679;
wire n_220;
wire n_663;
wire n_443;
wire n_528;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_385;
wire n_917;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1064;
wire n_633;
wire n_900;
wire n_1093;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_835;
wire n_446;
wire n_1076;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_291;
wire n_822;
wire n_1094;
wire n_840;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_188;
wire n_323;
wire n_550;
wire n_997;
wire n_635;
wire n_694;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1236;
wire n_228;
wire n_671;
wire n_1148;
wire n_654;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_658;
wire n_630;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_196;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1229;
wire n_415;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_195;
wire n_938;
wire n_895;
wire n_304;
wire n_583;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_265;
wire n_208;
wire n_275;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_963;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1001;
wire n_1115;
wire n_1002;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_548;
wire n_289;
wire n_523;
wire n_457;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_484;
wire n_411;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_573;
wire n_796;
wire n_531;
wire n_675;

INVx1_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_60),
.Y(n_181)
);

BUFx10_ASAP7_75t_L g182 ( 
.A(n_33),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_80),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_125),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_179),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_150),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_133),
.Y(n_187)
);

INVxp33_ASAP7_75t_SL g188 ( 
.A(n_146),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_51),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_120),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_177),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_102),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_48),
.Y(n_193)
);

INVxp33_ASAP7_75t_SL g194 ( 
.A(n_61),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_43),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_178),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_68),
.Y(n_197)
);

BUFx10_ASAP7_75t_L g198 ( 
.A(n_83),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_153),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_99),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_97),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_67),
.Y(n_202)
);

BUFx5_ASAP7_75t_L g203 ( 
.A(n_53),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_111),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_40),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_43),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_168),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_154),
.Y(n_208)
);

BUFx10_ASAP7_75t_L g209 ( 
.A(n_18),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_58),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_138),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_38),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_157),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_107),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_122),
.Y(n_215)
);

BUFx10_ASAP7_75t_L g216 ( 
.A(n_73),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_115),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_72),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_79),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_63),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_9),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_170),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_40),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_7),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_117),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_20),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_32),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g228 ( 
.A(n_59),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_20),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_149),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_94),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_148),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_62),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_147),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_2),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_139),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_64),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_19),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_27),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_130),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_34),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_162),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_95),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_176),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g245 ( 
.A(n_134),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_39),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_143),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_16),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_169),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_132),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_23),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g252 ( 
.A(n_105),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_65),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_29),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_151),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_22),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_9),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_108),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_74),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_11),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_135),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_45),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_8),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_14),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_57),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_152),
.Y(n_266)
);

BUFx10_ASAP7_75t_L g267 ( 
.A(n_165),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_82),
.Y(n_268)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_124),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_140),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_69),
.Y(n_271)
);

BUFx8_ASAP7_75t_SL g272 ( 
.A(n_16),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_45),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_78),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_113),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_121),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_163),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_5),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_35),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_144),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_19),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_52),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_171),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_98),
.Y(n_284)
);

BUFx10_ASAP7_75t_L g285 ( 
.A(n_100),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_34),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_88),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_75),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_160),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_24),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_32),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_155),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_141),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_13),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_156),
.Y(n_295)
);

BUFx10_ASAP7_75t_L g296 ( 
.A(n_5),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_114),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_142),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_91),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_47),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_212),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_272),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_203),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_269),
.B(n_227),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_203),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_203),
.Y(n_306)
);

INVxp67_ASAP7_75t_SL g307 ( 
.A(n_189),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_293),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_203),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_198),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_203),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_203),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_195),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_203),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_196),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_198),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_198),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_216),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_203),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_216),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_180),
.B(n_0),
.Y(n_321)
);

NOR2xp67_ASAP7_75t_L g322 ( 
.A(n_235),
.B(n_0),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_199),
.Y(n_323)
);

INVxp67_ASAP7_75t_SL g324 ( 
.A(n_193),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_205),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_251),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_256),
.Y(n_327)
);

INVxp67_ASAP7_75t_SL g328 ( 
.A(n_260),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_222),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_264),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_278),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g332 ( 
.A(n_286),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_216),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_255),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_267),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_267),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_266),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_284),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_267),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_246),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_285),
.Y(n_341)
);

OR2x2_ASAP7_75t_L g342 ( 
.A(n_229),
.B(n_1),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_285),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_285),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_181),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_182),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_191),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_257),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_195),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_182),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_181),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_182),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_186),
.B(n_1),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_209),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_262),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_191),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g357 ( 
.A(n_209),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_209),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_183),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_183),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_296),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_294),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g363 ( 
.A(n_296),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_236),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_296),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_184),
.Y(n_366)
);

INVxp67_ASAP7_75t_SL g367 ( 
.A(n_236),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_184),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_192),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_291),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_204),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_185),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_208),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_185),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_294),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_187),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_211),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_187),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_215),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_300),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_190),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_300),
.Y(n_382)
);

OR2x2_ASAP7_75t_L g383 ( 
.A(n_281),
.B(n_2),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_237),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_247),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_250),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_253),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_190),
.Y(n_388)
);

BUFx6f_ASAP7_75t_SL g389 ( 
.A(n_228),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_240),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_276),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_303),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_347),
.B(n_277),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_305),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_342),
.A2(n_282),
.B1(n_254),
.B2(n_206),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_306),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_309),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_309),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_311),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_312),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_314),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_319),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_347),
.B(n_364),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_369),
.Y(n_404)
);

AND2x4_ASAP7_75t_L g405 ( 
.A(n_371),
.B(n_228),
.Y(n_405)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_375),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_356),
.Y(n_407)
);

INVx6_ASAP7_75t_L g408 ( 
.A(n_356),
.Y(n_408)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_356),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_356),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_373),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_356),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_377),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_379),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_364),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_384),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_385),
.Y(n_417)
);

BUFx3_ASAP7_75t_L g418 ( 
.A(n_386),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_387),
.B(n_240),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_391),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_353),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_325),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_307),
.B(n_245),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_326),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_367),
.B(n_292),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_327),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_324),
.B(n_292),
.Y(n_427)
);

INVx5_ASAP7_75t_L g428 ( 
.A(n_389),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_330),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_331),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_328),
.B(n_295),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_321),
.Y(n_432)
);

OAI21x1_ASAP7_75t_L g433 ( 
.A1(n_335),
.A2(n_242),
.B(n_233),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_313),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_332),
.B(n_295),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_336),
.B(n_245),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_339),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_346),
.B(n_297),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_352),
.B(n_233),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_322),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_389),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_354),
.B(n_297),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_389),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_358),
.Y(n_444)
);

AND2x4_ASAP7_75t_L g445 ( 
.A(n_361),
.B(n_242),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_365),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_383),
.Y(n_447)
);

BUFx8_ASAP7_75t_L g448 ( 
.A(n_357),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_382),
.Y(n_449)
);

INVx6_ASAP7_75t_L g450 ( 
.A(n_301),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_349),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_304),
.B(n_188),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_310),
.B(n_299),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_350),
.B(n_261),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_362),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_345),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_310),
.B(n_299),
.Y(n_457)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_345),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_316),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g460 ( 
.A(n_380),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_351),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_397),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_397),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_397),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_397),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_452),
.B(n_308),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_452),
.B(n_308),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_459),
.B(n_351),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_398),
.Y(n_469)
);

INVx4_ASAP7_75t_L g470 ( 
.A(n_428),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_398),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_398),
.Y(n_472)
);

NOR3xp33_ASAP7_75t_L g473 ( 
.A(n_395),
.B(n_360),
.C(n_359),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g474 ( 
.A(n_459),
.B(n_359),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_398),
.Y(n_475)
);

INVx5_ASAP7_75t_L g476 ( 
.A(n_428),
.Y(n_476)
);

OR2x2_ASAP7_75t_L g477 ( 
.A(n_447),
.B(n_363),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_400),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_407),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_461),
.B(n_360),
.Y(n_480)
);

INVxp67_ASAP7_75t_SL g481 ( 
.A(n_403),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_407),
.Y(n_482)
);

OR2x2_ASAP7_75t_L g483 ( 
.A(n_447),
.B(n_366),
.Y(n_483)
);

INVx6_ASAP7_75t_L g484 ( 
.A(n_408),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_407),
.Y(n_485)
);

NAND2x1p5_ASAP7_75t_L g486 ( 
.A(n_433),
.B(n_244),
.Y(n_486)
);

INVx4_ASAP7_75t_L g487 ( 
.A(n_428),
.Y(n_487)
);

AND2x4_ASAP7_75t_L g488 ( 
.A(n_437),
.B(n_316),
.Y(n_488)
);

NAND3xp33_ASAP7_75t_L g489 ( 
.A(n_395),
.B(n_368),
.C(n_366),
.Y(n_489)
);

AND2x6_ASAP7_75t_L g490 ( 
.A(n_441),
.B(n_261),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_459),
.B(n_368),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_400),
.Y(n_492)
);

NOR3xp33_ASAP7_75t_L g493 ( 
.A(n_434),
.B(n_374),
.C(n_372),
.Y(n_493)
);

BUFx2_ASAP7_75t_L g494 ( 
.A(n_434),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_400),
.Y(n_495)
);

INVx4_ASAP7_75t_L g496 ( 
.A(n_428),
.Y(n_496)
);

AND2x6_ASAP7_75t_L g497 ( 
.A(n_441),
.B(n_298),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_400),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_402),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_402),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_421),
.B(n_317),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_402),
.Y(n_502)
);

INVx5_ASAP7_75t_L g503 ( 
.A(n_428),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_407),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_461),
.B(n_372),
.Y(n_505)
);

INVxp67_ASAP7_75t_SL g506 ( 
.A(n_403),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_402),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_392),
.Y(n_508)
);

AND3x1_ASAP7_75t_L g509 ( 
.A(n_453),
.B(n_376),
.C(n_374),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_415),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_461),
.B(n_376),
.Y(n_511)
);

INVx5_ASAP7_75t_L g512 ( 
.A(n_428),
.Y(n_512)
);

OAI22xp33_ASAP7_75t_L g513 ( 
.A1(n_447),
.A2(n_333),
.B1(n_317),
.B2(n_318),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_415),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_461),
.B(n_378),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_459),
.B(n_378),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_457),
.B(n_381),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_459),
.B(n_381),
.Y(n_518)
);

NAND2xp33_ASAP7_75t_SL g519 ( 
.A(n_459),
.B(n_388),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_415),
.Y(n_520)
);

INVx4_ASAP7_75t_L g521 ( 
.A(n_428),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_457),
.B(n_388),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_415),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_L g524 ( 
.A1(n_447),
.A2(n_188),
.B1(n_194),
.B2(n_318),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_392),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_449),
.B(n_390),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_448),
.Y(n_527)
);

BUFx10_ASAP7_75t_L g528 ( 
.A(n_450),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_447),
.A2(n_194),
.B1(n_320),
.B2(n_333),
.Y(n_529)
);

NOR2x1p5_ASAP7_75t_L g530 ( 
.A(n_456),
.B(n_458),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_459),
.B(n_390),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_394),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_480),
.A2(n_458),
.B1(n_459),
.B2(n_456),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_532),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_505),
.B(n_458),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_511),
.B(n_458),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_515),
.B(n_458),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_494),
.B(n_453),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_494),
.B(n_453),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_526),
.B(n_421),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_501),
.B(n_449),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_517),
.B(n_449),
.Y(n_542)
);

NAND2xp33_ASAP7_75t_L g543 ( 
.A(n_530),
.B(n_441),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_532),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_522),
.B(n_449),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_508),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_481),
.B(n_444),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_L g548 ( 
.A1(n_508),
.A2(n_432),
.B1(n_423),
.B2(n_405),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_525),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_525),
.Y(n_550)
);

NAND2xp33_ASAP7_75t_L g551 ( 
.A(n_530),
.B(n_441),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_495),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_506),
.B(n_444),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_520),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_466),
.B(n_444),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_483),
.B(n_437),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_528),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_495),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_467),
.B(n_444),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_488),
.B(n_394),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_488),
.B(n_396),
.Y(n_561)
);

AND2x4_ASAP7_75t_L g562 ( 
.A(n_488),
.B(n_437),
.Y(n_562)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_524),
.A2(n_432),
.B1(n_423),
.B2(n_442),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_520),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_483),
.B(n_437),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_520),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_498),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_477),
.B(n_444),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_498),
.Y(n_569)
);

OR2x6_ASAP7_75t_L g570 ( 
.A(n_489),
.B(n_450),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_477),
.B(n_425),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_528),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_513),
.B(n_423),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_499),
.B(n_425),
.Y(n_574)
);

AO221x1_ASAP7_75t_L g575 ( 
.A1(n_509),
.A2(n_455),
.B1(n_451),
.B2(n_443),
.C(n_448),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_499),
.B(n_427),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_468),
.B(n_446),
.Y(n_577)
);

NAND2xp33_ASAP7_75t_L g578 ( 
.A(n_519),
.B(n_443),
.Y(n_578)
);

INVx4_ASAP7_75t_SL g579 ( 
.A(n_490),
.Y(n_579)
);

NAND2x1_ASAP7_75t_L g580 ( 
.A(n_479),
.B(n_408),
.Y(n_580)
);

AOI21xp5_ASAP7_75t_L g581 ( 
.A1(n_502),
.A2(n_399),
.B(n_396),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_528),
.B(n_399),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_502),
.B(n_427),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_473),
.A2(n_442),
.B1(n_436),
.B2(n_446),
.Y(n_584)
);

INVx8_ASAP7_75t_L g585 ( 
.A(n_527),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_507),
.Y(n_586)
);

AND2x4_ASAP7_75t_L g587 ( 
.A(n_527),
.B(n_442),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_507),
.Y(n_588)
);

A2O1A1Ixp33_ASAP7_75t_L g589 ( 
.A1(n_529),
.A2(n_416),
.B(n_424),
.C(n_422),
.Y(n_589)
);

NOR3xp33_ASAP7_75t_L g590 ( 
.A(n_493),
.B(n_460),
.C(n_406),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_474),
.B(n_401),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_463),
.B(n_431),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_463),
.B(n_431),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_465),
.B(n_435),
.Y(n_594)
);

INVx8_ASAP7_75t_L g595 ( 
.A(n_490),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_465),
.B(n_435),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_462),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g598 ( 
.A(n_491),
.B(n_438),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_462),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_472),
.B(n_418),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_L g601 ( 
.A1(n_478),
.A2(n_405),
.B1(n_416),
.B2(n_422),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_472),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_475),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_485),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_475),
.B(n_418),
.Y(n_605)
);

INVxp67_ASAP7_75t_L g606 ( 
.A(n_531),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_484),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_464),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_510),
.Y(n_609)
);

NOR2xp67_ASAP7_75t_L g610 ( 
.A(n_516),
.B(n_320),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_518),
.B(n_438),
.Y(n_611)
);

AOI22xp33_ASAP7_75t_L g612 ( 
.A1(n_478),
.A2(n_405),
.B1(n_416),
.B2(n_422),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_464),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_479),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_492),
.B(n_401),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g616 ( 
.A1(n_479),
.A2(n_419),
.B(n_433),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_510),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_469),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_492),
.B(n_428),
.Y(n_619)
);

AOI22xp33_ASAP7_75t_L g620 ( 
.A1(n_500),
.A2(n_405),
.B1(n_416),
.B2(n_422),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_500),
.B(n_418),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_514),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_485),
.B(n_436),
.Y(n_623)
);

NAND3xp33_ASAP7_75t_L g624 ( 
.A(n_514),
.B(n_455),
.C(n_451),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_469),
.B(n_418),
.Y(n_625)
);

AOI22xp5_ASAP7_75t_L g626 ( 
.A1(n_490),
.A2(n_436),
.B1(n_454),
.B2(n_450),
.Y(n_626)
);

OAI221xp5_ASAP7_75t_L g627 ( 
.A1(n_523),
.A2(n_419),
.B1(n_440),
.B2(n_430),
.C(n_426),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_471),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_523),
.Y(n_629)
);

BUFx6f_ASAP7_75t_SL g630 ( 
.A(n_490),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_597),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_571),
.B(n_436),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_545),
.A2(n_315),
.B1(n_329),
.B2(n_323),
.Y(n_633)
);

OAI22xp5_ASAP7_75t_L g634 ( 
.A1(n_545),
.A2(n_411),
.B1(n_413),
.B2(n_404),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_604),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_571),
.B(n_541),
.Y(n_636)
);

OAI21xp5_ASAP7_75t_L g637 ( 
.A1(n_616),
.A2(n_589),
.B(n_581),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_541),
.B(n_436),
.Y(n_638)
);

OAI21xp5_ASAP7_75t_L g639 ( 
.A1(n_589),
.A2(n_433),
.B(n_486),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_540),
.B(n_334),
.Y(n_640)
);

NOR2xp67_ASAP7_75t_L g641 ( 
.A(n_542),
.B(n_406),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_535),
.A2(n_487),
.B(n_470),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_536),
.A2(n_487),
.B(n_470),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_534),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_538),
.B(n_337),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_556),
.B(n_454),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_599),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_608),
.Y(n_648)
);

AND2x4_ASAP7_75t_L g649 ( 
.A(n_562),
.B(n_404),
.Y(n_649)
);

OR2x4_ASAP7_75t_L g650 ( 
.A(n_556),
.B(n_440),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_613),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_565),
.B(n_548),
.Y(n_652)
);

NOR2xp67_ASAP7_75t_L g653 ( 
.A(n_624),
.B(n_460),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_539),
.B(n_450),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_565),
.B(n_454),
.Y(n_655)
);

AND2x4_ASAP7_75t_L g656 ( 
.A(n_562),
.B(n_411),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g657 ( 
.A1(n_547),
.A2(n_487),
.B(n_470),
.Y(n_657)
);

HB1xp67_ASAP7_75t_L g658 ( 
.A(n_587),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_548),
.B(n_454),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_544),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_553),
.A2(n_521),
.B(n_496),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_587),
.B(n_450),
.Y(n_662)
);

OAI21xp5_ASAP7_75t_L g663 ( 
.A1(n_592),
.A2(n_486),
.B(n_471),
.Y(n_663)
);

AOI21xp5_ASAP7_75t_L g664 ( 
.A1(n_537),
.A2(n_521),
.B(n_496),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_604),
.Y(n_665)
);

AOI21x1_ASAP7_75t_L g666 ( 
.A1(n_619),
.A2(n_393),
.B(n_410),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_563),
.B(n_454),
.Y(n_667)
);

A2O1A1Ixp33_ASAP7_75t_L g668 ( 
.A1(n_598),
.A2(n_405),
.B(n_504),
.C(n_482),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_606),
.B(n_338),
.Y(n_669)
);

A2O1A1Ixp33_ASAP7_75t_L g670 ( 
.A1(n_598),
.A2(n_504),
.B(n_482),
.C(n_417),
.Y(n_670)
);

O2A1O1Ixp33_ASAP7_75t_L g671 ( 
.A1(n_573),
.A2(n_426),
.B(n_430),
.C(n_429),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g672 ( 
.A1(n_537),
.A2(n_521),
.B(n_496),
.Y(n_672)
);

O2A1O1Ixp33_ASAP7_75t_L g673 ( 
.A1(n_568),
.A2(n_429),
.B(n_413),
.C(n_420),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_557),
.B(n_485),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_555),
.B(n_341),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g676 ( 
.A1(n_574),
.A2(n_504),
.B(n_482),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_559),
.B(n_341),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_611),
.B(n_343),
.Y(n_678)
);

AOI22xp5_ASAP7_75t_L g679 ( 
.A1(n_560),
.A2(n_450),
.B1(n_343),
.B2(n_344),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_593),
.A2(n_503),
.B(n_476),
.Y(n_680)
);

O2A1O1Ixp33_ASAP7_75t_L g681 ( 
.A1(n_560),
.A2(n_417),
.B(n_414),
.C(n_420),
.Y(n_681)
);

A2O1A1Ixp33_ASAP7_75t_L g682 ( 
.A1(n_611),
.A2(n_414),
.B(n_424),
.C(n_445),
.Y(n_682)
);

NOR3xp33_ASAP7_75t_L g683 ( 
.A(n_561),
.B(n_223),
.C(n_221),
.Y(n_683)
);

NOR2xp67_ASAP7_75t_L g684 ( 
.A(n_584),
.B(n_344),
.Y(n_684)
);

AOI21xp5_ASAP7_75t_L g685 ( 
.A1(n_594),
.A2(n_596),
.B(n_583),
.Y(n_685)
);

INVx4_ASAP7_75t_L g686 ( 
.A(n_585),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_576),
.B(n_439),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_557),
.B(n_485),
.Y(n_688)
);

AND2x4_ASAP7_75t_SL g689 ( 
.A(n_570),
.B(n_340),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_585),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_561),
.B(n_348),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_585),
.B(n_355),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_557),
.B(n_485),
.Y(n_693)
);

OR2x6_ASAP7_75t_L g694 ( 
.A(n_595),
.B(n_448),
.Y(n_694)
);

OR2x6_ASAP7_75t_L g695 ( 
.A(n_595),
.B(n_448),
.Y(n_695)
);

O2A1O1Ixp5_ASAP7_75t_L g696 ( 
.A1(n_591),
.A2(n_424),
.B(n_409),
.C(n_439),
.Y(n_696)
);

O2A1O1Ixp33_ASAP7_75t_L g697 ( 
.A1(n_623),
.A2(n_627),
.B(n_558),
.C(n_567),
.Y(n_697)
);

AOI21xp5_ASAP7_75t_L g698 ( 
.A1(n_600),
.A2(n_503),
.B(n_476),
.Y(n_698)
);

HB1xp67_ASAP7_75t_L g699 ( 
.A(n_570),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_575),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_557),
.B(n_533),
.Y(n_701)
);

AOI21xp5_ASAP7_75t_L g702 ( 
.A1(n_605),
.A2(n_503),
.B(n_476),
.Y(n_702)
);

O2A1O1Ixp33_ASAP7_75t_L g703 ( 
.A1(n_623),
.A2(n_424),
.B(n_280),
.C(n_393),
.Y(n_703)
);

AOI21xp5_ASAP7_75t_L g704 ( 
.A1(n_543),
.A2(n_551),
.B(n_572),
.Y(n_704)
);

AOI21xp5_ASAP7_75t_L g705 ( 
.A1(n_591),
.A2(n_615),
.B(n_621),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_577),
.B(n_439),
.Y(n_706)
);

OAI22xp5_ASAP7_75t_L g707 ( 
.A1(n_601),
.A2(n_486),
.B1(n_224),
.B2(n_226),
.Y(n_707)
);

OAI22xp5_ASAP7_75t_L g708 ( 
.A1(n_577),
.A2(n_263),
.B1(n_238),
.B2(n_279),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_546),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_570),
.B(n_370),
.Y(n_710)
);

AOI21xp5_ASAP7_75t_L g711 ( 
.A1(n_615),
.A2(n_625),
.B(n_564),
.Y(n_711)
);

AOI21xp5_ASAP7_75t_L g712 ( 
.A1(n_554),
.A2(n_503),
.B(n_476),
.Y(n_712)
);

OAI22xp5_ASAP7_75t_L g713 ( 
.A1(n_601),
.A2(n_290),
.B1(n_239),
.B2(n_241),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_595),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_612),
.B(n_439),
.Y(n_715)
);

AOI21xp5_ASAP7_75t_L g716 ( 
.A1(n_566),
.A2(n_503),
.B(n_476),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_549),
.Y(n_717)
);

OAI22x1_ASAP7_75t_L g718 ( 
.A1(n_626),
.A2(n_445),
.B1(n_439),
.B2(n_448),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_618),
.Y(n_719)
);

AOI21xp5_ASAP7_75t_L g720 ( 
.A1(n_582),
.A2(n_512),
.B(n_412),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_612),
.B(n_445),
.Y(n_721)
);

OAI321xp33_ASAP7_75t_L g722 ( 
.A1(n_620),
.A2(n_410),
.A3(n_412),
.B1(n_298),
.B2(n_273),
.C(n_248),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_590),
.B(n_445),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_620),
.B(n_445),
.Y(n_724)
);

NOR2xp67_ASAP7_75t_L g725 ( 
.A(n_610),
.B(n_409),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_614),
.B(n_409),
.Y(n_726)
);

AOI22xp5_ASAP7_75t_L g727 ( 
.A1(n_550),
.A2(n_497),
.B1(n_490),
.B2(n_484),
.Y(n_727)
);

BUFx6f_ASAP7_75t_L g728 ( 
.A(n_580),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_636),
.B(n_552),
.Y(n_729)
);

O2A1O1Ixp33_ASAP7_75t_L g730 ( 
.A1(n_678),
.A2(n_588),
.B(n_586),
.C(n_569),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_692),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_640),
.B(n_602),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_691),
.B(n_614),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_644),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_SL g735 ( 
.A(n_652),
.B(n_603),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_632),
.B(n_609),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_631),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_649),
.B(n_656),
.Y(n_738)
);

A2O1A1Ixp33_ASAP7_75t_L g739 ( 
.A1(n_685),
.A2(n_629),
.B(n_622),
.C(n_617),
.Y(n_739)
);

HB1xp67_ASAP7_75t_L g740 ( 
.A(n_658),
.Y(n_740)
);

BUFx2_ASAP7_75t_L g741 ( 
.A(n_633),
.Y(n_741)
);

OAI22xp5_ASAP7_75t_L g742 ( 
.A1(n_646),
.A2(n_655),
.B1(n_638),
.B2(n_650),
.Y(n_742)
);

O2A1O1Ixp33_ASAP7_75t_L g743 ( 
.A1(n_675),
.A2(n_578),
.B(n_582),
.C(n_607),
.Y(n_743)
);

NOR3xp33_ASAP7_75t_SL g744 ( 
.A(n_645),
.B(n_200),
.C(n_197),
.Y(n_744)
);

INVx4_ASAP7_75t_L g745 ( 
.A(n_686),
.Y(n_745)
);

AOI21xp5_ASAP7_75t_L g746 ( 
.A1(n_642),
.A2(n_619),
.B(n_512),
.Y(n_746)
);

NAND2xp33_ASAP7_75t_SL g747 ( 
.A(n_686),
.B(n_630),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_724),
.A2(n_628),
.B1(n_630),
.B2(n_497),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_L g749 ( 
.A1(n_667),
.A2(n_497),
.B1(n_490),
.B2(n_409),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_660),
.Y(n_750)
);

INVx4_ASAP7_75t_L g751 ( 
.A(n_714),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_689),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_SL g753 ( 
.A1(n_710),
.A2(n_302),
.B1(n_287),
.B2(n_252),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_677),
.B(n_484),
.Y(n_754)
);

AOI21xp5_ASAP7_75t_L g755 ( 
.A1(n_643),
.A2(n_512),
.B(n_412),
.Y(n_755)
);

O2A1O1Ixp33_ASAP7_75t_L g756 ( 
.A1(n_708),
.A2(n_409),
.B(n_410),
.C(n_6),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_649),
.B(n_497),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_656),
.B(n_497),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_669),
.Y(n_759)
);

O2A1O1Ixp33_ASAP7_75t_L g760 ( 
.A1(n_634),
.A2(n_3),
.B(n_4),
.C(n_6),
.Y(n_760)
);

AOI21xp5_ASAP7_75t_L g761 ( 
.A1(n_701),
.A2(n_512),
.B(n_202),
.Y(n_761)
);

O2A1O1Ixp33_ASAP7_75t_L g762 ( 
.A1(n_634),
.A2(n_3),
.B(n_4),
.C(n_7),
.Y(n_762)
);

AND2x4_ASAP7_75t_L g763 ( 
.A(n_662),
.B(n_579),
.Y(n_763)
);

A2O1A1Ixp33_ASAP7_75t_L g764 ( 
.A1(n_697),
.A2(n_243),
.B(n_207),
.C(n_289),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_676),
.A2(n_512),
.B(n_258),
.Y(n_765)
);

NOR2xp67_ASAP7_75t_L g766 ( 
.A(n_690),
.B(n_201),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_657),
.A2(n_249),
.B(n_213),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_709),
.Y(n_768)
);

NOR2xp67_ASAP7_75t_L g769 ( 
.A(n_679),
.B(n_210),
.Y(n_769)
);

INVxp67_ASAP7_75t_L g770 ( 
.A(n_653),
.Y(n_770)
);

BUFx3_ASAP7_75t_L g771 ( 
.A(n_635),
.Y(n_771)
);

A2O1A1Ixp33_ASAP7_75t_L g772 ( 
.A1(n_684),
.A2(n_265),
.B(n_217),
.C(n_218),
.Y(n_772)
);

O2A1O1Ixp33_ASAP7_75t_L g773 ( 
.A1(n_671),
.A2(n_8),
.B(n_10),
.C(n_11),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_650),
.B(n_484),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_L g775 ( 
.A1(n_687),
.A2(n_408),
.B1(n_259),
.B2(n_288),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_661),
.A2(n_268),
.B(n_219),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_647),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_R g778 ( 
.A(n_714),
.B(n_497),
.Y(n_778)
);

AOI21xp5_ASAP7_75t_L g779 ( 
.A1(n_711),
.A2(n_234),
.B(n_220),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_705),
.A2(n_270),
.B(n_225),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_714),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_648),
.Y(n_782)
);

OAI22xp5_ASAP7_75t_L g783 ( 
.A1(n_706),
.A2(n_408),
.B1(n_271),
.B2(n_283),
.Y(n_783)
);

OR2x2_ASAP7_75t_L g784 ( 
.A(n_654),
.B(n_10),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_651),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_659),
.B(n_579),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_707),
.A2(n_579),
.B1(n_408),
.B2(n_275),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_635),
.B(n_214),
.Y(n_788)
);

INVx3_ASAP7_75t_L g789 ( 
.A(n_635),
.Y(n_789)
);

INVx1_ASAP7_75t_SL g790 ( 
.A(n_699),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_723),
.B(n_408),
.Y(n_791)
);

BUFx2_ASAP7_75t_L g792 ( 
.A(n_665),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_704),
.A2(n_274),
.B(n_232),
.Y(n_793)
);

AOI22xp5_ASAP7_75t_L g794 ( 
.A1(n_641),
.A2(n_683),
.B1(n_713),
.B2(n_707),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_713),
.A2(n_230),
.B1(n_231),
.B2(n_14),
.Y(n_795)
);

AOI21xp5_ASAP7_75t_L g796 ( 
.A1(n_729),
.A2(n_637),
.B(n_663),
.Y(n_796)
);

AO21x1_ASAP7_75t_L g797 ( 
.A1(n_742),
.A2(n_663),
.B(n_673),
.Y(n_797)
);

OAI22xp5_ASAP7_75t_L g798 ( 
.A1(n_794),
.A2(n_721),
.B1(n_715),
.B2(n_682),
.Y(n_798)
);

A2O1A1Ixp33_ASAP7_75t_L g799 ( 
.A1(n_733),
.A2(n_681),
.B(n_722),
.C(n_703),
.Y(n_799)
);

OR2x2_ASAP7_75t_L g800 ( 
.A(n_741),
.B(n_717),
.Y(n_800)
);

A2O1A1Ixp33_ASAP7_75t_L g801 ( 
.A1(n_733),
.A2(n_722),
.B(n_700),
.C(n_725),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_759),
.B(n_694),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_736),
.A2(n_637),
.B(n_668),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_735),
.B(n_665),
.Y(n_804)
);

OAI21xp5_ASAP7_75t_L g805 ( 
.A1(n_735),
.A2(n_670),
.B(n_696),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_739),
.A2(n_639),
.B(n_672),
.Y(n_806)
);

OAI21xp5_ASAP7_75t_L g807 ( 
.A1(n_739),
.A2(n_639),
.B(n_666),
.Y(n_807)
);

OAI21x1_ASAP7_75t_L g808 ( 
.A1(n_755),
.A2(n_746),
.B(n_720),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_737),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_777),
.Y(n_810)
);

BUFx12f_ASAP7_75t_L g811 ( 
.A(n_752),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_781),
.Y(n_812)
);

OAI21x1_ASAP7_75t_L g813 ( 
.A1(n_786),
.A2(n_664),
.B(n_698),
.Y(n_813)
);

NAND3xp33_ASAP7_75t_L g814 ( 
.A(n_795),
.B(n_726),
.C(n_665),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_734),
.Y(n_815)
);

OAI22xp5_ASAP7_75t_L g816 ( 
.A1(n_732),
.A2(n_694),
.B1(n_695),
.B2(n_727),
.Y(n_816)
);

O2A1O1Ixp5_ASAP7_75t_L g817 ( 
.A1(n_764),
.A2(n_674),
.B(n_688),
.C(n_693),
.Y(n_817)
);

BUFx12f_ASAP7_75t_L g818 ( 
.A(n_731),
.Y(n_818)
);

OAI22xp5_ASAP7_75t_L g819 ( 
.A1(n_787),
.A2(n_784),
.B1(n_764),
.B2(n_750),
.Y(n_819)
);

BUFx2_ASAP7_75t_L g820 ( 
.A(n_792),
.Y(n_820)
);

HB1xp67_ASAP7_75t_L g821 ( 
.A(n_740),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_738),
.Y(n_822)
);

OAI21xp5_ASAP7_75t_L g823 ( 
.A1(n_730),
.A2(n_680),
.B(n_702),
.Y(n_823)
);

OAI21xp5_ASAP7_75t_L g824 ( 
.A1(n_743),
.A2(n_716),
.B(n_712),
.Y(n_824)
);

A2O1A1Ixp33_ASAP7_75t_L g825 ( 
.A1(n_756),
.A2(n_773),
.B(n_787),
.C(n_760),
.Y(n_825)
);

AO31x2_ASAP7_75t_L g826 ( 
.A1(n_768),
.A2(n_718),
.A3(n_719),
.B(n_728),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_774),
.B(n_728),
.Y(n_827)
);

A2O1A1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_762),
.A2(n_728),
.B(n_695),
.C(n_694),
.Y(n_828)
);

INVxp67_ASAP7_75t_SL g829 ( 
.A(n_771),
.Y(n_829)
);

OAI21x1_ASAP7_75t_L g830 ( 
.A1(n_765),
.A2(n_695),
.B(n_89),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_782),
.Y(n_831)
);

OAI21xp5_ASAP7_75t_L g832 ( 
.A1(n_754),
.A2(n_12),
.B(n_13),
.Y(n_832)
);

AO31x2_ASAP7_75t_L g833 ( 
.A1(n_754),
.A2(n_90),
.A3(n_175),
.B(n_174),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_783),
.A2(n_86),
.B(n_173),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_SL g835 ( 
.A(n_753),
.B(n_56),
.Y(n_835)
);

AO31x2_ASAP7_75t_L g836 ( 
.A1(n_785),
.A2(n_87),
.A3(n_172),
.B(n_166),
.Y(n_836)
);

NAND2x1p5_ASAP7_75t_L g837 ( 
.A(n_771),
.B(n_66),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_769),
.B(n_781),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_780),
.A2(n_85),
.B(n_164),
.Y(n_839)
);

AO31x2_ASAP7_75t_L g840 ( 
.A1(n_775),
.A2(n_84),
.A3(n_161),
.B(n_159),
.Y(n_840)
);

INVxp67_ASAP7_75t_SL g841 ( 
.A(n_789),
.Y(n_841)
);

BUFx8_ASAP7_75t_L g842 ( 
.A(n_781),
.Y(n_842)
);

AOI21xp33_ASAP7_75t_L g843 ( 
.A1(n_791),
.A2(n_748),
.B(n_790),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_744),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_789),
.Y(n_845)
);

OAI21x1_ASAP7_75t_L g846 ( 
.A1(n_761),
.A2(n_77),
.B(n_158),
.Y(n_846)
);

INVx8_ASAP7_75t_L g847 ( 
.A(n_763),
.Y(n_847)
);

A2O1A1Ixp33_ASAP7_75t_L g848 ( 
.A1(n_774),
.A2(n_12),
.B(n_15),
.C(n_17),
.Y(n_848)
);

NOR2xp67_ASAP7_75t_L g849 ( 
.A(n_751),
.B(n_70),
.Y(n_849)
);

NAND2x1p5_ASAP7_75t_L g850 ( 
.A(n_763),
.B(n_71),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_757),
.Y(n_851)
);

AOI221x1_ASAP7_75t_L g852 ( 
.A1(n_779),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.C(n_21),
.Y(n_852)
);

AOI22xp33_ASAP7_75t_L g853 ( 
.A1(n_835),
.A2(n_770),
.B1(n_748),
.B2(n_788),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_815),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_L g855 ( 
.A1(n_798),
.A2(n_788),
.B1(n_758),
.B2(n_749),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_831),
.Y(n_856)
);

INVx6_ASAP7_75t_L g857 ( 
.A(n_842),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_L g858 ( 
.A1(n_798),
.A2(n_749),
.B1(n_766),
.B2(n_747),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_L g859 ( 
.A1(n_819),
.A2(n_778),
.B1(n_781),
.B2(n_751),
.Y(n_859)
);

AOI22xp33_ASAP7_75t_L g860 ( 
.A1(n_819),
.A2(n_778),
.B1(n_776),
.B2(n_767),
.Y(n_860)
);

INVx1_ASAP7_75t_SL g861 ( 
.A(n_818),
.Y(n_861)
);

AOI22xp33_ASAP7_75t_L g862 ( 
.A1(n_800),
.A2(n_793),
.B1(n_745),
.B2(n_772),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_832),
.A2(n_843),
.B1(n_797),
.B2(n_822),
.Y(n_863)
);

AOI22xp33_ASAP7_75t_L g864 ( 
.A1(n_832),
.A2(n_745),
.B1(n_22),
.B2(n_23),
.Y(n_864)
);

AOI22xp33_ASAP7_75t_L g865 ( 
.A1(n_843),
.A2(n_21),
.B1(n_24),
.B2(n_25),
.Y(n_865)
);

AOI22xp33_ASAP7_75t_L g866 ( 
.A1(n_809),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_866)
);

AOI22xp33_ASAP7_75t_L g867 ( 
.A1(n_816),
.A2(n_26),
.B1(n_28),
.B2(n_29),
.Y(n_867)
);

AOI22xp33_ASAP7_75t_SL g868 ( 
.A1(n_816),
.A2(n_28),
.B1(n_30),
.B2(n_31),
.Y(n_868)
);

AOI22xp33_ASAP7_75t_L g869 ( 
.A1(n_851),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_869)
);

BUFx10_ASAP7_75t_L g870 ( 
.A(n_844),
.Y(n_870)
);

AOI22xp33_ASAP7_75t_L g871 ( 
.A1(n_810),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_811),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_827),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_873)
);

BUFx2_ASAP7_75t_L g874 ( 
.A(n_820),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_821),
.B(n_39),
.Y(n_875)
);

AOI22xp33_ASAP7_75t_SL g876 ( 
.A1(n_802),
.A2(n_41),
.B1(n_42),
.B2(n_44),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_829),
.B(n_41),
.Y(n_877)
);

CKINVDCx20_ASAP7_75t_R g878 ( 
.A(n_842),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_847),
.Y(n_879)
);

INVx6_ASAP7_75t_L g880 ( 
.A(n_847),
.Y(n_880)
);

INVx3_ASAP7_75t_SL g881 ( 
.A(n_847),
.Y(n_881)
);

INVx3_ASAP7_75t_SL g882 ( 
.A(n_812),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_804),
.Y(n_883)
);

INVx3_ASAP7_75t_SL g884 ( 
.A(n_812),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_804),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_841),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_826),
.Y(n_887)
);

HB1xp67_ASAP7_75t_L g888 ( 
.A(n_812),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_826),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_826),
.Y(n_890)
);

CKINVDCx11_ASAP7_75t_R g891 ( 
.A(n_838),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_845),
.B(n_796),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_833),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_SL g894 ( 
.A1(n_850),
.A2(n_42),
.B1(n_44),
.B2(n_46),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_833),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_833),
.Y(n_896)
);

AOI22xp33_ASAP7_75t_SL g897 ( 
.A1(n_850),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_897)
);

AOI22xp33_ASAP7_75t_L g898 ( 
.A1(n_803),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_898)
);

BUFx8_ASAP7_75t_L g899 ( 
.A(n_828),
.Y(n_899)
);

AOI22xp5_ASAP7_75t_L g900 ( 
.A1(n_825),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_900)
);

BUFx12f_ASAP7_75t_L g901 ( 
.A(n_837),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_836),
.Y(n_902)
);

OAI22xp5_ASAP7_75t_L g903 ( 
.A1(n_799),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_903)
);

INVxp67_ASAP7_75t_L g904 ( 
.A(n_814),
.Y(n_904)
);

AOI22xp5_ASAP7_75t_L g905 ( 
.A1(n_801),
.A2(n_848),
.B1(n_849),
.B2(n_837),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_836),
.Y(n_906)
);

NAND2xp33_ASAP7_75t_SL g907 ( 
.A(n_805),
.B(n_54),
.Y(n_907)
);

AOI22xp33_ASAP7_75t_SL g908 ( 
.A1(n_807),
.A2(n_55),
.B1(n_76),
.B2(n_81),
.Y(n_908)
);

OAI22xp33_ASAP7_75t_R g909 ( 
.A1(n_852),
.A2(n_92),
.B1(n_93),
.B2(n_96),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_805),
.Y(n_910)
);

OR2x2_ASAP7_75t_L g911 ( 
.A(n_883),
.B(n_807),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_885),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_910),
.B(n_806),
.Y(n_913)
);

INVx3_ASAP7_75t_L g914 ( 
.A(n_892),
.Y(n_914)
);

BUFx2_ASAP7_75t_L g915 ( 
.A(n_893),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_902),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_854),
.B(n_806),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_895),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_887),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_906),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_889),
.B(n_840),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_890),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_904),
.B(n_840),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_896),
.Y(n_924)
);

AND2x4_ASAP7_75t_L g925 ( 
.A(n_886),
.B(n_813),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_856),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_901),
.Y(n_927)
);

AOI21x1_ASAP7_75t_L g928 ( 
.A1(n_888),
.A2(n_808),
.B(n_823),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_863),
.Y(n_929)
);

OR2x6_ASAP7_75t_L g930 ( 
.A(n_880),
.B(n_823),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_863),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_882),
.Y(n_932)
);

HB1xp67_ASAP7_75t_L g933 ( 
.A(n_874),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_882),
.Y(n_934)
);

HB1xp67_ASAP7_75t_L g935 ( 
.A(n_884),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_884),
.Y(n_936)
);

INVx3_ASAP7_75t_L g937 ( 
.A(n_857),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_907),
.Y(n_938)
);

AOI22xp33_ASAP7_75t_SL g939 ( 
.A1(n_899),
.A2(n_903),
.B1(n_909),
.B2(n_877),
.Y(n_939)
);

OR2x6_ASAP7_75t_L g940 ( 
.A(n_880),
.B(n_830),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_905),
.Y(n_941)
);

CKINVDCx20_ASAP7_75t_R g942 ( 
.A(n_878),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_899),
.Y(n_943)
);

OAI21x1_ASAP7_75t_L g944 ( 
.A1(n_860),
.A2(n_824),
.B(n_817),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_859),
.Y(n_945)
);

BUFx2_ASAP7_75t_SL g946 ( 
.A(n_879),
.Y(n_946)
);

HB1xp67_ASAP7_75t_L g947 ( 
.A(n_875),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_879),
.Y(n_948)
);

INVx3_ASAP7_75t_L g949 ( 
.A(n_925),
.Y(n_949)
);

AND2x4_ASAP7_75t_L g950 ( 
.A(n_925),
.B(n_859),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_917),
.B(n_913),
.Y(n_951)
);

OAI22xp5_ASAP7_75t_L g952 ( 
.A1(n_939),
.A2(n_864),
.B1(n_867),
.B2(n_898),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_916),
.Y(n_953)
);

BUFx6f_ASAP7_75t_L g954 ( 
.A(n_944),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_917),
.B(n_913),
.Y(n_955)
);

OAI211xp5_ASAP7_75t_L g956 ( 
.A1(n_939),
.A2(n_864),
.B(n_900),
.C(n_898),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_917),
.B(n_867),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_942),
.Y(n_958)
);

OR2x2_ASAP7_75t_L g959 ( 
.A(n_914),
.B(n_840),
.Y(n_959)
);

AND2x4_ASAP7_75t_SL g960 ( 
.A(n_930),
.B(n_936),
.Y(n_960)
);

BUFx12f_ASAP7_75t_L g961 ( 
.A(n_927),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_913),
.B(n_855),
.Y(n_962)
);

O2A1O1Ixp33_ASAP7_75t_SL g963 ( 
.A1(n_942),
.A2(n_861),
.B(n_873),
.C(n_870),
.Y(n_963)
);

AND4x1_ASAP7_75t_L g964 ( 
.A(n_938),
.B(n_871),
.C(n_869),
.D(n_858),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_914),
.B(n_855),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_926),
.Y(n_966)
);

OAI211xp5_ASAP7_75t_L g967 ( 
.A1(n_938),
.A2(n_876),
.B(n_897),
.C(n_894),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_914),
.B(n_908),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_926),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_914),
.B(n_868),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_914),
.B(n_871),
.Y(n_971)
);

BUFx3_ASAP7_75t_L g972 ( 
.A(n_936),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_925),
.B(n_869),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_925),
.B(n_911),
.Y(n_974)
);

OAI21xp5_ASAP7_75t_L g975 ( 
.A1(n_941),
.A2(n_865),
.B(n_858),
.Y(n_975)
);

INVx3_ASAP7_75t_L g976 ( 
.A(n_925),
.Y(n_976)
);

AOI22xp5_ASAP7_75t_L g977 ( 
.A1(n_941),
.A2(n_929),
.B1(n_931),
.B2(n_945),
.Y(n_977)
);

AND2x2_ASAP7_75t_L g978 ( 
.A(n_925),
.B(n_860),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_947),
.B(n_870),
.Y(n_979)
);

INVx2_ASAP7_75t_SL g980 ( 
.A(n_932),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_926),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_911),
.B(n_824),
.Y(n_982)
);

INVxp67_ASAP7_75t_L g983 ( 
.A(n_933),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_929),
.B(n_853),
.Y(n_984)
);

OR2x6_ASAP7_75t_L g985 ( 
.A(n_930),
.B(n_857),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_931),
.B(n_853),
.Y(n_986)
);

OA21x2_ASAP7_75t_L g987 ( 
.A1(n_944),
.A2(n_923),
.B(n_918),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_926),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_L g989 ( 
.A1(n_938),
.A2(n_866),
.B1(n_862),
.B2(n_857),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_951),
.B(n_911),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_966),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_954),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_953),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_951),
.B(n_944),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_951),
.B(n_955),
.Y(n_995)
);

AND2x2_ASAP7_75t_L g996 ( 
.A(n_955),
.B(n_930),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_982),
.B(n_933),
.Y(n_997)
);

AOI22xp33_ASAP7_75t_L g998 ( 
.A1(n_952),
.A2(n_923),
.B1(n_945),
.B2(n_947),
.Y(n_998)
);

OR2x2_ASAP7_75t_L g999 ( 
.A(n_955),
.B(n_915),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_953),
.Y(n_1000)
);

HB1xp67_ASAP7_75t_L g1001 ( 
.A(n_983),
.Y(n_1001)
);

INVx3_ASAP7_75t_L g1002 ( 
.A(n_949),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_966),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_974),
.B(n_930),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_974),
.B(n_930),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_982),
.B(n_915),
.Y(n_1006)
);

BUFx2_ASAP7_75t_L g1007 ( 
.A(n_976),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_974),
.B(n_930),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_978),
.B(n_930),
.Y(n_1009)
);

HB1xp67_ASAP7_75t_L g1010 ( 
.A(n_983),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_969),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_949),
.B(n_928),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_953),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_969),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_981),
.Y(n_1015)
);

OAI221xp5_ASAP7_75t_L g1016 ( 
.A1(n_998),
.A2(n_952),
.B1(n_956),
.B2(n_964),
.C(n_967),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_1006),
.B(n_982),
.Y(n_1017)
);

BUFx2_ASAP7_75t_L g1018 ( 
.A(n_1001),
.Y(n_1018)
);

AND2x4_ASAP7_75t_L g1019 ( 
.A(n_996),
.B(n_949),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_997),
.B(n_958),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_998),
.A2(n_956),
.B(n_975),
.Y(n_1021)
);

AOI31xp33_ASAP7_75t_L g1022 ( 
.A1(n_1006),
.A2(n_963),
.A3(n_968),
.B(n_979),
.Y(n_1022)
);

OR2x2_ASAP7_75t_L g1023 ( 
.A(n_999),
.B(n_987),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_995),
.B(n_978),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_1014),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_1014),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_995),
.B(n_978),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_993),
.Y(n_1028)
);

OR2x6_ASAP7_75t_L g1029 ( 
.A(n_992),
.B(n_985),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_995),
.B(n_949),
.Y(n_1030)
);

AND2x4_ASAP7_75t_L g1031 ( 
.A(n_996),
.B(n_949),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_991),
.Y(n_1032)
);

BUFx2_ASAP7_75t_SL g1033 ( 
.A(n_992),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_996),
.B(n_976),
.Y(n_1034)
);

BUFx3_ASAP7_75t_L g1035 ( 
.A(n_1001),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_994),
.B(n_976),
.Y(n_1036)
);

OR2x2_ASAP7_75t_L g1037 ( 
.A(n_999),
.B(n_987),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_1032),
.Y(n_1038)
);

NOR2xp67_ASAP7_75t_L g1039 ( 
.A(n_1023),
.B(n_1002),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_1017),
.B(n_997),
.Y(n_1040)
);

AND2x2_ASAP7_75t_L g1041 ( 
.A(n_1024),
.B(n_990),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_1017),
.B(n_1010),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_1022),
.B(n_1010),
.Y(n_1043)
);

HB1xp67_ASAP7_75t_L g1044 ( 
.A(n_1018),
.Y(n_1044)
);

INVx2_ASAP7_75t_SL g1045 ( 
.A(n_1035),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_1032),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_1025),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_1024),
.B(n_990),
.Y(n_1048)
);

BUFx2_ASAP7_75t_L g1049 ( 
.A(n_1035),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_1041),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_1044),
.B(n_1022),
.Y(n_1051)
);

AND2x4_ASAP7_75t_L g1052 ( 
.A(n_1041),
.B(n_1024),
.Y(n_1052)
);

OR2x2_ASAP7_75t_L g1053 ( 
.A(n_1040),
.B(n_1023),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_1048),
.B(n_1021),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1038),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_1048),
.B(n_1021),
.Y(n_1056)
);

INVx1_ASAP7_75t_SL g1057 ( 
.A(n_1049),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_1055),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1057),
.Y(n_1059)
);

BUFx3_ASAP7_75t_L g1060 ( 
.A(n_1057),
.Y(n_1060)
);

BUFx2_ASAP7_75t_L g1061 ( 
.A(n_1051),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_1052),
.B(n_1049),
.Y(n_1062)
);

INVxp67_ASAP7_75t_L g1063 ( 
.A(n_1060),
.Y(n_1063)
);

OAI322xp33_ASAP7_75t_L g1064 ( 
.A1(n_1059),
.A2(n_1016),
.A3(n_1054),
.B1(n_1056),
.B2(n_1043),
.C1(n_1053),
.C2(n_1037),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_1058),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_1061),
.A2(n_1016),
.B1(n_1052),
.B2(n_1050),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1058),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1060),
.Y(n_1068)
);

OR4x1_ASAP7_75t_L g1069 ( 
.A(n_1059),
.B(n_1045),
.C(n_1047),
.D(n_1046),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_1060),
.Y(n_1070)
);

OAI211xp5_ASAP7_75t_L g1071 ( 
.A1(n_1061),
.A2(n_1045),
.B(n_1039),
.C(n_1018),
.Y(n_1071)
);

OR2x6_ASAP7_75t_L g1072 ( 
.A(n_1060),
.B(n_927),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_1062),
.Y(n_1073)
);

OR2x2_ASAP7_75t_L g1074 ( 
.A(n_1061),
.B(n_1042),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_1063),
.B(n_1062),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_1068),
.B(n_1062),
.Y(n_1076)
);

OAI211xp5_ASAP7_75t_L g1077 ( 
.A1(n_1071),
.A2(n_1039),
.B(n_1035),
.C(n_967),
.Y(n_1077)
);

OAI31xp33_ASAP7_75t_L g1078 ( 
.A1(n_1066),
.A2(n_1037),
.A3(n_989),
.B(n_970),
.Y(n_1078)
);

INVxp67_ASAP7_75t_L g1079 ( 
.A(n_1070),
.Y(n_1079)
);

OR2x2_ASAP7_75t_L g1080 ( 
.A(n_1074),
.B(n_1047),
.Y(n_1080)
);

INVx3_ASAP7_75t_L g1081 ( 
.A(n_1073),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_1072),
.Y(n_1082)
);

INVxp67_ASAP7_75t_L g1083 ( 
.A(n_1072),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_1072),
.Y(n_1084)
);

OA21x2_ASAP7_75t_L g1085 ( 
.A1(n_1065),
.A2(n_1038),
.B(n_1046),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_1067),
.B(n_1025),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1069),
.Y(n_1087)
);

AOI321xp33_ASAP7_75t_L g1088 ( 
.A1(n_1064),
.A2(n_989),
.A3(n_977),
.B1(n_970),
.B2(n_986),
.C(n_984),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_1064),
.A2(n_872),
.B(n_1020),
.Y(n_1089)
);

AND2x4_ASAP7_75t_SL g1090 ( 
.A(n_1073),
.B(n_1027),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1063),
.B(n_1026),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1075),
.Y(n_1092)
);

OAI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_1087),
.A2(n_1026),
.B1(n_992),
.B2(n_1033),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1075),
.Y(n_1094)
);

INVx1_ASAP7_75t_SL g1095 ( 
.A(n_1076),
.Y(n_1095)
);

INVx1_ASAP7_75t_SL g1096 ( 
.A(n_1076),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_SL g1097 ( 
.A1(n_1088),
.A2(n_992),
.B1(n_954),
.B2(n_973),
.Y(n_1097)
);

OAI32xp33_ASAP7_75t_L g1098 ( 
.A1(n_1081),
.A2(n_1027),
.A3(n_968),
.B1(n_999),
.B2(n_935),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1081),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1091),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1079),
.B(n_1027),
.Y(n_1101)
);

OR2x2_ASAP7_75t_L g1102 ( 
.A(n_1080),
.B(n_990),
.Y(n_1102)
);

O2A1O1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_1077),
.A2(n_975),
.B(n_968),
.C(n_970),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1083),
.B(n_1036),
.Y(n_1104)
);

NAND2xp33_ASAP7_75t_L g1105 ( 
.A(n_1089),
.B(n_1036),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_1091),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1085),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_1085),
.Y(n_1108)
);

OAI321xp33_ASAP7_75t_L g1109 ( 
.A1(n_1082),
.A2(n_977),
.A3(n_986),
.B1(n_984),
.B2(n_1029),
.C(n_959),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1086),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1095),
.B(n_1090),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_1096),
.B(n_1084),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_1099),
.B(n_1086),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_1107),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_1092),
.B(n_1030),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1094),
.B(n_1078),
.Y(n_1116)
);

AOI211xp5_ASAP7_75t_L g1117 ( 
.A1(n_1103),
.A2(n_927),
.B(n_992),
.C(n_994),
.Y(n_1117)
);

NOR3xp33_ASAP7_75t_SL g1118 ( 
.A(n_1100),
.B(n_1106),
.C(n_1098),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_1101),
.B(n_1033),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_1101),
.B(n_1030),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1108),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1110),
.B(n_1036),
.Y(n_1122)
);

OAI21xp5_ASAP7_75t_L g1123 ( 
.A1(n_1097),
.A2(n_964),
.B(n_935),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1102),
.B(n_994),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_1104),
.B(n_1019),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1093),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_1093),
.A2(n_1105),
.B1(n_1031),
.B2(n_1019),
.Y(n_1127)
);

NAND5xp2_ASAP7_75t_L g1128 ( 
.A(n_1118),
.B(n_1109),
.C(n_862),
.D(n_1034),
.E(n_973),
.Y(n_1128)
);

O2A1O1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_1121),
.A2(n_834),
.B(n_839),
.C(n_959),
.Y(n_1129)
);

AOI221xp5_ASAP7_75t_L g1130 ( 
.A1(n_1114),
.A2(n_954),
.B1(n_992),
.B2(n_973),
.C(n_957),
.Y(n_1130)
);

NAND4xp25_ASAP7_75t_L g1131 ( 
.A(n_1111),
.B(n_937),
.C(n_1007),
.D(n_972),
.Y(n_1131)
);

AOI21xp33_ASAP7_75t_L g1132 ( 
.A1(n_1112),
.A2(n_1028),
.B(n_959),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1113),
.B(n_1019),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_1111),
.B(n_937),
.Y(n_1134)
);

AOI221xp5_ASAP7_75t_L g1135 ( 
.A1(n_1116),
.A2(n_954),
.B1(n_992),
.B2(n_957),
.C(n_1012),
.Y(n_1135)
);

NAND3xp33_ASAP7_75t_L g1136 ( 
.A(n_1126),
.B(n_992),
.C(n_954),
.Y(n_1136)
);

AOI222xp33_ASAP7_75t_L g1137 ( 
.A1(n_1123),
.A2(n_1122),
.B1(n_1115),
.B2(n_1119),
.C1(n_1125),
.C2(n_1120),
.Y(n_1137)
);

NAND3xp33_ASAP7_75t_SL g1138 ( 
.A(n_1117),
.B(n_943),
.C(n_1034),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_1127),
.B(n_1019),
.Y(n_1139)
);

OAI21xp33_ASAP7_75t_L g1140 ( 
.A1(n_1124),
.A2(n_1031),
.B(n_1012),
.Y(n_1140)
);

OAI31xp33_ASAP7_75t_L g1141 ( 
.A1(n_1121),
.A2(n_971),
.A3(n_957),
.B(n_943),
.Y(n_1141)
);

AOI322xp5_ASAP7_75t_L g1142 ( 
.A1(n_1118),
.A2(n_971),
.A3(n_1009),
.B1(n_965),
.B2(n_962),
.C1(n_943),
.C2(n_921),
.Y(n_1142)
);

INVx1_ASAP7_75t_SL g1143 ( 
.A(n_1111),
.Y(n_1143)
);

AOI32xp33_ASAP7_75t_L g1144 ( 
.A1(n_1112),
.A2(n_1012),
.A3(n_971),
.B1(n_937),
.B2(n_1031),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1121),
.Y(n_1145)
);

NAND4xp25_ASAP7_75t_L g1146 ( 
.A(n_1111),
.B(n_937),
.C(n_1007),
.D(n_972),
.Y(n_1146)
);

NOR4xp25_ASAP7_75t_L g1147 ( 
.A(n_1121),
.B(n_1028),
.C(n_1011),
.D(n_1015),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1112),
.B(n_1031),
.Y(n_1148)
);

AOI221xp5_ASAP7_75t_L g1149 ( 
.A1(n_1118),
.A2(n_954),
.B1(n_1012),
.B2(n_921),
.C(n_1028),
.Y(n_1149)
);

NOR3xp33_ASAP7_75t_SL g1150 ( 
.A(n_1112),
.B(n_1003),
.C(n_1015),
.Y(n_1150)
);

AOI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_1112),
.A2(n_891),
.B1(n_927),
.B2(n_937),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1143),
.Y(n_1152)
);

OAI22x1_ASAP7_75t_L g1153 ( 
.A1(n_1145),
.A2(n_881),
.B1(n_943),
.B2(n_1007),
.Y(n_1153)
);

AOI221xp5_ASAP7_75t_L g1154 ( 
.A1(n_1149),
.A2(n_1128),
.B1(n_1147),
.B2(n_1150),
.C(n_1135),
.Y(n_1154)
);

OAI22xp5_ASAP7_75t_L g1155 ( 
.A1(n_1148),
.A2(n_954),
.B1(n_1012),
.B2(n_927),
.Y(n_1155)
);

BUFx2_ASAP7_75t_L g1156 ( 
.A(n_1133),
.Y(n_1156)
);

AOI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_1151),
.A2(n_927),
.B1(n_1012),
.B2(n_1029),
.Y(n_1157)
);

AOI221xp5_ASAP7_75t_L g1158 ( 
.A1(n_1132),
.A2(n_991),
.B1(n_1015),
.B2(n_1011),
.C(n_1003),
.Y(n_1158)
);

AO22x2_ASAP7_75t_L g1159 ( 
.A1(n_1142),
.A2(n_948),
.B1(n_1009),
.B2(n_1011),
.Y(n_1159)
);

INVx2_ASAP7_75t_SL g1160 ( 
.A(n_1134),
.Y(n_1160)
);

AOI221xp5_ASAP7_75t_L g1161 ( 
.A1(n_1141),
.A2(n_991),
.B1(n_1003),
.B2(n_921),
.C(n_1009),
.Y(n_1161)
);

AOI322xp5_ASAP7_75t_L g1162 ( 
.A1(n_1130),
.A2(n_965),
.A3(n_962),
.B1(n_950),
.B2(n_1005),
.C1(n_1004),
.C2(n_1008),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_SL g1163 ( 
.A(n_1137),
.B(n_927),
.Y(n_1163)
);

AOI222xp33_ASAP7_75t_L g1164 ( 
.A1(n_1136),
.A2(n_965),
.B1(n_962),
.B2(n_915),
.C1(n_927),
.C2(n_918),
.Y(n_1164)
);

OAI221xp5_ASAP7_75t_L g1165 ( 
.A1(n_1144),
.A2(n_940),
.B1(n_1029),
.B2(n_881),
.C(n_985),
.Y(n_1165)
);

OA22x2_ASAP7_75t_L g1166 ( 
.A1(n_1139),
.A2(n_1002),
.B1(n_1029),
.B2(n_980),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_1140),
.A2(n_1029),
.B1(n_972),
.B2(n_1002),
.Y(n_1167)
);

NOR2xp33_ASAP7_75t_L g1168 ( 
.A(n_1131),
.B(n_1146),
.Y(n_1168)
);

AOI211xp5_ASAP7_75t_L g1169 ( 
.A1(n_1138),
.A2(n_1008),
.B(n_1005),
.C(n_1004),
.Y(n_1169)
);

AOI221xp5_ASAP7_75t_L g1170 ( 
.A1(n_1129),
.A2(n_1008),
.B1(n_1005),
.B2(n_1004),
.C(n_950),
.Y(n_1170)
);

AO22x2_ASAP7_75t_L g1171 ( 
.A1(n_1145),
.A2(n_948),
.B1(n_934),
.B2(n_932),
.Y(n_1171)
);

AOI22xp5_ASAP7_75t_L g1172 ( 
.A1(n_1149),
.A2(n_1029),
.B1(n_940),
.B2(n_948),
.Y(n_1172)
);

AOI211xp5_ASAP7_75t_L g1173 ( 
.A1(n_1149),
.A2(n_936),
.B(n_879),
.C(n_948),
.Y(n_1173)
);

OA22x2_ASAP7_75t_L g1174 ( 
.A1(n_1143),
.A2(n_1002),
.B1(n_980),
.B2(n_946),
.Y(n_1174)
);

OAI211xp5_ASAP7_75t_L g1175 ( 
.A1(n_1143),
.A2(n_1002),
.B(n_976),
.C(n_936),
.Y(n_1175)
);

AND2x4_ASAP7_75t_L g1176 ( 
.A(n_1152),
.B(n_1002),
.Y(n_1176)
);

NOR2x1_ASAP7_75t_L g1177 ( 
.A(n_1156),
.B(n_946),
.Y(n_1177)
);

NOR2x1_ASAP7_75t_L g1178 ( 
.A(n_1163),
.B(n_946),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1171),
.Y(n_1179)
);

NAND4xp75_ASAP7_75t_L g1180 ( 
.A(n_1160),
.B(n_987),
.C(n_980),
.D(n_934),
.Y(n_1180)
);

OR2x2_ASAP7_75t_L g1181 ( 
.A(n_1153),
.B(n_987),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1154),
.B(n_987),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1168),
.A2(n_934),
.B(n_932),
.Y(n_1183)
);

NAND2xp33_ASAP7_75t_L g1184 ( 
.A(n_1155),
.B(n_936),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_1171),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1159),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1159),
.Y(n_1187)
);

NOR2x1_ASAP7_75t_L g1188 ( 
.A(n_1175),
.B(n_936),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1174),
.Y(n_1189)
);

NOR2x1_ASAP7_75t_L g1190 ( 
.A(n_1165),
.B(n_936),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1166),
.Y(n_1191)
);

AOI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1157),
.A2(n_940),
.B1(n_961),
.B2(n_985),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1164),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1169),
.Y(n_1194)
);

AND3x4_ASAP7_75t_L g1195 ( 
.A(n_1162),
.B(n_934),
.C(n_932),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1161),
.Y(n_1196)
);

NOR2x1p5_ASAP7_75t_L g1197 ( 
.A(n_1173),
.B(n_961),
.Y(n_1197)
);

AND2x4_ASAP7_75t_L g1198 ( 
.A(n_1191),
.B(n_1172),
.Y(n_1198)
);

OAI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1189),
.A2(n_1158),
.B(n_1170),
.Y(n_1199)
);

OAI21x1_ASAP7_75t_L g1200 ( 
.A1(n_1179),
.A2(n_1167),
.B(n_846),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_SL g1201 ( 
.A(n_1193),
.B(n_961),
.Y(n_1201)
);

AOI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1195),
.A2(n_1182),
.B1(n_1186),
.B2(n_1187),
.Y(n_1202)
);

OAI211xp5_ASAP7_75t_SL g1203 ( 
.A1(n_1178),
.A2(n_1013),
.B(n_1000),
.C(n_993),
.Y(n_1203)
);

A2O1A1Ixp33_ASAP7_75t_L g1204 ( 
.A1(n_1194),
.A2(n_1013),
.B(n_1000),
.C(n_993),
.Y(n_1204)
);

OR4x1_ASAP7_75t_L g1205 ( 
.A(n_1196),
.B(n_988),
.C(n_981),
.D(n_918),
.Y(n_1205)
);

NAND3xp33_ASAP7_75t_L g1206 ( 
.A(n_1185),
.B(n_879),
.C(n_936),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1177),
.A2(n_940),
.B(n_985),
.Y(n_1207)
);

NAND3xp33_ASAP7_75t_L g1208 ( 
.A(n_1176),
.B(n_1000),
.C(n_993),
.Y(n_1208)
);

XOR2xp5_ASAP7_75t_L g1209 ( 
.A(n_1176),
.B(n_101),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1181),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1188),
.Y(n_1211)
);

NAND3xp33_ASAP7_75t_SL g1212 ( 
.A(n_1183),
.B(n_1013),
.C(n_1000),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1211),
.Y(n_1213)
);

XNOR2x1_ASAP7_75t_L g1214 ( 
.A(n_1198),
.B(n_1190),
.Y(n_1214)
);

INVx2_ASAP7_75t_SL g1215 ( 
.A(n_1209),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1210),
.A2(n_1184),
.B(n_1192),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1201),
.B(n_1197),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1199),
.A2(n_1180),
.B(n_940),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1202),
.B(n_985),
.Y(n_1219)
);

AOI211xp5_ASAP7_75t_L g1220 ( 
.A1(n_1206),
.A2(n_1013),
.B(n_950),
.C(n_988),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1204),
.A2(n_1208),
.B1(n_1207),
.B2(n_1205),
.Y(n_1221)
);

AOI211xp5_ASAP7_75t_L g1222 ( 
.A1(n_1203),
.A2(n_950),
.B(n_912),
.C(n_922),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1212),
.Y(n_1223)
);

OAI31xp33_ASAP7_75t_SL g1224 ( 
.A1(n_1200),
.A2(n_950),
.A3(n_880),
.B(n_985),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1199),
.B(n_960),
.Y(n_1225)
);

OAI211xp5_ASAP7_75t_L g1226 ( 
.A1(n_1202),
.A2(n_928),
.B(n_104),
.C(n_106),
.Y(n_1226)
);

XOR2xp5_ASAP7_75t_L g1227 ( 
.A(n_1209),
.B(n_103),
.Y(n_1227)
);

INVxp67_ASAP7_75t_SL g1228 ( 
.A(n_1214),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1213),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1215),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1227),
.Y(n_1231)
);

AOI22xp33_ASAP7_75t_SL g1232 ( 
.A1(n_1225),
.A2(n_940),
.B1(n_960),
.B2(n_912),
.Y(n_1232)
);

OAI22x1_ASAP7_75t_L g1233 ( 
.A1(n_1223),
.A2(n_928),
.B1(n_922),
.B2(n_919),
.Y(n_1233)
);

INVx4_ASAP7_75t_L g1234 ( 
.A(n_1219),
.Y(n_1234)
);

AOI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1221),
.A2(n_940),
.B1(n_960),
.B2(n_919),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1217),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1216),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1229),
.A2(n_1218),
.B1(n_1220),
.B2(n_1226),
.Y(n_1238)
);

HB1xp67_ASAP7_75t_L g1239 ( 
.A(n_1237),
.Y(n_1239)
);

AO22x2_ASAP7_75t_L g1240 ( 
.A1(n_1228),
.A2(n_1224),
.B1(n_1222),
.B2(n_920),
.Y(n_1240)
);

INVxp67_ASAP7_75t_SL g1241 ( 
.A(n_1236),
.Y(n_1241)
);

XOR2xp5_ASAP7_75t_L g1242 ( 
.A(n_1231),
.B(n_109),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_SL g1243 ( 
.A1(n_1230),
.A2(n_110),
.B1(n_112),
.B2(n_116),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_SL g1244 ( 
.A1(n_1241),
.A2(n_1234),
.B1(n_1235),
.B2(n_1232),
.Y(n_1244)
);

AOI221xp5_ASAP7_75t_L g1245 ( 
.A1(n_1238),
.A2(n_1233),
.B1(n_920),
.B2(n_916),
.C(n_924),
.Y(n_1245)
);

XNOR2x1_ASAP7_75t_L g1246 ( 
.A(n_1242),
.B(n_118),
.Y(n_1246)
);

XNOR2xp5_ASAP7_75t_L g1247 ( 
.A(n_1239),
.B(n_119),
.Y(n_1247)
);

AO21x2_ASAP7_75t_L g1248 ( 
.A1(n_1247),
.A2(n_1243),
.B(n_1240),
.Y(n_1248)
);

OR2x2_ASAP7_75t_L g1249 ( 
.A(n_1248),
.B(n_1246),
.Y(n_1249)
);

AOI21xp33_ASAP7_75t_L g1250 ( 
.A1(n_1249),
.A2(n_1244),
.B(n_1245),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1250),
.A2(n_123),
.B(n_126),
.Y(n_1251)
);

AOI221xp5_ASAP7_75t_L g1252 ( 
.A1(n_1251),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.C(n_131),
.Y(n_1252)
);

AOI211xp5_ASAP7_75t_L g1253 ( 
.A1(n_1252),
.A2(n_136),
.B(n_137),
.C(n_145),
.Y(n_1253)
);


endmodule