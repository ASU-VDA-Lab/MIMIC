module fake_jpeg_2803_n_508 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_508);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_508;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

CKINVDCx14_ASAP7_75t_R g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_49),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_53),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_20),
.B(n_9),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_54),
.B(n_80),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_55),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_56),
.Y(n_154)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_59),
.Y(n_108)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_60),
.Y(n_112)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_62),
.Y(n_147)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g134 ( 
.A(n_63),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_64),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx8_ASAP7_75t_L g141 ( 
.A(n_65),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_66),
.Y(n_130)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_67),
.Y(n_145)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_68),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_69),
.Y(n_109)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_71),
.Y(n_129)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_20),
.Y(n_72)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

INVx3_ASAP7_75t_SL g73 ( 
.A(n_36),
.Y(n_73)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_36),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_96),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_75),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_76),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_78),
.Y(n_117)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_40),
.B(n_8),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_82),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_47),
.B(n_8),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_85),
.B(n_45),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_86),
.Y(n_127)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_87),
.Y(n_135)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_88),
.Y(n_152)
);

INVx4_ASAP7_75t_SL g89 ( 
.A(n_23),
.Y(n_89)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_89),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_90),
.B(n_95),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_91),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_24),
.Y(n_92)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_92),
.Y(n_126)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

NAND2xp33_ASAP7_75t_SL g131 ( 
.A(n_93),
.B(n_94),
.Y(n_131)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_23),
.Y(n_94)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_36),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_48),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_113),
.B(n_132),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_L g124 ( 
.A1(n_68),
.A2(n_36),
.B1(n_33),
.B2(n_25),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_124),
.A2(n_128),
.B1(n_137),
.B2(n_138),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_75),
.A2(n_29),
.B1(n_33),
.B2(n_37),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_73),
.B(n_47),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_48),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_136),
.B(n_149),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_65),
.A2(n_29),
.B1(n_35),
.B2(n_44),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_49),
.A2(n_29),
.B1(n_34),
.B2(n_38),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_50),
.A2(n_34),
.B1(n_27),
.B2(n_41),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_139),
.A2(n_140),
.B1(n_109),
.B2(n_134),
.Y(n_165)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_60),
.Y(n_142)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_142),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_77),
.A2(n_25),
.B1(n_37),
.B2(n_45),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_143),
.A2(n_28),
.B1(n_38),
.B2(n_19),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_65),
.A2(n_34),
.B1(n_36),
.B2(n_41),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_144),
.A2(n_90),
.B1(n_156),
.B2(n_140),
.Y(n_163)
);

AND2x2_ASAP7_75t_SL g146 ( 
.A(n_96),
.B(n_46),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_146),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_148),
.B(n_155),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_69),
.B(n_18),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_81),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_150),
.B(n_153),
.Y(n_179)
);

NOR2x1_ASAP7_75t_L g151 ( 
.A(n_67),
.B(n_26),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g186 ( 
.A(n_151),
.B(n_28),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_69),
.B(n_18),
.Y(n_153)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_110),
.Y(n_157)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_157),
.Y(n_217)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_99),
.Y(n_158)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_158),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_106),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_159),
.B(n_203),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_160),
.A2(n_194),
.B1(n_214),
.B2(n_3),
.Y(n_264)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_97),
.Y(n_162)
);

INVx2_ASAP7_75t_SL g229 ( 
.A(n_162),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_163),
.Y(n_239)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_100),
.Y(n_164)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_164),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_165),
.A2(n_130),
.B1(n_122),
.B2(n_108),
.Y(n_238)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_98),
.Y(n_166)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_166),
.Y(n_232)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_104),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_167),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_117),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_168),
.Y(n_251)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_141),
.Y(n_169)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_169),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_118),
.B(n_26),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_170),
.B(n_183),
.Y(n_215)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_119),
.Y(n_172)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_172),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_128),
.A2(n_19),
.B1(n_83),
.B2(n_91),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_174),
.A2(n_187),
.B1(n_154),
.B2(n_101),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_90),
.Y(n_175)
);

OAI21xp33_ASAP7_75t_L g245 ( 
.A1(n_175),
.A2(n_186),
.B(n_193),
.Y(n_245)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_176),
.Y(n_223)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_101),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_177),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g178 ( 
.A(n_109),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_178),
.Y(n_241)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_115),
.Y(n_180)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_180),
.Y(n_222)
);

FAx1_ASAP7_75t_SL g181 ( 
.A(n_146),
.B(n_151),
.CI(n_131),
.CON(n_181),
.SN(n_181)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_181),
.B(n_196),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_135),
.B(n_92),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_182),
.B(n_208),
.C(n_107),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_124),
.B(n_31),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_116),
.Y(n_184)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_184),
.Y(n_236)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_126),
.Y(n_185)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_185),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_143),
.A2(n_84),
.B1(n_86),
.B2(n_58),
.Y(n_187)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_111),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_188),
.Y(n_261)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_112),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_189),
.B(n_192),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_120),
.B(n_31),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_190),
.B(n_0),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_144),
.A2(n_28),
.B(n_71),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_191),
.A2(n_108),
.B(n_147),
.Y(n_224)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_121),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_114),
.A2(n_27),
.B1(n_41),
.B2(n_46),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_137),
.A2(n_56),
.B1(n_53),
.B2(n_66),
.Y(n_194)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_112),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_195),
.B(n_197),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_134),
.B(n_95),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_129),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_123),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_198),
.B(n_204),
.Y(n_246)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_111),
.Y(n_199)
);

INVx8_ASAP7_75t_L g230 ( 
.A(n_199),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_114),
.B(n_70),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_201),
.B(n_202),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_130),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_127),
.Y(n_204)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_145),
.Y(n_205)
);

INVx8_ASAP7_75t_L g259 ( 
.A(n_205),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_152),
.B(n_46),
.Y(n_206)
);

OAI21xp33_ASAP7_75t_L g247 ( 
.A1(n_206),
.A2(n_210),
.B(n_213),
.Y(n_247)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_129),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_207),
.B(n_209),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_105),
.B(n_64),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_133),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_155),
.A2(n_46),
.B1(n_41),
.B2(n_27),
.Y(n_210)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_145),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g248 ( 
.A(n_212),
.B(n_30),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_107),
.A2(n_27),
.B1(n_41),
.B2(n_46),
.Y(n_213)
);

OAI22xp33_ASAP7_75t_L g214 ( 
.A1(n_133),
.A2(n_62),
.B1(n_59),
.B2(n_27),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g286 ( 
.A1(n_216),
.A2(n_204),
.B1(n_198),
.B2(n_192),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_224),
.A2(n_256),
.B(n_14),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_173),
.A2(n_105),
.B1(n_147),
.B2(n_103),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_226),
.A2(n_252),
.B1(n_255),
.B2(n_178),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_227),
.B(n_228),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_186),
.A2(n_154),
.B1(n_125),
.B2(n_102),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_231),
.A2(n_243),
.B1(n_5),
.B2(n_6),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_182),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_235),
.B(n_240),
.Y(n_270)
);

INVx6_ASAP7_75t_L g237 ( 
.A(n_177),
.Y(n_237)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_237),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_238),
.B(n_264),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_190),
.B(n_103),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_183),
.A2(n_125),
.B1(n_102),
.B2(n_122),
.Y(n_243)
);

NAND2xp33_ASAP7_75t_SL g244 ( 
.A(n_175),
.B(n_181),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_244),
.A2(n_164),
.B(n_209),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g291 ( 
.A(n_248),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_200),
.A2(n_30),
.B1(n_1),
.B2(n_2),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_250),
.A2(n_205),
.B1(n_176),
.B2(n_169),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_165),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_179),
.B(n_0),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_254),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_170),
.B(n_1),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_181),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_191),
.A2(n_175),
.B(n_194),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_171),
.B(n_3),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_258),
.B(n_254),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_211),
.B(n_11),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_260),
.B(n_12),
.C(n_5),
.Y(n_290)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_222),
.Y(n_267)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_267),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_239),
.A2(n_160),
.B1(n_195),
.B2(n_188),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_268),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_235),
.B(n_180),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_269),
.B(n_273),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_256),
.A2(n_214),
.B1(n_172),
.B2(n_167),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_271),
.A2(n_287),
.B1(n_292),
.B2(n_297),
.Y(n_318)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_222),
.Y(n_272)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_272),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_242),
.B(n_157),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_229),
.Y(n_275)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_275),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_227),
.B(n_158),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g347 ( 
.A(n_276),
.B(n_277),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_242),
.B(n_161),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_239),
.A2(n_199),
.B1(n_212),
.B2(n_189),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_278),
.Y(n_352)
);

NOR3xp33_ASAP7_75t_L g279 ( 
.A(n_220),
.B(n_215),
.C(n_240),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_279),
.B(n_281),
.Y(n_317)
);

HB1xp67_ASAP7_75t_L g351 ( 
.A(n_280),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_232),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_282),
.A2(n_296),
.B(n_303),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_285),
.B(n_290),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_L g320 ( 
.A1(n_286),
.A2(n_295),
.B1(n_221),
.B2(n_236),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_220),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_288),
.B(n_298),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_228),
.B(n_184),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_289),
.B(n_294),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_215),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_244),
.B(n_17),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_293),
.B(n_302),
.C(n_308),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_253),
.B(n_4),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_238),
.A2(n_5),
.B1(n_7),
.B2(n_10),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_264),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_233),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_224),
.A2(n_7),
.B1(n_10),
.B2(n_11),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_299),
.A2(n_300),
.B1(n_305),
.B2(n_311),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_248),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_251),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_301),
.B(n_304),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_SL g302 ( 
.A(n_255),
.B(n_245),
.C(n_260),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_226),
.B(n_13),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_246),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_248),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_229),
.Y(n_306)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_306),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_307),
.A2(n_280),
.B(n_303),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_249),
.B(n_17),
.C(n_258),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_229),
.Y(n_309)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_309),
.Y(n_335)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_217),
.Y(n_310)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_310),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_247),
.A2(n_17),
.B1(n_252),
.B2(n_217),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g312 ( 
.A1(n_261),
.A2(n_17),
.B1(n_263),
.B2(n_219),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_312),
.A2(n_236),
.B1(n_265),
.B2(n_225),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_283),
.A2(n_261),
.B1(n_237),
.B2(n_263),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_314),
.A2(n_337),
.B1(n_287),
.B2(n_281),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_307),
.A2(n_262),
.B(n_234),
.Y(n_315)
);

AO21x1_ASAP7_75t_L g368 ( 
.A1(n_315),
.A2(n_319),
.B(n_322),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_291),
.A2(n_234),
.B(n_230),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_320),
.A2(n_330),
.B1(n_338),
.B2(n_346),
.Y(n_373)
);

XNOR2x2_ASAP7_75t_L g322 ( 
.A(n_270),
.B(n_221),
.Y(n_322)
);

OAI32xp33_ASAP7_75t_L g326 ( 
.A1(n_270),
.A2(n_273),
.A3(n_279),
.B1(n_277),
.B2(n_303),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_326),
.B(n_340),
.Y(n_382)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_267),
.Y(n_328)
);

INVx2_ASAP7_75t_SL g380 ( 
.A(n_328),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_266),
.B(n_234),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_SL g372 ( 
.A(n_332),
.B(n_343),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_291),
.A2(n_230),
.B(n_218),
.Y(n_333)
);

AOI21x1_ASAP7_75t_L g375 ( 
.A1(n_333),
.A2(n_344),
.B(n_353),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_283),
.A2(n_257),
.B1(n_218),
.B2(n_259),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_283),
.A2(n_289),
.B1(n_271),
.B2(n_266),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_269),
.B(n_225),
.Y(n_340)
);

AO22x1_ASAP7_75t_SL g341 ( 
.A1(n_283),
.A2(n_265),
.B1(n_257),
.B2(n_223),
.Y(n_341)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_341),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_285),
.B(n_223),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_282),
.A2(n_259),
.B(n_241),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_304),
.B(n_293),
.C(n_302),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_345),
.B(n_308),
.C(n_301),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_311),
.A2(n_223),
.B1(n_257),
.B2(n_299),
.Y(n_346)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_272),
.Y(n_349)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_349),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_284),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_350),
.B(n_284),
.Y(n_365)
);

OAI32xp33_ASAP7_75t_L g354 ( 
.A1(n_317),
.A2(n_303),
.A3(n_310),
.B1(n_275),
.B2(n_309),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_354),
.B(n_357),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_332),
.B(n_274),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_355),
.B(n_359),
.C(n_360),
.Y(n_390)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_321),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_356),
.B(n_361),
.Y(n_405)
);

OAI32xp33_ASAP7_75t_L g357 ( 
.A1(n_322),
.A2(n_306),
.A3(n_274),
.B1(n_295),
.B2(n_294),
.Y(n_357)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_358),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_316),
.B(n_276),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_324),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_316),
.B(n_298),
.C(n_290),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_362),
.B(n_369),
.C(n_374),
.Y(n_398)
);

AO22x1_ASAP7_75t_L g363 ( 
.A1(n_314),
.A2(n_297),
.B1(n_300),
.B2(n_305),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_363),
.B(n_371),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_338),
.A2(n_351),
.B1(n_318),
.B2(n_353),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_364),
.A2(n_381),
.B1(n_383),
.B2(n_384),
.Y(n_407)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_365),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_322),
.B(n_292),
.Y(n_369)
);

AOI322xp5_ASAP7_75t_L g370 ( 
.A1(n_326),
.A2(n_284),
.A3(n_286),
.B1(n_312),
.B2(n_324),
.C1(n_340),
.C2(n_342),
.Y(n_370)
);

BUFx24_ASAP7_75t_SL g388 ( 
.A(n_370),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_330),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_345),
.B(n_331),
.Y(n_374)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_328),
.Y(n_376)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_376),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_331),
.B(n_343),
.C(n_319),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_377),
.B(n_379),
.C(n_372),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_327),
.A2(n_352),
.B1(n_337),
.B2(n_348),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_378),
.A2(n_375),
.B(n_368),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_315),
.B(n_333),
.C(n_344),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_318),
.A2(n_346),
.B1(n_336),
.B2(n_327),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_336),
.A2(n_341),
.B1(n_339),
.B2(n_325),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_341),
.A2(n_313),
.B1(n_339),
.B2(n_325),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_349),
.Y(n_385)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_385),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_347),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_386),
.Y(n_395)
);

NOR2x1_ASAP7_75t_R g387 ( 
.A(n_313),
.B(n_323),
.Y(n_387)
);

AO21x1_ASAP7_75t_L g397 ( 
.A1(n_387),
.A2(n_347),
.B(n_334),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_361),
.A2(n_352),
.B1(n_348),
.B2(n_350),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_389),
.B(n_394),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_375),
.A2(n_368),
.B(n_382),
.Y(n_392)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_392),
.A2(n_406),
.B(n_412),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_366),
.A2(n_329),
.B1(n_334),
.B2(n_335),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_374),
.B(n_323),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_396),
.B(n_414),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_397),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_SL g400 ( 
.A(n_372),
.B(n_329),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_400),
.B(n_397),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_366),
.A2(n_335),
.B1(n_382),
.B2(n_371),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_401),
.B(n_403),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_378),
.A2(n_358),
.B1(n_364),
.B2(n_381),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_383),
.A2(n_373),
.B1(n_384),
.B2(n_369),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g425 ( 
.A1(n_408),
.A2(n_411),
.B1(n_407),
.B2(n_393),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_377),
.B(n_355),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_409),
.B(n_410),
.C(n_362),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_379),
.A2(n_359),
.B1(n_354),
.B2(n_357),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_387),
.A2(n_380),
.B(n_367),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_380),
.A2(n_367),
.B(n_376),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_385),
.Y(n_415)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_415),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_380),
.A2(n_363),
.B(n_360),
.Y(n_416)
);

CKINVDCx16_ASAP7_75t_R g439 ( 
.A(n_416),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_405),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_417),
.B(n_426),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_421),
.B(n_433),
.Y(n_444)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_405),
.Y(n_422)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_422),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_395),
.B(n_363),
.Y(n_423)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_423),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_409),
.B(n_410),
.C(n_398),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_424),
.B(n_427),
.C(n_411),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_425),
.A2(n_430),
.B1(n_431),
.B2(n_432),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_395),
.B(n_414),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_398),
.B(n_390),
.C(n_396),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_402),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_428),
.B(n_434),
.Y(n_449)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_394),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_402),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_413),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_399),
.B(n_401),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_399),
.Y(n_434)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_413),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_437),
.B(n_412),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_390),
.B(n_416),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_438),
.B(n_400),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_SL g454 ( 
.A(n_440),
.B(n_408),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_425),
.A2(n_403),
.B1(n_433),
.B2(n_404),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_441),
.A2(n_420),
.B1(n_435),
.B2(n_419),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_SL g461 ( 
.A(n_442),
.B(n_454),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_443),
.B(n_446),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_438),
.B(n_427),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_445),
.B(n_447),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_421),
.B(n_392),
.C(n_406),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_424),
.B(n_391),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g450 ( 
.A(n_417),
.B(n_397),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_450),
.B(n_456),
.Y(n_467)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_451),
.Y(n_472)
);

AO21x1_ASAP7_75t_L g452 ( 
.A1(n_429),
.A2(n_391),
.B(n_404),
.Y(n_452)
);

CKINVDCx16_ASAP7_75t_R g473 ( 
.A(n_452),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_439),
.B(n_389),
.C(n_393),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_455),
.B(n_457),
.C(n_426),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_422),
.B(n_388),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_439),
.B(n_407),
.C(n_415),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_434),
.B(n_436),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_459),
.B(n_434),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_462),
.A2(n_465),
.B1(n_475),
.B2(n_466),
.Y(n_484)
);

XNOR2x1_ASAP7_75t_L g463 ( 
.A(n_454),
.B(n_436),
.Y(n_463)
);

MAJx2_ASAP7_75t_L g479 ( 
.A(n_463),
.B(n_446),
.C(n_442),
.Y(n_479)
);

AND2x2_ASAP7_75t_L g478 ( 
.A(n_464),
.B(n_457),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_441),
.A2(n_423),
.B1(n_420),
.B2(n_419),
.Y(n_465)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_466),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_445),
.B(n_430),
.C(n_429),
.Y(n_469)
);

NOR2xp67_ASAP7_75t_SL g486 ( 
.A(n_469),
.B(n_470),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_444),
.B(n_440),
.C(n_428),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_444),
.B(n_418),
.C(n_431),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_474),
.B(n_448),
.C(n_458),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g475 ( 
.A1(n_460),
.A2(n_418),
.B1(n_432),
.B2(n_437),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_464),
.B(n_443),
.C(n_447),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_476),
.B(n_478),
.Y(n_488)
);

XOR2xp5_ASAP7_75t_L g492 ( 
.A(n_479),
.B(n_461),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_471),
.B(n_455),
.C(n_453),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_480),
.B(n_482),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_472),
.A2(n_460),
.B(n_452),
.Y(n_481)
);

NOR3xp33_ASAP7_75t_L g489 ( 
.A(n_481),
.B(n_472),
.C(n_469),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_467),
.A2(n_449),
.B1(n_458),
.B2(n_473),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_483),
.B(n_484),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_471),
.B(n_468),
.C(n_474),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_485),
.B(n_463),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_485),
.B(n_470),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_487),
.B(n_489),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_492),
.B(n_493),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_SL g494 ( 
.A1(n_488),
.A2(n_478),
.B(n_477),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_494),
.A2(n_491),
.B(n_475),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_490),
.B(n_476),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_495),
.B(n_486),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_491),
.B(n_480),
.Y(n_496)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_496),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g503 ( 
.A(n_499),
.Y(n_503)
);

O2A1O1Ixp33_ASAP7_75t_SL g502 ( 
.A1(n_500),
.A2(n_501),
.B(n_498),
.C(n_497),
.Y(n_502)
);

AOI21xp5_ASAP7_75t_SL g504 ( 
.A1(n_502),
.A2(n_462),
.B(n_465),
.Y(n_504)
);

HB1xp67_ASAP7_75t_L g505 ( 
.A(n_504),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_505),
.A2(n_503),
.B(n_479),
.Y(n_506)
);

NAND2x1p5_ASAP7_75t_L g507 ( 
.A(n_506),
.B(n_461),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_507),
.Y(n_508)
);


endmodule