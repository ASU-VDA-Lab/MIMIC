module fake_jpeg_25232_n_137 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_137);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_34),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_15),
.B(n_35),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_26),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_21),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_32),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_18),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_27),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_22),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_23),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_29),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_39),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_62),
.Y(n_73)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx4f_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

BUFx2_ASAP7_75t_R g65 ( 
.A(n_52),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_52),
.Y(n_75)
);

CKINVDCx11_ASAP7_75t_R g70 ( 
.A(n_65),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_70),
.B(n_72),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_60),
.A2(n_49),
.B1(n_40),
.B2(n_55),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_74),
.A2(n_50),
.B1(n_48),
.B2(n_45),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_75),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_62),
.B(n_43),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_76),
.B(n_0),
.Y(n_82)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_62),
.B(n_57),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_78),
.B(n_43),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_61),
.A2(n_56),
.B1(n_53),
.B2(n_51),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_79),
.A2(n_46),
.B1(n_44),
.B2(n_68),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_80),
.B(n_82),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_L g81 ( 
.A1(n_67),
.A2(n_41),
.B1(n_42),
.B2(n_47),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_81),
.A2(n_90),
.B1(n_83),
.B2(n_92),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_73),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_85),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_73),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_86),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_0),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_93),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_71),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_69),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_92),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_1),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_1),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_94),
.B(n_2),
.Y(n_102)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_98),
.A2(n_84),
.B1(n_88),
.B2(n_4),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_99),
.Y(n_110)
);

NOR3xp33_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_81),
.C(n_87),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_102),
.B(n_3),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_105),
.B(n_107),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_109),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_24),
.C(n_5),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_25),
.C(n_12),
.Y(n_122)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_96),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_103),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_95),
.Y(n_121)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_110),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_114),
.Y(n_124)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_106),
.B(n_98),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_116),
.B(n_120),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_110),
.A2(n_28),
.B(n_7),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_118),
.Y(n_123)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_111),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_119),
.Y(n_127)
);

BUFx24_ASAP7_75t_SL g120 ( 
.A(n_111),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_121),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_112),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_128),
.B(n_129),
.C(n_127),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_125),
.B(n_115),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_130),
.B(n_123),
.C(n_126),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_131),
.B(n_122),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_132),
.A2(n_31),
.B(n_13),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_122),
.B(n_14),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_134),
.B(n_33),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_135),
.A2(n_30),
.B(n_17),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_19),
.Y(n_137)
);


endmodule