module fake_jpeg_21778_n_26 (n_3, n_2, n_1, n_0, n_4, n_5, n_26);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_26;

wire n_13;
wire n_21;
wire n_10;
wire n_23;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

BUFx3_ASAP7_75t_L g6 ( 
.A(n_5),
.Y(n_6)
);

INVx2_ASAP7_75t_R g7 ( 
.A(n_1),
.Y(n_7)
);

INVx5_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

BUFx12f_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

OA22x2_ASAP7_75t_L g12 ( 
.A1(n_7),
.A2(n_3),
.B1(n_4),
.B2(n_9),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_12),
.A2(n_17),
.B1(n_13),
.B2(n_16),
.Y(n_20)
);

INVx13_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

OR2x2_ASAP7_75t_SL g14 ( 
.A(n_9),
.B(n_6),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_14),
.A2(n_18),
.B(n_12),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_11),
.B(n_8),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_15),
.B(n_16),
.Y(n_21)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

OA22x2_ASAP7_75t_L g17 ( 
.A1(n_10),
.A2(n_7),
.B1(n_9),
.B2(n_6),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_6),
.A2(n_10),
.B(n_7),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_19),
.B(n_20),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_22),
.B(n_21),
.C(n_19),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g24 ( 
.A(n_23),
.B(n_20),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_24),
.Y(n_25)
);

BUFx24_ASAP7_75t_SL g26 ( 
.A(n_25),
.Y(n_26)
);


endmodule