module fake_jpeg_30920_n_484 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_484);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_484;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx5_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_51),
.Y(n_130)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_53),
.Y(n_144)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_54),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_41),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_55),
.B(n_61),
.Y(n_111)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_58),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_22),
.B(n_16),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_59),
.B(n_63),
.Y(n_123)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_60),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_41),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_62),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_22),
.B(n_15),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_64),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_39),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_65),
.B(n_73),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_66),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

BUFx2_ASAP7_75t_L g153 ( 
.A(n_67),
.Y(n_153)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_69),
.Y(n_150)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_71),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_72),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_39),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_17),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_75),
.A2(n_28),
.B1(n_27),
.B2(n_38),
.Y(n_129)
);

BUFx24_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g138 ( 
.A(n_76),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_77),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_78),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_79),
.Y(n_152)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_80),
.Y(n_135)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_81),
.Y(n_141)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_82),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_48),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_83),
.B(n_88),
.Y(n_128)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_84),
.Y(n_146)
);

BUFx10_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_85),
.Y(n_139)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_87),
.Y(n_121)
);

INVx6_ASAP7_75t_SL g88 ( 
.A(n_17),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_24),
.B(n_15),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_94),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_39),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_90),
.B(n_92),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_91),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_39),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_30),
.Y(n_93)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_93),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_24),
.B(n_40),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_17),
.Y(n_95)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_95),
.Y(n_142)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_46),
.Y(n_96)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_96),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_20),
.Y(n_97)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_97),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_33),
.B(n_13),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_98),
.B(n_33),
.Y(n_114)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_23),
.Y(n_99)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_99),
.Y(n_156)
);

HAxp5_ASAP7_75t_SL g101 ( 
.A(n_76),
.B(n_23),
.CON(n_101),
.SN(n_101)
);

OR2x4_ASAP7_75t_L g180 ( 
.A(n_101),
.B(n_34),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_88),
.A2(n_45),
.B1(n_20),
.B2(n_31),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_104),
.A2(n_148),
.B1(n_51),
.B2(n_91),
.Y(n_158)
);

AND2x2_ASAP7_75t_SL g105 ( 
.A(n_81),
.B(n_45),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_105),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_95),
.A2(n_43),
.B1(n_31),
.B2(n_18),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_112),
.A2(n_115),
.B1(n_122),
.B2(n_125),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_114),
.B(n_11),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_84),
.A2(n_40),
.B1(n_43),
.B2(n_31),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_75),
.B(n_47),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_117),
.B(n_118),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_64),
.B(n_47),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_57),
.A2(n_18),
.B1(n_43),
.B2(n_42),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_58),
.A2(n_18),
.B1(n_23),
.B2(n_44),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_129),
.A2(n_37),
.B1(n_34),
.B2(n_76),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_83),
.B(n_38),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_136),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_52),
.B(n_28),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_60),
.B(n_44),
.C(n_23),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_155),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_72),
.A2(n_27),
.B1(n_34),
.B2(n_39),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_74),
.A2(n_37),
.B1(n_34),
.B2(n_13),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_133),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_157),
.B(n_164),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_158),
.A2(n_159),
.B1(n_183),
.B2(n_199),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_101),
.A2(n_97),
.B1(n_96),
.B2(n_87),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_128),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_160),
.Y(n_224)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_116),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_163),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_103),
.Y(n_164)
);

A2O1A1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_106),
.A2(n_123),
.B(n_100),
.C(n_107),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_165),
.B(n_85),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_109),
.B(n_99),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_166),
.B(n_174),
.Y(n_214)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_144),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_167),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_111),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_168),
.B(n_175),
.Y(n_213)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_126),
.Y(n_169)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_169),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_170),
.B(n_180),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_130),
.Y(n_171)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_171),
.Y(n_242)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_149),
.Y(n_173)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_173),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_123),
.B(n_62),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_128),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_120),
.B(n_66),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_176),
.B(n_200),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_153),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_177),
.B(n_179),
.Y(n_229)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_156),
.Y(n_178)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_178),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_145),
.Y(n_179)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_113),
.Y(n_181)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_181),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_131),
.A2(n_11),
.B1(n_10),
.B2(n_29),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g223 ( 
.A(n_182),
.B(n_196),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_153),
.A2(n_93),
.B1(n_67),
.B2(n_69),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_105),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_184),
.B(n_190),
.Y(n_233)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_147),
.Y(n_185)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_185),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_119),
.Y(n_186)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_186),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_116),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_188),
.Y(n_217)
);

AO22x2_ASAP7_75t_SL g189 ( 
.A1(n_125),
.A2(n_79),
.B1(n_78),
.B2(n_77),
.Y(n_189)
);

OA22x2_ASAP7_75t_L g212 ( 
.A1(n_189),
.A2(n_112),
.B1(n_142),
.B2(n_121),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_148),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_191),
.B(n_192),
.Y(n_244)
);

BUFx12f_ASAP7_75t_L g192 ( 
.A(n_144),
.Y(n_192)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_130),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_193),
.Y(n_219)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_108),
.Y(n_194)
);

HB1xp67_ASAP7_75t_L g237 ( 
.A(n_194),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_151),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g225 ( 
.A(n_195),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_132),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_119),
.Y(n_197)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_197),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_132),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_198),
.B(n_207),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g199 ( 
.A(n_138),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_146),
.Y(n_200)
);

INVx11_ASAP7_75t_L g201 ( 
.A(n_150),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_201),
.A2(n_204),
.B1(n_150),
.B2(n_154),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_104),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_202),
.B(n_203),
.Y(n_231)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_146),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_108),
.Y(n_204)
);

AOI21xp33_ASAP7_75t_SL g206 ( 
.A1(n_138),
.A2(n_85),
.B(n_53),
.Y(n_206)
);

AOI21xp33_ASAP7_75t_L g230 ( 
.A1(n_206),
.A2(n_135),
.B(n_29),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_139),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_212),
.B(n_230),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_141),
.C(n_110),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_215),
.B(n_235),
.C(n_193),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_191),
.A2(n_140),
.B1(n_152),
.B2(n_124),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_218),
.A2(n_220),
.B1(n_247),
.B2(n_172),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_161),
.A2(n_152),
.B1(n_124),
.B2(n_143),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_162),
.B(n_110),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_222),
.B(n_181),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_161),
.A2(n_139),
.B(n_135),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_226),
.A2(n_204),
.B(n_194),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_227),
.B(n_239),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_187),
.B(n_141),
.C(n_102),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_236),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_162),
.B(n_205),
.Y(n_239)
);

OA22x2_ASAP7_75t_L g241 ( 
.A1(n_172),
.A2(n_102),
.B1(n_143),
.B2(n_127),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_241),
.Y(n_263)
);

OAI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_202),
.A2(n_189),
.B1(n_161),
.B2(n_180),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_246),
.A2(n_160),
.B1(n_170),
.B2(n_166),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_189),
.A2(n_154),
.B1(n_127),
.B2(n_80),
.Y(n_247)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_221),
.Y(n_249)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_249),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_250),
.A2(n_256),
.B1(n_269),
.B2(n_284),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_211),
.B(n_174),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_251),
.B(n_270),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_252),
.A2(n_265),
.B1(n_267),
.B2(n_257),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_229),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_253),
.B(n_266),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_210),
.A2(n_176),
.B1(n_178),
.B2(n_173),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_254),
.A2(n_218),
.B1(n_224),
.B2(n_212),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_255),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_247),
.A2(n_214),
.B1(n_223),
.B2(n_228),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_210),
.A2(n_182),
.B(n_165),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_257),
.A2(n_261),
.B(n_267),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_258),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_210),
.A2(n_203),
.B(n_200),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_221),
.Y(n_262)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_262),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_264),
.B(n_243),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_239),
.B(n_185),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_223),
.A2(n_231),
.B(n_226),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_209),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_268),
.B(n_283),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_228),
.A2(n_163),
.B1(n_188),
.B2(n_169),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_225),
.B(n_199),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_231),
.A2(n_199),
.B(n_167),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_271),
.B(n_243),
.Y(n_301)
);

XNOR2x2_ASAP7_75t_L g272 ( 
.A(n_227),
.B(n_214),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_272),
.B(n_275),
.Y(n_310)
);

INVx4_ASAP7_75t_L g273 ( 
.A(n_242),
.Y(n_273)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_273),
.Y(n_287)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_232),
.Y(n_274)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_274),
.Y(n_318)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_232),
.Y(n_276)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_276),
.Y(n_294)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_238),
.Y(n_277)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_277),
.Y(n_296)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_238),
.Y(n_278)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_278),
.Y(n_300)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_248),
.Y(n_279)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_279),
.Y(n_302)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_248),
.Y(n_280)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_280),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_235),
.B(n_215),
.C(n_222),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_224),
.C(n_241),
.Y(n_288)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_245),
.Y(n_282)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_282),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_209),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_208),
.A2(n_241),
.B1(n_220),
.B2(n_212),
.Y(n_284)
);

OAI32xp33_ASAP7_75t_L g285 ( 
.A1(n_272),
.A2(n_244),
.A3(n_233),
.B1(n_213),
.B2(n_241),
.Y(n_285)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_285),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_288),
.B(n_292),
.C(n_297),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_289),
.B(n_303),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_290),
.A2(n_291),
.B1(n_265),
.B2(n_263),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_245),
.C(n_219),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_260),
.B(n_234),
.C(n_237),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_301),
.A2(n_279),
.B(n_276),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_264),
.B(n_212),
.Y(n_303)
);

BUFx24_ASAP7_75t_L g307 ( 
.A(n_271),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_307),
.Y(n_338)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_249),
.Y(n_308)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_308),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_268),
.B(n_243),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_311),
.B(n_315),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_281),
.B(n_255),
.C(n_265),
.Y(n_313)
);

MAJx2_ASAP7_75t_L g328 ( 
.A(n_313),
.B(n_261),
.C(n_275),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_284),
.A2(n_216),
.B1(n_234),
.B2(n_240),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_314),
.A2(n_263),
.B1(n_254),
.B2(n_259),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_283),
.B(n_240),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_262),
.Y(n_316)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_316),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_295),
.B(n_253),
.Y(n_319)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_319),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_320),
.B(n_325),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_317),
.B(n_306),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_322),
.B(n_323),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_311),
.B(n_256),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g327 ( 
.A(n_303),
.B(n_252),
.Y(n_327)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_327),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_328),
.B(n_310),
.C(n_314),
.Y(n_350)
);

NOR3xp33_ASAP7_75t_SL g329 ( 
.A(n_285),
.B(n_259),
.C(n_250),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_329),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_297),
.B(n_282),
.Y(n_330)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_330),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_315),
.B(n_280),
.Y(n_332)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_332),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_289),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_333),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_298),
.A2(n_269),
.B1(n_278),
.B2(n_277),
.Y(n_335)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_335),
.Y(n_356)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_337),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_288),
.B(n_273),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_339),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_298),
.A2(n_274),
.B1(n_216),
.B2(n_217),
.Y(n_340)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_340),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_307),
.A2(n_192),
.B(n_216),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g370 ( 
.A1(n_341),
.A2(n_345),
.B(n_321),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_299),
.B(n_171),
.Y(n_342)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_342),
.Y(n_373)
);

MAJx2_ASAP7_75t_L g343 ( 
.A(n_292),
.B(n_313),
.C(n_309),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_343),
.B(n_347),
.Y(n_375)
);

NAND3xp33_ASAP7_75t_L g344 ( 
.A(n_299),
.B(n_0),
.C(n_2),
.Y(n_344)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_344),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_309),
.B(n_2),
.Y(n_345)
);

INVxp33_ASAP7_75t_L g346 ( 
.A(n_290),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_346),
.A2(n_349),
.B(n_304),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_286),
.B(n_312),
.Y(n_347)
);

OAI21x1_ASAP7_75t_SL g348 ( 
.A1(n_307),
.A2(n_192),
.B(n_217),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_348),
.A2(n_287),
.B(n_302),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_310),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_SL g381 ( 
.A(n_350),
.B(n_354),
.Y(n_381)
);

XNOR2x2_ASAP7_75t_L g354 ( 
.A(n_338),
.B(n_293),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_343),
.B(n_305),
.C(n_318),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_357),
.B(n_371),
.C(n_342),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_326),
.B(n_305),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_359),
.B(n_361),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_326),
.B(n_316),
.Y(n_361)
);

NOR2x1_ASAP7_75t_SL g362 ( 
.A(n_348),
.B(n_308),
.Y(n_362)
);

CKINVDCx14_ASAP7_75t_R g384 ( 
.A(n_362),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_363),
.B(n_377),
.Y(n_387)
);

OAI22xp33_ASAP7_75t_L g391 ( 
.A1(n_364),
.A2(n_333),
.B1(n_341),
.B2(n_337),
.Y(n_391)
);

XOR2x2_ASAP7_75t_L g366 ( 
.A(n_343),
.B(n_304),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_366),
.B(n_331),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_370),
.B(n_376),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_328),
.B(n_286),
.C(n_300),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_327),
.A2(n_302),
.B(n_300),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_328),
.B(n_296),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_367),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_378),
.B(n_390),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_382),
.B(n_399),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_368),
.B(n_322),
.Y(n_383)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_383),
.Y(n_411)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_376),
.Y(n_385)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_385),
.Y(n_414)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_374),
.Y(n_386)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_386),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_359),
.B(n_325),
.C(n_324),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_388),
.B(n_394),
.C(n_401),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_353),
.B(n_319),
.Y(n_389)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_389),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_358),
.A2(n_324),
.B1(n_327),
.B2(n_331),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g403 ( 
.A(n_391),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_392),
.B(n_354),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_356),
.A2(n_335),
.B1(n_340),
.B2(n_323),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_393),
.A2(n_396),
.B1(n_397),
.B2(n_400),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_361),
.B(n_321),
.C(n_332),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_358),
.B(n_334),
.Y(n_395)
);

INVxp67_ASAP7_75t_SL g412 ( 
.A(n_395),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_351),
.A2(n_329),
.B1(n_334),
.B2(n_320),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_356),
.A2(n_345),
.B1(n_336),
.B2(n_296),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_362),
.A2(n_360),
.B1(n_369),
.B2(n_355),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_398),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_371),
.B(n_294),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_360),
.A2(n_336),
.B1(n_294),
.B2(n_287),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_357),
.B(n_366),
.C(n_375),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_382),
.B(n_375),
.C(n_350),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_404),
.B(n_409),
.C(n_417),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_399),
.B(n_377),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_405),
.B(n_420),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g426 ( 
.A(n_406),
.B(n_381),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_379),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_408),
.B(n_418),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_380),
.B(n_372),
.C(n_373),
.Y(n_409)
);

BUFx5_ASAP7_75t_L g416 ( 
.A(n_384),
.Y(n_416)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_416),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_380),
.B(n_373),
.C(n_363),
.Y(n_417)
);

NOR3xp33_ASAP7_75t_SL g420 ( 
.A(n_381),
.B(n_365),
.C(n_370),
.Y(n_420)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_422),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_411),
.B(n_394),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_424),
.B(n_425),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_402),
.B(n_413),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_SL g449 ( 
.A(n_426),
.B(n_417),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_403),
.A2(n_393),
.B1(n_355),
.B2(n_397),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_427),
.A2(n_406),
.B1(n_387),
.B2(n_364),
.Y(n_439)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_415),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_428),
.B(n_433),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_410),
.A2(n_388),
.B1(n_400),
.B2(n_352),
.Y(n_429)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_429),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_407),
.B(n_416),
.Y(n_430)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_430),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_412),
.B(n_392),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_431),
.B(n_435),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_402),
.B(n_401),
.Y(n_433)
);

INVx1_ASAP7_75t_SL g434 ( 
.A(n_414),
.Y(n_434)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_434),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_403),
.B(n_352),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_419),
.Y(n_436)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_436),
.Y(n_448)
);

OR2x2_ASAP7_75t_L g437 ( 
.A(n_434),
.B(n_391),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_437),
.A2(n_446),
.B1(n_4),
.B2(n_5),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_439),
.B(n_449),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_SL g443 ( 
.A(n_423),
.B(n_409),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_443),
.B(n_430),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_427),
.A2(n_387),
.B1(n_420),
.B2(n_413),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_426),
.B(n_404),
.Y(n_450)
);

XNOR2x1_ASAP7_75t_L g457 ( 
.A(n_450),
.B(n_29),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_450),
.B(n_433),
.C(n_425),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_451),
.B(n_454),
.Y(n_463)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_452),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_440),
.B(n_432),
.Y(n_453)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_453),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_445),
.B(n_432),
.Y(n_454)
);

INVxp67_ASAP7_75t_SL g455 ( 
.A(n_441),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_455),
.B(n_444),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_L g456 ( 
.A1(n_448),
.A2(n_421),
.B(n_201),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_456),
.A2(n_447),
.B(n_439),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_457),
.B(n_446),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_441),
.B(n_29),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_458),
.B(n_459),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_442),
.B(n_4),
.C(n_6),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_460),
.B(n_461),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_437),
.B(n_6),
.Y(n_461)
);

AO21x1_ASAP7_75t_L g476 ( 
.A1(n_466),
.A2(n_468),
.B(n_7),
.Y(n_476)
);

OAI21x1_ASAP7_75t_L g468 ( 
.A1(n_455),
.A2(n_438),
.B(n_449),
.Y(n_468)
);

INVxp33_ASAP7_75t_L g472 ( 
.A(n_470),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_471),
.B(n_462),
.C(n_7),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_463),
.A2(n_462),
.B(n_457),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_473),
.B(n_476),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g479 ( 
.A(n_474),
.B(n_475),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_469),
.B(n_6),
.C(n_7),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_L g478 ( 
.A1(n_472),
.A2(n_467),
.B1(n_466),
.B2(n_464),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_478),
.A2(n_465),
.B(n_8),
.Y(n_480)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_480),
.A2(n_481),
.B(n_479),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_477),
.Y(n_481)
);

OAI21x1_ASAP7_75t_SL g483 ( 
.A1(n_482),
.A2(n_9),
.B(n_481),
.Y(n_483)
);

OR2x2_ASAP7_75t_L g484 ( 
.A(n_483),
.B(n_9),
.Y(n_484)
);


endmodule