module real_jpeg_2152_n_9 (n_59, n_5, n_4, n_8, n_0, n_57, n_1, n_2, n_56, n_60, n_61, n_6, n_7, n_55, n_3, n_58, n_62, n_9);

input n_59;
input n_5;
input n_4;
input n_8;
input n_0;
input n_57;
input n_1;
input n_2;
input n_56;
input n_60;
input n_61;
input n_6;
input n_7;
input n_55;
input n_3;
input n_58;
input n_62;

output n_9;

wire n_17;
wire n_43;
wire n_37;
wire n_21;
wire n_38;
wire n_35;
wire n_50;
wire n_33;
wire n_29;
wire n_49;
wire n_10;
wire n_31;
wire n_52;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_11;
wire n_14;
wire n_51;
wire n_47;
wire n_45;
wire n_25;
wire n_42;
wire n_22;
wire n_53;
wire n_18;
wire n_36;
wire n_39;
wire n_40;
wire n_41;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_27;
wire n_48;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_0),
.B(n_20),
.C(n_46),
.Y(n_19)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx4f_ASAP7_75t_SL g34 ( 
.A(n_1),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_2),
.B(n_29),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_3),
.A2(n_28),
.B(n_32),
.Y(n_27)
);

AO22x1_ASAP7_75t_L g22 ( 
.A1(n_4),
.A2(n_23),
.B1(n_26),
.B2(n_37),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_5),
.B(n_22),
.C(n_38),
.Y(n_21)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g10 ( 
.A1(n_8),
.A2(n_11),
.B1(n_12),
.B2(n_16),
.Y(n_10)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_17),
.Y(n_9)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_14),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_14),
.B(n_53),
.Y(n_52)
);

INVx8_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx6_ASAP7_75t_SL g40 ( 
.A(n_15),
.Y(n_40)
);

INVx4_ASAP7_75t_SL g45 ( 
.A(n_15),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_50),
.C(n_51),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_41),
.C(n_42),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_25),
.Y(n_23)
);

CKINVDCx6p67_ASAP7_75t_R g49 ( 
.A(n_25),
.Y(n_49)
);

NAND3xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_35),
.C(n_36),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_35),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_32),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_34),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_40),
.Y(n_38)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_48),
.Y(n_46)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_55),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_56),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_57),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_58),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_59),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_60),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_61),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_62),
.Y(n_53)
);


endmodule