module fake_jpeg_26588_n_250 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_250);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_250;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_19),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_29),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_31),
.Y(n_34)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_0),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_30),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_11),
.B(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

HAxp5_ASAP7_75t_SL g36 ( 
.A(n_32),
.B(n_11),
.CON(n_36),
.SN(n_36)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_36),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_29),
.A2(n_20),
.B1(n_13),
.B2(n_16),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_38),
.A2(n_31),
.B1(n_16),
.B2(n_21),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_44),
.A2(n_52),
.B1(n_46),
.B2(n_55),
.Y(n_73)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_53),
.Y(n_60)
);

AND2x2_ASAP7_75t_SL g48 ( 
.A(n_41),
.B(n_30),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_51),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_30),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_49),
.B(n_54),
.Y(n_68)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_39),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g52 ( 
.A1(n_34),
.A2(n_32),
.B1(n_27),
.B2(n_28),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_34),
.B(n_30),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_35),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_55),
.Y(n_63)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_56),
.Y(n_74)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_41),
.A2(n_30),
.B1(n_29),
.B2(n_25),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_58),
.A2(n_29),
.B1(n_25),
.B2(n_35),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_41),
.C(n_34),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_72),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_65),
.A2(n_56),
.B1(n_50),
.B2(n_57),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_47),
.A2(n_32),
.B1(n_27),
.B2(n_42),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_67),
.A2(n_73),
.B1(n_76),
.B2(n_39),
.Y(n_81)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_47),
.A2(n_36),
.B(n_30),
.C(n_28),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_69),
.A2(n_48),
.B(n_58),
.Y(n_79)
);

OAI32xp33_ASAP7_75t_L g71 ( 
.A1(n_49),
.A2(n_35),
.A3(n_31),
.B1(n_38),
.B2(n_20),
.Y(n_71)
);

AOI32xp33_ASAP7_75t_L g88 ( 
.A1(n_71),
.A2(n_45),
.A3(n_22),
.B1(n_24),
.B2(n_12),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_13),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_48),
.C(n_58),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_26),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_44),
.A2(n_39),
.B1(n_21),
.B2(n_40),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_63),
.A2(n_45),
.B1(n_40),
.B2(n_39),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_77),
.A2(n_62),
.B1(n_70),
.B2(n_40),
.Y(n_94)
);

INVxp33_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_78),
.B(n_80),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_79),
.A2(n_84),
.B(n_89),
.Y(n_111)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_81),
.B(n_86),
.Y(n_96)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_82),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_83),
.A2(n_85),
.B1(n_87),
.B2(n_91),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_60),
.A2(n_48),
.B(n_57),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_65),
.A2(n_48),
.B1(n_50),
.B2(n_56),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_74),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_73),
.A2(n_39),
.B1(n_51),
.B2(n_45),
.Y(n_87)
);

NAND2xp67_ASAP7_75t_SL g102 ( 
.A(n_88),
.B(n_89),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_61),
.A2(n_51),
.B(n_10),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_61),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_61),
.A2(n_63),
.B1(n_71),
.B2(n_76),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_74),
.Y(n_93)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_94),
.A2(n_22),
.B1(n_37),
.B2(n_23),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_80),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_95),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_91),
.A2(n_61),
.B(n_69),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_97),
.A2(n_102),
.B(n_113),
.Y(n_133)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_101),
.Y(n_117)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_68),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_85),
.B(n_72),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_106),
.Y(n_122)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_86),
.B(n_81),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_107),
.B(n_108),
.Y(n_135)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_90),
.B(n_68),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_109),
.B(n_24),
.Y(n_137)
);

BUFx24_ASAP7_75t_SL g110 ( 
.A(n_92),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_92),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_79),
.A2(n_69),
.B(n_75),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_114),
.B(n_126),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_113),
.B(n_64),
.C(n_84),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_115),
.B(n_120),
.C(n_134),
.Y(n_148)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_112),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_124),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_118),
.B(n_123),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_88),
.C(n_62),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_66),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_108),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_103),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_96),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_125),
.B(n_128),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_82),
.Y(n_126)
);

OAI21xp33_ASAP7_75t_L g127 ( 
.A1(n_97),
.A2(n_102),
.B(n_105),
.Y(n_127)
);

AOI21xp33_ASAP7_75t_L g153 ( 
.A1(n_127),
.A2(n_14),
.B(n_12),
.Y(n_153)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_100),
.B(n_82),
.Y(n_129)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_100),
.B(n_80),
.Y(n_130)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_130),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_98),
.B(n_93),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_131),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_101),
.A2(n_40),
.B1(n_66),
.B2(n_43),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_132),
.A2(n_137),
.B1(n_37),
.B2(n_33),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_111),
.B(n_24),
.C(n_43),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_99),
.B(n_24),
.C(n_26),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_136),
.B(n_139),
.C(n_140),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_138),
.A2(n_37),
.B1(n_22),
.B2(n_23),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_94),
.B(n_24),
.C(n_26),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_24),
.C(n_33),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_118),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_124),
.A2(n_23),
.B1(n_17),
.B2(n_15),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_142),
.A2(n_23),
.B1(n_17),
.B2(n_15),
.Y(n_175)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_144),
.Y(n_171)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_117),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_140),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_147),
.Y(n_167)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_135),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_SL g176 ( 
.A(n_153),
.B(n_156),
.C(n_160),
.Y(n_176)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_122),
.Y(n_154)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_154),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_115),
.B(n_33),
.C(n_37),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_163),
.C(n_134),
.Y(n_173)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_122),
.Y(n_159)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_159),
.Y(n_180)
);

AOI21xp33_ASAP7_75t_L g160 ( 
.A1(n_133),
.A2(n_14),
.B(n_12),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_136),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_161),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_162),
.A2(n_119),
.B1(n_116),
.B2(n_125),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_120),
.B(n_33),
.C(n_37),
.Y(n_163)
);

XOR2x2_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_133),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_165),
.A2(n_158),
.B(n_146),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_166),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_157),
.A2(n_119),
.B1(n_139),
.B2(n_128),
.Y(n_168)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_168),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_121),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_172),
.C(n_173),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_155),
.C(n_163),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_174),
.B(n_178),
.C(n_152),
.Y(n_192)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_175),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_149),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_177),
.B(n_182),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_37),
.C(n_17),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_164),
.A2(n_18),
.B1(n_17),
.B2(n_15),
.Y(n_181)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_181),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_145),
.B(n_6),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_176),
.A2(n_147),
.B1(n_150),
.B2(n_149),
.Y(n_188)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_188),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_169),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_151),
.Y(n_190)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_190),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_165),
.A2(n_143),
.B1(n_144),
.B2(n_154),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_191),
.A2(n_194),
.B(n_18),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_195),
.C(n_197),
.Y(n_207)
);

FAx1_ASAP7_75t_L g194 ( 
.A(n_171),
.B(n_159),
.CI(n_158),
.CON(n_194),
.SN(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_170),
.C(n_173),
.Y(n_195)
);

NAND3xp33_ASAP7_75t_L g196 ( 
.A(n_176),
.B(n_180),
.C(n_179),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_196),
.B(n_175),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_172),
.B(n_142),
.C(n_162),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_184),
.B(n_178),
.Y(n_198)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_198),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_199),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_169),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_200),
.B(n_203),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_202),
.A2(n_4),
.B(n_8),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_197),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_187),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_6),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_206),
.B(n_208),
.Y(n_215)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_14),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_192),
.B(n_18),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_209),
.B(n_186),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_4),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_4),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_207),
.B(n_186),
.C(n_189),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_211),
.B(n_217),
.Y(n_222)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_213),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_209),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_207),
.B(n_194),
.C(n_193),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_218),
.B(n_220),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_216),
.A2(n_201),
.B(n_204),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_221),
.A2(n_225),
.B(n_228),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_223),
.B(n_2),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_211),
.A2(n_205),
.B(n_208),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_199),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_227),
.B(n_229),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_4),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_2),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_219),
.C(n_213),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_230),
.B(n_232),
.C(n_235),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_2),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_236),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_226),
.A2(n_228),
.B(n_223),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_222),
.A2(n_2),
.B(n_3),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_3),
.Y(n_237)
);

BUFx24_ASAP7_75t_SL g240 ( 
.A(n_237),
.Y(n_240)
);

NOR2xp67_ASAP7_75t_L g238 ( 
.A(n_233),
.B(n_3),
.Y(n_238)
);

O2A1O1Ixp33_ASAP7_75t_SL g243 ( 
.A1(n_238),
.A2(n_5),
.B(n_7),
.C(n_9),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_234),
.B(n_5),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_239),
.B(n_7),
.Y(n_245)
);

OAI32xp33_ASAP7_75t_L g246 ( 
.A1(n_243),
.A2(n_244),
.A3(n_245),
.B1(n_240),
.B2(n_1),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_242),
.B(n_5),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_246),
.B(n_247),
.Y(n_248)
);

MAJx2_ASAP7_75t_L g247 ( 
.A(n_244),
.B(n_241),
.C(n_7),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_248),
.A2(n_7),
.B1(n_9),
.B2(n_0),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_9),
.Y(n_250)
);


endmodule