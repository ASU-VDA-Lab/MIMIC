module fake_jpeg_26860_n_60 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_60);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_60;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

INVx1_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

BUFx24_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g19 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_19),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_14),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_22),
.Y(n_26)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_11),
.B(n_1),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_23),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_9),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_28),
.B(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_31),
.Y(n_41)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_29),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_34),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_26),
.A2(n_20),
.B(n_19),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_25),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_28),
.B(n_10),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_18),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_32),
.B(n_7),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_40),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_32),
.B(n_7),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_39),
.A2(n_18),
.B(n_12),
.Y(n_43)
);

MAJx2_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_5),
.C(n_6),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_41),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_44),
.Y(n_48)
);

INVxp33_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_46),
.B(n_1),
.C(n_3),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_45),
.Y(n_51)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_47),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_53),
.Y(n_54)
);

AOI31xp67_ASAP7_75t_L g56 ( 
.A1(n_55),
.A2(n_50),
.A3(n_49),
.B(n_46),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_56),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_54),
.B(n_8),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_54),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_57),
.Y(n_60)
);


endmodule