module fake_netlist_1_5544_n_505 (n_20, n_12, n_56, n_47, n_52, n_67, n_50, n_7, n_1, n_60, n_16, n_22, n_3, n_19, n_10, n_34, n_40, n_68, n_25, n_30, n_36, n_9, n_13, n_75, n_53, n_26, n_11, n_64, n_72, n_69, n_39, n_43, n_73, n_62, n_38, n_23, n_0, n_33, n_4, n_59, n_24, n_35, n_6, n_32, n_8, n_15, n_74, n_57, n_61, n_51, n_44, n_71, n_66, n_70, n_46, n_45, n_42, n_21, n_2, n_37, n_48, n_27, n_63, n_18, n_17, n_54, n_28, n_41, n_58, n_65, n_55, n_49, n_5, n_29, n_14, n_31, n_505, n_449);
input n_20;
input n_12;
input n_56;
input n_47;
input n_52;
input n_67;
input n_50;
input n_7;
input n_1;
input n_60;
input n_16;
input n_22;
input n_3;
input n_19;
input n_10;
input n_34;
input n_40;
input n_68;
input n_25;
input n_30;
input n_36;
input n_9;
input n_13;
input n_75;
input n_53;
input n_26;
input n_11;
input n_64;
input n_72;
input n_69;
input n_39;
input n_43;
input n_73;
input n_62;
input n_38;
input n_23;
input n_0;
input n_33;
input n_4;
input n_59;
input n_24;
input n_35;
input n_6;
input n_32;
input n_8;
input n_15;
input n_74;
input n_57;
input n_61;
input n_51;
input n_44;
input n_71;
input n_66;
input n_70;
input n_46;
input n_45;
input n_42;
input n_21;
input n_2;
input n_37;
input n_48;
input n_27;
input n_63;
input n_18;
input n_17;
input n_54;
input n_28;
input n_41;
input n_58;
input n_65;
input n_55;
input n_49;
input n_5;
input n_29;
input n_14;
input n_31;
output n_505;
output n_449;
wire n_107;
wire n_156;
wire n_154;
wire n_239;
wire n_7;
wire n_309;
wire n_356;
wire n_327;
wire n_25;
wire n_204;
wire n_169;
wire n_384;
wire n_370;
wire n_439;
wire n_180;
wire n_99;
wire n_43;
wire n_73;
wire n_440;
wire n_199;
wire n_279;
wire n_357;
wire n_74;
wire n_308;
wire n_44;
wire n_394;
wire n_189;
wire n_226;
wire n_352;
wire n_447;
wire n_66;
wire n_379;
wire n_316;
wire n_285;
wire n_471;
wire n_47;
wire n_475;
wire n_281;
wire n_497;
wire n_399;
wire n_11;
wire n_295;
wire n_371;
wire n_368;
wire n_373;
wire n_139;
wire n_342;
wire n_151;
wire n_71;
wire n_288;
wire n_176;
wire n_436;
wire n_438;
wire n_359;
wire n_195;
wire n_300;
wire n_487;
wire n_461;
wire n_223;
wire n_405;
wire n_19;
wire n_409;
wire n_482;
wire n_261;
wire n_423;
wire n_483;
wire n_220;
wire n_353;
wire n_410;
wire n_104;
wire n_303;
wire n_502;
wire n_468;
wire n_159;
wire n_91;
wire n_301;
wire n_340;
wire n_148;
wire n_149;
wire n_378;
wire n_246;
wire n_191;
wire n_143;
wire n_446;
wire n_63;
wire n_402;
wire n_54;
wire n_387;
wire n_125;
wire n_145;
wire n_166;
wire n_492;
wire n_181;
wire n_123;
wire n_219;
wire n_343;
wire n_494;
wire n_135;
wire n_481;
wire n_315;
wire n_397;
wire n_53;
wire n_213;
wire n_196;
wire n_293;
wire n_127;
wire n_312;
wire n_424;
wire n_23;
wire n_110;
wire n_182;
wire n_269;
wire n_186;
wire n_137;
wire n_334;
wire n_164;
wire n_433;
wire n_120;
wire n_392;
wire n_155;
wire n_162;
wire n_114;
wire n_50;
wire n_3;
wire n_331;
wire n_330;
wire n_231;
wire n_9;
wire n_428;
wire n_178;
wire n_478;
wire n_229;
wire n_97;
wire n_133;
wire n_324;
wire n_442;
wire n_422;
wire n_192;
wire n_329;
wire n_6;
wire n_8;
wire n_187;
wire n_188;
wire n_443;
wire n_304;
wire n_18;
wire n_441;
wire n_425;
wire n_314;
wire n_307;
wire n_215;
wire n_172;
wire n_109;
wire n_332;
wire n_198;
wire n_386;
wire n_351;
wire n_1;
wire n_16;
wire n_95;
wire n_40;
wire n_210;
wire n_426;
wire n_228;
wire n_278;
wire n_115;
wire n_270;
wire n_476;
wire n_404;
wire n_289;
wire n_179;
wire n_366;
wire n_362;
wire n_485;
wire n_396;
wire n_354;
wire n_152;
wire n_70;
wire n_458;
wire n_375;
wire n_17;
wire n_322;
wire n_317;
wire n_221;
wire n_328;
wire n_491;
wire n_388;
wire n_266;
wire n_80;
wire n_326;
wire n_275;
wire n_493;
wire n_274;
wire n_150;
wire n_235;
wire n_38;
wire n_272;
wire n_299;
wire n_100;
wire n_280;
wire n_141;
wire n_160;
wire n_499;
wire n_377;
wire n_263;
wire n_193;
wire n_232;
wire n_344;
wire n_147;
wire n_185;
wire n_367;
wire n_267;
wire n_171;
wire n_450;
wire n_140;
wire n_111;
wire n_212;
wire n_30;
wire n_13;
wire n_254;
wire n_435;
wire n_64;
wire n_69;
wire n_248;
wire n_407;
wire n_83;
wire n_200;
wire n_262;
wire n_119;
wire n_503;
wire n_339;
wire n_347;
wire n_124;
wire n_79;
wire n_129;
wire n_157;
wire n_103;
wire n_421;
wire n_52;
wire n_253;
wire n_434;
wire n_273;
wire n_325;
wire n_163;
wire n_348;
wire n_96;
wire n_72;
wire n_77;
wire n_90;
wire n_214;
wire n_167;
wire n_364;
wire n_33;
wire n_464;
wire n_76;
wire n_470;
wire n_61;
wire n_463;
wire n_216;
wire n_153;
wire n_355;
wire n_121;
wire n_286;
wire n_408;
wire n_247;
wire n_431;
wire n_161;
wire n_224;
wire n_484;
wire n_165;
wire n_413;
wire n_65;
wire n_5;
wire n_496;
wire n_393;
wire n_211;
wire n_85;
wire n_320;
wire n_264;
wire n_102;
wire n_283;
wire n_290;
wire n_217;
wire n_201;
wire n_277;
wire n_259;
wire n_244;
wire n_276;
wire n_297;
wire n_225;
wire n_350;
wire n_208;
wire n_419;
wire n_252;
wire n_168;
wire n_271;
wire n_94;
wire n_194;
wire n_282;
wire n_58;
wire n_113;
wire n_242;
wire n_498;
wire n_501;
wire n_284;
wire n_321;
wire n_302;
wire n_116;
wire n_292;
wire n_118;
wire n_233;
wire n_257;
wire n_26;
wire n_203;
wire n_477;
wire n_460;
wire n_243;
wire n_318;
wire n_346;
wire n_98;
wire n_345;
wire n_230;
wire n_452;
wire n_337;
wire n_146;
wire n_32;
wire n_93;
wire n_406;
wire n_372;
wire n_467;
wire n_41;
wire n_417;
wire n_451;
wire n_445;
wire n_500;
wire n_10;
wire n_390;
wire n_75;
wire n_82;
wire n_183;
wire n_132;
wire n_170;
wire n_205;
wire n_158;
wire n_126;
wire n_473;
wire n_249;
wire n_389;
wire n_360;
wire n_363;
wire n_427;
wire n_106;
wire n_296;
wire n_42;
wire n_21;
wire n_437;
wire n_89;
wire n_480;
wire n_130;
wire n_310;
wire n_341;
wire n_14;
wire n_236;
wire n_136;
wire n_260;
wire n_222;
wire n_381;
wire n_34;
wire n_142;
wire n_385;
wire n_227;
wire n_395;
wire n_454;
wire n_453;
wire n_250;
wire n_268;
wire n_190;
wire n_62;
wire n_4;
wire n_59;
wire n_323;
wire n_376;
wire n_240;
wire n_459;
wire n_88;
wire n_46;
wire n_174;
wire n_108;
wire n_335;
wire n_37;
wire n_122;
wire n_374;
wire n_380;
wire n_87;
wire n_466;
wire n_349;
wire n_207;
wire n_197;
wire n_81;
wire n_298;
wire n_112;
wire n_78;
wire n_68;
wire n_444;
wire n_105;
wire n_251;
wire n_36;
wire n_416;
wire n_432;
wire n_465;
wire n_414;
wire n_369;
wire n_469;
wire n_361;
wire n_237;
wire n_15;
wire n_429;
wire n_256;
wire n_398;
wire n_117;
wire n_238;
wire n_365;
wire n_294;
wire n_2;
wire n_338;
wire n_391;
wire n_209;
wire n_241;
wire n_20;
wire n_84;
wire n_449;
wire n_12;
wire n_56;
wire n_412;
wire n_455;
wire n_67;
wire n_504;
wire n_456;
wire n_22;
wire n_479;
wire n_311;
wire n_383;
wire n_202;
wire n_319;
wire n_39;
wire n_101;
wire n_291;
wire n_489;
wire n_245;
wire n_486;
wire n_24;
wire n_35;
wire n_490;
wire n_472;
wire n_400;
wire n_457;
wire n_134;
wire n_48;
wire n_255;
wire n_55;
wire n_336;
wire n_29;
wire n_218;
wire n_173;
wire n_488;
wire n_382;
wire n_138;
wire n_60;
wire n_462;
wire n_474;
wire n_305;
wire n_495;
wire n_430;
wire n_418;
wire n_92;
wire n_313;
wire n_333;
wire n_358;
wire n_175;
wire n_128;
wire n_306;
wire n_415;
wire n_0;
wire n_258;
wire n_234;
wire n_184;
wire n_265;
wire n_57;
wire n_51;
wire n_411;
wire n_287;
wire n_144;
wire n_403;
wire n_45;
wire n_131;
wire n_420;
wire n_86;
wire n_27;
wire n_177;
wire n_28;
wire n_448;
wire n_49;
wire n_206;
wire n_31;
INVx1_ASAP7_75t_L g76 ( .A(n_30), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_65), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_54), .Y(n_78) );
CKINVDCx5p33_ASAP7_75t_R g79 ( .A(n_44), .Y(n_79) );
INVxp33_ASAP7_75t_L g80 ( .A(n_72), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_26), .Y(n_81) );
HB1xp67_ASAP7_75t_L g82 ( .A(n_3), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_69), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_68), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_74), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_62), .Y(n_86) );
INVxp67_ASAP7_75t_SL g87 ( .A(n_48), .Y(n_87) );
CKINVDCx16_ASAP7_75t_R g88 ( .A(n_11), .Y(n_88) );
OR2x2_ASAP7_75t_L g89 ( .A(n_50), .B(n_37), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_66), .Y(n_90) );
INVxp33_ASAP7_75t_L g91 ( .A(n_71), .Y(n_91) );
BUFx3_ASAP7_75t_L g92 ( .A(n_29), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_39), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_61), .Y(n_94) );
HB1xp67_ASAP7_75t_L g95 ( .A(n_75), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_45), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_20), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_73), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_8), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_70), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_3), .Y(n_101) );
CKINVDCx5p33_ASAP7_75t_R g102 ( .A(n_38), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_5), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_19), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_6), .Y(n_105) );
INVxp33_ASAP7_75t_SL g106 ( .A(n_58), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_13), .Y(n_107) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_10), .Y(n_108) );
BUFx3_ASAP7_75t_L g109 ( .A(n_41), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_31), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_35), .Y(n_111) );
INVxp67_ASAP7_75t_L g112 ( .A(n_34), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_76), .Y(n_113) );
OA21x2_ASAP7_75t_L g114 ( .A1(n_76), .A2(n_25), .B(n_64), .Y(n_114) );
NOR2xp33_ASAP7_75t_L g115 ( .A(n_95), .B(n_0), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_95), .B(n_0), .Y(n_116) );
AND2x2_ASAP7_75t_L g117 ( .A(n_82), .B(n_1), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_77), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_92), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_77), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_92), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_78), .Y(n_122) );
AND2x2_ASAP7_75t_L g123 ( .A(n_82), .B(n_1), .Y(n_123) );
INVxp67_ASAP7_75t_L g124 ( .A(n_108), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_78), .Y(n_125) );
AND2x6_ASAP7_75t_L g126 ( .A(n_92), .B(n_27), .Y(n_126) );
INVxp67_ASAP7_75t_L g127 ( .A(n_108), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_83), .Y(n_128) );
AND2x4_ASAP7_75t_L g129 ( .A(n_109), .B(n_2), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_83), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_97), .B(n_2), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_97), .B(n_4), .Y(n_132) );
AND2x2_ASAP7_75t_L g133 ( .A(n_80), .B(n_4), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_88), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g135 ( .A(n_80), .B(n_5), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_119), .Y(n_136) );
AND2x2_ASAP7_75t_L g137 ( .A(n_124), .B(n_91), .Y(n_137) );
AND2x4_ASAP7_75t_L g138 ( .A(n_129), .B(n_109), .Y(n_138) );
BUFx3_ASAP7_75t_L g139 ( .A(n_129), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_113), .B(n_91), .Y(n_140) );
AND2x4_ASAP7_75t_L g141 ( .A(n_129), .B(n_109), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_129), .Y(n_142) );
INVx3_ASAP7_75t_L g143 ( .A(n_129), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_119), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_119), .Y(n_145) );
INVx2_ASAP7_75t_L g146 ( .A(n_121), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_121), .Y(n_147) );
NAND3xp33_ASAP7_75t_L g148 ( .A(n_113), .B(n_98), .C(n_111), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_114), .Y(n_149) );
AND2x2_ASAP7_75t_L g150 ( .A(n_124), .B(n_88), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_121), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_118), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g153 ( .A(n_127), .B(n_118), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_120), .Y(n_154) );
BUFx3_ASAP7_75t_L g155 ( .A(n_126), .Y(n_155) );
AOI22xp33_ASAP7_75t_L g156 ( .A1(n_120), .A2(n_99), .B1(n_101), .B2(n_103), .Y(n_156) );
OR2x2_ASAP7_75t_L g157 ( .A(n_127), .B(n_117), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_114), .Y(n_158) );
HB1xp67_ASAP7_75t_L g159 ( .A(n_133), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_122), .B(n_112), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_143), .Y(n_161) );
AO22x1_ASAP7_75t_L g162 ( .A1(n_138), .A2(n_126), .B1(n_87), .B2(n_133), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_143), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_153), .B(n_133), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_157), .B(n_134), .Y(n_165) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_157), .B(n_116), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_143), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_143), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_136), .Y(n_169) );
AOI22xp33_ASAP7_75t_L g170 ( .A1(n_139), .A2(n_117), .B1(n_123), .B2(n_115), .Y(n_170) );
CKINVDCx5p33_ASAP7_75t_R g171 ( .A(n_150), .Y(n_171) );
BUFx4f_ASAP7_75t_L g172 ( .A(n_138), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_143), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_153), .B(n_117), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_140), .B(n_123), .Y(n_175) );
NAND2x2_ASAP7_75t_L g176 ( .A(n_157), .B(n_116), .Y(n_176) );
INVx5_ASAP7_75t_L g177 ( .A(n_138), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_139), .Y(n_178) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_155), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_139), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_139), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_142), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g183 ( .A(n_137), .B(n_123), .Y(n_183) );
INVx5_ASAP7_75t_L g184 ( .A(n_138), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_142), .Y(n_185) );
AND2x2_ASAP7_75t_L g186 ( .A(n_159), .B(n_137), .Y(n_186) );
BUFx3_ASAP7_75t_L g187 ( .A(n_155), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_140), .B(n_135), .Y(n_188) );
INVx4_ASAP7_75t_L g189 ( .A(n_138), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_137), .B(n_135), .Y(n_190) );
AND2x2_ASAP7_75t_L g191 ( .A(n_159), .B(n_115), .Y(n_191) );
CKINVDCx6p67_ASAP7_75t_R g192 ( .A(n_150), .Y(n_192) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_150), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_161), .Y(n_194) );
AOI221x1_ASAP7_75t_L g195 ( .A1(n_182), .A2(n_149), .B1(n_158), .B2(n_96), .C(n_94), .Y(n_195) );
OAI22xp5_ASAP7_75t_L g196 ( .A1(n_176), .A2(n_182), .B1(n_185), .B2(n_172), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_166), .B(n_160), .Y(n_197) );
OAI22x1_ASAP7_75t_L g198 ( .A1(n_171), .A2(n_138), .B1(n_141), .B2(n_158), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_161), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_163), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_163), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_167), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_192), .Y(n_203) );
INVx3_ASAP7_75t_L g204 ( .A(n_189), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_167), .A2(n_158), .B(n_141), .Y(n_205) );
AOI22xp33_ASAP7_75t_SL g206 ( .A1(n_176), .A2(n_160), .B1(n_141), .B2(n_107), .Y(n_206) );
OAI22xp5_ASAP7_75t_L g207 ( .A1(n_176), .A2(n_156), .B1(n_152), .B2(n_154), .Y(n_207) );
BUFx8_ASAP7_75t_L g208 ( .A(n_186), .Y(n_208) );
BUFx3_ASAP7_75t_L g209 ( .A(n_172), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_168), .Y(n_210) );
BUFx3_ASAP7_75t_L g211 ( .A(n_172), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_192), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_168), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_169), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_173), .Y(n_215) );
AO22x1_ASAP7_75t_L g216 ( .A1(n_177), .A2(n_141), .B1(n_126), .B2(n_87), .Y(n_216) );
OAI22xp5_ASAP7_75t_L g217 ( .A1(n_185), .A2(n_156), .B1(n_152), .B2(n_154), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_173), .Y(n_218) );
BUFx2_ASAP7_75t_L g219 ( .A(n_189), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g220 ( .A(n_165), .B(n_141), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_175), .B(n_141), .Y(n_221) );
BUFx6f_ASAP7_75t_L g222 ( .A(n_187), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_169), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_178), .Y(n_224) );
AND2x2_ASAP7_75t_L g225 ( .A(n_186), .B(n_122), .Y(n_225) );
OAI21x1_ASAP7_75t_L g226 ( .A1(n_195), .A2(n_158), .B(n_114), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_214), .Y(n_227) );
INVxp33_ASAP7_75t_SL g228 ( .A(n_203), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_214), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_214), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g231 ( .A(n_208), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_197), .B(n_183), .Y(n_232) );
AOI22xp33_ASAP7_75t_L g233 ( .A1(n_207), .A2(n_190), .B1(n_191), .B2(n_188), .Y(n_233) );
INVx3_ASAP7_75t_L g234 ( .A(n_222), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_223), .Y(n_235) );
INVx4_ASAP7_75t_L g236 ( .A(n_222), .Y(n_236) );
OAI22xp5_ASAP7_75t_L g237 ( .A1(n_196), .A2(n_170), .B1(n_125), .B2(n_130), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_221), .B(n_164), .Y(n_238) );
AO21x2_ASAP7_75t_L g239 ( .A1(n_196), .A2(n_86), .B(n_90), .Y(n_239) );
OAI22xp5_ASAP7_75t_L g240 ( .A1(n_206), .A2(n_125), .B1(n_130), .B2(n_128), .Y(n_240) );
AND2x2_ASAP7_75t_SL g241 ( .A(n_208), .B(n_189), .Y(n_241) );
AND2x4_ASAP7_75t_L g242 ( .A(n_209), .B(n_189), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_220), .B(n_193), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_223), .Y(n_244) );
OAI22xp5_ASAP7_75t_L g245 ( .A1(n_217), .A2(n_128), .B1(n_177), .B2(n_184), .Y(n_245) );
OAI22xp33_ASAP7_75t_L g246 ( .A1(n_207), .A2(n_131), .B1(n_132), .B2(n_174), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g247 ( .A1(n_225), .A2(n_191), .B1(n_184), .B2(n_177), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_223), .Y(n_248) );
CKINVDCx5p33_ASAP7_75t_R g249 ( .A(n_208), .Y(n_249) );
AOI22xp33_ASAP7_75t_L g250 ( .A1(n_225), .A2(n_177), .B1(n_184), .B2(n_148), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_224), .Y(n_251) );
OAI22xp5_ASAP7_75t_L g252 ( .A1(n_217), .A2(n_184), .B1(n_177), .B2(n_148), .Y(n_252) );
AND2x2_ASAP7_75t_L g253 ( .A(n_241), .B(n_224), .Y(n_253) );
OR2x2_ASAP7_75t_L g254 ( .A(n_251), .B(n_224), .Y(n_254) );
AND2x2_ASAP7_75t_SL g255 ( .A(n_241), .B(n_208), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_233), .B(n_194), .Y(n_256) );
AND2x2_ASAP7_75t_L g257 ( .A(n_241), .B(n_194), .Y(n_257) );
NAND4xp25_ASAP7_75t_L g258 ( .A(n_232), .B(n_132), .C(n_131), .D(n_103), .Y(n_258) );
OAI221xp5_ASAP7_75t_L g259 ( .A1(n_233), .A2(n_212), .B1(n_219), .B2(n_105), .C(n_104), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_251), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_238), .B(n_199), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g262 ( .A(n_243), .B(n_209), .Y(n_262) );
BUFx4f_ASAP7_75t_SL g263 ( .A(n_231), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_238), .B(n_232), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_227), .Y(n_265) );
OR2x2_ASAP7_75t_L g266 ( .A(n_229), .B(n_198), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_229), .Y(n_267) );
AOI22xp33_ASAP7_75t_L g268 ( .A1(n_237), .A2(n_246), .B1(n_240), .B2(n_241), .Y(n_268) );
BUFx2_ASAP7_75t_L g269 ( .A(n_227), .Y(n_269) );
BUFx12f_ASAP7_75t_L g270 ( .A(n_249), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g271 ( .A1(n_243), .A2(n_219), .B1(n_198), .B2(n_211), .Y(n_271) );
INVx4_ASAP7_75t_L g272 ( .A(n_236), .Y(n_272) );
OR2x2_ASAP7_75t_L g273 ( .A(n_248), .B(n_199), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_248), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_260), .Y(n_275) );
INVx2_ASAP7_75t_SL g276 ( .A(n_255), .Y(n_276) );
AOI222xp33_ASAP7_75t_L g277 ( .A1(n_264), .A2(n_237), .B1(n_240), .B2(n_246), .C1(n_231), .C2(n_104), .Y(n_277) );
OR2x2_ASAP7_75t_L g278 ( .A(n_264), .B(n_239), .Y(n_278) );
OAI22xp5_ASAP7_75t_L g279 ( .A1(n_268), .A2(n_255), .B1(n_259), .B2(n_261), .Y(n_279) );
OAI22xp5_ASAP7_75t_L g280 ( .A1(n_268), .A2(n_245), .B1(n_247), .B2(n_235), .Y(n_280) );
OAI321xp33_ASAP7_75t_L g281 ( .A1(n_258), .A2(n_245), .A3(n_252), .B1(n_89), .B2(n_247), .C(n_99), .Y(n_281) );
OAI221xp5_ASAP7_75t_SL g282 ( .A1(n_258), .A2(n_101), .B1(n_105), .B2(n_250), .C(n_110), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_260), .B(n_227), .Y(n_283) );
OR2x6_ASAP7_75t_L g284 ( .A(n_272), .B(n_236), .Y(n_284) );
OAI321xp33_ASAP7_75t_L g285 ( .A1(n_259), .A2(n_252), .A3(n_89), .B1(n_112), .B2(n_250), .C(n_96), .Y(n_285) );
NAND4xp25_ASAP7_75t_L g286 ( .A(n_271), .B(n_98), .C(n_94), .D(n_111), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_263), .B(n_228), .Y(n_287) );
OR2x6_ASAP7_75t_L g288 ( .A(n_272), .B(n_236), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_267), .B(n_230), .Y(n_289) );
BUFx2_ASAP7_75t_L g290 ( .A(n_269), .Y(n_290) );
INVx2_ASAP7_75t_SL g291 ( .A(n_255), .Y(n_291) );
AND2x2_ASAP7_75t_SL g292 ( .A(n_272), .B(n_236), .Y(n_292) );
OAI221xp5_ASAP7_75t_SL g293 ( .A1(n_261), .A2(n_85), .B1(n_86), .B2(n_90), .C(n_110), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_267), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_274), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_274), .B(n_230), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_275), .Y(n_297) );
AND2x2_ASAP7_75t_L g298 ( .A(n_283), .B(n_269), .Y(n_298) );
OAI22xp5_ASAP7_75t_L g299 ( .A1(n_282), .A2(n_257), .B1(n_253), .B2(n_254), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_294), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_295), .B(n_254), .Y(n_301) );
OAI21xp33_ASAP7_75t_L g302 ( .A1(n_286), .A2(n_85), .B(n_89), .Y(n_302) );
NAND3xp33_ASAP7_75t_L g303 ( .A(n_277), .B(n_272), .C(n_262), .Y(n_303) );
OAI33xp33_ASAP7_75t_L g304 ( .A1(n_279), .A2(n_256), .A3(n_266), .B1(n_273), .B2(n_144), .B3(n_147), .Y(n_304) );
INVx1_ASAP7_75t_SL g305 ( .A(n_287), .Y(n_305) );
BUFx2_ASAP7_75t_L g306 ( .A(n_290), .Y(n_306) );
AOI22xp33_ASAP7_75t_L g307 ( .A1(n_276), .A2(n_257), .B1(n_253), .B2(n_239), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_283), .Y(n_308) );
OAI22xp5_ASAP7_75t_L g309 ( .A1(n_293), .A2(n_257), .B1(n_253), .B2(n_256), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_289), .Y(n_310) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_290), .Y(n_311) );
AOI22xp5_ASAP7_75t_L g312 ( .A1(n_280), .A2(n_263), .B1(n_242), .B2(n_239), .Y(n_312) );
INVx2_ASAP7_75t_L g313 ( .A(n_289), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g314 ( .A1(n_276), .A2(n_273), .B1(n_266), .B2(n_265), .Y(n_314) );
OAI221xp5_ASAP7_75t_L g315 ( .A1(n_278), .A2(n_209), .B1(n_211), .B2(n_204), .C(n_265), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_296), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_296), .B(n_265), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_278), .Y(n_318) );
AND4x1_ASAP7_75t_L g319 ( .A(n_281), .B(n_270), .C(n_7), .D(n_8), .Y(n_319) );
AOI211xp5_ASAP7_75t_L g320 ( .A1(n_285), .A2(n_162), .B(n_216), .C(n_242), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_292), .B(n_239), .Y(n_321) );
OR2x2_ASAP7_75t_L g322 ( .A(n_284), .B(n_239), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_292), .Y(n_323) );
OR2x2_ASAP7_75t_L g324 ( .A(n_284), .B(n_230), .Y(n_324) );
INVx1_ASAP7_75t_SL g325 ( .A(n_305), .Y(n_325) );
AOI331xp33_ASAP7_75t_L g326 ( .A1(n_307), .A2(n_6), .A3(n_7), .B1(n_9), .B2(n_10), .B3(n_11), .C1(n_12), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_297), .Y(n_327) );
INVx1_ASAP7_75t_SL g328 ( .A(n_298), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_297), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_318), .B(n_284), .Y(n_330) );
INVx2_ASAP7_75t_SL g331 ( .A(n_324), .Y(n_331) );
NAND4xp25_ASAP7_75t_L g332 ( .A(n_312), .B(n_106), .C(n_195), .D(n_242), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_308), .B(n_291), .Y(n_333) );
NAND5xp2_ASAP7_75t_L g334 ( .A(n_320), .B(n_291), .C(n_270), .D(n_205), .E(n_288), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_319), .B(n_270), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_318), .B(n_288), .Y(n_336) );
INVx3_ASAP7_75t_L g337 ( .A(n_324), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_313), .B(n_288), .Y(n_338) );
OR2x2_ASAP7_75t_L g339 ( .A(n_306), .B(n_288), .Y(n_339) );
A2O1A1Ixp33_ASAP7_75t_L g340 ( .A1(n_302), .A2(n_244), .B(n_235), .C(n_242), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_310), .B(n_244), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_303), .B(n_9), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_300), .Y(n_343) );
AOI221xp5_ASAP7_75t_L g344 ( .A1(n_304), .A2(n_162), .B1(n_216), .B2(n_242), .C(n_79), .Y(n_344) );
AND2x4_ASAP7_75t_L g345 ( .A(n_323), .B(n_236), .Y(n_345) );
OR2x2_ASAP7_75t_L g346 ( .A(n_306), .B(n_311), .Y(n_346) );
OR2x2_ASAP7_75t_L g347 ( .A(n_298), .B(n_244), .Y(n_347) );
NOR3xp33_ASAP7_75t_SL g348 ( .A(n_315), .B(n_81), .C(n_84), .Y(n_348) );
AND2x4_ASAP7_75t_L g349 ( .A(n_323), .B(n_234), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_313), .Y(n_350) );
OAI31xp33_ASAP7_75t_L g351 ( .A1(n_321), .A2(n_211), .A3(n_204), .B(n_144), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_316), .B(n_12), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_316), .B(n_114), .Y(n_353) );
AOI31xp33_ASAP7_75t_L g354 ( .A1(n_321), .A2(n_322), .A3(n_299), .B(n_314), .Y(n_354) );
OR2x2_ASAP7_75t_L g355 ( .A(n_322), .B(n_13), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_317), .Y(n_356) );
NOR3xp33_ASAP7_75t_L g357 ( .A(n_309), .B(n_204), .C(n_234), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_317), .B(n_114), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_301), .B(n_14), .Y(n_359) );
OA21x2_ASAP7_75t_L g360 ( .A1(n_312), .A2(n_226), .B(n_144), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_318), .B(n_234), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_297), .Y(n_362) );
NAND4xp25_ASAP7_75t_L g363 ( .A(n_312), .B(n_204), .C(n_151), .D(n_147), .Y(n_363) );
INVx4_ASAP7_75t_L g364 ( .A(n_324), .Y(n_364) );
INVx1_ASAP7_75t_SL g365 ( .A(n_305), .Y(n_365) );
INVx1_ASAP7_75t_SL g366 ( .A(n_325), .Y(n_366) );
INVx2_ASAP7_75t_SL g367 ( .A(n_339), .Y(n_367) );
AND2x4_ASAP7_75t_L g368 ( .A(n_337), .B(n_234), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_328), .B(n_14), .Y(n_369) );
A2O1A1Ixp33_ASAP7_75t_L g370 ( .A1(n_354), .A2(n_234), .B(n_226), .C(n_93), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_356), .B(n_15), .Y(n_371) );
NAND2x1_ASAP7_75t_L g372 ( .A(n_364), .B(n_126), .Y(n_372) );
OAI21xp5_ASAP7_75t_L g373 ( .A1(n_342), .A2(n_126), .B(n_226), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_356), .B(n_15), .Y(n_374) );
NAND4xp75_ASAP7_75t_L g375 ( .A(n_335), .B(n_16), .C(n_17), .D(n_18), .Y(n_375) );
OAI31xp33_ASAP7_75t_L g376 ( .A1(n_334), .A2(n_17), .A3(n_18), .B(n_19), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_343), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_365), .B(n_21), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_350), .B(n_21), .Y(n_379) );
OAI32xp33_ASAP7_75t_L g380 ( .A1(n_355), .A2(n_22), .A3(n_23), .B1(n_100), .B2(n_102), .Y(n_380) );
NAND2x1_ASAP7_75t_L g381 ( .A(n_364), .B(n_126), .Y(n_381) );
OR2x6_ASAP7_75t_L g382 ( .A(n_364), .B(n_149), .Y(n_382) );
OR2x2_ASAP7_75t_L g383 ( .A(n_346), .B(n_22), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_362), .Y(n_384) );
NOR2x1_ASAP7_75t_L g385 ( .A(n_355), .B(n_23), .Y(n_385) );
OAI32xp33_ASAP7_75t_L g386 ( .A1(n_339), .A2(n_145), .A3(n_151), .B1(n_146), .B2(n_136), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_327), .Y(n_387) );
NOR3xp33_ASAP7_75t_L g388 ( .A(n_359), .B(n_146), .C(n_136), .Y(n_388) );
NAND3xp33_ASAP7_75t_SL g389 ( .A(n_351), .B(n_145), .C(n_136), .Y(n_389) );
XNOR2xp5_ASAP7_75t_L g390 ( .A(n_330), .B(n_24), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_330), .B(n_28), .Y(n_391) );
OAI31xp33_ASAP7_75t_L g392 ( .A1(n_340), .A2(n_218), .A3(n_215), .B(n_213), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_336), .B(n_32), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_346), .B(n_33), .Y(n_394) );
OR2x2_ASAP7_75t_L g395 ( .A(n_331), .B(n_36), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_336), .B(n_40), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_327), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_337), .B(n_42), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_352), .B(n_43), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_337), .B(n_46), .Y(n_400) );
O2A1O1Ixp33_ASAP7_75t_L g401 ( .A1(n_332), .A2(n_200), .B(n_218), .C(n_215), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_338), .B(n_47), .Y(n_402) );
OR2x2_ASAP7_75t_L g403 ( .A(n_331), .B(n_347), .Y(n_403) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_347), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_329), .B(n_361), .Y(n_405) );
OAI31xp33_ASAP7_75t_L g406 ( .A1(n_363), .A2(n_202), .A3(n_201), .B(n_200), .Y(n_406) );
INVxp67_ASAP7_75t_L g407 ( .A(n_338), .Y(n_407) );
INVxp67_ASAP7_75t_L g408 ( .A(n_333), .Y(n_408) );
OR2x2_ASAP7_75t_L g409 ( .A(n_404), .B(n_360), .Y(n_409) );
OR2x2_ASAP7_75t_L g410 ( .A(n_403), .B(n_360), .Y(n_410) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_384), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_366), .B(n_345), .Y(n_412) );
NAND2xp33_ASAP7_75t_SL g413 ( .A(n_390), .B(n_348), .Y(n_413) );
INVx2_ASAP7_75t_SL g414 ( .A(n_382), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_408), .B(n_345), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_378), .B(n_349), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_370), .A2(n_357), .B1(n_341), .B2(n_349), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_387), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_397), .Y(n_419) );
INVx2_ASAP7_75t_SL g420 ( .A(n_382), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_407), .B(n_358), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_367), .B(n_358), .Y(n_422) );
NOR2x1_ASAP7_75t_SL g423 ( .A(n_382), .B(n_353), .Y(n_423) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_370), .A2(n_326), .B1(n_344), .B2(n_353), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_367), .B(n_49), .Y(n_425) );
AOI21xp33_ASAP7_75t_SL g426 ( .A1(n_378), .A2(n_51), .B(n_52), .Y(n_426) );
OAI21xp33_ASAP7_75t_L g427 ( .A1(n_385), .A2(n_149), .B(n_213), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g428 ( .A1(n_375), .A2(n_126), .B1(n_210), .B2(n_202), .Y(n_428) );
XOR2x2_ASAP7_75t_L g429 ( .A(n_383), .B(n_53), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_368), .B(n_55), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_379), .Y(n_431) );
OAI21xp33_ASAP7_75t_SL g432 ( .A1(n_382), .A2(n_201), .B(n_210), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_379), .Y(n_433) );
NOR2xp33_ASAP7_75t_SL g434 ( .A(n_406), .B(n_126), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_371), .B(n_56), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_374), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_368), .B(n_57), .Y(n_437) );
NOR2x1_ASAP7_75t_SL g438 ( .A(n_394), .B(n_184), .Y(n_438) );
INVx1_ASAP7_75t_SL g439 ( .A(n_402), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_369), .Y(n_440) );
XNOR2x1_ASAP7_75t_L g441 ( .A(n_391), .B(n_59), .Y(n_441) );
INVx3_ASAP7_75t_L g442 ( .A(n_368), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_391), .B(n_60), .Y(n_443) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_380), .B(n_399), .Y(n_444) );
AOI222xp33_ASAP7_75t_L g445 ( .A1(n_389), .A2(n_184), .B1(n_177), .B2(n_178), .C1(n_181), .C2(n_180), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_393), .B(n_63), .Y(n_446) );
NAND3xp33_ASAP7_75t_L g447 ( .A(n_376), .B(n_222), .C(n_180), .Y(n_447) );
OAI321xp33_ASAP7_75t_L g448 ( .A1(n_373), .A2(n_222), .A3(n_67), .B1(n_181), .B2(n_179), .C(n_155), .Y(n_448) );
UNKNOWN g449 ( );
INVx1_ASAP7_75t_SL g450 ( .A(n_402), .Y(n_450) );
INVx1_ASAP7_75t_SL g451 ( .A(n_393), .Y(n_451) );
AOI211xp5_ASAP7_75t_L g452 ( .A1(n_392), .A2(n_222), .B(n_155), .C(n_179), .Y(n_452) );
AOI221xp5_ASAP7_75t_L g453 ( .A1(n_388), .A2(n_399), .B1(n_396), .B2(n_398), .C(n_400), .Y(n_453) );
AOI221xp5_ASAP7_75t_L g454 ( .A1(n_396), .A2(n_179), .B1(n_187), .B2(n_222), .C(n_400), .Y(n_454) );
INVx2_ASAP7_75t_SL g455 ( .A(n_395), .Y(n_455) );
OAI211xp5_ASAP7_75t_SL g456 ( .A1(n_372), .A2(n_179), .B(n_187), .C(n_381), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_386), .Y(n_457) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_404), .Y(n_458) );
INVx1_ASAP7_75t_SL g459 ( .A(n_366), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g460 ( .A1(n_376), .A2(n_334), .B1(n_357), .B2(n_342), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_377), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_404), .B(n_403), .Y(n_462) );
INVx1_ASAP7_75t_SL g463 ( .A(n_366), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_404), .B(n_405), .Y(n_464) );
XNOR2x1_ASAP7_75t_L g465 ( .A(n_390), .B(n_325), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_461), .B(n_458), .Y(n_466) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_458), .Y(n_467) );
NAND4xp25_ASAP7_75t_L g468 ( .A(n_460), .B(n_444), .C(n_413), .D(n_453), .Y(n_468) );
XOR2xp5_ASAP7_75t_L g469 ( .A(n_465), .B(n_441), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_464), .Y(n_470) );
XNOR2xp5_ASAP7_75t_L g471 ( .A(n_465), .B(n_429), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_462), .B(n_422), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_411), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_423), .A2(n_432), .B(n_441), .Y(n_474) );
NAND2x1p5_ASAP7_75t_L g475 ( .A(n_420), .B(n_414), .Y(n_475) );
OAI211xp5_ASAP7_75t_SL g476 ( .A1(n_460), .A2(n_440), .B(n_463), .C(n_459), .Y(n_476) );
AOI31xp33_ASAP7_75t_L g477 ( .A1(n_444), .A2(n_413), .A3(n_417), .B(n_420), .Y(n_477) );
INVxp67_ASAP7_75t_L g478 ( .A(n_412), .Y(n_478) );
OAI211xp5_ASAP7_75t_SL g479 ( .A1(n_436), .A2(n_427), .B(n_416), .C(n_428), .Y(n_479) );
XNOR2xp5_ASAP7_75t_L g480 ( .A(n_429), .B(n_451), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_416), .A2(n_415), .B1(n_414), .B2(n_412), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_410), .B(n_409), .Y(n_482) );
AOI211xp5_ASAP7_75t_L g483 ( .A1(n_468), .A2(n_424), .B(n_426), .C(n_447), .Y(n_483) );
OAI211xp5_ASAP7_75t_L g484 ( .A1(n_474), .A2(n_452), .B(n_415), .C(n_445), .Y(n_484) );
NAND3xp33_ASAP7_75t_L g485 ( .A(n_477), .B(n_434), .C(n_457), .Y(n_485) );
AOI211xp5_ASAP7_75t_L g486 ( .A1(n_476), .A2(n_456), .B(n_439), .C(n_450), .Y(n_486) );
AOI211xp5_ASAP7_75t_SL g487 ( .A1(n_477), .A2(n_448), .B(n_446), .C(n_443), .Y(n_487) );
AO22x1_ASAP7_75t_L g488 ( .A1(n_467), .A2(n_425), .B1(n_437), .B2(n_430), .Y(n_488) );
OAI22xp5_ASAP7_75t_SL g489 ( .A1(n_469), .A2(n_455), .B1(n_438), .B2(n_442), .Y(n_489) );
AOI21xp5_ASAP7_75t_SL g490 ( .A1(n_471), .A2(n_425), .B(n_454), .Y(n_490) );
AOI222xp33_ASAP7_75t_L g491 ( .A1(n_480), .A2(n_433), .B1(n_431), .B2(n_421), .C1(n_419), .C2(n_418), .Y(n_491) );
OAI211xp5_ASAP7_75t_L g492 ( .A1(n_483), .A2(n_485), .B(n_484), .C(n_490), .Y(n_492) );
AOI22xp33_ASAP7_75t_SL g493 ( .A1(n_489), .A2(n_475), .B1(n_470), .B2(n_478), .Y(n_493) );
AOI22xp5_ASAP7_75t_L g494 ( .A1(n_491), .A2(n_481), .B1(n_479), .B2(n_475), .Y(n_494) );
NOR3x1_ASAP7_75t_SL g495 ( .A(n_487), .B(n_449), .C(n_411), .Y(n_495) );
O2A1O1Ixp33_ASAP7_75t_L g496 ( .A1(n_486), .A2(n_466), .B(n_482), .C(n_435), .Y(n_496) );
XNOR2xp5_ASAP7_75t_L g497 ( .A(n_492), .B(n_494), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_495), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_493), .A2(n_472), .B1(n_466), .B2(n_473), .Y(n_499) );
INVx2_ASAP7_75t_L g500 ( .A(n_497), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_499), .Y(n_501) );
XNOR2xp5_ASAP7_75t_L g502 ( .A(n_500), .B(n_498), .Y(n_502) );
NOR3xp33_ASAP7_75t_SL g503 ( .A(n_502), .B(n_501), .C(n_500), .Y(n_503) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_503), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g505 ( .A1(n_504), .A2(n_496), .B(n_488), .Y(n_505) );
endmodule