module fake_jpeg_24689_n_301 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_301);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_301;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_288;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_125;
wire n_80;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_41),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

BUFx24_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_39),
.Y(n_48)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

AND2x2_ASAP7_75t_SL g42 ( 
.A(n_18),
.B(n_1),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_1),
.Y(n_47)
);

INVx3_ASAP7_75t_SL g43 ( 
.A(n_20),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_43),
.A2(n_22),
.B1(n_18),
.B2(n_30),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_44),
.Y(n_46)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_47),
.B(n_48),
.Y(n_100)
);

OA22x2_ASAP7_75t_L g103 ( 
.A1(n_50),
.A2(n_40),
.B1(n_39),
.B2(n_38),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_26),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_51),
.B(n_19),
.C(n_21),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_45),
.A2(n_18),
.B1(n_22),
.B2(n_30),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_53),
.A2(n_55),
.B1(n_56),
.B2(n_70),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_1),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_54),
.A2(n_59),
.B(n_57),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_45),
.A2(n_18),
.B1(n_30),
.B2(n_31),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_45),
.A2(n_31),
.B1(n_27),
.B2(n_23),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_31),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_59),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_27),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_64),
.Y(n_80)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_61),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_42),
.A2(n_35),
.B1(n_34),
.B2(n_17),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_21),
.B1(n_19),
.B2(n_23),
.Y(n_75)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_63),
.Y(n_84)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_69),
.B(n_71),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_43),
.A2(n_27),
.B1(n_19),
.B2(n_21),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_36),
.B(n_28),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_51),
.B(n_29),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_74),
.B(n_79),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_75),
.A2(n_17),
.B1(n_34),
.B2(n_35),
.Y(n_111)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_77),
.B(n_78),
.Y(n_110)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_28),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_47),
.B(n_33),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_81),
.B(n_82),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_54),
.B(n_33),
.Y(n_82)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_83),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_52),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_86),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g109 ( 
.A1(n_87),
.A2(n_38),
.B(n_23),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_32),
.Y(n_88)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_97),
.Y(n_117)
);

AND2x2_ASAP7_75t_SL g90 ( 
.A(n_54),
.B(n_38),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_90),
.B(n_96),
.C(n_85),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_48),
.A2(n_36),
.B(n_37),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_92),
.A2(n_102),
.B(n_90),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_32),
.Y(n_94)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_49),
.B(n_63),
.Y(n_95)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_48),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_99),
.A2(n_103),
.B1(n_43),
.B2(n_58),
.Y(n_113)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_101),
.B(n_58),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_67),
.B(n_25),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_46),
.Y(n_116)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_49),
.Y(n_104)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_104),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_61),
.B(n_29),
.Y(n_106)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_106),
.Y(n_134)
);

AO21x1_ASAP7_75t_L g146 ( 
.A1(n_109),
.A2(n_103),
.B(n_76),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_111),
.B(n_98),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_113),
.A2(n_114),
.B1(n_126),
.B2(n_133),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_97),
.A2(n_85),
.B1(n_105),
.B2(n_92),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_115),
.A2(n_124),
.B(n_127),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_116),
.B(n_44),
.Y(n_166)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_121),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_100),
.C(n_87),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_100),
.A2(n_25),
.B(n_17),
.C(n_34),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_73),
.B(n_69),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_125),
.B(n_131),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_96),
.A2(n_43),
.B1(n_40),
.B2(n_37),
.Y(n_126)
);

O2A1O1Ixp33_ASAP7_75t_L g127 ( 
.A1(n_103),
.A2(n_40),
.B(n_43),
.C(n_44),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_40),
.Y(n_128)
);

XNOR2x1_ASAP7_75t_SL g142 ( 
.A(n_128),
.B(n_115),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_91),
.B(n_79),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_100),
.A2(n_67),
.B1(n_44),
.B2(n_25),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_91),
.B(n_35),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_135),
.B(n_76),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_137),
.B(n_144),
.C(n_129),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_110),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_138),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_125),
.B(n_75),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_143),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_142),
.A2(n_2),
.B(n_3),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_135),
.B(n_131),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_114),
.C(n_109),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_145),
.B(n_147),
.Y(n_175)
);

OAI21xp33_ASAP7_75t_SL g196 ( 
.A1(n_146),
.A2(n_16),
.B(n_3),
.Y(n_196)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_110),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_104),
.Y(n_148)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_148),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_128),
.A2(n_83),
.B1(n_103),
.B2(n_99),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_149),
.A2(n_152),
.B1(n_157),
.B2(n_151),
.Y(n_189)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_150),
.B(n_151),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_117),
.Y(n_151)
);

OAI22x1_ASAP7_75t_SL g152 ( 
.A1(n_128),
.A2(n_127),
.B1(n_124),
.B2(n_133),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_119),
.B(n_84),
.Y(n_153)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_153),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_117),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_154),
.B(n_155),
.Y(n_195)
);

BUFx5_ASAP7_75t_L g155 ( 
.A(n_120),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_132),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_127),
.A2(n_89),
.B1(n_101),
.B2(n_80),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_120),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_160),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_84),
.Y(n_159)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_159),
.Y(n_192)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_124),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_162),
.B(n_112),
.Y(n_167)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_126),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_163),
.B(n_165),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_112),
.B(n_107),
.Y(n_164)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_164),
.Y(n_177)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_111),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_108),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_167),
.B(n_193),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_144),
.B(n_132),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_169),
.B(n_180),
.C(n_186),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_136),
.A2(n_123),
.B1(n_108),
.B2(n_77),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_170),
.A2(n_182),
.B1(n_185),
.B2(n_173),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_152),
.A2(n_118),
.B1(n_123),
.B2(n_134),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_172),
.A2(n_182),
.B1(n_183),
.B2(n_157),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_174),
.B(n_4),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_129),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_176),
.B(n_165),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_166),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_155),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_179),
.B(n_189),
.Y(n_217)
);

AOI22x1_ASAP7_75t_L g182 ( 
.A1(n_146),
.A2(n_72),
.B1(n_78),
.B2(n_107),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_161),
.A2(n_130),
.B1(n_118),
.B2(n_134),
.Y(n_183)
);

AND2x4_ASAP7_75t_L g185 ( 
.A(n_146),
.B(n_72),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_185),
.A2(n_188),
.B(n_194),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_137),
.B(n_130),
.C(n_93),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_138),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_190),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_139),
.B(n_2),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_136),
.A2(n_93),
.B(n_3),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_196),
.B(n_2),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_197),
.A2(n_201),
.B1(n_209),
.B2(n_170),
.Y(n_222)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_191),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_198),
.B(n_200),
.Y(n_229)
);

BUFx4f_ASAP7_75t_SL g199 ( 
.A(n_182),
.Y(n_199)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_199),
.Y(n_230)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_175),
.Y(n_200)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_178),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_204),
.B(n_207),
.Y(n_233)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_205),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_185),
.A2(n_160),
.B1(n_163),
.B2(n_145),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_195),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_210),
.A2(n_216),
.B1(n_219),
.B2(n_5),
.Y(n_237)
);

A2O1A1O1Ixp25_ASAP7_75t_L g211 ( 
.A1(n_185),
.A2(n_156),
.B(n_161),
.C(n_154),
.D(n_139),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_211),
.B(n_6),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_212),
.B(n_221),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_169),
.B(n_147),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_186),
.C(n_180),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_171),
.B(n_150),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_214),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_168),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_215),
.Y(n_224)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_171),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_187),
.B(n_162),
.Y(n_218)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_218),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_177),
.B(n_140),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_172),
.B(n_140),
.Y(n_220)
);

AOI321xp33_ASAP7_75t_L g231 ( 
.A1(n_220),
.A2(n_188),
.A3(n_184),
.B1(n_177),
.B2(n_181),
.C(n_192),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_222),
.A2(n_236),
.B(n_203),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_220),
.A2(n_173),
.B1(n_183),
.B2(n_194),
.Y(n_225)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_225),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_226),
.B(n_228),
.C(n_232),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_202),
.B(n_176),
.C(n_174),
.Y(n_228)
);

XNOR2x1_ASAP7_75t_L g250 ( 
.A(n_231),
.B(n_207),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_202),
.B(n_158),
.C(n_179),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_4),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_234),
.B(n_238),
.C(n_239),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_214),
.A2(n_5),
.B(n_6),
.Y(n_236)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_237),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_212),
.B(n_5),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_217),
.A2(n_199),
.B1(n_208),
.B2(n_203),
.Y(n_241)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_241),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_199),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_242)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_242),
.Y(n_248)
);

XOR2x2_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_211),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_244),
.A2(n_257),
.B(n_233),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_224),
.B(n_200),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_249),
.B(n_253),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_250),
.A2(n_252),
.B1(n_239),
.B2(n_230),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_223),
.B(n_205),
.Y(n_251)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_251),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_204),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_209),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_256),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_235),
.B(n_206),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_210),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_201),
.C(n_221),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_258),
.B(n_226),
.C(n_228),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_259),
.B(n_262),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_263),
.C(n_266),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_247),
.B(n_229),
.C(n_227),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_244),
.Y(n_265)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_265),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_227),
.C(n_238),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_231),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_267),
.B(n_271),
.Y(n_272)
);

BUFx24_ASAP7_75t_SL g269 ( 
.A(n_245),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_257),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_243),
.A2(n_224),
.B1(n_234),
.B2(n_10),
.Y(n_270)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_270),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_246),
.B(n_8),
.C(n_9),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_264),
.A2(n_255),
.B1(n_252),
.B2(n_251),
.Y(n_273)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_273),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_261),
.B(n_253),
.Y(n_276)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_276),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_268),
.B(n_248),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_280),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_254),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_281),
.A2(n_16),
.B(n_13),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_260),
.A2(n_250),
.B1(n_254),
.B2(n_12),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_282),
.B(n_8),
.C(n_9),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_279),
.B(n_266),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_283),
.B(n_288),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_284),
.A2(n_285),
.B(n_275),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_12),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_290),
.B(n_292),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_287),
.B(n_273),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_276),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_293),
.A2(n_294),
.B1(n_272),
.B2(n_284),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_274),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_277),
.C(n_279),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_296),
.A2(n_14),
.B(n_295),
.Y(n_299)
);

AOI221xp5_ASAP7_75t_L g298 ( 
.A1(n_297),
.A2(n_283),
.B1(n_282),
.B2(n_15),
.C(n_14),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_298),
.B(n_299),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_296),
.Y(n_301)
);


endmodule