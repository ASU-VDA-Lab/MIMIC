module fake_aes_9012_n_682 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_682);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_682;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVxp33_ASAP7_75t_SL g79 ( .A(n_42), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_77), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_27), .Y(n_81) );
INVxp67_ASAP7_75t_SL g82 ( .A(n_53), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_16), .Y(n_83) );
HB1xp67_ASAP7_75t_L g84 ( .A(n_51), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_33), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_21), .Y(n_86) );
INVxp33_ASAP7_75t_L g87 ( .A(n_16), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_39), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_69), .Y(n_89) );
INVxp33_ASAP7_75t_SL g90 ( .A(n_76), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_55), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_45), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_25), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_65), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_20), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_75), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_62), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_58), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_64), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_63), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_78), .Y(n_101) );
HB1xp67_ASAP7_75t_L g102 ( .A(n_41), .Y(n_102) );
NOR2xp67_ASAP7_75t_L g103 ( .A(n_73), .B(n_74), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_29), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_28), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_2), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_66), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_46), .Y(n_108) );
INVx2_ASAP7_75t_L g109 ( .A(n_72), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_4), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_47), .Y(n_111) );
INVxp67_ASAP7_75t_SL g112 ( .A(n_3), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g113 ( .A(n_14), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_38), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_70), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_34), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_60), .Y(n_117) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_61), .Y(n_118) );
INVxp67_ASAP7_75t_SL g119 ( .A(n_50), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_31), .Y(n_120) );
INVxp67_ASAP7_75t_L g121 ( .A(n_11), .Y(n_121) );
INVxp67_ASAP7_75t_SL g122 ( .A(n_40), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_13), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_59), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_15), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_35), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_44), .Y(n_127) );
CKINVDCx16_ASAP7_75t_R g128 ( .A(n_17), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_84), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_102), .B(n_0), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_83), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_128), .B(n_0), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_108), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_118), .Y(n_134) );
AND2x2_ASAP7_75t_L g135 ( .A(n_87), .B(n_1), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_118), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g137 ( .A(n_113), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_125), .Y(n_138) );
HB1xp67_ASAP7_75t_L g139 ( .A(n_106), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_121), .B(n_1), .Y(n_140) );
BUFx2_ASAP7_75t_L g141 ( .A(n_106), .Y(n_141) );
CKINVDCx5p33_ASAP7_75t_R g142 ( .A(n_110), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_110), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_108), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_127), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_85), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g147 ( .A(n_123), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_109), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_86), .Y(n_149) );
INVx1_ASAP7_75t_SL g150 ( .A(n_115), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_86), .Y(n_151) );
CKINVDCx5p33_ASAP7_75t_R g152 ( .A(n_85), .Y(n_152) );
HB1xp67_ASAP7_75t_L g153 ( .A(n_112), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_88), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_96), .Y(n_155) );
INVx4_ASAP7_75t_L g156 ( .A(n_118), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_118), .Y(n_157) );
BUFx2_ASAP7_75t_L g158 ( .A(n_96), .Y(n_158) );
OA21x2_ASAP7_75t_L g159 ( .A1(n_88), .A2(n_23), .B(n_68), .Y(n_159) );
OAI22xp5_ASAP7_75t_L g160 ( .A1(n_79), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_160) );
CKINVDCx20_ASAP7_75t_R g161 ( .A(n_126), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_126), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_127), .Y(n_163) );
CKINVDCx20_ASAP7_75t_R g164 ( .A(n_89), .Y(n_164) );
AND2x2_ASAP7_75t_L g165 ( .A(n_89), .B(n_5), .Y(n_165) );
INVx4_ASAP7_75t_L g166 ( .A(n_118), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g167 ( .A(n_79), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_91), .Y(n_168) );
INVx6_ASAP7_75t_L g169 ( .A(n_90), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_109), .Y(n_170) );
CKINVDCx5p33_ASAP7_75t_R g171 ( .A(n_90), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_80), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_91), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_156), .Y(n_174) );
NAND2x1p5_ASAP7_75t_L g175 ( .A(n_165), .B(n_92), .Y(n_175) );
AOI22xp5_ASAP7_75t_L g176 ( .A1(n_167), .A2(n_82), .B1(n_122), .B2(n_119), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_156), .Y(n_177) );
AND2x4_ASAP7_75t_L g178 ( .A(n_129), .B(n_101), .Y(n_178) );
AND2x4_ASAP7_75t_L g179 ( .A(n_172), .B(n_101), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_165), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_151), .Y(n_181) );
INVx2_ASAP7_75t_SL g182 ( .A(n_158), .Y(n_182) );
INVx3_ASAP7_75t_L g183 ( .A(n_156), .Y(n_183) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_134), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_151), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_166), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_166), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_166), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_158), .B(n_81), .Y(n_189) );
AND2x4_ASAP7_75t_L g190 ( .A(n_172), .B(n_92), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_169), .B(n_124), .Y(n_191) );
BUFx2_ASAP7_75t_L g192 ( .A(n_141), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_133), .Y(n_193) );
CKINVDCx5p33_ASAP7_75t_R g194 ( .A(n_161), .Y(n_194) );
NAND3x1_ASAP7_75t_L g195 ( .A(n_132), .B(n_93), .C(n_94), .Y(n_195) );
AND2x4_ASAP7_75t_L g196 ( .A(n_141), .B(n_93), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_134), .Y(n_197) );
INVx4_ASAP7_75t_L g198 ( .A(n_159), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_169), .B(n_120), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_173), .Y(n_200) );
BUFx6f_ASAP7_75t_L g201 ( .A(n_134), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_173), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_133), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_146), .B(n_117), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_144), .Y(n_205) );
CKINVDCx5p33_ASAP7_75t_R g206 ( .A(n_146), .Y(n_206) );
INVxp67_ASAP7_75t_L g207 ( .A(n_139), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_144), .Y(n_208) );
BUFx4f_ASAP7_75t_L g209 ( .A(n_145), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_148), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_148), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_170), .Y(n_212) );
BUFx6f_ASAP7_75t_L g213 ( .A(n_134), .Y(n_213) );
INVx3_ASAP7_75t_L g214 ( .A(n_170), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_131), .Y(n_215) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_134), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_135), .B(n_94), .Y(n_217) );
BUFx3_ASAP7_75t_L g218 ( .A(n_169), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g219 ( .A(n_137), .Y(n_219) );
NAND2xp33_ASAP7_75t_L g220 ( .A(n_167), .B(n_95), .Y(n_220) );
HB1xp67_ASAP7_75t_L g221 ( .A(n_142), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_138), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_152), .B(n_116), .Y(n_223) );
INVx2_ASAP7_75t_SL g224 ( .A(n_169), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_136), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_149), .Y(n_226) );
BUFx3_ASAP7_75t_L g227 ( .A(n_152), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_154), .Y(n_228) );
INVxp67_ASAP7_75t_L g229 ( .A(n_142), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_136), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_163), .Y(n_231) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_155), .Y(n_232) );
BUFx2_ASAP7_75t_L g233 ( .A(n_143), .Y(n_233) );
BUFx6f_ASAP7_75t_L g234 ( .A(n_136), .Y(n_234) );
BUFx3_ASAP7_75t_L g235 ( .A(n_155), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_136), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_168), .B(n_104), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_162), .B(n_114), .Y(n_238) );
BUFx3_ASAP7_75t_L g239 ( .A(n_162), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_209), .B(n_171), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_214), .Y(n_241) );
INVx2_ASAP7_75t_L g242 ( .A(n_214), .Y(n_242) );
AND2x2_ASAP7_75t_L g243 ( .A(n_192), .B(n_143), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_178), .B(n_171), .Y(n_244) );
BUFx4f_ASAP7_75t_L g245 ( .A(n_175), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_178), .B(n_135), .Y(n_246) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_198), .Y(n_247) );
AOI22xp33_ASAP7_75t_L g248 ( .A1(n_231), .A2(n_153), .B1(n_95), .B2(n_160), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_178), .B(n_130), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_193), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_193), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_238), .B(n_140), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_209), .B(n_107), .Y(n_253) );
NOR2xp33_ASAP7_75t_L g254 ( .A(n_189), .B(n_105), .Y(n_254) );
BUFx2_ASAP7_75t_L g255 ( .A(n_192), .Y(n_255) );
BUFx3_ASAP7_75t_L g256 ( .A(n_233), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_175), .Y(n_257) );
NAND2xp33_ASAP7_75t_SL g258 ( .A(n_206), .B(n_164), .Y(n_258) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_179), .A2(n_150), .B1(n_97), .B2(n_111), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_175), .Y(n_260) );
CKINVDCx5p33_ASAP7_75t_R g261 ( .A(n_219), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_214), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_203), .Y(n_263) );
HB1xp67_ASAP7_75t_L g264 ( .A(n_182), .Y(n_264) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_198), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_217), .B(n_100), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_205), .Y(n_267) );
INVx1_ASAP7_75t_SL g268 ( .A(n_233), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_224), .B(n_99), .Y(n_269) );
O2A1O1Ixp33_ASAP7_75t_L g270 ( .A1(n_180), .A2(n_98), .B(n_159), .C(n_103), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_224), .B(n_159), .Y(n_271) );
CKINVDCx20_ASAP7_75t_R g272 ( .A(n_219), .Y(n_272) );
INVx4_ASAP7_75t_L g273 ( .A(n_209), .Y(n_273) );
NOR3xp33_ASAP7_75t_SL g274 ( .A(n_206), .B(n_147), .C(n_6), .Y(n_274) );
BUFx2_ASAP7_75t_L g275 ( .A(n_227), .Y(n_275) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_182), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_217), .B(n_159), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_196), .B(n_157), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_196), .B(n_5), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_208), .Y(n_280) );
NOR3xp33_ASAP7_75t_L g281 ( .A(n_220), .B(n_6), .C(n_7), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_210), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_196), .B(n_157), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_211), .Y(n_284) );
NAND2xp5_ASAP7_75t_SL g285 ( .A(n_181), .B(n_157), .Y(n_285) );
INVx2_ASAP7_75t_SL g286 ( .A(n_227), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_212), .Y(n_287) );
NOR2xp33_ASAP7_75t_R g288 ( .A(n_232), .B(n_7), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g289 ( .A(n_191), .B(n_157), .Y(n_289) );
NOR2xp33_ASAP7_75t_L g290 ( .A(n_199), .B(n_157), .Y(n_290) );
BUFx6f_ASAP7_75t_L g291 ( .A(n_198), .Y(n_291) );
INVxp67_ASAP7_75t_SL g292 ( .A(n_207), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_231), .B(n_136), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_226), .B(n_8), .Y(n_294) );
CKINVDCx5p33_ASAP7_75t_R g295 ( .A(n_194), .Y(n_295) );
INVx5_ASAP7_75t_L g296 ( .A(n_183), .Y(n_296) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_174), .Y(n_297) );
NOR3xp33_ASAP7_75t_SL g298 ( .A(n_232), .B(n_8), .C(n_9), .Y(n_298) );
NOR3xp33_ASAP7_75t_L g299 ( .A(n_220), .B(n_9), .C(n_10), .Y(n_299) );
INVx1_ASAP7_75t_SL g300 ( .A(n_235), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_183), .Y(n_301) );
OR2x2_ASAP7_75t_L g302 ( .A(n_221), .B(n_194), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_228), .B(n_10), .Y(n_303) );
BUFx3_ASAP7_75t_L g304 ( .A(n_218), .Y(n_304) );
INVxp67_ASAP7_75t_L g305 ( .A(n_235), .Y(n_305) );
BUFx6f_ASAP7_75t_L g306 ( .A(n_174), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_215), .Y(n_307) );
CKINVDCx11_ASAP7_75t_R g308 ( .A(n_239), .Y(n_308) );
BUFx3_ASAP7_75t_L g309 ( .A(n_218), .Y(n_309) );
INVx4_ASAP7_75t_L g310 ( .A(n_183), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_252), .B(n_190), .Y(n_311) );
AND2x4_ASAP7_75t_L g312 ( .A(n_257), .B(n_239), .Y(n_312) );
CKINVDCx20_ASAP7_75t_R g313 ( .A(n_272), .Y(n_313) );
OAI21xp5_ASAP7_75t_L g314 ( .A1(n_271), .A2(n_195), .B(n_202), .Y(n_314) );
AOI22xp33_ASAP7_75t_L g315 ( .A1(n_279), .A2(n_179), .B1(n_190), .B2(n_204), .Y(n_315) );
BUFx2_ASAP7_75t_L g316 ( .A(n_256), .Y(n_316) );
BUFx2_ASAP7_75t_L g317 ( .A(n_255), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_244), .B(n_229), .Y(n_318) );
INVx1_ASAP7_75t_SL g319 ( .A(n_268), .Y(n_319) );
OAI22xp5_ASAP7_75t_L g320 ( .A1(n_245), .A2(n_179), .B1(n_190), .B2(n_176), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_260), .B(n_222), .Y(n_321) );
INVx5_ASAP7_75t_L g322 ( .A(n_247), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_245), .B(n_200), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_247), .Y(n_324) );
NOR2xp67_ASAP7_75t_SL g325 ( .A(n_273), .B(n_185), .Y(n_325) );
BUFx6f_ASAP7_75t_L g326 ( .A(n_247), .Y(n_326) );
BUFx8_ASAP7_75t_SL g327 ( .A(n_261), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_250), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_243), .B(n_237), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_247), .Y(n_330) );
INVx3_ASAP7_75t_L g331 ( .A(n_310), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_251), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_265), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_280), .Y(n_334) );
AOI22xp5_ASAP7_75t_L g335 ( .A1(n_252), .A2(n_195), .B1(n_223), .B2(n_187), .Y(n_335) );
BUFx6f_ASAP7_75t_L g336 ( .A(n_265), .Y(n_336) );
AOI222xp33_ASAP7_75t_L g337 ( .A1(n_258), .A2(n_177), .B1(n_186), .B2(n_187), .C1(n_188), .C2(n_15), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_265), .Y(n_338) );
INVx3_ASAP7_75t_L g339 ( .A(n_310), .Y(n_339) );
INVx3_ASAP7_75t_L g340 ( .A(n_296), .Y(n_340) );
INVx5_ASAP7_75t_L g341 ( .A(n_265), .Y(n_341) );
CKINVDCx11_ASAP7_75t_R g342 ( .A(n_308), .Y(n_342) );
CKINVDCx8_ASAP7_75t_R g343 ( .A(n_295), .Y(n_343) );
OAI22xp5_ASAP7_75t_L g344 ( .A1(n_249), .A2(n_188), .B1(n_186), .B2(n_177), .Y(n_344) );
CKINVDCx11_ASAP7_75t_R g345 ( .A(n_300), .Y(n_345) );
BUFx3_ASAP7_75t_L g346 ( .A(n_304), .Y(n_346) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_292), .B(n_11), .Y(n_347) );
CKINVDCx6p67_ASAP7_75t_R g348 ( .A(n_275), .Y(n_348) );
INVx3_ASAP7_75t_L g349 ( .A(n_296), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_282), .Y(n_350) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_264), .Y(n_351) );
BUFx6f_ASAP7_75t_L g352 ( .A(n_291), .Y(n_352) );
BUFx2_ASAP7_75t_L g353 ( .A(n_264), .Y(n_353) );
BUFx2_ASAP7_75t_R g354 ( .A(n_302), .Y(n_354) );
BUFx2_ASAP7_75t_L g355 ( .A(n_276), .Y(n_355) );
OAI21x1_ASAP7_75t_L g356 ( .A1(n_270), .A2(n_236), .B(n_197), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_287), .Y(n_357) );
OAI221xp5_ASAP7_75t_L g358 ( .A1(n_248), .A2(n_236), .B1(n_230), .B2(n_225), .C(n_197), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_246), .B(n_12), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_276), .B(n_307), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_281), .A2(n_230), .B1(n_225), .B2(n_234), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_254), .B(n_12), .Y(n_362) );
AND2x4_ASAP7_75t_L g363 ( .A(n_286), .B(n_13), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_291), .Y(n_364) );
OAI22xp5_ASAP7_75t_L g365 ( .A1(n_266), .A2(n_14), .B1(n_17), .B2(n_234), .Y(n_365) );
BUFx6f_ASAP7_75t_L g366 ( .A(n_326), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_329), .B(n_248), .Y(n_367) );
OAI22xp5_ASAP7_75t_L g368 ( .A1(n_311), .A2(n_305), .B1(n_273), .B2(n_259), .Y(n_368) );
BUFx2_ASAP7_75t_SL g369 ( .A(n_313), .Y(n_369) );
OAI22xp5_ASAP7_75t_L g370 ( .A1(n_353), .A2(n_263), .B1(n_267), .B2(n_284), .Y(n_370) );
AOI22xp5_ASAP7_75t_L g371 ( .A1(n_319), .A2(n_299), .B1(n_240), .B2(n_254), .Y(n_371) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_327), .Y(n_372) );
AOI22xp33_ASAP7_75t_SL g373 ( .A1(n_353), .A2(n_288), .B1(n_269), .B2(n_274), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_329), .B(n_240), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_321), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_360), .B(n_269), .Y(n_376) );
BUFx10_ASAP7_75t_L g377 ( .A(n_312), .Y(n_377) );
OAI22xp5_ASAP7_75t_L g378 ( .A1(n_355), .A2(n_277), .B1(n_283), .B2(n_278), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_360), .B(n_274), .Y(n_379) );
BUFx2_ASAP7_75t_L g380 ( .A(n_317), .Y(n_380) );
OAI22xp33_ASAP7_75t_L g381 ( .A1(n_317), .A2(n_303), .B1(n_294), .B2(n_288), .Y(n_381) );
BUFx2_ASAP7_75t_L g382 ( .A(n_316), .Y(n_382) );
O2A1O1Ixp5_ASAP7_75t_L g383 ( .A1(n_314), .A2(n_271), .B(n_253), .C(n_290), .Y(n_383) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_337), .A2(n_309), .B1(n_304), .B2(n_253), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_316), .B(n_241), .Y(n_385) );
CKINVDCx8_ASAP7_75t_R g386 ( .A(n_355), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_328), .A2(n_309), .B1(n_291), .B2(n_242), .Y(n_387) );
BUFx4f_ASAP7_75t_SL g388 ( .A(n_313), .Y(n_388) );
AOI22xp5_ASAP7_75t_L g389 ( .A1(n_318), .A2(n_298), .B1(n_301), .B2(n_291), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_328), .A2(n_262), .B1(n_306), .B2(n_297), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_321), .B(n_298), .Y(n_391) );
AOI22xp33_ASAP7_75t_SL g392 ( .A1(n_320), .A2(n_296), .B1(n_289), .B2(n_290), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_351), .Y(n_393) );
CKINVDCx20_ASAP7_75t_R g394 ( .A(n_345), .Y(n_394) );
NAND2xp5_ASAP7_75t_SL g395 ( .A(n_341), .B(n_306), .Y(n_395) );
NAND3xp33_ASAP7_75t_SL g396 ( .A(n_343), .B(n_315), .C(n_335), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_326), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_332), .A2(n_306), .B1(n_297), .B2(n_296), .Y(n_398) );
NAND2x1_ASAP7_75t_L g399 ( .A(n_325), .B(n_306), .Y(n_399) );
CKINVDCx8_ASAP7_75t_R g400 ( .A(n_342), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_396), .A2(n_363), .B1(n_347), .B2(n_362), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_366), .Y(n_402) );
AOI22xp33_ASAP7_75t_SL g403 ( .A1(n_388), .A2(n_363), .B1(n_312), .B2(n_354), .Y(n_403) );
BUFx3_ASAP7_75t_L g404 ( .A(n_377), .Y(n_404) );
OR2x2_ASAP7_75t_L g405 ( .A(n_375), .B(n_348), .Y(n_405) );
AOI22xp5_ASAP7_75t_L g406 ( .A1(n_367), .A2(n_335), .B1(n_363), .B2(n_359), .Y(n_406) );
OAI22xp33_ASAP7_75t_L g407 ( .A1(n_386), .A2(n_348), .B1(n_343), .B2(n_332), .Y(n_407) );
OAI21xp5_ASAP7_75t_L g408 ( .A1(n_383), .A2(n_356), .B(n_357), .Y(n_408) );
AO31x2_ASAP7_75t_L g409 ( .A1(n_378), .A2(n_365), .A3(n_364), .B(n_324), .Y(n_409) );
AO21x2_ASAP7_75t_L g410 ( .A1(n_389), .A2(n_356), .B(n_338), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_374), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_392), .A2(n_334), .B1(n_357), .B2(n_350), .Y(n_412) );
AOI222xp33_ASAP7_75t_L g413 ( .A1(n_388), .A2(n_379), .B1(n_391), .B2(n_376), .C1(n_380), .C2(n_393), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_373), .A2(n_312), .B1(n_323), .B2(n_350), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_369), .A2(n_323), .B1(n_334), .B2(n_349), .Y(n_415) );
OAI22xp33_ASAP7_75t_L g416 ( .A1(n_370), .A2(n_339), .B1(n_331), .B2(n_341), .Y(n_416) );
OAI21xp5_ASAP7_75t_L g417 ( .A1(n_371), .A2(n_361), .B(n_293), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_381), .B(n_322), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_368), .A2(n_340), .B1(n_349), .B2(n_346), .Y(n_419) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_382), .Y(n_420) );
BUFx6f_ASAP7_75t_SL g421 ( .A(n_400), .Y(n_421) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_385), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_397), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_377), .B(n_322), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_377), .B(n_341), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_397), .B(n_341), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_384), .B(n_322), .Y(n_427) );
AOI22xp33_ASAP7_75t_SL g428 ( .A1(n_394), .A2(n_341), .B1(n_322), .B2(n_349), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_395), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_384), .A2(n_340), .B1(n_346), .B2(n_331), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_402), .Y(n_431) );
INVx3_ASAP7_75t_L g432 ( .A(n_404), .Y(n_432) );
AOI21xp5_ASAP7_75t_L g433 ( .A1(n_412), .A2(n_395), .B(n_399), .Y(n_433) );
OAI33xp33_ASAP7_75t_L g434 ( .A1(n_407), .A2(n_344), .A3(n_372), .B1(n_285), .B2(n_364), .B3(n_324), .Y(n_434) );
BUFx2_ASAP7_75t_L g435 ( .A(n_429), .Y(n_435) );
NOR4xp25_ASAP7_75t_SL g436 ( .A(n_429), .B(n_394), .C(n_358), .D(n_285), .Y(n_436) );
AND2x6_ASAP7_75t_L g437 ( .A(n_406), .B(n_366), .Y(n_437) );
AO21x2_ASAP7_75t_L g438 ( .A1(n_408), .A2(n_338), .B(n_330), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_423), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_402), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_423), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_411), .B(n_341), .Y(n_442) );
NOR2x1_ASAP7_75t_L g443 ( .A(n_418), .B(n_404), .Y(n_443) );
OAI21x1_ASAP7_75t_L g444 ( .A1(n_408), .A2(n_390), .B(n_398), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_411), .Y(n_445) );
OAI22xp5_ASAP7_75t_L g446 ( .A1(n_406), .A2(n_390), .B1(n_387), .B2(n_398), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_410), .Y(n_447) );
OR2x6_ASAP7_75t_L g448 ( .A(n_427), .B(n_366), .Y(n_448) );
INVx3_ASAP7_75t_L g449 ( .A(n_404), .Y(n_449) );
INVx5_ASAP7_75t_L g450 ( .A(n_425), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_413), .B(n_322), .Y(n_451) );
INVx2_ASAP7_75t_SL g452 ( .A(n_425), .Y(n_452) );
AOI221xp5_ASAP7_75t_L g453 ( .A1(n_401), .A2(n_289), .B1(n_325), .B2(n_387), .C(n_340), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_410), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_410), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_413), .B(n_366), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_422), .B(n_326), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_409), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_426), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_426), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_409), .Y(n_461) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_403), .A2(n_339), .B1(n_331), .B2(n_330), .Y(n_462) );
NAND4xp25_ASAP7_75t_SL g463 ( .A(n_414), .B(n_333), .C(n_19), .D(n_22), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_409), .Y(n_464) );
NOR5xp2_ASAP7_75t_SL g465 ( .A(n_416), .B(n_18), .C(n_24), .D(n_26), .E(n_30), .Y(n_465) );
INVx3_ASAP7_75t_L g466 ( .A(n_409), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_441), .Y(n_467) );
AND2x4_ASAP7_75t_L g468 ( .A(n_448), .B(n_409), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_441), .B(n_420), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_441), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_459), .B(n_405), .Y(n_471) );
INVx4_ASAP7_75t_L g472 ( .A(n_432), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_439), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_445), .Y(n_474) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_457), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_459), .B(n_405), .Y(n_476) );
INVx1_ASAP7_75t_SL g477 ( .A(n_450), .Y(n_477) );
AOI221x1_ASAP7_75t_SL g478 ( .A1(n_445), .A2(n_421), .B1(n_424), .B2(n_415), .C(n_428), .Y(n_478) );
INVx4_ASAP7_75t_L g479 ( .A(n_432), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_435), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_435), .Y(n_481) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_457), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_460), .B(n_430), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_460), .B(n_419), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_456), .B(n_417), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_458), .Y(n_486) );
CKINVDCx5p33_ASAP7_75t_R g487 ( .A(n_450), .Y(n_487) );
OAI22xp33_ASAP7_75t_L g488 ( .A1(n_450), .A2(n_417), .B1(n_336), .B2(n_352), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_458), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_431), .B(n_352), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_458), .Y(n_491) );
INVx2_ASAP7_75t_SL g492 ( .A(n_432), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_461), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_431), .B(n_440), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_431), .Y(n_495) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_432), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_440), .B(n_352), .Y(n_497) );
AND2x4_ASAP7_75t_L g498 ( .A(n_448), .B(n_333), .Y(n_498) );
INVx1_ASAP7_75t_SL g499 ( .A(n_450), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_461), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_461), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_466), .B(n_352), .Y(n_502) );
INVx1_ASAP7_75t_SL g503 ( .A(n_450), .Y(n_503) );
BUFx2_ASAP7_75t_L g504 ( .A(n_437), .Y(n_504) );
INVx4_ASAP7_75t_L g505 ( .A(n_449), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_464), .Y(n_506) );
INVx4_ASAP7_75t_L g507 ( .A(n_449), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_464), .Y(n_508) );
BUFx2_ASAP7_75t_L g509 ( .A(n_437), .Y(n_509) );
INVx2_ASAP7_75t_L g510 ( .A(n_464), .Y(n_510) );
OA21x2_ASAP7_75t_L g511 ( .A1(n_447), .A2(n_352), .B(n_336), .Y(n_511) );
O2A1O1Ixp33_ASAP7_75t_L g512 ( .A1(n_434), .A2(n_339), .B(n_421), .C(n_297), .Y(n_512) );
OAI221xp5_ASAP7_75t_L g513 ( .A1(n_462), .A2(n_421), .B1(n_297), .B2(n_326), .C(n_336), .Y(n_513) );
INVxp67_ASAP7_75t_L g514 ( .A(n_449), .Y(n_514) );
INVx4_ASAP7_75t_L g515 ( .A(n_449), .Y(n_515) );
NAND3xp33_ASAP7_75t_L g516 ( .A(n_512), .B(n_443), .C(n_451), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_469), .B(n_450), .Y(n_517) );
INVx1_ASAP7_75t_SL g518 ( .A(n_487), .Y(n_518) );
INVx1_ASAP7_75t_SL g519 ( .A(n_487), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_467), .Y(n_520) );
NOR2xp33_ASAP7_75t_R g521 ( .A(n_477), .B(n_463), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_475), .B(n_452), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_473), .Y(n_523) );
NAND3xp33_ASAP7_75t_SL g524 ( .A(n_499), .B(n_436), .C(n_451), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_482), .B(n_450), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_471), .B(n_442), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_471), .B(n_476), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_472), .B(n_443), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_470), .B(n_448), .Y(n_529) );
NOR2x1_ASAP7_75t_L g530 ( .A(n_472), .B(n_463), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_474), .B(n_437), .Y(n_531) );
INVxp67_ASAP7_75t_L g532 ( .A(n_496), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_484), .B(n_437), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_503), .B(n_437), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_467), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_485), .B(n_437), .Y(n_536) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_495), .Y(n_537) );
NAND2xp33_ASAP7_75t_SL g538 ( .A(n_472), .B(n_436), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_483), .B(n_437), .Y(n_539) );
OA21x2_ASAP7_75t_L g540 ( .A1(n_486), .A2(n_447), .B(n_455), .Y(n_540) );
INVx2_ASAP7_75t_SL g541 ( .A(n_507), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_483), .B(n_437), .Y(n_542) );
NOR3xp33_ASAP7_75t_SL g543 ( .A(n_513), .B(n_446), .C(n_433), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_480), .Y(n_544) );
INVx2_ASAP7_75t_SL g545 ( .A(n_507), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_494), .B(n_466), .Y(n_546) );
NAND5xp2_ASAP7_75t_SL g547 ( .A(n_478), .B(n_453), .C(n_465), .D(n_433), .E(n_43), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_485), .B(n_448), .Y(n_548) );
INVxp67_ASAP7_75t_L g549 ( .A(n_481), .Y(n_549) );
NAND4xp25_ASAP7_75t_L g550 ( .A(n_468), .B(n_453), .C(n_466), .D(n_446), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_494), .B(n_466), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_495), .B(n_454), .Y(n_552) );
NOR2xp67_ASAP7_75t_SL g553 ( .A(n_507), .B(n_465), .Y(n_553) );
INVx1_ASAP7_75t_SL g554 ( .A(n_479), .Y(n_554) );
NOR2xp33_ASAP7_75t_SL g555 ( .A(n_479), .B(n_448), .Y(n_555) );
CKINVDCx5p33_ASAP7_75t_R g556 ( .A(n_479), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_481), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_486), .B(n_447), .Y(n_558) );
INVx2_ASAP7_75t_SL g559 ( .A(n_479), .Y(n_559) );
INVxp67_ASAP7_75t_L g560 ( .A(n_511), .Y(n_560) );
NOR2x1_ASAP7_75t_L g561 ( .A(n_505), .B(n_438), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_489), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_492), .B(n_444), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_527), .B(n_501), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_547), .A2(n_509), .B1(n_504), .B2(n_468), .Y(n_565) );
NAND2xp33_ASAP7_75t_R g566 ( .A(n_556), .B(n_465), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g567 ( .A1(n_530), .A2(n_504), .B1(n_509), .B2(n_514), .Y(n_567) );
AND2x2_ASAP7_75t_L g568 ( .A(n_517), .B(n_515), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_548), .B(n_515), .Y(n_569) );
AOI311xp33_ASAP7_75t_L g570 ( .A1(n_544), .A2(n_500), .A3(n_506), .B(n_491), .C(n_493), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_523), .Y(n_571) );
NAND4xp25_ASAP7_75t_L g572 ( .A(n_550), .B(n_468), .C(n_505), .D(n_515), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_525), .B(n_505), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_537), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_518), .B(n_515), .Y(n_575) );
INVxp67_ASAP7_75t_SL g576 ( .A(n_560), .Y(n_576) );
XNOR2xp5_ASAP7_75t_L g577 ( .A(n_526), .B(n_498), .Y(n_577) );
AOI21x1_ASAP7_75t_SL g578 ( .A1(n_531), .A2(n_468), .B(n_498), .Y(n_578) );
O2A1O1Ixp33_ASAP7_75t_L g579 ( .A1(n_524), .A2(n_488), .B(n_498), .C(n_502), .Y(n_579) );
OAI21xp5_ASAP7_75t_L g580 ( .A1(n_516), .A2(n_505), .B(n_502), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_557), .B(n_500), .Y(n_581) );
INVxp67_ASAP7_75t_L g582 ( .A(n_541), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_549), .B(n_506), .Y(n_583) );
NOR2xp33_ASAP7_75t_SL g584 ( .A(n_556), .B(n_498), .Y(n_584) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_538), .A2(n_511), .B(n_491), .Y(n_585) );
OAI31xp33_ASAP7_75t_L g586 ( .A1(n_538), .A2(n_510), .A3(n_508), .B(n_497), .Y(n_586) );
OAI22xp33_ASAP7_75t_SL g587 ( .A1(n_528), .A2(n_511), .B1(n_490), .B2(n_444), .Y(n_587) );
INVxp67_ASAP7_75t_L g588 ( .A(n_553), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_536), .B(n_438), .Y(n_589) );
INVx1_ASAP7_75t_SL g590 ( .A(n_519), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_520), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_520), .Y(n_592) );
OAI22xp33_ASAP7_75t_L g593 ( .A1(n_555), .A2(n_559), .B1(n_522), .B2(n_545), .Y(n_593) );
OAI322xp33_ASAP7_75t_L g594 ( .A1(n_549), .A2(n_234), .A3(n_201), .B1(n_213), .B2(n_216), .C1(n_184), .C2(n_326), .Y(n_594) );
OAI22xp33_ASAP7_75t_L g595 ( .A1(n_559), .A2(n_336), .B1(n_444), .B2(n_438), .Y(n_595) );
OA21x2_ASAP7_75t_L g596 ( .A1(n_560), .A2(n_438), .B(n_36), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_535), .Y(n_597) );
INVxp67_ASAP7_75t_L g598 ( .A(n_528), .Y(n_598) );
CKINVDCx14_ASAP7_75t_R g599 ( .A(n_521), .Y(n_599) );
AOI221xp5_ASAP7_75t_L g600 ( .A1(n_532), .A2(n_234), .B1(n_216), .B2(n_213), .C(n_201), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_562), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g602 ( .A(n_529), .B(n_32), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_546), .B(n_37), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_551), .B(n_48), .Y(n_604) );
OAI21xp5_ASAP7_75t_L g605 ( .A1(n_543), .A2(n_49), .B(n_52), .Y(n_605) );
AOI21xp5_ASAP7_75t_L g606 ( .A1(n_561), .A2(n_336), .B(n_234), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_589), .B(n_563), .Y(n_607) );
NAND3xp33_ASAP7_75t_L g608 ( .A(n_598), .B(n_543), .C(n_533), .Y(n_608) );
HB1xp67_ASAP7_75t_SL g609 ( .A(n_599), .Y(n_609) );
NAND4xp25_ASAP7_75t_SL g610 ( .A(n_590), .B(n_554), .C(n_539), .D(n_542), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_564), .B(n_535), .Y(n_611) );
AOI21xp33_ASAP7_75t_SL g612 ( .A1(n_593), .A2(n_566), .B(n_582), .Y(n_612) );
OAI21xp33_ASAP7_75t_L g613 ( .A1(n_572), .A2(n_521), .B(n_534), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_571), .Y(n_614) );
XOR2x2_ASAP7_75t_L g615 ( .A(n_577), .B(n_558), .Y(n_615) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_582), .B(n_552), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_573), .B(n_540), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_565), .A2(n_540), .B1(n_216), .B2(n_213), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_601), .Y(n_619) );
INVx1_ASAP7_75t_SL g620 ( .A(n_568), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g621 ( .A(n_593), .B(n_540), .Y(n_621) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_574), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_591), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_583), .Y(n_624) );
INVx1_ASAP7_75t_SL g625 ( .A(n_569), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_576), .B(n_54), .Y(n_626) );
NOR3xp33_ASAP7_75t_SL g627 ( .A(n_580), .B(n_56), .C(n_57), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_581), .Y(n_628) );
OAI21xp33_ASAP7_75t_L g629 ( .A1(n_567), .A2(n_184), .B(n_201), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_576), .Y(n_630) );
AND2x2_ASAP7_75t_L g631 ( .A(n_592), .B(n_67), .Y(n_631) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_597), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_588), .B(n_71), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_614), .Y(n_634) );
AOI32xp33_ASAP7_75t_L g635 ( .A1(n_620), .A2(n_584), .A3(n_570), .B1(n_575), .B2(n_604), .Y(n_635) );
NAND4xp75_ASAP7_75t_L g636 ( .A(n_621), .B(n_586), .C(n_585), .D(n_605), .Y(n_636) );
INVxp67_ASAP7_75t_L g637 ( .A(n_609), .Y(n_637) );
AOI22xp5_ASAP7_75t_L g638 ( .A1(n_613), .A2(n_588), .B1(n_602), .B2(n_603), .Y(n_638) );
INVx2_ASAP7_75t_SL g639 ( .A(n_625), .Y(n_639) );
OAI21xp5_ASAP7_75t_L g640 ( .A1(n_612), .A2(n_579), .B(n_585), .Y(n_640) );
AOI21xp33_ASAP7_75t_L g641 ( .A1(n_608), .A2(n_579), .B(n_587), .Y(n_641) );
INVxp67_ASAP7_75t_L g642 ( .A(n_622), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_624), .B(n_606), .Y(n_643) );
AOI21xp33_ASAP7_75t_L g644 ( .A1(n_621), .A2(n_596), .B(n_606), .Y(n_644) );
INVx3_ASAP7_75t_L g645 ( .A(n_617), .Y(n_645) );
OAI221xp5_ASAP7_75t_L g646 ( .A1(n_615), .A2(n_596), .B1(n_600), .B2(n_578), .C(n_594), .Y(n_646) );
XNOR2x2_ASAP7_75t_L g647 ( .A(n_615), .B(n_578), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_617), .Y(n_648) );
OAI211xp5_ASAP7_75t_L g649 ( .A1(n_618), .A2(n_595), .B(n_201), .C(n_213), .Y(n_649) );
INVx1_ASAP7_75t_SL g650 ( .A(n_632), .Y(n_650) );
NAND2xp33_ASAP7_75t_SL g651 ( .A(n_627), .B(n_184), .Y(n_651) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_641), .A2(n_628), .B1(n_616), .B2(n_619), .C(n_630), .Y(n_652) );
INVxp67_ASAP7_75t_L g653 ( .A(n_637), .Y(n_653) );
INVx1_ASAP7_75t_SL g654 ( .A(n_650), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_634), .Y(n_655) );
NOR2x1_ASAP7_75t_L g656 ( .A(n_636), .B(n_626), .Y(n_656) );
NAND2xp33_ASAP7_75t_L g657 ( .A(n_635), .B(n_618), .Y(n_657) );
INVx1_ASAP7_75t_SL g658 ( .A(n_639), .Y(n_658) );
NOR2x1_ASAP7_75t_L g659 ( .A(n_640), .B(n_633), .Y(n_659) );
XNOR2xp5_ASAP7_75t_L g660 ( .A(n_647), .B(n_607), .Y(n_660) );
OAI21xp33_ASAP7_75t_L g661 ( .A1(n_640), .A2(n_616), .B(n_610), .Y(n_661) );
AOI21xp5_ASAP7_75t_L g662 ( .A1(n_646), .A2(n_629), .B(n_611), .Y(n_662) );
BUFx2_ASAP7_75t_L g663 ( .A(n_642), .Y(n_663) );
OAI211xp5_ASAP7_75t_SL g664 ( .A1(n_644), .A2(n_633), .B(n_623), .C(n_607), .Y(n_664) );
AOI211xp5_ASAP7_75t_L g665 ( .A1(n_649), .A2(n_631), .B(n_184), .C(n_216), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g666 ( .A1(n_645), .A2(n_648), .B1(n_638), .B2(n_643), .Y(n_666) );
AOI211xp5_ASAP7_75t_L g667 ( .A1(n_651), .A2(n_641), .B(n_640), .C(n_612), .Y(n_667) );
OAI211xp5_ASAP7_75t_L g668 ( .A1(n_635), .A2(n_637), .B(n_641), .C(n_640), .Y(n_668) );
CKINVDCx20_ASAP7_75t_R g669 ( .A(n_653), .Y(n_669) );
OAI221xp5_ASAP7_75t_L g670 ( .A1(n_668), .A2(n_667), .B1(n_657), .B2(n_661), .C(n_660), .Y(n_670) );
INVx2_ASAP7_75t_L g671 ( .A(n_663), .Y(n_671) );
CKINVDCx20_ASAP7_75t_R g672 ( .A(n_658), .Y(n_672) );
AND2x4_ASAP7_75t_L g673 ( .A(n_654), .B(n_659), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_669), .Y(n_674) );
NOR4xp25_ASAP7_75t_L g675 ( .A(n_670), .B(n_652), .C(n_666), .D(n_664), .Y(n_675) );
AND3x2_ASAP7_75t_L g676 ( .A(n_673), .B(n_665), .C(n_655), .Y(n_676) );
INVx1_ASAP7_75t_L g677 ( .A(n_674), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_676), .Y(n_678) );
INVxp67_ASAP7_75t_SL g679 ( .A(n_677), .Y(n_679) );
INVxp67_ASAP7_75t_L g680 ( .A(n_678), .Y(n_680) );
AOI222xp33_ASAP7_75t_L g681 ( .A1(n_680), .A2(n_673), .B1(n_671), .B2(n_672), .C1(n_675), .C2(n_656), .Y(n_681) );
AOI21xp5_ASAP7_75t_L g682 ( .A1(n_681), .A2(n_679), .B(n_662), .Y(n_682) );
endmodule