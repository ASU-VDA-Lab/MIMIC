module fake_jpeg_24252_n_317 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_317);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_145;
wire n_18;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

INVx4_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_6),
.B(n_11),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_12),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_32),
.B(n_37),
.Y(n_56)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx3_ASAP7_75t_SL g40 ( 
.A(n_34),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_16),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_36),
.B(n_39),
.Y(n_51)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_54),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_26),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_49),
.B(n_27),
.Y(n_64)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_29),
.A2(n_15),
.B1(n_14),
.B2(n_33),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_52),
.A2(n_33),
.B1(n_14),
.B2(n_15),
.Y(n_71)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_25),
.Y(n_67)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_60),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_66),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_35),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_67),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_39),
.Y(n_68)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_71),
.A2(n_50),
.B1(n_44),
.B2(n_37),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_39),
.Y(n_72)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_35),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_46),
.Y(n_95)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_76),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_41),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_58),
.A2(n_33),
.B1(n_15),
.B2(n_14),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_77),
.A2(n_79),
.B1(n_45),
.B2(n_57),
.Y(n_87)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_59),
.Y(n_78)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_42),
.A2(n_14),
.B1(n_15),
.B2(n_32),
.Y(n_79)
);

AND2x2_ASAP7_75t_SL g80 ( 
.A(n_45),
.B(n_37),
.Y(n_80)
);

AND2x2_ASAP7_75t_SL g85 ( 
.A(n_80),
.B(n_53),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_82),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_36),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_83),
.B(n_96),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_85),
.A2(n_80),
.B(n_67),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_87),
.A2(n_71),
.B1(n_77),
.B2(n_79),
.Y(n_123)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_73),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_94),
.B(n_98),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_95),
.B(n_97),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_36),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_55),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_62),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_99),
.B(n_100),
.Y(n_117)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_103),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_64),
.B(n_47),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_105),
.A2(n_65),
.B1(n_70),
.B2(n_60),
.Y(n_129)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_60),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_96),
.B(n_21),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_107),
.B(n_109),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_108),
.A2(n_63),
.B(n_76),
.Y(n_147)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_96),
.B(n_21),
.Y(n_110)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_116),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_83),
.B(n_28),
.Y(n_115)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_115),
.Y(n_142)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_91),
.Y(n_116)
);

AND2x6_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_80),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_118),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_89),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_120),
.Y(n_136)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_124),
.Y(n_157)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_93),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_122),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_123),
.A2(n_129),
.B1(n_106),
.B2(n_102),
.Y(n_141)
);

FAx1_ASAP7_75t_SL g124 ( 
.A(n_90),
.B(n_80),
.CI(n_32),
.CON(n_124),
.SN(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_125),
.B(n_126),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_83),
.B(n_85),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_94),
.B(n_30),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_87),
.Y(n_138)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_86),
.A2(n_16),
.B(n_28),
.C(n_23),
.Y(n_128)
);

OAI32xp33_ASAP7_75t_L g137 ( 
.A1(n_128),
.A2(n_88),
.A3(n_92),
.B1(n_99),
.B2(n_98),
.Y(n_137)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_130),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_119),
.A2(n_40),
.B1(n_65),
.B2(n_84),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_132),
.A2(n_84),
.B1(n_119),
.B2(n_153),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_137),
.B(n_146),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_138),
.B(n_143),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_111),
.B(n_92),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_152),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_141),
.A2(n_145),
.B1(n_40),
.B2(n_61),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_108),
.B(n_88),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_112),
.B(n_127),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_144),
.A2(n_126),
.B(n_124),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_123),
.A2(n_100),
.B1(n_44),
.B2(n_30),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_130),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_147),
.A2(n_115),
.B(n_26),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_151),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_124),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_149),
.B(n_150),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_113),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_112),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_111),
.B(n_93),
.Y(n_152)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_114),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g194 ( 
.A1(n_159),
.A2(n_175),
.B1(n_179),
.B2(n_24),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_156),
.B(n_125),
.C(n_135),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_160),
.B(n_176),
.C(n_154),
.Y(n_189)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_164),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_162),
.B(n_166),
.Y(n_185)
);

BUFx12f_ASAP7_75t_L g163 ( 
.A(n_156),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_163),
.Y(n_187)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_178),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_142),
.B(n_120),
.Y(n_166)
);

NOR2x1_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_126),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_167),
.B(n_23),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_135),
.A2(n_118),
.B1(n_121),
.B2(n_109),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_168),
.A2(n_172),
.B1(n_182),
.B2(n_43),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_169),
.B(n_170),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_157),
.B(n_131),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_151),
.A2(n_128),
.B1(n_61),
.B2(n_116),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_122),
.C(n_110),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_107),
.Y(n_177)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_177),
.Y(n_203)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_145),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_136),
.B(n_101),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_183),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_134),
.A2(n_61),
.B1(n_48),
.B2(n_91),
.Y(n_182)
);

AOI32xp33_ASAP7_75t_L g183 ( 
.A1(n_149),
.A2(n_75),
.A3(n_104),
.B1(n_48),
.B2(n_78),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_134),
.Y(n_184)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_184),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_189),
.A2(n_190),
.B(n_195),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_163),
.A2(n_144),
.B(n_148),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_160),
.A2(n_144),
.B1(n_141),
.B2(n_138),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_191),
.A2(n_209),
.B1(n_172),
.B2(n_173),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_171),
.B(n_139),
.Y(n_193)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_193),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_196),
.Y(n_213)
);

XOR2x2_ASAP7_75t_L g195 ( 
.A(n_167),
.B(n_143),
.Y(n_195)
);

OA21x2_ASAP7_75t_L g196 ( 
.A1(n_163),
.A2(n_18),
.B(n_28),
.Y(n_196)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_197),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_174),
.B(n_43),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_174),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_161),
.B(n_104),
.Y(n_200)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_200),
.Y(n_218)
);

OAI21xp33_ASAP7_75t_L g201 ( 
.A1(n_169),
.A2(n_11),
.B(n_13),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_12),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_171),
.B(n_25),
.Y(n_202)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_202),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_205),
.B(n_206),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_177),
.B(n_23),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_158),
.B(n_74),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_207),
.B(n_208),
.Y(n_220)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_168),
.A2(n_26),
.B1(n_18),
.B2(n_24),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_189),
.B(n_190),
.C(n_191),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_212),
.B(n_216),
.C(n_219),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_226),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_215),
.A2(n_227),
.B1(n_209),
.B2(n_193),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_188),
.B(n_187),
.C(n_208),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_188),
.B(n_170),
.C(n_176),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_195),
.Y(n_221)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_221),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g224 ( 
.A(n_204),
.Y(n_224)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_224),
.Y(n_240)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_204),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_229),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_179),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_187),
.A2(n_175),
.B1(n_182),
.B2(n_24),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_69),
.C(n_38),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_185),
.C(n_206),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_197),
.B(n_69),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_205),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_220),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_0),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_233),
.B(n_245),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_211),
.A2(n_192),
.B1(n_203),
.B2(n_199),
.Y(n_235)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_235),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_216),
.A2(n_210),
.B1(n_212),
.B2(n_224),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_236),
.A2(n_238),
.B1(n_20),
.B2(n_27),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_218),
.Y(n_237)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_237),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_223),
.A2(n_196),
.B1(n_202),
.B2(n_186),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_241),
.B(n_242),
.C(n_226),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_185),
.C(n_196),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_250),
.Y(n_259)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_228),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_213),
.B(n_25),
.Y(n_246)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_246),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_230),
.A2(n_18),
.B1(n_27),
.B2(n_19),
.Y(n_247)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_247),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_229),
.B(n_25),
.Y(n_248)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_248),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_222),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_249),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_38),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_234),
.Y(n_270)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_253),
.Y(n_269)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_9),
.Y(n_255)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_255),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_236),
.B(n_239),
.C(n_231),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_82),
.C(n_20),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_239),
.B(n_38),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_250),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_244),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_262),
.A2(n_265),
.B1(n_241),
.B2(n_234),
.Y(n_271)
);

BUFx12_ASAP7_75t_L g264 ( 
.A(n_240),
.Y(n_264)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_264),
.Y(n_280)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_243),
.Y(n_265)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_266),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_257),
.A2(n_232),
.B(n_242),
.Y(n_268)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_268),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_272),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_271),
.B(n_274),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_251),
.B(n_38),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_277),
.C(n_278),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_17),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_264),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_82),
.C(n_20),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_7),
.Y(n_278)
);

XNOR2x1_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_0),
.Y(n_279)
);

XNOR2x1_ASAP7_75t_L g284 ( 
.A(n_279),
.B(n_255),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_282),
.B(n_290),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_284),
.A2(n_13),
.B(n_11),
.Y(n_301)
);

NAND2xp33_ASAP7_75t_SL g285 ( 
.A(n_279),
.B(n_252),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_285),
.A2(n_288),
.B(n_291),
.Y(n_299)
);

BUFx24_ASAP7_75t_SL g287 ( 
.A(n_280),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_8),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_275),
.A2(n_254),
.B(n_260),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_253),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_273),
.A2(n_267),
.B(n_264),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_281),
.A2(n_258),
.B1(n_256),
.B2(n_263),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_292),
.A2(n_269),
.B1(n_278),
.B2(n_27),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_289),
.B(n_272),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_300),
.C(n_283),
.Y(n_303)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_295),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_286),
.A2(n_19),
.B1(n_17),
.B2(n_6),
.Y(n_296)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_296),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_293),
.B(n_19),
.Y(n_298)
);

AOI322xp5_ASAP7_75t_L g305 ( 
.A1(n_298),
.A2(n_301),
.A3(n_302),
.B1(n_7),
.B2(n_1),
.C1(n_2),
.C2(n_3),
.Y(n_305)
);

AOI21xp33_ASAP7_75t_L g300 ( 
.A1(n_284),
.A2(n_6),
.B(n_13),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_303),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_289),
.C(n_297),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_306),
.C(n_301),
.Y(n_310)
);

BUFx24_ASAP7_75t_SL g309 ( 
.A(n_305),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_299),
.A2(n_283),
.B1(n_19),
.B2(n_7),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_310),
.A2(n_308),
.B1(n_307),
.B2(n_2),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_312),
.B(n_309),
.Y(n_313)
);

AOI322xp5_ASAP7_75t_L g314 ( 
.A1(n_313),
.A2(n_311),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_314),
.A2(n_0),
.B(n_1),
.Y(n_315)
);

OAI211xp5_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_4),
.B(n_5),
.C(n_284),
.Y(n_316)
);

AO31x2_ASAP7_75t_SL g317 ( 
.A1(n_316),
.A2(n_4),
.A3(n_5),
.B(n_284),
.Y(n_317)
);


endmodule