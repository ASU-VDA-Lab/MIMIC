module fake_jpeg_7295_n_250 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_250);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_250;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx24_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

HB1xp67_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_34),
.Y(n_43)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_22),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_22),
.B1(n_18),
.B2(n_37),
.Y(n_49)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_7),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_38),
.B(n_11),
.Y(n_64)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_42),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_24),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_46),
.A2(n_57),
.B(n_60),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_33),
.A2(n_22),
.B1(n_24),
.B2(n_18),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_47),
.A2(n_49),
.B1(n_61),
.B2(n_60),
.Y(n_71)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_51),
.B(n_52),
.Y(n_66)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_26),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_53),
.B(n_54),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_26),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g81 ( 
.A(n_55),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_36),
.A2(n_16),
.B1(n_21),
.B2(n_29),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_64),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_42),
.A2(n_16),
.B1(n_21),
.B2(n_25),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_42),
.A2(n_25),
.B1(n_23),
.B2(n_15),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_34),
.B(n_28),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_62),
.B(n_27),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_31),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_63),
.B(n_65),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_28),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_67),
.B(n_72),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_54),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_69),
.A2(n_50),
.B1(n_56),
.B2(n_58),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_57),
.A2(n_41),
.B1(n_40),
.B2(n_25),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_70),
.A2(n_84),
.B1(n_65),
.B2(n_56),
.Y(n_102)
);

OA22x2_ASAP7_75t_L g94 ( 
.A1(n_71),
.A2(n_47),
.B1(n_23),
.B2(n_56),
.Y(n_94)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

OAI21xp33_ASAP7_75t_L g98 ( 
.A1(n_74),
.A2(n_75),
.B(n_50),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_41),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_76),
.B(n_82),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_40),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_85),
.Y(n_87)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_79),
.Y(n_93)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_44),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_51),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_83),
.B(n_52),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_61),
.A2(n_23),
.B1(n_20),
.B2(n_40),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_28),
.Y(n_85)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_86),
.Y(n_129)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_88),
.Y(n_112)
);

AND2x4_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_46),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_90),
.A2(n_98),
.B(n_105),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g91 ( 
.A(n_66),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_91),
.B(n_96),
.Y(n_111)
);

AND2x6_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_46),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_92),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_94),
.A2(n_95),
.B1(n_102),
.B2(n_70),
.Y(n_109)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_67),
.B(n_51),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_99),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_81),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_101),
.B(n_103),
.Y(n_116)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

INVx13_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_104),
.B(n_107),
.Y(n_124)
);

AOI32xp33_ASAP7_75t_L g105 ( 
.A1(n_77),
.A2(n_63),
.A3(n_59),
.B1(n_45),
.B2(n_53),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_85),
.B(n_64),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_73),
.C(n_82),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_81),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_72),
.A2(n_58),
.B1(n_48),
.B2(n_45),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_108),
.A2(n_68),
.B(n_77),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_109),
.A2(n_94),
.B1(n_69),
.B2(n_105),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_110),
.A2(n_115),
.B(n_118),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_85),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_119),
.Y(n_134)
);

XNOR2x1_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_120),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_87),
.A2(n_68),
.B(n_73),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_90),
.A2(n_68),
.B(n_74),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_78),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_106),
.B(n_70),
.C(n_80),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_78),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_125),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_91),
.B(n_80),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_90),
.B(n_71),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g132 ( 
.A(n_126),
.B(n_92),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_96),
.B(n_75),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_128),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_90),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_55),
.Y(n_130)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_130),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_132),
.B(n_144),
.C(n_117),
.Y(n_166)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_116),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_141),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_135),
.A2(n_146),
.B1(n_154),
.B2(n_114),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_93),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_136),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_119),
.B(n_95),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_138),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_88),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_127),
.B(n_94),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_140),
.A2(n_142),
.B(n_149),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_93),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_110),
.A2(n_84),
.B(n_103),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_122),
.B(n_94),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_126),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_109),
.A2(n_48),
.B1(n_101),
.B2(n_107),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_116),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_147),
.B(n_152),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_122),
.A2(n_27),
.B(n_17),
.Y(n_149)
);

O2A1O1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_111),
.A2(n_55),
.B(n_104),
.C(n_27),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_151),
.A2(n_111),
.B1(n_124),
.B2(n_131),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_79),
.Y(n_152)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_0),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_153),
.A2(n_121),
.B(n_124),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_117),
.A2(n_79),
.B1(n_55),
.B2(n_81),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_138),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_160),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_158),
.B(n_153),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_159),
.B(n_162),
.Y(n_180)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_151),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_134),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_165),
.Y(n_188)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_146),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_172),
.C(n_149),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_143),
.A2(n_130),
.B1(n_128),
.B2(n_115),
.Y(n_167)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_167),
.Y(n_178)
);

INVxp33_ASAP7_75t_L g168 ( 
.A(n_145),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_168),
.B(n_173),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_143),
.A2(n_126),
.B1(n_118),
.B2(n_120),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_169),
.A2(n_150),
.B1(n_114),
.B2(n_113),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_170),
.A2(n_132),
.B1(n_135),
.B2(n_148),
.Y(n_176)
);

BUFx12f_ASAP7_75t_L g171 ( 
.A(n_133),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_171),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_145),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_147),
.B(n_131),
.Y(n_174)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_174),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_176),
.B(n_186),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_170),
.A2(n_142),
.B1(n_137),
.B2(n_154),
.Y(n_177)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_165),
.A2(n_140),
.B1(n_148),
.B2(n_139),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_182),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_160),
.A2(n_140),
.B1(n_139),
.B2(n_120),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_185),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_164),
.Y(n_198)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_171),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_162),
.A2(n_150),
.B1(n_112),
.B2(n_153),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_187),
.A2(n_171),
.B(n_20),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_166),
.C(n_172),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_192),
.C(n_184),
.Y(n_197)
);

AO22x1_ASAP7_75t_L g200 ( 
.A1(n_191),
.A2(n_159),
.B1(n_161),
.B2(n_157),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_163),
.B(n_112),
.C(n_20),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_179),
.A2(n_175),
.B(n_156),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_194),
.B(n_204),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_190),
.A2(n_155),
.B1(n_175),
.B2(n_158),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_195),
.A2(n_180),
.B1(n_178),
.B2(n_188),
.Y(n_209)
);

NOR2x1_ASAP7_75t_L g196 ( 
.A(n_191),
.B(n_164),
.Y(n_196)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_196),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_197),
.B(n_198),
.C(n_202),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g212 ( 
.A(n_200),
.B(n_203),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_171),
.C(n_20),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_17),
.C(n_1),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_176),
.B(n_186),
.C(n_183),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_206),
.B(n_208),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_177),
.B(n_17),
.C(n_1),
.Y(n_208)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_209),
.Y(n_225)
);

INVxp33_ASAP7_75t_L g211 ( 
.A(n_196),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_211),
.A2(n_217),
.B1(n_7),
.B2(n_14),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_201),
.A2(n_180),
.B1(n_188),
.B2(n_193),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_213),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_207),
.B(n_181),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_214),
.B(n_219),
.Y(n_224)
);

INVxp33_ASAP7_75t_L g217 ( 
.A(n_200),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_208),
.B(n_192),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_202),
.B(n_185),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_220),
.Y(n_222)
);

NOR3xp33_ASAP7_75t_L g223 ( 
.A(n_211),
.B(n_204),
.C(n_206),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_226),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_210),
.A2(n_205),
.B(n_198),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_216),
.B(n_197),
.C(n_199),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_227),
.B(n_228),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_217),
.A2(n_199),
.B(n_187),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_229),
.B(n_11),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_232),
.B(n_233),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_221),
.A2(n_212),
.B1(n_218),
.B2(n_215),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_218),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_234),
.A2(n_236),
.B(n_225),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_222),
.B(n_215),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_235),
.B(n_223),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_229),
.B(n_216),
.Y(n_236)
);

AOI322xp5_ASAP7_75t_L g242 ( 
.A1(n_237),
.A2(n_240),
.A3(n_231),
.B1(n_233),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_239),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_230),
.B(n_212),
.C(n_9),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_6),
.C(n_14),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_241),
.A2(n_11),
.B(n_13),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_244),
.Y(n_246)
);

AOI322xp5_ASAP7_75t_L g244 ( 
.A1(n_240),
.A2(n_10),
.A3(n_14),
.B1(n_13),
.B2(n_3),
.C1(n_6),
.C2(n_12),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_245),
.A2(n_10),
.B(n_12),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_247),
.A2(n_243),
.B(n_17),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_248),
.A2(n_246),
.B1(n_10),
.B2(n_2),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_0),
.Y(n_250)
);


endmodule