module real_jpeg_8950_n_6 (n_5, n_4, n_0, n_1, n_2, n_3, n_6);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_3;

output n_6;

wire n_17;
wire n_8;
wire n_43;
wire n_37;
wire n_21;
wire n_38;
wire n_35;
wire n_33;
wire n_29;
wire n_10;
wire n_31;
wire n_9;
wire n_12;
wire n_24;
wire n_34;
wire n_44;
wire n_28;
wire n_46;
wire n_23;
wire n_11;
wire n_14;
wire n_45;
wire n_25;
wire n_42;
wire n_7;
wire n_22;
wire n_18;
wire n_40;
wire n_36;
wire n_39;
wire n_41;
wire n_26;
wire n_27;
wire n_20;
wire n_19;
wire n_32;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

OR2x2_ASAP7_75t_SL g29 ( 
.A(n_1),
.B(n_30),
.Y(n_29)
);

OR2x2_ASAP7_75t_SL g37 ( 
.A(n_1),
.B(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_2),
.B(n_4),
.Y(n_13)
);

OR2x2_ASAP7_75t_L g18 ( 
.A(n_3),
.B(n_19),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

OA21x2_ASAP7_75t_L g22 ( 
.A1(n_5),
.A2(n_9),
.B(n_13),
.Y(n_22)
);

OAI211xp5_ASAP7_75t_L g6 ( 
.A1(n_7),
.A2(n_14),
.B(n_20),
.C(n_40),
.Y(n_6)
);

AOI221xp5_ASAP7_75t_L g20 ( 
.A1(n_7),
.A2(n_21),
.B1(n_23),
.B2(n_26),
.C(n_31),
.Y(n_20)
);

OA21x2_ASAP7_75t_L g7 ( 
.A1(n_8),
.A2(n_9),
.B(n_13),
.Y(n_7)
);

AO21x1_ASAP7_75t_L g33 ( 
.A1(n_8),
.A2(n_16),
.B(n_34),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_8),
.B(n_16),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_8),
.B(n_17),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g9 ( 
.A(n_10),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_12),
.Y(n_10)
);

AOI221xp5_ASAP7_75t_L g40 ( 
.A1(n_11),
.A2(n_22),
.B1(n_41),
.B2(n_42),
.C(n_44),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_11),
.B(n_17),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_18),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_16),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_16),
.B(n_28),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_16),
.A2(n_36),
.B(n_38),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_16),
.B(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_16),
.B(n_29),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

OR2x2_ASAP7_75t_SL g39 ( 
.A(n_19),
.B(n_30),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_35),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);


endmodule