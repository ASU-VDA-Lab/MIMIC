module fake_netlist_6_2441_n_1747 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1747);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1747;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1605;
wire n_1413;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_91),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_36),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_141),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_23),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_112),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_38),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_61),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_118),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_115),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_104),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_74),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_53),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_121),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_101),
.Y(n_169)
);

BUFx10_ASAP7_75t_L g170 ( 
.A(n_66),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_108),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_146),
.Y(n_172)
);

BUFx10_ASAP7_75t_L g173 ( 
.A(n_94),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_144),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_151),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_49),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_50),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_18),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_39),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_133),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_150),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_129),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_99),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_149),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_90),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_154),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_50),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_127),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_54),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_29),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_75),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_68),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_116),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_4),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_24),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_131),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_95),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_136),
.Y(n_198)
);

BUFx10_ASAP7_75t_L g199 ( 
.A(n_142),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g200 ( 
.A(n_51),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_13),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_58),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_3),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_31),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_78),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_62),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_135),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_15),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_12),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g210 ( 
.A(n_79),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_132),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_9),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_96),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_92),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_21),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_155),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_111),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_81),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_123),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_49),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_86),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_67),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_117),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_42),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_31),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_113),
.Y(n_226)
);

INVx2_ASAP7_75t_SL g227 ( 
.A(n_36),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_53),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_72),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_143),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_11),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_82),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_57),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_105),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_93),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_32),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_84),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_110),
.Y(n_238)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_120),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_6),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_138),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_51),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_45),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_23),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_59),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_114),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_76),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_15),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_77),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_148),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_45),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_57),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_60),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_28),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_7),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_7),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_55),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_107),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_152),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_126),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_52),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_109),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_83),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_28),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_63),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_125),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_19),
.Y(n_267)
);

INVx2_ASAP7_75t_SL g268 ( 
.A(n_97),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_119),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_106),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_6),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_33),
.Y(n_272)
);

BUFx2_ASAP7_75t_L g273 ( 
.A(n_140),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_22),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_44),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_1),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_14),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_73),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_18),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_29),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_153),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_33),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_54),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_103),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_38),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_3),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_134),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_64),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_87),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_98),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_24),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_69),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_71),
.Y(n_293)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_89),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_32),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_48),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_137),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_30),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_102),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_46),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_37),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_39),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_14),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_27),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_4),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_43),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_5),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_19),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_5),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_200),
.Y(n_310)
);

INVxp33_ASAP7_75t_L g311 ( 
.A(n_264),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_156),
.Y(n_312)
);

INVxp67_ASAP7_75t_SL g313 ( 
.A(n_168),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_158),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_200),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_163),
.Y(n_316)
);

CKINVDCx14_ASAP7_75t_R g317 ( 
.A(n_210),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_175),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_200),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_241),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_200),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_194),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_166),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_290),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_258),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_200),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_200),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_169),
.Y(n_328)
);

BUFx6f_ASAP7_75t_L g329 ( 
.A(n_258),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_200),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_172),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_174),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_200),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_185),
.Y(n_334)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_205),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_200),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_180),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_215),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_215),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_182),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_183),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_184),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_194),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_188),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_192),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_193),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_167),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_215),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_196),
.Y(n_349)
);

INVxp33_ASAP7_75t_SL g350 ( 
.A(n_157),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_215),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_197),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_215),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_251),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_206),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_207),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_211),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_216),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_258),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_217),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_251),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_218),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_221),
.Y(n_363)
);

INVxp33_ASAP7_75t_SL g364 ( 
.A(n_161),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_177),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_251),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_222),
.Y(n_367)
);

INVxp33_ASAP7_75t_SL g368 ( 
.A(n_201),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_251),
.Y(n_369)
);

BUFx2_ASAP7_75t_L g370 ( 
.A(n_236),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_226),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_251),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_298),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_232),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_298),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_258),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_234),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_298),
.Y(n_378)
);

BUFx2_ASAP7_75t_L g379 ( 
.A(n_236),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_237),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_238),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_326),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_338),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_338),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_339),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_339),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_325),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_348),
.B(n_210),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_318),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_348),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_326),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_350),
.B(n_273),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_351),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_317),
.B(n_273),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_351),
.B(n_278),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_353),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_326),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_364),
.B(n_278),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_353),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_325),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_325),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_325),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_354),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_347),
.B(n_195),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_321),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_354),
.B(n_268),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_370),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_361),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_321),
.Y(n_409)
);

AND2x4_ASAP7_75t_L g410 ( 
.A(n_373),
.B(n_205),
.Y(n_410)
);

OA21x2_ASAP7_75t_L g411 ( 
.A1(n_359),
.A2(n_277),
.B(n_231),
.Y(n_411)
);

CKINVDCx6p67_ASAP7_75t_R g412 ( 
.A(n_334),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_361),
.B(n_268),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_366),
.Y(n_414)
);

NAND2xp33_ASAP7_75t_L g415 ( 
.A(n_325),
.B(n_227),
.Y(n_415)
);

INVx4_ASAP7_75t_L g416 ( 
.A(n_325),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_329),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_329),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_366),
.Y(n_419)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_329),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_329),
.Y(n_421)
);

NAND2xp33_ASAP7_75t_SL g422 ( 
.A(n_311),
.B(n_227),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_335),
.B(n_294),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_329),
.Y(n_424)
);

BUFx2_ASAP7_75t_L g425 ( 
.A(n_370),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_369),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_369),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_329),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_372),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_372),
.B(n_245),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_359),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_376),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_373),
.B(n_249),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_359),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_335),
.B(n_294),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_368),
.B(n_313),
.Y(n_436)
);

OR2x6_ASAP7_75t_L g437 ( 
.A(n_375),
.B(n_162),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_342),
.Y(n_438)
);

AND2x4_ASAP7_75t_L g439 ( 
.A(n_375),
.B(n_378),
.Y(n_439)
);

NAND3xp33_ASAP7_75t_L g440 ( 
.A(n_343),
.B(n_176),
.C(n_159),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_376),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_335),
.B(n_160),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_310),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_376),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_310),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_378),
.B(n_250),
.Y(n_446)
);

INVx4_ASAP7_75t_L g447 ( 
.A(n_411),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_382),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_430),
.B(n_312),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_411),
.Y(n_450)
);

INVx1_ASAP7_75t_SL g451 ( 
.A(n_389),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_382),
.Y(n_452)
);

NAND2xp33_ASAP7_75t_L g453 ( 
.A(n_433),
.B(n_314),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_382),
.Y(n_454)
);

BUFx10_ASAP7_75t_L g455 ( 
.A(n_436),
.Y(n_455)
);

OR2x6_ASAP7_75t_L g456 ( 
.A(n_437),
.B(n_160),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_387),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_411),
.Y(n_458)
);

BUFx3_ASAP7_75t_L g459 ( 
.A(n_411),
.Y(n_459)
);

NAND3xp33_ASAP7_75t_L g460 ( 
.A(n_398),
.B(n_365),
.C(n_323),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_411),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_430),
.B(n_316),
.Y(n_462)
);

AND2x4_ASAP7_75t_L g463 ( 
.A(n_410),
.B(n_164),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_382),
.Y(n_464)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_398),
.A2(n_224),
.B1(n_280),
.B2(n_306),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_436),
.B(n_328),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_392),
.B(n_331),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_391),
.Y(n_468)
);

AOI22xp33_ASAP7_75t_L g469 ( 
.A1(n_442),
.A2(n_322),
.B1(n_231),
.B2(n_283),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_387),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_411),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_443),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_387),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_387),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_443),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_445),
.Y(n_476)
);

INVx4_ASAP7_75t_L g477 ( 
.A(n_387),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_392),
.B(n_332),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_391),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_404),
.A2(n_248),
.B1(n_244),
.B2(n_225),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_387),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_445),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_394),
.B(n_337),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_423),
.B(n_340),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_394),
.B(n_341),
.Y(n_485)
);

AOI22xp33_ASAP7_75t_L g486 ( 
.A1(n_442),
.A2(n_190),
.B1(n_242),
.B2(n_240),
.Y(n_486)
);

INVx4_ASAP7_75t_L g487 ( 
.A(n_387),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_383),
.Y(n_488)
);

INVx2_ASAP7_75t_SL g489 ( 
.A(n_423),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_423),
.B(n_379),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_435),
.B(n_379),
.Y(n_491)
);

INVx2_ASAP7_75t_SL g492 ( 
.A(n_435),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_435),
.B(n_344),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_383),
.Y(n_494)
);

AOI22xp33_ASAP7_75t_L g495 ( 
.A1(n_410),
.A2(n_187),
.B1(n_243),
.B2(n_240),
.Y(n_495)
);

AO22x2_ASAP7_75t_L g496 ( 
.A1(n_440),
.A2(n_257),
.B1(n_300),
.B2(n_261),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_391),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_387),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_391),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_400),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_397),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_397),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_384),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_407),
.B(n_345),
.Y(n_504)
);

NAND2xp33_ASAP7_75t_SL g505 ( 
.A(n_425),
.B(n_346),
.Y(n_505)
);

AND2x2_ASAP7_75t_SL g506 ( 
.A(n_404),
.B(n_162),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_397),
.Y(n_507)
);

OR2x2_ASAP7_75t_L g508 ( 
.A(n_425),
.B(n_349),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_407),
.B(n_355),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_433),
.B(n_371),
.Y(n_510)
);

AOI22xp33_ASAP7_75t_L g511 ( 
.A1(n_410),
.A2(n_439),
.B1(n_440),
.B2(n_395),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_384),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_385),
.Y(n_513)
);

AND2x6_ASAP7_75t_L g514 ( 
.A(n_410),
.B(n_186),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_400),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_446),
.B(n_374),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_397),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_385),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_446),
.B(n_377),
.Y(n_519)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_425),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_386),
.Y(n_521)
);

INVxp33_ASAP7_75t_L g522 ( 
.A(n_388),
.Y(n_522)
);

INVx4_ASAP7_75t_L g523 ( 
.A(n_400),
.Y(n_523)
);

OR2x6_ASAP7_75t_L g524 ( 
.A(n_437),
.B(n_388),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_405),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_405),
.Y(n_526)
);

BUFx10_ASAP7_75t_L g527 ( 
.A(n_438),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_386),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_405),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_395),
.B(n_380),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_390),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g532 ( 
.A(n_400),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_390),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_393),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_422),
.B(n_381),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_439),
.B(n_315),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_422),
.B(n_352),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_439),
.B(n_315),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_400),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_410),
.B(n_356),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_439),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_439),
.B(n_319),
.Y(n_542)
);

INVxp33_ASAP7_75t_L g543 ( 
.A(n_406),
.Y(n_543)
);

NAND2xp33_ASAP7_75t_SL g544 ( 
.A(n_406),
.B(n_357),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_438),
.B(n_358),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_405),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_400),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_393),
.B(n_319),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_400),
.Y(n_549)
);

CKINVDCx16_ASAP7_75t_R g550 ( 
.A(n_389),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_413),
.B(n_360),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_412),
.Y(n_552)
);

BUFx6f_ASAP7_75t_SL g553 ( 
.A(n_437),
.Y(n_553)
);

AND2x6_ASAP7_75t_L g554 ( 
.A(n_409),
.B(n_186),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_396),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_409),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_396),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_409),
.Y(n_558)
);

INVx2_ASAP7_75t_SL g559 ( 
.A(n_437),
.Y(n_559)
);

INVx2_ASAP7_75t_SL g560 ( 
.A(n_437),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_399),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_399),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_403),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_403),
.B(n_327),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_409),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_431),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_431),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_408),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_408),
.B(n_327),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_419),
.B(n_362),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_400),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_414),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_419),
.B(n_363),
.Y(n_573)
);

INVx4_ASAP7_75t_L g574 ( 
.A(n_401),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_401),
.Y(n_575)
);

BUFx6f_ASAP7_75t_SL g576 ( 
.A(n_437),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_426),
.B(n_427),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_401),
.Y(n_578)
);

INVx2_ASAP7_75t_SL g579 ( 
.A(n_413),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_426),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_427),
.B(n_330),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_429),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_434),
.Y(n_583)
);

BUFx10_ASAP7_75t_L g584 ( 
.A(n_429),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_414),
.B(n_330),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_414),
.B(n_367),
.Y(n_586)
);

INVx4_ASAP7_75t_L g587 ( 
.A(n_401),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_434),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_416),
.B(n_170),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_401),
.Y(n_590)
);

INVx4_ASAP7_75t_L g591 ( 
.A(n_401),
.Y(n_591)
);

INVx8_ASAP7_75t_L g592 ( 
.A(n_524),
.Y(n_592)
);

INVx8_ASAP7_75t_L g593 ( 
.A(n_524),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_541),
.Y(n_594)
);

O2A1O1Ixp33_ASAP7_75t_L g595 ( 
.A1(n_579),
.A2(n_415),
.B(n_252),
.C(n_178),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_541),
.B(n_258),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_579),
.B(n_416),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_541),
.B(n_223),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_489),
.B(n_164),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_506),
.B(n_223),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_506),
.B(n_266),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_SL g602 ( 
.A1(n_480),
.A2(n_320),
.B1(n_324),
.B2(n_254),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_572),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_530),
.B(n_416),
.Y(n_604)
);

BUFx6f_ASAP7_75t_SL g605 ( 
.A(n_527),
.Y(n_605)
);

INVx8_ASAP7_75t_L g606 ( 
.A(n_524),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_519),
.B(n_416),
.Y(n_607)
);

INVxp67_ASAP7_75t_L g608 ( 
.A(n_508),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_489),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_506),
.B(n_266),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_L g611 ( 
.A1(n_492),
.A2(n_297),
.B1(n_292),
.B2(n_239),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_522),
.B(n_412),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_492),
.B(n_416),
.Y(n_613)
);

A2O1A1Ixp33_ASAP7_75t_L g614 ( 
.A1(n_536),
.A2(n_333),
.B(n_336),
.C(n_219),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_475),
.B(n_418),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_536),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_538),
.B(n_213),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_538),
.B(n_253),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_543),
.B(n_202),
.Y(n_619)
);

AND2x4_ASAP7_75t_SL g620 ( 
.A(n_527),
.B(n_412),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_475),
.B(n_418),
.Y(n_621)
);

INVx2_ASAP7_75t_SL g622 ( 
.A(n_490),
.Y(n_622)
);

AOI22xp5_ASAP7_75t_L g623 ( 
.A1(n_453),
.A2(n_544),
.B1(n_540),
.B2(n_516),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_510),
.B(n_203),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_572),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_490),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_542),
.B(n_260),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_476),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_476),
.B(n_418),
.Y(n_629)
);

BUFx5_ASAP7_75t_L g630 ( 
.A(n_459),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_484),
.B(n_204),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_482),
.B(n_418),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_482),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_542),
.A2(n_288),
.B1(n_230),
.B2(n_259),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_488),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_491),
.B(n_208),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_488),
.Y(n_637)
);

OA22x2_ASAP7_75t_L g638 ( 
.A1(n_480),
.A2(n_212),
.B1(n_220),
.B2(n_190),
.Y(n_638)
);

AOI22xp33_ASAP7_75t_SL g639 ( 
.A1(n_455),
.A2(n_199),
.B1(n_173),
.B2(n_170),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_493),
.B(n_466),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_SL g641 ( 
.A(n_552),
.B(n_170),
.Y(n_641)
);

INVxp67_ASAP7_75t_L g642 ( 
.A(n_508),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_449),
.B(n_462),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_570),
.B(n_262),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_494),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_472),
.Y(n_646)
);

AOI22xp5_ASAP7_75t_L g647 ( 
.A1(n_524),
.A2(n_270),
.B1(n_265),
.B2(n_269),
.Y(n_647)
);

CKINVDCx14_ASAP7_75t_R g648 ( 
.A(n_505),
.Y(n_648)
);

O2A1O1Ixp33_ASAP7_75t_L g649 ( 
.A1(n_450),
.A2(n_415),
.B(n_212),
.C(n_179),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_494),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_559),
.B(n_287),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_491),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_511),
.B(n_428),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_472),
.B(n_428),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_460),
.B(n_209),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_566),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_566),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_472),
.B(n_428),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_463),
.B(n_428),
.Y(n_659)
);

NAND3x1_ASAP7_75t_L g660 ( 
.A(n_465),
.B(n_243),
.C(n_309),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_463),
.B(n_428),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_527),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_551),
.B(n_228),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_503),
.Y(n_664)
);

BUFx3_ASAP7_75t_L g665 ( 
.A(n_584),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_455),
.B(n_233),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_566),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_567),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_573),
.B(n_289),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_463),
.B(n_165),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_503),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_527),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_455),
.B(n_255),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_567),
.Y(n_674)
);

OR2x2_ASAP7_75t_L g675 ( 
.A(n_520),
.B(n_256),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_463),
.B(n_450),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_512),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_512),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_483),
.B(n_267),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_458),
.B(n_165),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_458),
.B(n_461),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_485),
.B(n_271),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_SL g683 ( 
.A1(n_455),
.A2(n_173),
.B1(n_199),
.B2(n_181),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_461),
.B(n_171),
.Y(n_684)
);

OAI22xp33_ASAP7_75t_L g685 ( 
.A1(n_524),
.A2(n_214),
.B1(n_171),
.B2(n_259),
.Y(n_685)
);

OAI22xp33_ASAP7_75t_SL g686 ( 
.A1(n_467),
.A2(n_181),
.B1(n_191),
.B2(n_198),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_567),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_471),
.B(n_191),
.Y(n_688)
);

AOI22xp33_ASAP7_75t_L g689 ( 
.A1(n_514),
.A2(n_281),
.B1(n_198),
.B2(n_288),
.Y(n_689)
);

AOI22xp5_ASAP7_75t_L g690 ( 
.A1(n_559),
.A2(n_293),
.B1(n_247),
.B2(n_235),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_469),
.B(n_272),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_471),
.B(n_214),
.Y(n_692)
);

INVx2_ASAP7_75t_SL g693 ( 
.A(n_586),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_504),
.B(n_276),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_513),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_459),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_560),
.B(n_333),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_560),
.B(n_336),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_513),
.B(n_219),
.Y(n_699)
);

NAND3xp33_ASAP7_75t_L g700 ( 
.A(n_486),
.B(n_509),
.C(n_478),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_496),
.Y(n_701)
);

AND2x4_ASAP7_75t_SL g702 ( 
.A(n_584),
.B(n_173),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_518),
.B(n_229),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_459),
.B(n_229),
.Y(n_704)
);

AO22x1_ASAP7_75t_L g705 ( 
.A1(n_514),
.A2(n_309),
.B1(n_275),
.B2(n_274),
.Y(n_705)
);

A2O1A1Ixp33_ASAP7_75t_L g706 ( 
.A1(n_518),
.A2(n_284),
.B(n_299),
.C(n_281),
.Y(n_706)
);

NAND3xp33_ASAP7_75t_L g707 ( 
.A(n_495),
.B(n_291),
.C(n_302),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_496),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_521),
.B(n_230),
.Y(n_709)
);

AOI22xp33_ASAP7_75t_L g710 ( 
.A1(n_514),
.A2(n_247),
.B1(n_299),
.B2(n_263),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_521),
.B(n_235),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_583),
.Y(n_712)
);

INVx1_ASAP7_75t_SL g713 ( 
.A(n_451),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_528),
.B(n_246),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_465),
.B(n_279),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_528),
.B(n_246),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_447),
.B(n_263),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_584),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_535),
.B(n_282),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_531),
.B(n_284),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_583),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_531),
.Y(n_722)
);

INVx1_ASAP7_75t_SL g723 ( 
.A(n_550),
.Y(n_723)
);

BUFx2_ASAP7_75t_L g724 ( 
.A(n_550),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_533),
.B(n_417),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_447),
.B(n_285),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_447),
.B(n_401),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_533),
.Y(n_728)
);

OAI22xp33_ASAP7_75t_L g729 ( 
.A1(n_456),
.A2(n_303),
.B1(n_176),
.B2(n_179),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_447),
.B(n_401),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_496),
.Y(n_731)
);

NAND2xp33_ASAP7_75t_L g732 ( 
.A(n_514),
.B(n_534),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_514),
.A2(n_304),
.B1(n_187),
.B2(n_189),
.Y(n_733)
);

INVx3_ASAP7_75t_L g734 ( 
.A(n_584),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_534),
.B(n_417),
.Y(n_735)
);

AOI22xp5_ASAP7_75t_L g736 ( 
.A1(n_553),
.A2(n_199),
.B1(n_286),
.B2(n_295),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_555),
.B(n_301),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_555),
.B(n_417),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_537),
.B(n_305),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_564),
.B(n_402),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_583),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_557),
.B(n_307),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_564),
.B(n_402),
.Y(n_743)
);

HB1xp67_ASAP7_75t_L g744 ( 
.A(n_496),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_557),
.B(n_561),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_561),
.B(n_562),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_562),
.B(n_159),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_563),
.B(n_444),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_588),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_563),
.B(n_444),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_568),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_545),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_568),
.B(n_402),
.Y(n_753)
);

INVx8_ASAP7_75t_L g754 ( 
.A(n_553),
.Y(n_754)
);

NAND2xp33_ASAP7_75t_L g755 ( 
.A(n_514),
.B(n_376),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_588),
.Y(n_756)
);

NOR3xp33_ASAP7_75t_L g757 ( 
.A(n_589),
.B(n_308),
.C(n_220),
.Y(n_757)
);

A2O1A1Ixp33_ASAP7_75t_L g758 ( 
.A1(n_580),
.A2(n_189),
.B(n_257),
.C(n_275),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_580),
.B(n_444),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_582),
.B(n_402),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_582),
.B(n_444),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_577),
.Y(n_762)
);

OAI21xp33_ASAP7_75t_L g763 ( 
.A1(n_655),
.A2(n_303),
.B(n_296),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_628),
.Y(n_764)
);

INVx2_ASAP7_75t_SL g765 ( 
.A(n_693),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_676),
.A2(n_591),
.B(n_523),
.Y(n_766)
);

OAI21xp33_ASAP7_75t_L g767 ( 
.A1(n_655),
.A2(n_308),
.B(n_304),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_681),
.A2(n_591),
.B(n_523),
.Y(n_768)
);

AO21x1_ASAP7_75t_L g769 ( 
.A1(n_600),
.A2(n_610),
.B(n_601),
.Y(n_769)
);

INVx2_ASAP7_75t_SL g770 ( 
.A(n_713),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_727),
.A2(n_591),
.B(n_523),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_628),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_633),
.Y(n_773)
);

AOI21xp33_ASAP7_75t_L g774 ( 
.A1(n_663),
.A2(n_456),
.B(n_548),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_643),
.B(n_514),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_727),
.A2(n_591),
.B(n_477),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_633),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_730),
.A2(n_574),
.B(n_587),
.Y(n_778)
);

HB1xp67_ASAP7_75t_L g779 ( 
.A(n_622),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_616),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_762),
.B(n_457),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_730),
.A2(n_574),
.B(n_587),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_656),
.Y(n_783)
);

INVx4_ASAP7_75t_L g784 ( 
.A(n_754),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_732),
.A2(n_574),
.B(n_587),
.Y(n_785)
);

AND2x4_ASAP7_75t_L g786 ( 
.A(n_609),
.B(n_456),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_607),
.A2(n_574),
.B(n_587),
.Y(n_787)
);

OAI21xp5_ASAP7_75t_L g788 ( 
.A1(n_717),
.A2(n_501),
.B(n_502),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_640),
.B(n_457),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_755),
.A2(n_477),
.B(n_487),
.Y(n_790)
);

BUFx4f_ASAP7_75t_L g791 ( 
.A(n_754),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_696),
.A2(n_477),
.B(n_487),
.Y(n_792)
);

AOI22xp5_ASAP7_75t_L g793 ( 
.A1(n_640),
.A2(n_553),
.B1(n_576),
.B2(n_456),
.Y(n_793)
);

BUFx2_ASAP7_75t_L g794 ( 
.A(n_724),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_624),
.B(n_457),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_624),
.B(n_457),
.Y(n_796)
);

OAI22xp5_ASAP7_75t_L g797 ( 
.A1(n_623),
.A2(n_576),
.B1(n_553),
.B2(n_456),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_631),
.B(n_470),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_656),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_608),
.B(n_569),
.Y(n_800)
);

AOI22xp5_ASAP7_75t_L g801 ( 
.A1(n_726),
.A2(n_576),
.B1(n_581),
.B2(n_585),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_642),
.B(n_477),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_631),
.B(n_470),
.Y(n_803)
);

AOI22xp5_ASAP7_75t_L g804 ( 
.A1(n_726),
.A2(n_554),
.B1(n_470),
.B2(n_575),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_657),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_646),
.B(n_470),
.Y(n_806)
);

NOR2x1_ASAP7_75t_L g807 ( 
.A(n_665),
.B(n_487),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_646),
.B(n_473),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_635),
.B(n_473),
.Y(n_809)
);

A2O1A1Ixp33_ASAP7_75t_L g810 ( 
.A1(n_701),
.A2(n_296),
.B(n_565),
.C(n_546),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_696),
.A2(n_523),
.B(n_487),
.Y(n_811)
);

HB1xp67_ASAP7_75t_L g812 ( 
.A(n_626),
.Y(n_812)
);

INVx2_ASAP7_75t_SL g813 ( 
.A(n_675),
.Y(n_813)
);

AND2x4_ASAP7_75t_L g814 ( 
.A(n_652),
.B(n_590),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_637),
.B(n_473),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_645),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_619),
.B(n_473),
.Y(n_817)
);

OAI21xp5_ASAP7_75t_L g818 ( 
.A1(n_717),
.A2(n_501),
.B(n_452),
.Y(n_818)
);

NOR2x1_ASAP7_75t_L g819 ( 
.A(n_665),
.B(n_474),
.Y(n_819)
);

OAI21xp5_ASAP7_75t_L g820 ( 
.A1(n_704),
.A2(n_479),
.B(n_502),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_636),
.B(n_525),
.Y(n_821)
);

AOI21xp5_ASAP7_75t_L g822 ( 
.A1(n_653),
.A2(n_578),
.B(n_515),
.Y(n_822)
);

O2A1O1Ixp33_ASAP7_75t_L g823 ( 
.A1(n_600),
.A2(n_565),
.B(n_546),
.C(n_468),
.Y(n_823)
);

AND2x4_ASAP7_75t_L g824 ( 
.A(n_594),
.B(n_590),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_604),
.A2(n_743),
.B(n_740),
.Y(n_825)
);

OAI22xp5_ASAP7_75t_L g826 ( 
.A1(n_704),
.A2(n_590),
.B1(n_500),
.B2(n_575),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_740),
.A2(n_578),
.B(n_515),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_650),
.B(n_474),
.Y(n_828)
);

NAND2xp33_ASAP7_75t_L g829 ( 
.A(n_630),
.B(n_515),
.Y(n_829)
);

BUFx3_ASAP7_75t_L g830 ( 
.A(n_754),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_743),
.A2(n_578),
.B(n_515),
.Y(n_831)
);

BUFx6f_ASAP7_75t_L g832 ( 
.A(n_592),
.Y(n_832)
);

AOI22xp5_ASAP7_75t_L g833 ( 
.A1(n_651),
.A2(n_554),
.B1(n_575),
.B2(n_481),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_664),
.B(n_474),
.Y(n_834)
);

AO21x1_ASAP7_75t_L g835 ( 
.A1(n_601),
.A2(n_558),
.B(n_556),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_671),
.Y(n_836)
);

INVx2_ASAP7_75t_SL g837 ( 
.A(n_612),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_619),
.B(n_525),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_613),
.A2(n_578),
.B(n_515),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_677),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_678),
.B(n_474),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_695),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_659),
.A2(n_578),
.B(n_532),
.Y(n_843)
);

OAI21xp5_ASAP7_75t_L g844 ( 
.A1(n_610),
.A2(n_499),
.B(n_452),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_661),
.A2(n_578),
.B(n_515),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_654),
.A2(n_547),
.B(n_571),
.Y(n_846)
);

O2A1O1Ixp33_ASAP7_75t_SL g847 ( 
.A1(n_685),
.A2(n_546),
.B(n_565),
.C(n_468),
.Y(n_847)
);

AO21x1_ASAP7_75t_L g848 ( 
.A1(n_651),
.A2(n_558),
.B(n_556),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_658),
.A2(n_597),
.B(n_680),
.Y(n_849)
);

AOI21xp33_ASAP7_75t_L g850 ( 
.A1(n_663),
.A2(n_682),
.B(n_679),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_722),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_744),
.B(n_481),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_630),
.B(n_532),
.Y(n_853)
);

AO21x1_ASAP7_75t_L g854 ( 
.A1(n_684),
.A2(n_526),
.B(n_529),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_708),
.B(n_481),
.Y(n_855)
);

OAI21xp5_ASAP7_75t_L g856 ( 
.A1(n_688),
.A2(n_497),
.B(n_499),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_692),
.A2(n_532),
.B(n_571),
.Y(n_857)
);

AOI21x1_ASAP7_75t_L g858 ( 
.A1(n_753),
.A2(n_479),
.B(n_497),
.Y(n_858)
);

CKINVDCx20_ASAP7_75t_R g859 ( 
.A(n_602),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_697),
.A2(n_532),
.B(n_571),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_697),
.A2(n_532),
.B(n_571),
.Y(n_861)
);

OAI21xp5_ASAP7_75t_L g862 ( 
.A1(n_698),
.A2(n_746),
.B(n_745),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_728),
.B(n_751),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_599),
.B(n_481),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_731),
.B(n_498),
.Y(n_865)
);

O2A1O1Ixp5_ASAP7_75t_L g866 ( 
.A1(n_598),
.A2(n_529),
.B(n_526),
.C(n_464),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_749),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_715),
.B(n_498),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_L g869 ( 
.A(n_700),
.B(n_498),
.Y(n_869)
);

AOI21x1_ASAP7_75t_L g870 ( 
.A1(n_753),
.A2(n_464),
.B(n_454),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_698),
.A2(n_532),
.B(n_571),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_749),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_599),
.B(n_498),
.Y(n_873)
);

OAI321xp33_ASAP7_75t_L g874 ( 
.A1(n_679),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_8),
.C(n_9),
.Y(n_874)
);

INVx2_ASAP7_75t_L g875 ( 
.A(n_667),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_667),
.Y(n_876)
);

O2A1O1Ixp5_ASAP7_75t_L g877 ( 
.A1(n_598),
.A2(n_454),
.B(n_448),
.C(n_468),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_756),
.Y(n_878)
);

INVx4_ASAP7_75t_L g879 ( 
.A(n_718),
.Y(n_879)
);

INVx1_ASAP7_75t_SL g880 ( 
.A(n_723),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_615),
.A2(n_571),
.B(n_547),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_L g882 ( 
.A1(n_682),
.A2(n_554),
.B1(n_575),
.B2(n_549),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_666),
.B(n_517),
.Y(n_883)
);

HB1xp67_ASAP7_75t_L g884 ( 
.A(n_599),
.Y(n_884)
);

OAI321xp33_ASAP7_75t_L g885 ( 
.A1(n_729),
.A2(n_719),
.A3(n_736),
.B1(n_690),
.B2(n_691),
.C(n_739),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_621),
.A2(n_547),
.B(n_549),
.Y(n_886)
);

CKINVDCx5p33_ASAP7_75t_R g887 ( 
.A(n_662),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_673),
.B(n_517),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_756),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_603),
.Y(n_890)
);

OAI21xp5_ASAP7_75t_L g891 ( 
.A1(n_670),
.A2(n_448),
.B(n_517),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_737),
.B(n_549),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_617),
.B(n_549),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_603),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_629),
.A2(n_547),
.B(n_539),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_668),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_L g897 ( 
.A(n_617),
.B(n_539),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_625),
.Y(n_898)
);

AO21x2_ASAP7_75t_L g899 ( 
.A1(n_596),
.A2(n_448),
.B(n_507),
.Y(n_899)
);

OAI22xp5_ASAP7_75t_L g900 ( 
.A1(n_734),
.A2(n_500),
.B1(n_539),
.B2(n_547),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_668),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_737),
.B(n_539),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_674),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_742),
.B(n_500),
.Y(n_904)
);

CKINVDCx8_ASAP7_75t_R g905 ( 
.A(n_672),
.Y(n_905)
);

AOI22x1_ASAP7_75t_L g906 ( 
.A1(n_625),
.A2(n_721),
.B1(n_687),
.B2(n_712),
.Y(n_906)
);

AOI21x1_ASAP7_75t_L g907 ( 
.A1(n_760),
.A2(n_507),
.B(n_441),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_674),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_644),
.B(n_500),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_687),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_712),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_632),
.A2(n_547),
.B(n_402),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_742),
.B(n_507),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_725),
.A2(n_402),
.B(n_441),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_735),
.A2(n_402),
.B(n_441),
.Y(n_915)
);

NOR2xp67_ASAP7_75t_L g916 ( 
.A(n_611),
.B(n_147),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_738),
.A2(n_402),
.B(n_441),
.Y(n_917)
);

AOI21xp5_ASAP7_75t_L g918 ( 
.A1(n_748),
.A2(n_432),
.B(n_424),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_721),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_734),
.B(n_554),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_750),
.A2(n_432),
.B(n_424),
.Y(n_921)
);

INVx11_ASAP7_75t_L g922 ( 
.A(n_605),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_759),
.A2(n_432),
.B(n_424),
.Y(n_923)
);

AOI21x1_ASAP7_75t_L g924 ( 
.A1(n_760),
.A2(n_432),
.B(n_424),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_630),
.B(n_718),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_630),
.B(n_554),
.Y(n_926)
);

OAI21xp5_ASAP7_75t_L g927 ( 
.A1(n_741),
.A2(n_554),
.B(n_421),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_761),
.A2(n_596),
.B(n_627),
.Y(n_928)
);

AOI22xp33_ASAP7_75t_L g929 ( 
.A1(n_638),
.A2(n_630),
.B1(n_733),
.B2(n_741),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_630),
.B(n_376),
.Y(n_930)
);

OR2x2_ASAP7_75t_L g931 ( 
.A(n_752),
.B(n_0),
.Y(n_931)
);

BUFx2_ASAP7_75t_L g932 ( 
.A(n_660),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_618),
.A2(n_421),
.B(n_420),
.Y(n_933)
);

AND2x4_ASAP7_75t_L g934 ( 
.A(n_620),
.B(n_145),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_699),
.B(n_421),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_618),
.A2(n_420),
.B(n_417),
.Y(n_936)
);

O2A1O1Ixp5_ASAP7_75t_L g937 ( 
.A1(n_703),
.A2(n_420),
.B(n_376),
.C(n_10),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_592),
.Y(n_938)
);

AND2x4_ASAP7_75t_L g939 ( 
.A(n_620),
.B(n_100),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_647),
.A2(n_139),
.B1(n_130),
.B2(n_128),
.Y(n_940)
);

AOI21x1_ASAP7_75t_L g941 ( 
.A1(n_709),
.A2(n_124),
.B(n_122),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_627),
.A2(n_88),
.B(n_85),
.Y(n_942)
);

OAI22xp5_ASAP7_75t_L g943 ( 
.A1(n_634),
.A2(n_80),
.B1(n_70),
.B2(n_65),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_711),
.B(n_2),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_669),
.B(n_8),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_714),
.B(n_10),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_716),
.B(n_11),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_720),
.Y(n_948)
);

OAI21xp5_ASAP7_75t_L g949 ( 
.A1(n_614),
.A2(n_12),
.B(n_13),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_800),
.B(n_719),
.Y(n_950)
);

O2A1O1Ixp33_ASAP7_75t_SL g951 ( 
.A1(n_850),
.A2(n_706),
.B(n_747),
.C(n_649),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_R g952 ( 
.A(n_887),
.B(n_648),
.Y(n_952)
);

OAI22xp5_ASAP7_75t_L g953 ( 
.A1(n_868),
.A2(n_592),
.B1(n_593),
.B2(n_606),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_SL g954 ( 
.A(n_885),
.B(n_702),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_800),
.B(n_694),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_829),
.A2(n_593),
.B(n_606),
.Y(n_956)
);

INVx8_ASAP7_75t_L g957 ( 
.A(n_832),
.Y(n_957)
);

INVx3_ASAP7_75t_L g958 ( 
.A(n_832),
.Y(n_958)
);

O2A1O1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_945),
.A2(n_686),
.B(n_595),
.C(n_758),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_775),
.A2(n_593),
.B(n_606),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_948),
.B(n_702),
.Y(n_961)
);

AND2x2_ASAP7_75t_SL g962 ( 
.A(n_791),
.B(n_641),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_880),
.B(n_605),
.Y(n_963)
);

OAI22xp5_ASAP7_75t_SL g964 ( 
.A1(n_859),
.A2(n_639),
.B1(n_683),
.B2(n_707),
.Y(n_964)
);

O2A1O1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_949),
.A2(n_757),
.B(n_710),
.C(n_689),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_770),
.B(n_638),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_764),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_825),
.A2(n_705),
.B(n_17),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_813),
.B(n_16),
.Y(n_969)
);

OR2x6_ASAP7_75t_L g970 ( 
.A(n_794),
.B(n_16),
.Y(n_970)
);

OAI22xp5_ASAP7_75t_L g971 ( 
.A1(n_868),
.A2(n_17),
.B1(n_20),
.B2(n_21),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_799),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_779),
.B(n_20),
.Y(n_973)
);

BUFx2_ASAP7_75t_L g974 ( 
.A(n_932),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_821),
.B(n_884),
.Y(n_975)
);

OAI22xp5_ASAP7_75t_L g976 ( 
.A1(n_884),
.A2(n_793),
.B1(n_801),
.B2(n_817),
.Y(n_976)
);

AOI22xp5_ASAP7_75t_L g977 ( 
.A1(n_945),
.A2(n_22),
.B1(n_25),
.B2(n_26),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_849),
.A2(n_803),
.B(n_798),
.Y(n_978)
);

HB1xp67_ASAP7_75t_L g979 ( 
.A(n_779),
.Y(n_979)
);

BUFx12f_ASAP7_75t_L g980 ( 
.A(n_765),
.Y(n_980)
);

AOI22x1_ASAP7_75t_L g981 ( 
.A1(n_928),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_869),
.A2(n_30),
.B(n_34),
.C(n_35),
.Y(n_982)
);

AO22x1_ASAP7_75t_L g983 ( 
.A1(n_934),
.A2(n_58),
.B1(n_35),
.B2(n_37),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_L g984 ( 
.A1(n_817),
.A2(n_34),
.B1(n_40),
.B2(n_41),
.Y(n_984)
);

BUFx12f_ASAP7_75t_L g985 ( 
.A(n_837),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_786),
.B(n_40),
.Y(n_986)
);

CKINVDCx20_ASAP7_75t_R g987 ( 
.A(n_905),
.Y(n_987)
);

NOR3xp33_ASAP7_75t_L g988 ( 
.A(n_874),
.B(n_41),
.C(n_42),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_812),
.B(n_43),
.Y(n_989)
);

CKINVDCx20_ASAP7_75t_R g990 ( 
.A(n_830),
.Y(n_990)
);

NAND2x1p5_ASAP7_75t_L g991 ( 
.A(n_784),
.B(n_44),
.Y(n_991)
);

AO21x1_ASAP7_75t_L g992 ( 
.A1(n_869),
.A2(n_46),
.B(n_47),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_838),
.B(n_47),
.Y(n_993)
);

A2O1A1Ixp33_ASAP7_75t_L g994 ( 
.A1(n_893),
.A2(n_48),
.B(n_52),
.C(n_55),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_863),
.B(n_883),
.Y(n_995)
);

BUFx8_ASAP7_75t_SL g996 ( 
.A(n_791),
.Y(n_996)
);

AO21x2_ASAP7_75t_L g997 ( 
.A1(n_854),
.A2(n_56),
.B(n_774),
.Y(n_997)
);

BUFx4f_ASAP7_75t_L g998 ( 
.A(n_832),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_893),
.A2(n_897),
.B(n_862),
.C(n_767),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_799),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_R g1001 ( 
.A(n_830),
.B(n_56),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_922),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_929),
.A2(n_873),
.B1(n_864),
.B2(n_789),
.Y(n_1003)
);

A2O1A1Ixp33_ASAP7_75t_L g1004 ( 
.A1(n_897),
.A2(n_763),
.B(n_888),
.C(n_909),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_772),
.Y(n_1005)
);

HB1xp67_ASAP7_75t_L g1006 ( 
.A(n_812),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_931),
.B(n_802),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_802),
.B(n_816),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_773),
.Y(n_1009)
);

BUFx2_ASAP7_75t_L g1010 ( 
.A(n_934),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_836),
.B(n_840),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_784),
.B(n_786),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_879),
.B(n_939),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_777),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_842),
.B(n_851),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_780),
.B(n_814),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_867),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_814),
.B(n_852),
.Y(n_1018)
);

HB1xp67_ASAP7_75t_L g1019 ( 
.A(n_939),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_872),
.Y(n_1020)
);

OR2x2_ASAP7_75t_L g1021 ( 
.A(n_944),
.B(n_946),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_878),
.Y(n_1022)
);

NOR2xp33_ASAP7_75t_L g1023 ( 
.A(n_879),
.B(n_852),
.Y(n_1023)
);

AOI22xp33_ASAP7_75t_L g1024 ( 
.A1(n_916),
.A2(n_769),
.B1(n_947),
.B2(n_797),
.Y(n_1024)
);

OAI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_929),
.A2(n_795),
.B1(n_796),
.B2(n_892),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_902),
.A2(n_904),
.B(n_822),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_805),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_913),
.B(n_781),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_785),
.A2(n_857),
.B(n_787),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_R g1030 ( 
.A(n_832),
.B(n_938),
.Y(n_1030)
);

AOI22x1_ASAP7_75t_L g1031 ( 
.A1(n_933),
.A2(n_936),
.B1(n_910),
.B2(n_908),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_768),
.A2(n_853),
.B(n_790),
.Y(n_1032)
);

OR2x2_ASAP7_75t_L g1033 ( 
.A(n_889),
.B(n_890),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_855),
.B(n_865),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_SL g1035 ( 
.A(n_938),
.B(n_824),
.Y(n_1035)
);

INVx4_ASAP7_75t_L g1036 ( 
.A(n_938),
.Y(n_1036)
);

INVx2_ASAP7_75t_SL g1037 ( 
.A(n_938),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_853),
.A2(n_839),
.B(n_766),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_894),
.B(n_898),
.Y(n_1039)
);

NOR2xp67_ASAP7_75t_L g1040 ( 
.A(n_942),
.B(n_909),
.Y(n_1040)
);

O2A1O1Ixp33_ASAP7_75t_L g1041 ( 
.A1(n_810),
.A2(n_940),
.B(n_847),
.C(n_937),
.Y(n_1041)
);

NOR3xp33_ASAP7_75t_SL g1042 ( 
.A(n_810),
.B(n_943),
.C(n_925),
.Y(n_1042)
);

INVx4_ASAP7_75t_L g1043 ( 
.A(n_824),
.Y(n_1043)
);

NOR3xp33_ASAP7_75t_SL g1044 ( 
.A(n_809),
.B(n_834),
.C(n_815),
.Y(n_1044)
);

AOI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_819),
.A2(n_882),
.B1(n_833),
.B2(n_848),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_930),
.A2(n_843),
.B(n_845),
.Y(n_1046)
);

OR2x2_ASAP7_75t_L g1047 ( 
.A(n_783),
.B(n_911),
.Y(n_1047)
);

O2A1O1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_847),
.A2(n_937),
.B(n_828),
.C(n_841),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_919),
.Y(n_1049)
);

O2A1O1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_805),
.A2(n_875),
.B(n_903),
.C(n_901),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_930),
.A2(n_771),
.B(n_776),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_SL g1052 ( 
.A(n_807),
.B(n_876),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_875),
.B(n_876),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_778),
.A2(n_782),
.B(n_856),
.Y(n_1054)
);

OAI22x1_ASAP7_75t_L g1055 ( 
.A1(n_906),
.A2(n_903),
.B1(n_901),
.B2(n_896),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_896),
.Y(n_1056)
);

AOI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_926),
.A2(n_920),
.B1(n_804),
.B2(n_835),
.Y(n_1057)
);

A2O1A1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_823),
.A2(n_927),
.B(n_866),
.C(n_877),
.Y(n_1058)
);

INVx2_ASAP7_75t_SL g1059 ( 
.A(n_899),
.Y(n_1059)
);

O2A1O1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_826),
.A2(n_935),
.B(n_866),
.C(n_877),
.Y(n_1060)
);

BUFx6f_ASAP7_75t_L g1061 ( 
.A(n_941),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_846),
.A2(n_881),
.B(n_891),
.Y(n_1062)
);

OAI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_806),
.A2(n_808),
.B1(n_900),
.B2(n_827),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_860),
.B(n_861),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_858),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_918),
.Y(n_1066)
);

INVx4_ASAP7_75t_L g1067 ( 
.A(n_899),
.Y(n_1067)
);

O2A1O1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_844),
.A2(n_820),
.B(n_788),
.C(n_818),
.Y(n_1068)
);

BUFx3_ASAP7_75t_L g1069 ( 
.A(n_871),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_792),
.A2(n_811),
.B(n_895),
.Y(n_1070)
);

INVxp67_ASAP7_75t_L g1071 ( 
.A(n_831),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_886),
.A2(n_912),
.B(n_915),
.Y(n_1072)
);

AOI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_921),
.A2(n_923),
.B1(n_914),
.B2(n_917),
.Y(n_1073)
);

INVx6_ASAP7_75t_L g1074 ( 
.A(n_924),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_870),
.Y(n_1075)
);

INVx3_ASAP7_75t_L g1076 ( 
.A(n_907),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_SL g1077 ( 
.A(n_850),
.B(n_643),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_829),
.A2(n_775),
.B(n_825),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_887),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_764),
.Y(n_1080)
);

BUFx6f_ASAP7_75t_L g1081 ( 
.A(n_832),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_850),
.B(n_643),
.Y(n_1082)
);

OR2x2_ASAP7_75t_L g1083 ( 
.A(n_880),
.B(n_451),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_829),
.A2(n_775),
.B(n_825),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_800),
.B(n_643),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_764),
.Y(n_1086)
);

OAI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_850),
.A2(n_643),
.B1(n_868),
.B2(n_884),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_800),
.B(n_643),
.Y(n_1088)
);

BUFx2_ASAP7_75t_L g1089 ( 
.A(n_794),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_800),
.B(n_643),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_800),
.B(n_643),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_887),
.Y(n_1092)
);

OAI21x1_ASAP7_75t_L g1093 ( 
.A1(n_1029),
.A2(n_1070),
.B(n_1046),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_978),
.A2(n_1054),
.B(n_1026),
.Y(n_1094)
);

AOI221xp5_ASAP7_75t_L g1095 ( 
.A1(n_1082),
.A2(n_950),
.B1(n_955),
.B2(n_1091),
.C(n_1090),
.Y(n_1095)
);

AO21x1_ASAP7_75t_L g1096 ( 
.A1(n_1087),
.A2(n_954),
.B(n_1077),
.Y(n_1096)
);

AO22x2_ASAP7_75t_L g1097 ( 
.A1(n_988),
.A2(n_976),
.B1(n_971),
.B2(n_984),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_1007),
.B(n_1085),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_978),
.A2(n_1054),
.B(n_1026),
.Y(n_1099)
);

INVx5_ASAP7_75t_L g1100 ( 
.A(n_957),
.Y(n_1100)
);

NOR2x1_ASAP7_75t_L g1101 ( 
.A(n_1088),
.B(n_1034),
.Y(n_1101)
);

OAI21x1_ASAP7_75t_L g1102 ( 
.A1(n_1029),
.A2(n_1070),
.B(n_1046),
.Y(n_1102)
);

A2O1A1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_965),
.A2(n_959),
.B(n_999),
.C(n_1041),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_1015),
.Y(n_1104)
);

AO31x2_ASAP7_75t_L g1105 ( 
.A1(n_1025),
.A2(n_1062),
.A3(n_1067),
.B(n_1058),
.Y(n_1105)
);

AND2x4_ASAP7_75t_L g1106 ( 
.A(n_1012),
.B(n_1010),
.Y(n_1106)
);

OAI21x1_ASAP7_75t_L g1107 ( 
.A1(n_1038),
.A2(n_1032),
.B(n_1031),
.Y(n_1107)
);

OR2x2_ASAP7_75t_L g1108 ( 
.A(n_1083),
.B(n_1089),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_961),
.B(n_964),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_1078),
.A2(n_1084),
.B(n_1032),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1049),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1033),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_1079),
.Y(n_1113)
);

AO31x2_ASAP7_75t_L g1114 ( 
.A1(n_1078),
.A2(n_1084),
.A3(n_1072),
.B(n_1063),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_1051),
.A2(n_1072),
.B(n_960),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_1028),
.A2(n_1040),
.B(n_1051),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_960),
.A2(n_1076),
.B(n_1050),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_974),
.B(n_1021),
.Y(n_1118)
);

AND2x4_ASAP7_75t_L g1119 ( 
.A(n_1012),
.B(n_1019),
.Y(n_1119)
);

OR2x2_ASAP7_75t_L g1120 ( 
.A(n_975),
.B(n_979),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1017),
.Y(n_1121)
);

OR2x2_ASAP7_75t_L g1122 ( 
.A(n_1006),
.B(n_1016),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_1023),
.B(n_1011),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_1092),
.Y(n_1124)
);

CKINVDCx11_ASAP7_75t_R g1125 ( 
.A(n_987),
.Y(n_1125)
);

INVx3_ASAP7_75t_L g1126 ( 
.A(n_1081),
.Y(n_1126)
);

OA21x2_ASAP7_75t_L g1127 ( 
.A1(n_1004),
.A2(n_1024),
.B(n_968),
.Y(n_1127)
);

AND2x4_ASAP7_75t_L g1128 ( 
.A(n_1013),
.B(n_1036),
.Y(n_1128)
);

INVx3_ASAP7_75t_L g1129 ( 
.A(n_1081),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1020),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_962),
.B(n_986),
.Y(n_1131)
);

AO31x2_ASAP7_75t_L g1132 ( 
.A1(n_968),
.A2(n_1003),
.A3(n_992),
.B(n_1055),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_995),
.A2(n_1008),
.B1(n_965),
.B2(n_1018),
.Y(n_1133)
);

OAI21x1_ASAP7_75t_L g1134 ( 
.A1(n_1076),
.A2(n_1050),
.B(n_956),
.Y(n_1134)
);

AO31x2_ASAP7_75t_L g1135 ( 
.A1(n_1065),
.A2(n_1075),
.A3(n_953),
.B(n_994),
.Y(n_1135)
);

OAI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_1071),
.A2(n_1057),
.B(n_1048),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1068),
.A2(n_956),
.B(n_1064),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1060),
.A2(n_951),
.B(n_1066),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_989),
.B(n_966),
.Y(n_1139)
);

BUFx2_ASAP7_75t_L g1140 ( 
.A(n_990),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1069),
.A2(n_1045),
.B(n_1052),
.Y(n_1141)
);

AO21x1_ASAP7_75t_L g1142 ( 
.A1(n_993),
.A2(n_1039),
.B(n_977),
.Y(n_1142)
);

NAND3xp33_ASAP7_75t_L g1143 ( 
.A(n_982),
.B(n_981),
.C(n_969),
.Y(n_1143)
);

OAI21x1_ASAP7_75t_L g1144 ( 
.A1(n_1073),
.A2(n_1053),
.B(n_1056),
.Y(n_1144)
);

OR2x2_ASAP7_75t_L g1145 ( 
.A(n_1005),
.B(n_1014),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1035),
.A2(n_1059),
.B(n_998),
.Y(n_1146)
);

INVx2_ASAP7_75t_SL g1147 ( 
.A(n_980),
.Y(n_1147)
);

BUFx2_ASAP7_75t_L g1148 ( 
.A(n_985),
.Y(n_1148)
);

INVxp67_ASAP7_75t_L g1149 ( 
.A(n_973),
.Y(n_1149)
);

INVx5_ASAP7_75t_L g1150 ( 
.A(n_957),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1022),
.Y(n_1151)
);

BUFx2_ASAP7_75t_L g1152 ( 
.A(n_970),
.Y(n_1152)
);

OAI21x1_ASAP7_75t_L g1153 ( 
.A1(n_972),
.A2(n_1027),
.B(n_1000),
.Y(n_1153)
);

NOR2xp67_ASAP7_75t_L g1154 ( 
.A(n_1036),
.B(n_1043),
.Y(n_1154)
);

O2A1O1Ixp33_ASAP7_75t_SL g1155 ( 
.A1(n_1009),
.A2(n_1086),
.B(n_1080),
.C(n_1047),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1043),
.Y(n_1156)
);

OR2x2_ASAP7_75t_L g1157 ( 
.A(n_963),
.B(n_1037),
.Y(n_1157)
);

OAI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1042),
.A2(n_1044),
.B(n_998),
.Y(n_1158)
);

AO21x1_ASAP7_75t_L g1159 ( 
.A1(n_991),
.A2(n_997),
.B(n_1061),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1074),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_970),
.B(n_952),
.Y(n_1161)
);

AO31x2_ASAP7_75t_L g1162 ( 
.A1(n_997),
.A2(n_1061),
.A3(n_1074),
.B(n_983),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_958),
.A2(n_991),
.B(n_1074),
.Y(n_1163)
);

OAI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_958),
.A2(n_970),
.B(n_1061),
.Y(n_1164)
);

AO31x2_ASAP7_75t_L g1165 ( 
.A1(n_1030),
.A2(n_957),
.A3(n_1001),
.B(n_1081),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_L g1166 ( 
.A(n_996),
.B(n_1002),
.Y(n_1166)
);

AO31x2_ASAP7_75t_L g1167 ( 
.A1(n_999),
.A2(n_854),
.A3(n_1025),
.B(n_1054),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_1085),
.B(n_1088),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_978),
.A2(n_829),
.B(n_1054),
.Y(n_1169)
);

NAND3xp33_ASAP7_75t_SL g1170 ( 
.A(n_950),
.B(n_438),
.C(n_404),
.Y(n_1170)
);

BUFx3_ASAP7_75t_L g1171 ( 
.A(n_1089),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_1085),
.B(n_1088),
.Y(n_1172)
);

OR2x2_ASAP7_75t_L g1173 ( 
.A(n_955),
.B(n_451),
.Y(n_1173)
);

OAI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1082),
.A2(n_850),
.B(n_999),
.Y(n_1174)
);

BUFx3_ASAP7_75t_L g1175 ( 
.A(n_1089),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_978),
.A2(n_829),
.B(n_1054),
.Y(n_1176)
);

OR2x2_ASAP7_75t_L g1177 ( 
.A(n_955),
.B(n_451),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1029),
.A2(n_1070),
.B(n_1046),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_978),
.A2(n_829),
.B(n_1054),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_978),
.A2(n_829),
.B(n_1054),
.Y(n_1180)
);

A2O1A1Ixp33_ASAP7_75t_L g1181 ( 
.A1(n_1082),
.A2(n_850),
.B(n_950),
.C(n_1085),
.Y(n_1181)
);

OR2x2_ASAP7_75t_L g1182 ( 
.A(n_955),
.B(n_451),
.Y(n_1182)
);

AOI221x1_ASAP7_75t_L g1183 ( 
.A1(n_988),
.A2(n_850),
.B1(n_1082),
.B2(n_976),
.C(n_1087),
.Y(n_1183)
);

AOI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1082),
.A2(n_950),
.B1(n_850),
.B2(n_1085),
.Y(n_1184)
);

INVxp67_ASAP7_75t_L g1185 ( 
.A(n_1083),
.Y(n_1185)
);

INVxp67_ASAP7_75t_L g1186 ( 
.A(n_1083),
.Y(n_1186)
);

AND2x2_ASAP7_75t_L g1187 ( 
.A(n_1007),
.B(n_522),
.Y(n_1187)
);

AND2x2_ASAP7_75t_SL g1188 ( 
.A(n_988),
.B(n_506),
.Y(n_1188)
);

NAND2x1p5_ASAP7_75t_L g1189 ( 
.A(n_998),
.B(n_1036),
.Y(n_1189)
);

AND2x4_ASAP7_75t_L g1190 ( 
.A(n_1012),
.B(n_1010),
.Y(n_1190)
);

INVxp67_ASAP7_75t_SL g1191 ( 
.A(n_979),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1029),
.A2(n_1070),
.B(n_1046),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_978),
.A2(n_829),
.B(n_1054),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_978),
.A2(n_829),
.B(n_1054),
.Y(n_1194)
);

BUFx3_ASAP7_75t_L g1195 ( 
.A(n_1089),
.Y(n_1195)
);

INVx3_ASAP7_75t_L g1196 ( 
.A(n_1081),
.Y(n_1196)
);

BUFx8_ASAP7_75t_L g1197 ( 
.A(n_1089),
.Y(n_1197)
);

A2O1A1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_1082),
.A2(n_850),
.B(n_950),
.C(n_1085),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_978),
.A2(n_829),
.B(n_1054),
.Y(n_1199)
);

AOI221xp5_ASAP7_75t_SL g1200 ( 
.A1(n_1085),
.A2(n_1088),
.B1(n_1091),
.B2(n_1090),
.C(n_971),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1085),
.B(n_1088),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_978),
.A2(n_829),
.B(n_1054),
.Y(n_1202)
);

AO31x2_ASAP7_75t_L g1203 ( 
.A1(n_999),
.A2(n_854),
.A3(n_1025),
.B(n_1054),
.Y(n_1203)
);

AOI22xp5_ASAP7_75t_L g1204 ( 
.A1(n_1082),
.A2(n_950),
.B1(n_850),
.B2(n_1085),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_1029),
.A2(n_1070),
.B(n_1046),
.Y(n_1205)
);

INVx4_ASAP7_75t_L g1206 ( 
.A(n_957),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_978),
.A2(n_829),
.B(n_1054),
.Y(n_1207)
);

AOI221xp5_ASAP7_75t_SL g1208 ( 
.A1(n_1085),
.A2(n_1088),
.B1(n_1091),
.B2(n_1090),
.C(n_971),
.Y(n_1208)
);

AOI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1082),
.A2(n_950),
.B1(n_850),
.B2(n_1085),
.Y(n_1209)
);

AOI221x1_ASAP7_75t_L g1210 ( 
.A1(n_988),
.A2(n_850),
.B1(n_1082),
.B2(n_976),
.C(n_1087),
.Y(n_1210)
);

AOI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1082),
.A2(n_950),
.B1(n_850),
.B2(n_1085),
.Y(n_1211)
);

OAI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1082),
.A2(n_850),
.B(n_999),
.Y(n_1212)
);

AOI31xp67_ASAP7_75t_L g1213 ( 
.A1(n_1064),
.A2(n_1073),
.A3(n_1045),
.B(n_1077),
.Y(n_1213)
);

INVx5_ASAP7_75t_L g1214 ( 
.A(n_957),
.Y(n_1214)
);

AND2x2_ASAP7_75t_L g1215 ( 
.A(n_1007),
.B(n_522),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1015),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1029),
.A2(n_1070),
.B(n_1046),
.Y(n_1217)
);

AO31x2_ASAP7_75t_L g1218 ( 
.A1(n_999),
.A2(n_854),
.A3(n_1025),
.B(n_1054),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_978),
.A2(n_829),
.B(n_1054),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1085),
.B(n_1088),
.Y(n_1220)
);

BUFx12f_ASAP7_75t_L g1221 ( 
.A(n_1002),
.Y(n_1221)
);

AOI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1082),
.A2(n_950),
.B1(n_850),
.B2(n_1085),
.Y(n_1222)
);

AOI221x1_ASAP7_75t_L g1223 ( 
.A1(n_988),
.A2(n_850),
.B1(n_1082),
.B2(n_976),
.C(n_1087),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_967),
.Y(n_1224)
);

AOI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1082),
.A2(n_950),
.B1(n_850),
.B2(n_1085),
.Y(n_1225)
);

O2A1O1Ixp33_ASAP7_75t_L g1226 ( 
.A1(n_950),
.A2(n_850),
.B(n_1082),
.C(n_1085),
.Y(n_1226)
);

AO31x2_ASAP7_75t_L g1227 ( 
.A1(n_999),
.A2(n_854),
.A3(n_1025),
.B(n_1054),
.Y(n_1227)
);

NOR4xp25_ASAP7_75t_L g1228 ( 
.A(n_982),
.B(n_850),
.C(n_874),
.D(n_994),
.Y(n_1228)
);

BUFx6f_ASAP7_75t_L g1229 ( 
.A(n_1081),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_978),
.A2(n_829),
.B(n_1054),
.Y(n_1230)
);

OAI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1082),
.A2(n_850),
.B(n_999),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1085),
.B(n_1088),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_978),
.A2(n_829),
.B(n_1054),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_SL g1234 ( 
.A1(n_1109),
.A2(n_1123),
.B1(n_1188),
.B2(n_1097),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_SL g1235 ( 
.A1(n_1097),
.A2(n_1131),
.B1(n_1212),
.B2(n_1231),
.Y(n_1235)
);

BUFx8_ASAP7_75t_SL g1236 ( 
.A(n_1221),
.Y(n_1236)
);

INVx1_ASAP7_75t_SL g1237 ( 
.A(n_1108),
.Y(n_1237)
);

CKINVDCx11_ASAP7_75t_R g1238 ( 
.A(n_1125),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_SL g1239 ( 
.A1(n_1174),
.A2(n_1212),
.B1(n_1231),
.B2(n_1098),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_SL g1240 ( 
.A1(n_1174),
.A2(n_1232),
.B1(n_1143),
.B2(n_1152),
.Y(n_1240)
);

BUFx2_ASAP7_75t_L g1241 ( 
.A(n_1171),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1111),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1172),
.A2(n_1168),
.B1(n_1201),
.B2(n_1220),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1095),
.A2(n_1184),
.B1(n_1222),
.B2(n_1211),
.Y(n_1244)
);

INVx6_ASAP7_75t_L g1245 ( 
.A(n_1100),
.Y(n_1245)
);

CKINVDCx20_ASAP7_75t_R g1246 ( 
.A(n_1113),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_L g1247 ( 
.A1(n_1168),
.A2(n_1201),
.B1(n_1220),
.B2(n_1225),
.Y(n_1247)
);

BUFx3_ASAP7_75t_L g1248 ( 
.A(n_1197),
.Y(n_1248)
);

INVx1_ASAP7_75t_SL g1249 ( 
.A(n_1175),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1184),
.A2(n_1209),
.B1(n_1211),
.B2(n_1204),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1121),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_1124),
.Y(n_1252)
);

OAI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1204),
.A2(n_1222),
.B1(n_1225),
.B2(n_1209),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1130),
.Y(n_1254)
);

OAI22xp5_ASAP7_75t_L g1255 ( 
.A1(n_1149),
.A2(n_1118),
.B1(n_1187),
.B2(n_1215),
.Y(n_1255)
);

INVx3_ASAP7_75t_L g1256 ( 
.A(n_1206),
.Y(n_1256)
);

CKINVDCx11_ASAP7_75t_R g1257 ( 
.A(n_1140),
.Y(n_1257)
);

BUFx12f_ASAP7_75t_L g1258 ( 
.A(n_1197),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_SL g1259 ( 
.A1(n_1158),
.A2(n_1127),
.B1(n_1133),
.B2(n_1139),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1170),
.A2(n_1142),
.B1(n_1096),
.B2(n_1173),
.Y(n_1260)
);

BUFx3_ASAP7_75t_L g1261 ( 
.A(n_1195),
.Y(n_1261)
);

BUFx4f_ASAP7_75t_L g1262 ( 
.A(n_1189),
.Y(n_1262)
);

AOI22xp33_ASAP7_75t_L g1263 ( 
.A1(n_1133),
.A2(n_1101),
.B1(n_1136),
.B2(n_1104),
.Y(n_1263)
);

CKINVDCx20_ASAP7_75t_R g1264 ( 
.A(n_1166),
.Y(n_1264)
);

OAI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1183),
.A2(n_1210),
.B1(n_1223),
.B2(n_1182),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1181),
.B(n_1198),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1151),
.Y(n_1267)
);

BUFx2_ASAP7_75t_R g1268 ( 
.A(n_1148),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1101),
.A2(n_1136),
.B1(n_1216),
.B2(n_1177),
.Y(n_1269)
);

INVx1_ASAP7_75t_SL g1270 ( 
.A(n_1157),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_L g1271 ( 
.A1(n_1138),
.A2(n_1112),
.B1(n_1185),
.B2(n_1186),
.Y(n_1271)
);

INVx3_ASAP7_75t_L g1272 ( 
.A(n_1206),
.Y(n_1272)
);

CKINVDCx11_ASAP7_75t_R g1273 ( 
.A(n_1229),
.Y(n_1273)
);

BUFx4_ASAP7_75t_SL g1274 ( 
.A(n_1120),
.Y(n_1274)
);

CKINVDCx11_ASAP7_75t_R g1275 ( 
.A(n_1229),
.Y(n_1275)
);

BUFx6f_ASAP7_75t_L g1276 ( 
.A(n_1229),
.Y(n_1276)
);

BUFx4f_ASAP7_75t_SL g1277 ( 
.A(n_1147),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1164),
.A2(n_1122),
.B1(n_1141),
.B2(n_1191),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1164),
.A2(n_1161),
.B1(n_1228),
.B2(n_1224),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1228),
.A2(n_1119),
.B1(n_1159),
.B2(n_1190),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1103),
.A2(n_1226),
.B1(n_1119),
.B2(n_1190),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1153),
.Y(n_1282)
);

INVx8_ASAP7_75t_L g1283 ( 
.A(n_1150),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1106),
.A2(n_1128),
.B1(n_1156),
.B2(n_1099),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1106),
.A2(n_1128),
.B1(n_1094),
.B2(n_1233),
.Y(n_1285)
);

BUFx3_ASAP7_75t_L g1286 ( 
.A(n_1165),
.Y(n_1286)
);

OAI22xp33_ASAP7_75t_R g1287 ( 
.A1(n_1160),
.A2(n_1200),
.B1(n_1208),
.B2(n_1165),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1155),
.Y(n_1288)
);

OAI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1146),
.A2(n_1214),
.B1(n_1150),
.B2(n_1154),
.Y(n_1289)
);

OAI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1214),
.A2(n_1154),
.B1(n_1116),
.B2(n_1230),
.Y(n_1290)
);

INVxp67_ASAP7_75t_SL g1291 ( 
.A(n_1134),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1126),
.Y(n_1292)
);

CKINVDCx20_ASAP7_75t_R g1293 ( 
.A(n_1126),
.Y(n_1293)
);

CKINVDCx11_ASAP7_75t_R g1294 ( 
.A(n_1129),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_SL g1295 ( 
.A1(n_1163),
.A2(n_1219),
.B1(n_1169),
.B2(n_1207),
.Y(n_1295)
);

CKINVDCx6p67_ASAP7_75t_R g1296 ( 
.A(n_1196),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_L g1297 ( 
.A1(n_1176),
.A2(n_1179),
.B1(n_1180),
.B2(n_1202),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1137),
.A2(n_1199),
.B1(n_1194),
.B2(n_1193),
.Y(n_1298)
);

OAI22xp33_ASAP7_75t_L g1299 ( 
.A1(n_1200),
.A2(n_1208),
.B1(n_1196),
.B2(n_1110),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1135),
.B(n_1105),
.Y(n_1300)
);

OAI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1213),
.A2(n_1132),
.B1(n_1218),
.B2(n_1227),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1144),
.Y(n_1302)
);

BUFx8_ASAP7_75t_L g1303 ( 
.A(n_1162),
.Y(n_1303)
);

BUFx8_ASAP7_75t_SL g1304 ( 
.A(n_1162),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1135),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_SL g1306 ( 
.A1(n_1093),
.A2(n_1102),
.B1(n_1217),
.B2(n_1205),
.Y(n_1306)
);

BUFx6f_ASAP7_75t_L g1307 ( 
.A(n_1117),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1105),
.B(n_1132),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_SL g1309 ( 
.A1(n_1178),
.A2(n_1192),
.B1(n_1115),
.B2(n_1107),
.Y(n_1309)
);

OAI21xp5_ASAP7_75t_SL g1310 ( 
.A1(n_1167),
.A2(n_1203),
.B(n_1218),
.Y(n_1310)
);

INVx1_ASAP7_75t_SL g1311 ( 
.A(n_1105),
.Y(n_1311)
);

INVx6_ASAP7_75t_L g1312 ( 
.A(n_1114),
.Y(n_1312)
);

INVx2_ASAP7_75t_L g1313 ( 
.A(n_1114),
.Y(n_1313)
);

OAI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1167),
.A2(n_1203),
.B1(n_1218),
.B2(n_1227),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1167),
.A2(n_1203),
.B1(n_1227),
.B2(n_1114),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_SL g1316 ( 
.A1(n_1109),
.A2(n_404),
.B1(n_506),
.B2(n_641),
.Y(n_1316)
);

BUFx2_ASAP7_75t_SL g1317 ( 
.A(n_1100),
.Y(n_1317)
);

AOI22xp5_ASAP7_75t_SL g1318 ( 
.A1(n_1109),
.A2(n_859),
.B1(n_1123),
.B2(n_1131),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1174),
.A2(n_1082),
.B1(n_850),
.B2(n_988),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_1125),
.Y(n_1320)
);

OAI22xp5_ASAP7_75t_L g1321 ( 
.A1(n_1123),
.A2(n_1085),
.B1(n_1090),
.B2(n_1088),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1098),
.B(n_1232),
.Y(n_1322)
);

INVx5_ASAP7_75t_L g1323 ( 
.A(n_1100),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1145),
.Y(n_1324)
);

OAI22xp5_ASAP7_75t_L g1325 ( 
.A1(n_1123),
.A2(n_1085),
.B1(n_1090),
.B2(n_1088),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1145),
.Y(n_1326)
);

CKINVDCx11_ASAP7_75t_R g1327 ( 
.A(n_1125),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_1145),
.Y(n_1328)
);

OAI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1123),
.A2(n_1085),
.B1(n_1090),
.B2(n_1088),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1145),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_SL g1331 ( 
.A1(n_1109),
.A2(n_404),
.B1(n_506),
.B2(n_641),
.Y(n_1331)
);

INVx3_ASAP7_75t_L g1332 ( 
.A(n_1206),
.Y(n_1332)
);

BUFx2_ASAP7_75t_L g1333 ( 
.A(n_1171),
.Y(n_1333)
);

BUFx3_ASAP7_75t_L g1334 ( 
.A(n_1197),
.Y(n_1334)
);

BUFx10_ASAP7_75t_L g1335 ( 
.A(n_1113),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1145),
.Y(n_1336)
);

BUFx3_ASAP7_75t_L g1337 ( 
.A(n_1197),
.Y(n_1337)
);

INVx1_ASAP7_75t_SL g1338 ( 
.A(n_1108),
.Y(n_1338)
);

CKINVDCx14_ASAP7_75t_R g1339 ( 
.A(n_1125),
.Y(n_1339)
);

INVxp67_ASAP7_75t_L g1340 ( 
.A(n_1108),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1109),
.A2(n_850),
.B1(n_1082),
.B2(n_506),
.Y(n_1341)
);

OAI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1184),
.A2(n_950),
.B1(n_1088),
.B2(n_1085),
.Y(n_1342)
);

OAI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1184),
.A2(n_950),
.B1(n_1088),
.B2(n_1085),
.Y(n_1343)
);

AOI22xp33_ASAP7_75t_SL g1344 ( 
.A1(n_1109),
.A2(n_404),
.B1(n_506),
.B2(n_641),
.Y(n_1344)
);

CKINVDCx6p67_ASAP7_75t_R g1345 ( 
.A(n_1125),
.Y(n_1345)
);

AOI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1109),
.A2(n_438),
.B1(n_320),
.B2(n_324),
.Y(n_1346)
);

BUFx3_ASAP7_75t_L g1347 ( 
.A(n_1197),
.Y(n_1347)
);

CKINVDCx6p67_ASAP7_75t_R g1348 ( 
.A(n_1125),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1174),
.A2(n_1082),
.B1(n_850),
.B2(n_988),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_SL g1350 ( 
.A1(n_1109),
.A2(n_404),
.B1(n_506),
.B2(n_641),
.Y(n_1350)
);

CKINVDCx20_ASAP7_75t_R g1351 ( 
.A(n_1125),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1174),
.A2(n_1082),
.B1(n_850),
.B2(n_988),
.Y(n_1352)
);

OR2x2_ASAP7_75t_L g1353 ( 
.A(n_1310),
.B(n_1308),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1305),
.Y(n_1354)
);

OAI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1297),
.A2(n_1298),
.B(n_1302),
.Y(n_1355)
);

AND2x4_ASAP7_75t_L g1356 ( 
.A(n_1285),
.B(n_1286),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1235),
.B(n_1239),
.Y(n_1357)
);

OAI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1319),
.A2(n_1352),
.B(n_1349),
.Y(n_1358)
);

INVx1_ASAP7_75t_SL g1359 ( 
.A(n_1237),
.Y(n_1359)
);

HB1xp67_ASAP7_75t_L g1360 ( 
.A(n_1340),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1300),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1282),
.Y(n_1362)
);

INVx2_ASAP7_75t_SL g1363 ( 
.A(n_1245),
.Y(n_1363)
);

OAI222xp33_ASAP7_75t_L g1364 ( 
.A1(n_1316),
.A2(n_1350),
.B1(n_1344),
.B2(n_1331),
.C1(n_1341),
.C2(n_1234),
.Y(n_1364)
);

AOI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1288),
.A2(n_1266),
.B(n_1313),
.Y(n_1365)
);

BUFx3_ASAP7_75t_L g1366 ( 
.A(n_1303),
.Y(n_1366)
);

AOI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1247),
.A2(n_1281),
.B(n_1243),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1319),
.A2(n_1352),
.B1(n_1349),
.B2(n_1244),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1312),
.Y(n_1369)
);

OR2x2_ASAP7_75t_L g1370 ( 
.A(n_1315),
.B(n_1311),
.Y(n_1370)
);

BUFx3_ASAP7_75t_L g1371 ( 
.A(n_1303),
.Y(n_1371)
);

AND2x2_ASAP7_75t_L g1372 ( 
.A(n_1250),
.B(n_1259),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1322),
.B(n_1321),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1291),
.Y(n_1374)
);

BUFx2_ASAP7_75t_L g1375 ( 
.A(n_1304),
.Y(n_1375)
);

OAI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1244),
.A2(n_1325),
.B(n_1329),
.Y(n_1376)
);

HB1xp67_ASAP7_75t_L g1377 ( 
.A(n_1340),
.Y(n_1377)
);

AO21x1_ASAP7_75t_L g1378 ( 
.A1(n_1265),
.A2(n_1253),
.B(n_1343),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1314),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1314),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1250),
.A2(n_1253),
.B1(n_1240),
.B2(n_1265),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1242),
.Y(n_1382)
);

AOI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1251),
.A2(n_1254),
.B(n_1267),
.Y(n_1383)
);

OR2x2_ASAP7_75t_L g1384 ( 
.A(n_1315),
.B(n_1263),
.Y(n_1384)
);

BUFx6f_ASAP7_75t_L g1385 ( 
.A(n_1307),
.Y(n_1385)
);

OR2x2_ASAP7_75t_L g1386 ( 
.A(n_1263),
.B(n_1301),
.Y(n_1386)
);

BUFx3_ASAP7_75t_L g1387 ( 
.A(n_1283),
.Y(n_1387)
);

INVx1_ASAP7_75t_SL g1388 ( 
.A(n_1338),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1297),
.A2(n_1285),
.B(n_1284),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1307),
.Y(n_1390)
);

OR2x2_ASAP7_75t_L g1391 ( 
.A(n_1301),
.B(n_1269),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1307),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1287),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1299),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1299),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1284),
.A2(n_1260),
.B(n_1280),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1328),
.B(n_1279),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1295),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1306),
.Y(n_1399)
);

HB1xp67_ASAP7_75t_L g1400 ( 
.A(n_1324),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1309),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1326),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1330),
.Y(n_1403)
);

BUFx6f_ASAP7_75t_L g1404 ( 
.A(n_1323),
.Y(n_1404)
);

NAND2x1_ASAP7_75t_L g1405 ( 
.A(n_1245),
.B(n_1269),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1336),
.Y(n_1406)
);

AND2x4_ASAP7_75t_L g1407 ( 
.A(n_1280),
.B(n_1323),
.Y(n_1407)
);

OA21x2_ASAP7_75t_L g1408 ( 
.A1(n_1279),
.A2(n_1278),
.B(n_1271),
.Y(n_1408)
);

AO21x2_ASAP7_75t_L g1409 ( 
.A1(n_1290),
.A2(n_1343),
.B(n_1342),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1292),
.Y(n_1410)
);

HB1xp67_ASAP7_75t_L g1411 ( 
.A(n_1270),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1290),
.Y(n_1412)
);

BUFx3_ASAP7_75t_L g1413 ( 
.A(n_1283),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1342),
.Y(n_1414)
);

BUFx2_ASAP7_75t_L g1415 ( 
.A(n_1241),
.Y(n_1415)
);

HB1xp67_ASAP7_75t_L g1416 ( 
.A(n_1274),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1289),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1255),
.A2(n_1271),
.B1(n_1346),
.B2(n_1278),
.Y(n_1418)
);

INVx2_ASAP7_75t_SL g1419 ( 
.A(n_1283),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1317),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1318),
.B(n_1276),
.Y(n_1421)
);

INVx2_ASAP7_75t_SL g1422 ( 
.A(n_1274),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1333),
.Y(n_1423)
);

INVxp67_ASAP7_75t_L g1424 ( 
.A(n_1411),
.Y(n_1424)
);

OR2x2_ASAP7_75t_L g1425 ( 
.A(n_1353),
.B(n_1249),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1354),
.Y(n_1426)
);

AOI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1376),
.A2(n_1262),
.B(n_1332),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1361),
.B(n_1294),
.Y(n_1428)
);

AO32x2_ASAP7_75t_L g1429 ( 
.A1(n_1393),
.A2(n_1268),
.A3(n_1257),
.B1(n_1296),
.B2(n_1275),
.Y(n_1429)
);

OAI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1368),
.A2(n_1262),
.B1(n_1293),
.B2(n_1261),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1353),
.B(n_1348),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1358),
.A2(n_1332),
.B(n_1272),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1373),
.B(n_1339),
.Y(n_1433)
);

O2A1O1Ixp33_ASAP7_75t_SL g1434 ( 
.A1(n_1364),
.A2(n_1351),
.B(n_1246),
.C(n_1264),
.Y(n_1434)
);

BUFx3_ASAP7_75t_L g1435 ( 
.A(n_1366),
.Y(n_1435)
);

OAI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1381),
.A2(n_1272),
.B(n_1256),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1379),
.B(n_1345),
.Y(n_1437)
);

OA21x2_ASAP7_75t_L g1438 ( 
.A1(n_1355),
.A2(n_1365),
.B(n_1389),
.Y(n_1438)
);

OAI21xp33_ASAP7_75t_SL g1439 ( 
.A1(n_1357),
.A2(n_1273),
.B(n_1277),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1379),
.B(n_1347),
.Y(n_1440)
);

OAI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1418),
.A2(n_1320),
.B(n_1252),
.Y(n_1441)
);

NOR2x1_ASAP7_75t_SL g1442 ( 
.A(n_1409),
.B(n_1258),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1380),
.B(n_1337),
.Y(n_1443)
);

OR2x6_ASAP7_75t_L g1444 ( 
.A(n_1389),
.B(n_1248),
.Y(n_1444)
);

AND2x4_ASAP7_75t_L g1445 ( 
.A(n_1369),
.B(n_1334),
.Y(n_1445)
);

OAI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1357),
.A2(n_1277),
.B1(n_1335),
.B2(n_1327),
.Y(n_1446)
);

AO21x2_ASAP7_75t_L g1447 ( 
.A1(n_1365),
.A2(n_1335),
.B(n_1238),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1362),
.Y(n_1448)
);

NAND2xp5_ASAP7_75t_L g1449 ( 
.A(n_1360),
.B(n_1236),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1382),
.B(n_1406),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1370),
.B(n_1391),
.Y(n_1451)
);

O2A1O1Ixp33_ASAP7_75t_SL g1452 ( 
.A1(n_1422),
.A2(n_1416),
.B(n_1405),
.C(n_1393),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_L g1453 ( 
.A(n_1377),
.Y(n_1453)
);

OAI21xp5_ASAP7_75t_L g1454 ( 
.A1(n_1367),
.A2(n_1396),
.B(n_1372),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1397),
.B(n_1409),
.Y(n_1455)
);

OAI211xp5_ASAP7_75t_L g1456 ( 
.A1(n_1367),
.A2(n_1372),
.B(n_1408),
.C(n_1414),
.Y(n_1456)
);

NOR2x1_ASAP7_75t_SL g1457 ( 
.A(n_1409),
.B(n_1412),
.Y(n_1457)
);

OA21x2_ASAP7_75t_L g1458 ( 
.A1(n_1355),
.A2(n_1395),
.B(n_1394),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1397),
.B(n_1409),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1401),
.B(n_1362),
.Y(n_1460)
);

CKINVDCx10_ASAP7_75t_R g1461 ( 
.A(n_1422),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1401),
.B(n_1399),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1359),
.B(n_1388),
.Y(n_1463)
);

OA21x2_ASAP7_75t_L g1464 ( 
.A1(n_1394),
.A2(n_1395),
.B(n_1396),
.Y(n_1464)
);

OR2x6_ASAP7_75t_L g1465 ( 
.A(n_1356),
.B(n_1405),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1356),
.B(n_1410),
.Y(n_1466)
);

NOR2xp33_ASAP7_75t_L g1467 ( 
.A(n_1388),
.B(n_1423),
.Y(n_1467)
);

BUFx12f_ASAP7_75t_L g1468 ( 
.A(n_1415),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1356),
.B(n_1410),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1383),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1402),
.B(n_1403),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1402),
.B(n_1403),
.Y(n_1472)
);

OR2x6_ASAP7_75t_L g1473 ( 
.A(n_1407),
.B(n_1378),
.Y(n_1473)
);

OAI21xp5_ASAP7_75t_L g1474 ( 
.A1(n_1398),
.A2(n_1408),
.B(n_1417),
.Y(n_1474)
);

CKINVDCx20_ASAP7_75t_R g1475 ( 
.A(n_1415),
.Y(n_1475)
);

INVx3_ASAP7_75t_L g1476 ( 
.A(n_1385),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1458),
.B(n_1374),
.Y(n_1477)
);

BUFx12f_ASAP7_75t_L g1478 ( 
.A(n_1468),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1426),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1455),
.B(n_1400),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_SL g1481 ( 
.A1(n_1473),
.A2(n_1408),
.B1(n_1375),
.B2(n_1386),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1455),
.B(n_1412),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1448),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1448),
.Y(n_1484)
);

HB1xp67_ASAP7_75t_L g1485 ( 
.A(n_1470),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1466),
.B(n_1469),
.Y(n_1486)
);

OR2x2_ASAP7_75t_L g1487 ( 
.A(n_1458),
.B(n_1386),
.Y(n_1487)
);

CKINVDCx20_ASAP7_75t_R g1488 ( 
.A(n_1475),
.Y(n_1488)
);

NAND2xp5_ASAP7_75t_L g1489 ( 
.A(n_1459),
.B(n_1378),
.Y(n_1489)
);

INVx1_ASAP7_75t_SL g1490 ( 
.A(n_1425),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1470),
.Y(n_1491)
);

HB1xp67_ASAP7_75t_L g1492 ( 
.A(n_1470),
.Y(n_1492)
);

INVx3_ASAP7_75t_L g1493 ( 
.A(n_1476),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1459),
.B(n_1390),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1450),
.Y(n_1495)
);

INVxp67_ASAP7_75t_L g1496 ( 
.A(n_1450),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1430),
.A2(n_1408),
.B1(n_1384),
.B2(n_1407),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1460),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1471),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1471),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1438),
.B(n_1392),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1472),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1485),
.Y(n_1503)
);

OAI221xp5_ASAP7_75t_L g1504 ( 
.A1(n_1481),
.A2(n_1434),
.B1(n_1441),
.B2(n_1454),
.C(n_1439),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1483),
.Y(n_1505)
);

OAI211xp5_ASAP7_75t_L g1506 ( 
.A1(n_1481),
.A2(n_1439),
.B(n_1456),
.C(n_1474),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1489),
.B(n_1464),
.Y(n_1507)
);

OR2x2_ASAP7_75t_L g1508 ( 
.A(n_1487),
.B(n_1464),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1486),
.B(n_1457),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1487),
.B(n_1464),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1497),
.A2(n_1473),
.B1(n_1384),
.B2(n_1425),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1486),
.B(n_1457),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1486),
.B(n_1473),
.Y(n_1513)
);

INVx1_ASAP7_75t_SL g1514 ( 
.A(n_1490),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_1480),
.B(n_1433),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1494),
.B(n_1473),
.Y(n_1516)
);

BUFx3_ASAP7_75t_L g1517 ( 
.A(n_1493),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1494),
.B(n_1473),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1487),
.B(n_1464),
.Y(n_1519)
);

INVx3_ASAP7_75t_L g1520 ( 
.A(n_1491),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1483),
.Y(n_1521)
);

AO21x2_ASAP7_75t_L g1522 ( 
.A1(n_1489),
.A2(n_1442),
.B(n_1447),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1480),
.B(n_1451),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1483),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1494),
.B(n_1444),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1482),
.B(n_1453),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1482),
.B(n_1490),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1484),
.Y(n_1528)
);

NAND3xp33_ASAP7_75t_L g1529 ( 
.A(n_1497),
.B(n_1463),
.C(n_1467),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_1492),
.Y(n_1530)
);

INVxp67_ASAP7_75t_SL g1531 ( 
.A(n_1492),
.Y(n_1531)
);

INVxp67_ASAP7_75t_L g1532 ( 
.A(n_1479),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1498),
.B(n_1444),
.Y(n_1533)
);

AOI22xp33_ASAP7_75t_L g1534 ( 
.A1(n_1478),
.A2(n_1462),
.B1(n_1437),
.B2(n_1465),
.Y(n_1534)
);

INVx4_ASAP7_75t_L g1535 ( 
.A(n_1478),
.Y(n_1535)
);

OAI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1478),
.A2(n_1465),
.B1(n_1375),
.B2(n_1431),
.Y(n_1536)
);

INVx3_ASAP7_75t_L g1537 ( 
.A(n_1517),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1532),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1507),
.B(n_1508),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_1530),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1532),
.Y(n_1541)
);

HB1xp67_ASAP7_75t_L g1542 ( 
.A(n_1530),
.Y(n_1542)
);

BUFx2_ASAP7_75t_L g1543 ( 
.A(n_1535),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_L g1544 ( 
.A(n_1507),
.B(n_1523),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1505),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1509),
.B(n_1498),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1509),
.B(n_1498),
.Y(n_1547)
);

HB1xp67_ASAP7_75t_L g1548 ( 
.A(n_1503),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1505),
.Y(n_1549)
);

INVxp67_ASAP7_75t_L g1550 ( 
.A(n_1514),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1509),
.B(n_1495),
.Y(n_1551)
);

NAND2x1p5_ASAP7_75t_L g1552 ( 
.A(n_1514),
.B(n_1438),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1512),
.B(n_1495),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1520),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1508),
.B(n_1477),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1521),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1512),
.B(n_1495),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1512),
.B(n_1496),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1521),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1523),
.B(n_1499),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1524),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1513),
.B(n_1533),
.Y(n_1562)
);

AND2x4_ASAP7_75t_L g1563 ( 
.A(n_1533),
.B(n_1501),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1513),
.B(n_1496),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1513),
.B(n_1533),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1523),
.B(n_1499),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1520),
.Y(n_1567)
);

BUFx2_ASAP7_75t_L g1568 ( 
.A(n_1535),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1527),
.B(n_1500),
.Y(n_1569)
);

OR2x2_ASAP7_75t_L g1570 ( 
.A(n_1527),
.B(n_1500),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1524),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1528),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1526),
.B(n_1502),
.Y(n_1573)
);

INVx2_ASAP7_75t_L g1574 ( 
.A(n_1552),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1538),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1544),
.B(n_1508),
.Y(n_1576)
);

NOR2x1_ASAP7_75t_L g1577 ( 
.A(n_1543),
.B(n_1568),
.Y(n_1577)
);

INVx1_ASAP7_75t_SL g1578 ( 
.A(n_1543),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1562),
.B(n_1525),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1548),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1550),
.B(n_1515),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1550),
.B(n_1515),
.Y(n_1582)
);

INVx2_ASAP7_75t_L g1583 ( 
.A(n_1552),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1562),
.B(n_1525),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1562),
.B(n_1525),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1544),
.B(n_1510),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1566),
.B(n_1510),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1548),
.Y(n_1588)
);

AOI32xp33_ASAP7_75t_L g1589 ( 
.A1(n_1568),
.A2(n_1504),
.A3(n_1536),
.B1(n_1511),
.B2(n_1518),
.Y(n_1589)
);

AOI21xp5_ASAP7_75t_L g1590 ( 
.A1(n_1573),
.A2(n_1504),
.B(n_1506),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1545),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1545),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1549),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1565),
.B(n_1516),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1549),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1538),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1565),
.B(n_1516),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1541),
.Y(n_1598)
);

AND2x4_ASAP7_75t_L g1599 ( 
.A(n_1565),
.B(n_1535),
.Y(n_1599)
);

HB1xp67_ASAP7_75t_L g1600 ( 
.A(n_1540),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1556),
.Y(n_1601)
);

OR2x6_ASAP7_75t_L g1602 ( 
.A(n_1537),
.B(n_1535),
.Y(n_1602)
);

AND2x2_ASAP7_75t_SL g1603 ( 
.A(n_1540),
.B(n_1535),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1564),
.B(n_1516),
.Y(n_1604)
);

AOI33xp33_ASAP7_75t_L g1605 ( 
.A1(n_1541),
.A2(n_1511),
.A3(n_1536),
.B1(n_1534),
.B2(n_1437),
.B3(n_1440),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1556),
.Y(n_1606)
);

INVxp67_ASAP7_75t_SL g1607 ( 
.A(n_1542),
.Y(n_1607)
);

OAI221xp5_ASAP7_75t_SL g1608 ( 
.A1(n_1539),
.A2(n_1506),
.B1(n_1529),
.B2(n_1534),
.C(n_1519),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1559),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1564),
.B(n_1518),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1559),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1561),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1561),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1552),
.Y(n_1614)
);

OR2x6_ASAP7_75t_L g1615 ( 
.A(n_1537),
.B(n_1478),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1600),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1590),
.B(n_1564),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1591),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1591),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1579),
.B(n_1558),
.Y(n_1620)
);

AND2x4_ASAP7_75t_L g1621 ( 
.A(n_1577),
.B(n_1599),
.Y(n_1621)
);

NOR2xp33_ASAP7_75t_SL g1622 ( 
.A(n_1608),
.B(n_1603),
.Y(n_1622)
);

INVx3_ASAP7_75t_L g1623 ( 
.A(n_1599),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1581),
.B(n_1566),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1582),
.B(n_1573),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1592),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1592),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1594),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1578),
.B(n_1529),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1579),
.B(n_1584),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1593),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1605),
.B(n_1518),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1593),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1595),
.Y(n_1634)
);

AND2x4_ASAP7_75t_L g1635 ( 
.A(n_1599),
.B(n_1537),
.Y(n_1635)
);

AND3x2_ASAP7_75t_L g1636 ( 
.A(n_1607),
.B(n_1542),
.C(n_1428),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1595),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1584),
.B(n_1558),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1575),
.B(n_1539),
.Y(n_1639)
);

OR2x2_ASAP7_75t_L g1640 ( 
.A(n_1596),
.B(n_1539),
.Y(n_1640)
);

OR2x2_ASAP7_75t_L g1641 ( 
.A(n_1598),
.B(n_1560),
.Y(n_1641)
);

BUFx2_ASAP7_75t_L g1642 ( 
.A(n_1603),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1589),
.B(n_1569),
.Y(n_1643)
);

NOR2xp33_ASAP7_75t_L g1644 ( 
.A(n_1615),
.B(n_1488),
.Y(n_1644)
);

OAI21xp5_ASAP7_75t_L g1645 ( 
.A1(n_1615),
.A2(n_1446),
.B(n_1552),
.Y(n_1645)
);

OR2x2_ASAP7_75t_L g1646 ( 
.A(n_1585),
.B(n_1560),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1604),
.B(n_1569),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1585),
.B(n_1526),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1576),
.B(n_1570),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1601),
.Y(n_1650)
);

OAI22xp5_ASAP7_75t_L g1651 ( 
.A1(n_1643),
.A2(n_1615),
.B1(n_1602),
.B2(n_1488),
.Y(n_1651)
);

OAI221xp5_ASAP7_75t_SL g1652 ( 
.A1(n_1617),
.A2(n_1615),
.B1(n_1602),
.B2(n_1576),
.C(n_1586),
.Y(n_1652)
);

OAI221xp5_ASAP7_75t_L g1653 ( 
.A1(n_1622),
.A2(n_1602),
.B1(n_1431),
.B2(n_1588),
.C(n_1580),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1644),
.B(n_1604),
.Y(n_1654)
);

AOI21xp33_ASAP7_75t_L g1655 ( 
.A1(n_1642),
.A2(n_1602),
.B(n_1588),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1618),
.Y(n_1656)
);

AOI21xp5_ASAP7_75t_L g1657 ( 
.A1(n_1629),
.A2(n_1449),
.B(n_1580),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1624),
.B(n_1610),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1616),
.B(n_1610),
.Y(n_1659)
);

AOI322xp5_ASAP7_75t_L g1660 ( 
.A1(n_1632),
.A2(n_1597),
.A3(n_1594),
.B1(n_1558),
.B2(n_1563),
.C1(n_1557),
.C2(n_1551),
.Y(n_1660)
);

AOI221xp5_ASAP7_75t_L g1661 ( 
.A1(n_1625),
.A2(n_1614),
.B1(n_1574),
.B2(n_1583),
.C(n_1606),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1644),
.B(n_1597),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1630),
.B(n_1537),
.Y(n_1663)
);

OAI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1621),
.A2(n_1444),
.B1(n_1435),
.B2(n_1465),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1621),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1619),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1626),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1636),
.B(n_1551),
.Y(n_1668)
);

OAI22xp33_ASAP7_75t_L g1669 ( 
.A1(n_1645),
.A2(n_1444),
.B1(n_1465),
.B2(n_1371),
.Y(n_1669)
);

AOI322xp5_ASAP7_75t_L g1670 ( 
.A1(n_1630),
.A2(n_1563),
.A3(n_1553),
.B1(n_1551),
.B2(n_1557),
.C1(n_1547),
.C2(n_1546),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1627),
.Y(n_1671)
);

OAI22xp33_ASAP7_75t_L g1672 ( 
.A1(n_1628),
.A2(n_1465),
.B1(n_1371),
.B2(n_1366),
.Y(n_1672)
);

NOR3xp33_ASAP7_75t_L g1673 ( 
.A(n_1623),
.B(n_1583),
.C(n_1574),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1636),
.B(n_1553),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_SL g1675 ( 
.A(n_1621),
.B(n_1614),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1656),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1665),
.B(n_1628),
.Y(n_1677)
);

OAI221xp5_ASAP7_75t_L g1678 ( 
.A1(n_1652),
.A2(n_1623),
.B1(n_1647),
.B2(n_1639),
.C(n_1640),
.Y(n_1678)
);

OAI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1653),
.A2(n_1623),
.B1(n_1646),
.B2(n_1648),
.Y(n_1679)
);

HB1xp67_ASAP7_75t_L g1680 ( 
.A(n_1665),
.Y(n_1680)
);

OAI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1668),
.A2(n_1638),
.B1(n_1620),
.B2(n_1635),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1666),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1654),
.B(n_1620),
.Y(n_1683)
);

AOI22xp33_ASAP7_75t_L g1684 ( 
.A1(n_1651),
.A2(n_1650),
.B1(n_1631),
.B2(n_1633),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1657),
.B(n_1638),
.Y(n_1685)
);

NOR3xp33_ASAP7_75t_L g1686 ( 
.A(n_1655),
.B(n_1659),
.C(n_1662),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1667),
.Y(n_1687)
);

AOI21xp5_ASAP7_75t_L g1688 ( 
.A1(n_1675),
.A2(n_1635),
.B(n_1639),
.Y(n_1688)
);

INVxp67_ASAP7_75t_L g1689 ( 
.A(n_1675),
.Y(n_1689)
);

AOI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1669),
.A2(n_1635),
.B1(n_1522),
.B2(n_1637),
.Y(n_1690)
);

OAI211xp5_ASAP7_75t_L g1691 ( 
.A1(n_1660),
.A2(n_1634),
.B(n_1640),
.C(n_1649),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1671),
.B(n_1658),
.Y(n_1692)
);

NOR4xp25_ASAP7_75t_L g1693 ( 
.A(n_1661),
.B(n_1674),
.C(n_1669),
.D(n_1672),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1663),
.Y(n_1694)
);

AOI221xp5_ASAP7_75t_L g1695 ( 
.A1(n_1693),
.A2(n_1673),
.B1(n_1672),
.B2(n_1663),
.C(n_1664),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1694),
.B(n_1670),
.Y(n_1696)
);

INVx1_ASAP7_75t_SL g1697 ( 
.A(n_1688),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1680),
.Y(n_1698)
);

OAI21xp33_ASAP7_75t_L g1699 ( 
.A1(n_1684),
.A2(n_1641),
.B(n_1586),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1689),
.B(n_1641),
.Y(n_1700)
);

AOI211xp5_ASAP7_75t_SL g1701 ( 
.A1(n_1680),
.A2(n_1452),
.B(n_1429),
.C(n_1427),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1686),
.B(n_1601),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1683),
.B(n_1587),
.Y(n_1703)
);

NOR2xp33_ASAP7_75t_L g1704 ( 
.A(n_1692),
.B(n_1685),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1677),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_SL g1706 ( 
.A(n_1678),
.B(n_1468),
.Y(n_1706)
);

NOR3xp33_ASAP7_75t_L g1707 ( 
.A(n_1697),
.B(n_1682),
.C(n_1676),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1704),
.B(n_1684),
.Y(n_1708)
);

AOI22xp33_ASAP7_75t_SL g1709 ( 
.A1(n_1706),
.A2(n_1679),
.B1(n_1691),
.B2(n_1681),
.Y(n_1709)
);

A2O1A1Ixp33_ASAP7_75t_L g1710 ( 
.A1(n_1701),
.A2(n_1690),
.B(n_1687),
.C(n_1613),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_SL g1711 ( 
.A(n_1695),
.B(n_1609),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1696),
.B(n_1609),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1698),
.Y(n_1713)
);

NAND3xp33_ASAP7_75t_SL g1714 ( 
.A(n_1701),
.B(n_1428),
.C(n_1587),
.Y(n_1714)
);

O2A1O1Ixp33_ASAP7_75t_L g1715 ( 
.A1(n_1702),
.A2(n_1424),
.B(n_1613),
.C(n_1612),
.Y(n_1715)
);

OR2x2_ASAP7_75t_L g1716 ( 
.A(n_1712),
.B(n_1700),
.Y(n_1716)
);

OAI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1709),
.A2(n_1703),
.B1(n_1699),
.B2(n_1705),
.Y(n_1717)
);

OAI211xp5_ASAP7_75t_SL g1718 ( 
.A1(n_1708),
.A2(n_1612),
.B(n_1611),
.C(n_1429),
.Y(n_1718)
);

OAI22xp5_ASAP7_75t_L g1719 ( 
.A1(n_1711),
.A2(n_1611),
.B1(n_1563),
.B2(n_1555),
.Y(n_1719)
);

O2A1O1Ixp5_ASAP7_75t_L g1720 ( 
.A1(n_1710),
.A2(n_1555),
.B(n_1563),
.C(n_1420),
.Y(n_1720)
);

OAI21xp5_ASAP7_75t_L g1721 ( 
.A1(n_1717),
.A2(n_1707),
.B(n_1714),
.Y(n_1721)
);

NAND2xp33_ASAP7_75t_L g1722 ( 
.A(n_1716),
.B(n_1713),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1719),
.B(n_1715),
.Y(n_1723)
);

AOI322xp5_ASAP7_75t_L g1724 ( 
.A1(n_1718),
.A2(n_1563),
.A3(n_1531),
.B1(n_1553),
.B2(n_1557),
.C1(n_1440),
.C2(n_1443),
.Y(n_1724)
);

AOI221xp5_ASAP7_75t_SL g1725 ( 
.A1(n_1720),
.A2(n_1443),
.B1(n_1555),
.B2(n_1420),
.C(n_1429),
.Y(n_1725)
);

NOR2xp33_ASAP7_75t_L g1726 ( 
.A(n_1716),
.B(n_1461),
.Y(n_1726)
);

BUFx2_ASAP7_75t_L g1727 ( 
.A(n_1721),
.Y(n_1727)
);

AOI22xp33_ASAP7_75t_L g1728 ( 
.A1(n_1723),
.A2(n_1522),
.B1(n_1447),
.B2(n_1445),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1722),
.Y(n_1729)
);

NOR2xp67_ASAP7_75t_L g1730 ( 
.A(n_1726),
.B(n_1554),
.Y(n_1730)
);

OAI211xp5_ASAP7_75t_L g1731 ( 
.A1(n_1724),
.A2(n_1429),
.B(n_1461),
.C(n_1366),
.Y(n_1731)
);

OAI221xp5_ASAP7_75t_SL g1732 ( 
.A1(n_1731),
.A2(n_1725),
.B1(n_1429),
.B2(n_1435),
.C(n_1371),
.Y(n_1732)
);

AOI22xp5_ASAP7_75t_SL g1733 ( 
.A1(n_1729),
.A2(n_1429),
.B1(n_1435),
.B2(n_1413),
.Y(n_1733)
);

AND4x1_ASAP7_75t_L g1734 ( 
.A(n_1727),
.B(n_1421),
.C(n_1432),
.D(n_1436),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1733),
.Y(n_1735)
);

AOI211xp5_ASAP7_75t_L g1736 ( 
.A1(n_1735),
.A2(n_1732),
.B(n_1730),
.C(n_1734),
.Y(n_1736)
);

OAI22xp5_ASAP7_75t_L g1737 ( 
.A1(n_1736),
.A2(n_1728),
.B1(n_1567),
.B2(n_1554),
.Y(n_1737)
);

AOI22xp33_ASAP7_75t_L g1738 ( 
.A1(n_1737),
.A2(n_1728),
.B1(n_1522),
.B2(n_1445),
.Y(n_1738)
);

AOI22xp5_ASAP7_75t_L g1739 ( 
.A1(n_1738),
.A2(n_1522),
.B1(n_1554),
.B2(n_1567),
.Y(n_1739)
);

AOI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1739),
.A2(n_1419),
.B(n_1447),
.Y(n_1740)
);

XOR2xp5_ASAP7_75t_L g1741 ( 
.A(n_1739),
.B(n_1445),
.Y(n_1741)
);

AO21x2_ASAP7_75t_L g1742 ( 
.A1(n_1740),
.A2(n_1567),
.B(n_1572),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1741),
.B(n_1445),
.Y(n_1743)
);

AOI22x1_ASAP7_75t_L g1744 ( 
.A1(n_1742),
.A2(n_1419),
.B1(n_1363),
.B2(n_1404),
.Y(n_1744)
);

OAI22xp33_ASAP7_75t_L g1745 ( 
.A1(n_1743),
.A2(n_1570),
.B1(n_1571),
.B2(n_1572),
.Y(n_1745)
);

OAI221xp5_ASAP7_75t_R g1746 ( 
.A1(n_1744),
.A2(n_1522),
.B1(n_1531),
.B2(n_1442),
.C(n_1571),
.Y(n_1746)
);

AOI211xp5_ASAP7_75t_L g1747 ( 
.A1(n_1746),
.A2(n_1745),
.B(n_1387),
.C(n_1413),
.Y(n_1747)
);


endmodule