module real_aes_17482_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_831, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_831;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_815;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g112 ( .A(n_0), .B(n_113), .Y(n_112) );
AOI22xp5_ASAP7_75t_L g500 ( .A1(n_1), .A2(n_4), .B1(n_151), .B2(n_501), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g193 ( .A1(n_2), .A2(n_42), .B1(n_158), .B2(n_194), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_3), .A2(n_25), .B1(n_194), .B2(n_236), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g224 ( .A1(n_5), .A2(n_17), .B1(n_148), .B2(n_225), .Y(n_224) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_6), .A2(n_60), .B1(n_208), .B2(n_238), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g604 ( .A1(n_7), .A2(n_18), .B1(n_158), .B2(n_179), .Y(n_604) );
INVx1_ASAP7_75t_L g113 ( .A(n_8), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g517 ( .A(n_9), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_10), .A2(n_100), .B1(n_114), .B2(n_828), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g820 ( .A(n_11), .Y(n_820) );
CKINVDCx5p33_ASAP7_75t_R g178 ( .A(n_12), .Y(n_178) );
AOI22xp5_ASAP7_75t_L g206 ( .A1(n_13), .A2(n_19), .B1(n_207), .B2(n_210), .Y(n_206) );
OR2x2_ASAP7_75t_L g105 ( .A(n_14), .B(n_38), .Y(n_105) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_15), .Y(n_150) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_16), .Y(n_229) );
AOI22xp5_ASAP7_75t_L g147 ( .A1(n_20), .A2(n_97), .B1(n_148), .B2(n_151), .Y(n_147) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_21), .A2(n_39), .B1(n_183), .B2(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_22), .B(n_149), .Y(n_180) );
OAI21x1_ASAP7_75t_L g166 ( .A1(n_23), .A2(n_56), .B(n_167), .Y(n_166) );
CKINVDCx5p33_ASAP7_75t_R g496 ( .A(n_24), .Y(n_496) );
CKINVDCx5p33_ASAP7_75t_R g169 ( .A(n_26), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_27), .B(n_155), .Y(n_524) );
INVx4_ASAP7_75t_R g572 ( .A(n_28), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g195 ( .A1(n_29), .A2(n_46), .B1(n_196), .B2(n_197), .Y(n_195) );
AOI22xp33_ASAP7_75t_L g276 ( .A1(n_30), .A2(n_53), .B1(n_148), .B2(n_197), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g242 ( .A(n_31), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_32), .B(n_183), .Y(n_182) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_33), .Y(n_259) );
INVx1_ASAP7_75t_L g503 ( .A(n_34), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_35), .B(n_194), .Y(n_530) );
A2O1A1Ixp33_ASAP7_75t_SL g515 ( .A1(n_36), .A2(n_154), .B(n_158), .C(n_516), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g492 ( .A1(n_37), .A2(n_54), .B1(n_158), .B2(n_197), .Y(n_492) );
AOI22xp5_ASAP7_75t_L g234 ( .A1(n_40), .A2(n_85), .B1(n_158), .B2(n_235), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g211 ( .A1(n_41), .A2(n_45), .B1(n_158), .B2(n_179), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g512 ( .A(n_43), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g156 ( .A1(n_44), .A2(n_58), .B1(n_148), .B2(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g527 ( .A(n_47), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_48), .B(n_158), .Y(n_529) );
CKINVDCx5p33_ASAP7_75t_R g544 ( .A(n_49), .Y(n_544) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_50), .Y(n_116) );
INVx2_ASAP7_75t_L g128 ( .A(n_51), .Y(n_128) );
INVx1_ASAP7_75t_L g108 ( .A(n_52), .Y(n_108) );
BUFx3_ASAP7_75t_L g812 ( .A(n_52), .Y(n_812) );
CKINVDCx5p33_ASAP7_75t_R g573 ( .A(n_55), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_57), .A2(n_86), .B1(n_158), .B2(n_197), .Y(n_605) );
AOI22xp5_ASAP7_75t_L g130 ( .A1(n_59), .A2(n_131), .B1(n_471), .B2(n_472), .Y(n_130) );
INVx1_ASAP7_75t_L g471 ( .A(n_59), .Y(n_471) );
AOI22xp33_ASAP7_75t_L g275 ( .A1(n_61), .A2(n_74), .B1(n_157), .B2(n_196), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g607 ( .A(n_62), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g257 ( .A1(n_63), .A2(n_76), .B1(n_158), .B2(n_179), .Y(n_257) );
AOI22xp5_ASAP7_75t_L g256 ( .A1(n_64), .A2(n_96), .B1(n_148), .B2(n_210), .Y(n_256) );
AND2x4_ASAP7_75t_L g144 ( .A(n_65), .B(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g167 ( .A(n_66), .Y(n_167) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_67), .A2(n_88), .B1(n_196), .B2(n_197), .Y(n_499) );
AO22x1_ASAP7_75t_L g561 ( .A1(n_68), .A2(n_75), .B1(n_222), .B2(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g145 ( .A(n_69), .Y(n_145) );
OAI22xp5_ASAP7_75t_L g479 ( .A1(n_70), .A2(n_480), .B1(n_481), .B2(n_805), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_70), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g814 ( .A1(n_70), .A2(n_131), .B1(n_472), .B2(n_480), .Y(n_814) );
AND2x2_ASAP7_75t_L g519 ( .A(n_71), .B(n_189), .Y(n_519) );
CKINVDCx5p33_ASAP7_75t_R g510 ( .A(n_72), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_73), .B(n_238), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_77), .B(n_194), .Y(n_545) );
INVx2_ASAP7_75t_L g155 ( .A(n_78), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_79), .B(n_189), .Y(n_521) );
CKINVDCx5p33_ASAP7_75t_R g569 ( .A(n_80), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g237 ( .A1(n_81), .A2(n_95), .B1(n_197), .B2(n_238), .Y(n_237) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_82), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_83), .B(n_165), .Y(n_559) );
CKINVDCx5p33_ASAP7_75t_R g200 ( .A(n_84), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_87), .B(n_189), .Y(n_188) );
CKINVDCx5p33_ASAP7_75t_R g217 ( .A(n_89), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g541 ( .A(n_90), .B(n_189), .Y(n_541) );
INVx1_ASAP7_75t_L g111 ( .A(n_91), .Y(n_111) );
NOR2xp33_ASAP7_75t_L g120 ( .A(n_91), .B(n_121), .Y(n_120) );
NAND2xp33_ASAP7_75t_L g185 ( .A(n_92), .B(n_149), .Y(n_185) );
A2O1A1Ixp33_ASAP7_75t_L g567 ( .A1(n_93), .A2(n_213), .B(n_238), .C(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g574 ( .A(n_94), .B(n_575), .Y(n_574) );
NAND2xp33_ASAP7_75t_L g549 ( .A(n_98), .B(n_184), .Y(n_549) );
BUFx12f_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx6_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
INVx6_ASAP7_75t_L g829 ( .A(n_102), .Y(n_829) );
NAND2x2_ASAP7_75t_L g102 ( .A(n_103), .B(n_106), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
BUFx2_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g122 ( .A(n_105), .Y(n_122) );
NOR2x1_ASAP7_75t_L g827 ( .A(n_105), .B(n_812), .Y(n_827) );
NOR2x1p5_ASAP7_75t_L g106 ( .A(n_107), .B(n_109), .Y(n_106) );
AND3x2_ASAP7_75t_L g476 ( .A(n_107), .B(n_110), .C(n_122), .Y(n_476) );
HB1xp67_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g121 ( .A(n_108), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_110), .B(n_112), .Y(n_109) );
BUFx6f_ASAP7_75t_L g813 ( .A(n_110), .Y(n_813) );
BUFx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx2_ASAP7_75t_L g818 ( .A(n_111), .Y(n_818) );
OR2x6_ASAP7_75t_L g114 ( .A(n_115), .B(n_123), .Y(n_114) );
INVx1_ASAP7_75t_L g477 ( .A(n_115), .Y(n_477) );
NOR2xp67_ASAP7_75t_SL g115 ( .A(n_116), .B(n_117), .Y(n_115) );
BUFx12f_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx4_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
AND2x6_ASAP7_75t_SL g119 ( .A(n_120), .B(n_122), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_122), .B(n_811), .Y(n_810) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_124), .B(n_478), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_129), .Y(n_124) );
INVxp67_ASAP7_75t_SL g125 ( .A(n_126), .Y(n_125) );
BUFx8_ASAP7_75t_SL g126 ( .A(n_127), .Y(n_126) );
INVx3_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g809 ( .A(n_128), .Y(n_809) );
NOR2xp33_ASAP7_75t_L g824 ( .A(n_128), .B(n_825), .Y(n_824) );
OAI21xp5_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_474), .B(n_477), .Y(n_129) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx2_ASAP7_75t_L g473 ( .A(n_132), .Y(n_473) );
OR2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_374), .Y(n_132) );
NAND4xp25_ASAP7_75t_L g133 ( .A(n_134), .B(n_298), .C(n_329), .D(n_358), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g134 ( .A(n_135), .B(n_265), .Y(n_134) );
OAI322xp33_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_201), .A3(n_230), .B1(n_243), .B2(n_251), .C1(n_260), .C2(n_262), .Y(n_135) );
INVxp67_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_137), .B(n_455), .Y(n_454) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_171), .Y(n_137) );
AND2x2_ASAP7_75t_L g295 ( .A(n_138), .B(n_296), .Y(n_295) );
INVx4_ASAP7_75t_L g331 ( .A(n_138), .Y(n_331) );
INVx3_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x2_ASAP7_75t_L g306 ( .A(n_139), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g309 ( .A(n_139), .B(n_203), .Y(n_309) );
AND2x2_ASAP7_75t_L g326 ( .A(n_139), .B(n_219), .Y(n_326) );
AND2x2_ASAP7_75t_L g424 ( .A(n_139), .B(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx2_ASAP7_75t_L g247 ( .A(n_140), .Y(n_247) );
AND2x4_ASAP7_75t_L g430 ( .A(n_140), .B(n_425), .Y(n_430) );
AO31x2_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_146), .A3(n_162), .B(n_168), .Y(n_140) );
AO31x2_ASAP7_75t_L g254 ( .A1(n_141), .A2(n_214), .A3(n_255), .B(n_258), .Y(n_254) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AOI21xp5_ASAP7_75t_L g566 ( .A1(n_142), .A2(n_567), .B(n_570), .Y(n_566) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AO31x2_ASAP7_75t_L g191 ( .A1(n_143), .A2(n_192), .A3(n_198), .B(n_199), .Y(n_191) );
AO31x2_ASAP7_75t_L g204 ( .A1(n_143), .A2(n_205), .A3(n_214), .B(n_216), .Y(n_204) );
AO31x2_ASAP7_75t_L g219 ( .A1(n_143), .A2(n_220), .A3(n_227), .B(n_228), .Y(n_219) );
AO31x2_ASAP7_75t_L g602 ( .A1(n_143), .A2(n_170), .A3(n_603), .B(n_606), .Y(n_602) );
BUFx10_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g187 ( .A(n_144), .Y(n_187) );
BUFx10_ASAP7_75t_L g494 ( .A(n_144), .Y(n_494) );
INVx1_ASAP7_75t_L g518 ( .A(n_144), .Y(n_518) );
OAI22xp5_ASAP7_75t_L g146 ( .A1(n_147), .A2(n_153), .B1(n_156), .B2(n_159), .Y(n_146) );
INVx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVxp67_ASAP7_75t_SL g562 ( .A(n_149), .Y(n_562) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g152 ( .A(n_150), .Y(n_152) );
INVx3_ASAP7_75t_L g158 ( .A(n_150), .Y(n_158) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_150), .Y(n_184) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_150), .Y(n_194) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_150), .Y(n_197) );
INVx1_ASAP7_75t_L g209 ( .A(n_150), .Y(n_209) );
INVx1_ASAP7_75t_L g223 ( .A(n_150), .Y(n_223) );
INVx1_ASAP7_75t_L g226 ( .A(n_150), .Y(n_226) );
INVx2_ASAP7_75t_L g236 ( .A(n_150), .Y(n_236) );
INVx1_ASAP7_75t_L g238 ( .A(n_150), .Y(n_238) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g511 ( .A(n_152), .B(n_512), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g181 ( .A1(n_153), .A2(n_182), .B(n_185), .Y(n_181) );
OAI22xp5_ASAP7_75t_L g192 ( .A1(n_153), .A2(n_159), .B1(n_193), .B2(n_195), .Y(n_192) );
OAI22xp5_ASAP7_75t_L g205 ( .A1(n_153), .A2(n_206), .B1(n_211), .B2(n_212), .Y(n_205) );
OAI22xp5_ASAP7_75t_L g220 ( .A1(n_153), .A2(n_159), .B1(n_221), .B2(n_224), .Y(n_220) );
OAI22xp5_ASAP7_75t_L g233 ( .A1(n_153), .A2(n_234), .B1(n_237), .B2(n_239), .Y(n_233) );
OAI22xp5_ASAP7_75t_L g255 ( .A1(n_153), .A2(n_212), .B1(n_256), .B2(n_257), .Y(n_255) );
OAI22xp5_ASAP7_75t_L g274 ( .A1(n_153), .A2(n_159), .B1(n_275), .B2(n_276), .Y(n_274) );
OAI22xp5_ASAP7_75t_L g490 ( .A1(n_153), .A2(n_491), .B1(n_492), .B2(n_493), .Y(n_490) );
OAI22xp5_ASAP7_75t_L g498 ( .A1(n_153), .A2(n_239), .B1(n_499), .B2(n_500), .Y(n_498) );
OAI22x1_ASAP7_75t_L g603 ( .A1(n_153), .A2(n_239), .B1(n_604), .B2(n_605), .Y(n_603) );
INVx6_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
O2A1O1Ixp5_ASAP7_75t_L g177 ( .A1(n_154), .A2(n_178), .B(n_179), .C(n_180), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_154), .A2(n_549), .B(n_550), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_154), .B(n_561), .Y(n_560) );
A2O1A1Ixp33_ASAP7_75t_L g618 ( .A1(n_154), .A2(n_557), .B(n_561), .C(n_564), .Y(n_618) );
BUFx8_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g161 ( .A(n_155), .Y(n_161) );
INVx1_ASAP7_75t_L g213 ( .A(n_155), .Y(n_213) );
INVx1_ASAP7_75t_L g514 ( .A(n_155), .Y(n_514) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx4_ASAP7_75t_L g179 ( .A(n_158), .Y(n_179) );
INVx1_ASAP7_75t_L g210 ( .A(n_158), .Y(n_210) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g493 ( .A(n_160), .Y(n_493) );
BUFx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g547 ( .A(n_161), .Y(n_547) );
AO31x2_ASAP7_75t_L g273 ( .A1(n_162), .A2(n_240), .A3(n_274), .B(n_277), .Y(n_273) );
AO21x2_ASAP7_75t_L g565 ( .A1(n_162), .A2(n_566), .B(n_574), .Y(n_565) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
NOR2xp33_ASAP7_75t_SL g216 ( .A(n_164), .B(n_217), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g241 ( .A(n_164), .B(n_242), .Y(n_241) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g170 ( .A(n_165), .Y(n_170) );
INVx2_ASAP7_75t_L g215 ( .A(n_165), .Y(n_215) );
OAI21xp33_ASAP7_75t_L g564 ( .A1(n_165), .A2(n_518), .B(n_559), .Y(n_564) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_166), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g168 ( .A(n_169), .B(n_170), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_170), .B(n_278), .Y(n_277) );
AND2x4_ASAP7_75t_L g435 ( .A(n_171), .B(n_336), .Y(n_435) );
INVx1_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx1_ASAP7_75t_L g264 ( .A(n_172), .Y(n_264) );
INVxp67_ASAP7_75t_SL g422 ( .A(n_172), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_173), .B(n_190), .Y(n_172) );
AND2x2_ASAP7_75t_L g252 ( .A(n_173), .B(n_191), .Y(n_252) );
INVx1_ASAP7_75t_L g293 ( .A(n_173), .Y(n_293) );
OAI21x1_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_176), .B(n_188), .Y(n_173) );
OAI21x1_ASAP7_75t_L g288 ( .A1(n_174), .A2(n_176), .B(n_188), .Y(n_288) );
INVx2_ASAP7_75t_SL g174 ( .A(n_175), .Y(n_174) );
INVx4_ASAP7_75t_L g189 ( .A(n_175), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_175), .B(n_200), .Y(n_199) );
BUFx3_ASAP7_75t_L g227 ( .A(n_175), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_175), .B(n_229), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_175), .B(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g531 ( .A(n_175), .B(n_494), .Y(n_531) );
OAI21x1_ASAP7_75t_L g176 ( .A1(n_177), .A2(n_181), .B(n_186), .Y(n_176) );
O2A1O1Ixp33_ASAP7_75t_L g543 ( .A1(n_179), .A2(n_544), .B(n_545), .C(n_546), .Y(n_543) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g196 ( .A(n_184), .Y(n_196) );
OAI22xp33_ASAP7_75t_L g571 ( .A1(n_184), .A2(n_226), .B1(n_572), .B2(n_573), .Y(n_571) );
INVx2_ASAP7_75t_SL g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_SL g240 ( .A(n_187), .Y(n_240) );
INVx2_ASAP7_75t_L g198 ( .A(n_189), .Y(n_198) );
NOR2x1_ASAP7_75t_L g551 ( .A(n_189), .B(n_552), .Y(n_551) );
INVx2_ASAP7_75t_L g284 ( .A(n_190), .Y(n_284) );
AND2x2_ASAP7_75t_L g348 ( .A(n_190), .B(n_287), .Y(n_348) );
INVx2_ASAP7_75t_L g190 ( .A(n_191), .Y(n_190) );
INVx1_ASAP7_75t_L g302 ( .A(n_191), .Y(n_302) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_191), .Y(n_355) );
OR2x2_ASAP7_75t_L g426 ( .A(n_191), .B(n_232), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g509 ( .A(n_194), .B(n_510), .Y(n_509) );
INVx2_ASAP7_75t_L g501 ( .A(n_197), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_197), .B(n_526), .Y(n_525) );
AO31x2_ASAP7_75t_L g489 ( .A1(n_198), .A2(n_490), .A3(n_494), .B(n_495), .Y(n_489) );
NAND4xp25_ASAP7_75t_L g304 ( .A(n_201), .B(n_305), .C(n_308), .D(n_310), .Y(n_304) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
AND2x2_ASAP7_75t_L g442 ( .A(n_202), .B(n_430), .Y(n_442) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_218), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_203), .B(n_271), .Y(n_270) );
AND2x4_ASAP7_75t_L g296 ( .A(n_203), .B(n_297), .Y(n_296) );
INVx2_ASAP7_75t_L g316 ( .A(n_203), .Y(n_316) );
INVx1_ASAP7_75t_L g333 ( .A(n_203), .Y(n_333) );
INVx1_ASAP7_75t_L g341 ( .A(n_203), .Y(n_341) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_203), .Y(n_455) );
INVx4_ASAP7_75t_SL g203 ( .A(n_204), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_204), .B(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g373 ( .A(n_204), .B(n_273), .Y(n_373) );
AND2x2_ASAP7_75t_L g381 ( .A(n_204), .B(n_219), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_204), .B(n_404), .Y(n_403) );
BUFx2_ASAP7_75t_L g446 ( .A(n_204), .Y(n_446) );
INVx1_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_209), .B(n_569), .Y(n_568) );
INVx1_ASAP7_75t_SL g212 ( .A(n_213), .Y(n_212) );
INVx1_ASAP7_75t_L g239 ( .A(n_213), .Y(n_239) );
AO31x2_ASAP7_75t_L g497 ( .A1(n_214), .A2(n_240), .A3(n_498), .B(n_502), .Y(n_497) );
AOI21x1_ASAP7_75t_L g506 ( .A1(n_214), .A2(n_507), .B(n_519), .Y(n_506) );
BUFx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g495 ( .A(n_215), .B(n_496), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_215), .B(n_503), .Y(n_502) );
INVx2_ASAP7_75t_L g575 ( .A(n_215), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g606 ( .A(n_215), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g250 ( .A(n_219), .Y(n_250) );
OR2x2_ASAP7_75t_L g311 ( .A(n_219), .B(n_273), .Y(n_311) );
INVx2_ASAP7_75t_L g318 ( .A(n_219), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_219), .B(n_271), .Y(n_342) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_219), .Y(n_429) );
OAI21xp33_ASAP7_75t_SL g523 ( .A1(n_222), .A2(n_524), .B(n_525), .Y(n_523) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AO31x2_ASAP7_75t_L g232 ( .A1(n_227), .A2(n_233), .A3(n_240), .B(n_241), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_230), .B(n_401), .Y(n_400) );
BUFx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
AND2x2_ASAP7_75t_L g253 ( .A(n_232), .B(n_254), .Y(n_253) );
BUFx2_ASAP7_75t_L g263 ( .A(n_232), .Y(n_263) );
INVx2_ASAP7_75t_L g281 ( .A(n_232), .Y(n_281) );
AND2x4_ASAP7_75t_L g313 ( .A(n_232), .B(n_285), .Y(n_313) );
OR2x2_ASAP7_75t_L g393 ( .A(n_232), .B(n_293), .Y(n_393) );
INVx2_ASAP7_75t_SL g235 ( .A(n_236), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_236), .B(n_517), .Y(n_516) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_239), .B(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_244), .B(n_248), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_245), .B(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g310 ( .A(n_245), .B(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_245), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_246), .B(n_316), .Y(n_324) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx2_ASAP7_75t_L g269 ( .A(n_247), .Y(n_269) );
OR2x2_ASAP7_75t_L g362 ( .A(n_247), .B(n_272), .Y(n_362) );
INVx1_ASAP7_75t_L g289 ( .A(n_248), .Y(n_289) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g261 ( .A(n_249), .Y(n_261) );
INVx1_ASAP7_75t_L g297 ( .A(n_250), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_252), .B(n_253), .Y(n_251) );
OAI322xp33_ASAP7_75t_L g265 ( .A1(n_252), .A2(n_266), .A3(n_279), .B1(n_282), .B2(n_289), .C1(n_290), .C2(n_294), .Y(n_265) );
AND2x4_ASAP7_75t_L g312 ( .A(n_252), .B(n_313), .Y(n_312) );
AOI211xp5_ASAP7_75t_SL g343 ( .A1(n_252), .A2(n_344), .B(n_345), .C(n_349), .Y(n_343) );
AND2x2_ASAP7_75t_L g363 ( .A(n_252), .B(n_253), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_252), .B(n_280), .Y(n_369) );
AND2x4_ASAP7_75t_SL g291 ( .A(n_253), .B(n_292), .Y(n_291) );
NAND3xp33_ASAP7_75t_L g382 ( .A(n_253), .B(n_309), .C(n_337), .Y(n_382) );
AND2x2_ASAP7_75t_L g413 ( .A(n_253), .B(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g280 ( .A(n_254), .B(n_281), .Y(n_280) );
INVx3_ASAP7_75t_L g285 ( .A(n_254), .Y(n_285) );
BUFx2_ASAP7_75t_L g353 ( .A(n_254), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_263), .B(n_287), .Y(n_286) );
NAND2x1_ASAP7_75t_L g327 ( .A(n_263), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g346 ( .A(n_263), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_264), .B(n_280), .Y(n_411) );
OR2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_270), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g354 ( .A(n_269), .B(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_273), .Y(n_307) );
AND2x4_ASAP7_75t_L g317 ( .A(n_273), .B(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g404 ( .A(n_273), .Y(n_404) );
INVx2_ASAP7_75t_L g425 ( .A(n_273), .Y(n_425) );
OAI22xp33_ASAP7_75t_L g437 ( .A1(n_279), .A2(n_438), .B1(n_440), .B2(n_441), .Y(n_437) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g349 ( .A(n_280), .B(n_350), .Y(n_349) );
AND2x4_ASAP7_75t_L g303 ( .A(n_281), .B(n_287), .Y(n_303) );
OR2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_286), .Y(n_282) );
INVx1_ASAP7_75t_L g322 ( .A(n_283), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
AND2x4_ASAP7_75t_L g292 ( .A(n_284), .B(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g414 ( .A(n_284), .Y(n_414) );
INVx2_ASAP7_75t_L g300 ( .A(n_285), .Y(n_300) );
AND2x2_ASAP7_75t_L g328 ( .A(n_285), .B(n_287), .Y(n_328) );
INVx3_ASAP7_75t_L g336 ( .A(n_285), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_285), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g321 ( .A(n_286), .Y(n_321) );
INVx2_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
BUFx2_ASAP7_75t_L g337 ( .A(n_288), .Y(n_337) );
OAI222xp33_ASAP7_75t_L g460 ( .A1(n_290), .A2(n_450), .B1(n_461), .B2(n_464), .C1(n_466), .C2(n_468), .Y(n_460) );
INVx3_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g401 ( .A(n_292), .Y(n_401) );
AND2x2_ASAP7_75t_L g465 ( .A(n_292), .B(n_335), .Y(n_465) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_295), .B(n_386), .Y(n_385) );
AOI221xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_304), .B1(n_312), .B2(n_314), .C(n_319), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVx1_ASAP7_75t_L g387 ( .A(n_300), .Y(n_387) );
INVx2_ASAP7_75t_L g449 ( .A(n_301), .Y(n_449) );
AND2x4_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx2_ASAP7_75t_L g350 ( .A(n_302), .Y(n_350) );
AND2x2_ASAP7_75t_L g386 ( .A(n_302), .B(n_387), .Y(n_386) );
AND2x4_ASAP7_75t_L g352 ( .A(n_303), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g378 ( .A(n_303), .B(n_379), .Y(n_378) );
INVx1_ASAP7_75t_L g467 ( .A(n_303), .Y(n_467) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g416 ( .A(n_307), .Y(n_416) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
AND2x2_ASAP7_75t_L g439 ( .A(n_309), .B(n_317), .Y(n_439) );
AND2x2_ASAP7_75t_L g462 ( .A(n_309), .B(n_463), .Y(n_462) );
OR2x2_ASAP7_75t_L g323 ( .A(n_311), .B(n_324), .Y(n_323) );
INVx2_ASAP7_75t_L g458 ( .A(n_311), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g399 ( .A1(n_312), .A2(n_366), .B1(n_400), .B2(n_402), .Y(n_399) );
OAI21xp5_ASAP7_75t_L g427 ( .A1(n_312), .A2(n_428), .B(n_431), .Y(n_427) );
INVxp67_ASAP7_75t_L g344 ( .A(n_313), .Y(n_344) );
INVx2_ASAP7_75t_SL g448 ( .A(n_313), .Y(n_448) );
AND2x4_ASAP7_75t_L g314 ( .A(n_315), .B(n_317), .Y(n_314) );
OR2x2_ASAP7_75t_L g361 ( .A(n_315), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g459 ( .A(n_315), .B(n_458), .Y(n_459) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g332 ( .A(n_317), .B(n_333), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_317), .B(n_341), .Y(n_357) );
INVx2_ASAP7_75t_L g384 ( .A(n_317), .Y(n_384) );
OAI22xp33_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_323), .B1(n_325), .B2(n_327), .Y(n_319) );
NOR2xp33_ASAP7_75t_SL g320 ( .A(n_321), .B(n_322), .Y(n_320) );
AOI22xp5_ASAP7_75t_L g407 ( .A1(n_321), .A2(n_395), .B1(n_408), .B2(n_410), .Y(n_407) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g417 ( .A(n_326), .B(n_418), .Y(n_417) );
AOI21xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_334), .B(n_338), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
INVx1_ASAP7_75t_L g398 ( .A(n_331), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_331), .B(n_381), .Y(n_409) );
INVx1_ASAP7_75t_L g367 ( .A(n_333), .Y(n_367) );
AND2x2_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_335), .B(n_348), .Y(n_440) );
INVx2_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
OAI21xp33_ASAP7_75t_L g453 ( .A1(n_336), .A2(n_454), .B(n_456), .Y(n_453) );
OAI21xp5_ASAP7_75t_SL g338 ( .A1(n_339), .A2(n_343), .B(n_351), .Y(n_338) );
BUFx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
OR2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
INVx1_ASAP7_75t_L g397 ( .A(n_342), .Y(n_397) );
INVx1_ASAP7_75t_L g463 ( .A(n_342), .Y(n_463) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
INVx1_ASAP7_75t_L g436 ( .A(n_346), .Y(n_436) );
OR2x2_ASAP7_75t_L g447 ( .A(n_347), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND3xp33_ASAP7_75t_L g351 ( .A(n_352), .B(n_354), .C(n_356), .Y(n_351) );
AOI22xp5_ASAP7_75t_L g412 ( .A1(n_352), .A2(n_413), .B1(n_415), .B2(n_417), .Y(n_412) );
INVx1_ASAP7_75t_L g379 ( .A(n_353), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_354), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g392 ( .A(n_355), .Y(n_392) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_357), .B(n_361), .Y(n_360) );
OAI221xp5_ASAP7_75t_L g419 ( .A1(n_357), .A2(n_420), .B1(n_423), .B2(n_426), .C(n_427), .Y(n_419) );
AOI21xp5_ASAP7_75t_L g358 ( .A1(n_359), .A2(n_363), .B(n_364), .Y(n_358) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_L g368 ( .A(n_362), .Y(n_368) );
OAI22xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_369), .B1(n_370), .B2(n_831), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AND2x4_ASAP7_75t_L g366 ( .A(n_367), .B(n_368), .Y(n_366) );
INVxp67_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx2_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
AND2x4_ASAP7_75t_L g451 ( .A(n_373), .B(n_429), .Y(n_451) );
NAND4xp25_ASAP7_75t_L g374 ( .A(n_375), .B(n_405), .C(n_432), .D(n_452), .Y(n_374) );
NOR2xp33_ASAP7_75t_L g375 ( .A(n_376), .B(n_388), .Y(n_375) );
OAI221xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_380), .B1(n_382), .B2(n_383), .C(n_385), .Y(n_376) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_378), .A2(n_435), .B1(n_457), .B2(n_459), .Y(n_456) );
INVx1_ASAP7_75t_L g431 ( .A(n_380), .Y(n_431) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g415 ( .A(n_381), .B(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_381), .B(n_424), .Y(n_423) );
NAND2x1_ASAP7_75t_L g468 ( .A(n_381), .B(n_469), .Y(n_468) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_383), .B(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g390 ( .A(n_387), .B(n_391), .Y(n_390) );
OAI21xp33_ASAP7_75t_SL g388 ( .A1(n_389), .A2(n_394), .B(n_399), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
NOR2x1_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g418 ( .A(n_404), .Y(n_418) );
AOI211xp5_ASAP7_75t_L g432 ( .A1(n_404), .A2(n_433), .B(n_437), .C(n_443), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g405 ( .A(n_406), .B(n_419), .Y(n_405) );
NAND2xp5_ASAP7_75t_SL g406 ( .A(n_407), .B(n_412), .Y(n_406) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
OR2x2_ASAP7_75t_L g466 ( .A(n_414), .B(n_467), .Y(n_466) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AND2x4_ASAP7_75t_L g428 ( .A(n_429), .B(n_430), .Y(n_428) );
INVx3_ASAP7_75t_L g470 ( .A(n_430), .Y(n_470) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
NAND2x1p5_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
OAI22xp33_ASAP7_75t_R g443 ( .A1(n_444), .A2(n_447), .B1(n_449), .B2(n_450), .Y(n_443) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AND2x4_ASAP7_75t_L g457 ( .A(n_446), .B(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_453), .B(n_460), .Y(n_452) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx3_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx4_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AOI221xp5_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_806), .B1(n_814), .B2(n_815), .C(n_819), .Y(n_478) );
INVx1_ASAP7_75t_L g805 ( .A(n_481), .Y(n_805) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AND2x4_ASAP7_75t_L g482 ( .A(n_483), .B(n_697), .Y(n_482) );
NOR2xp67_ASAP7_75t_L g483 ( .A(n_484), .B(n_639), .Y(n_483) );
NAND3xp33_ASAP7_75t_SL g484 ( .A(n_485), .B(n_576), .C(n_621), .Y(n_484) );
OAI21xp5_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_532), .B(n_553), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g576 ( .A1(n_486), .A2(n_577), .B1(n_596), .B2(n_608), .Y(n_576) );
AOI22x1_ASAP7_75t_L g701 ( .A1(n_486), .A2(n_702), .B1(n_706), .B2(n_707), .Y(n_701) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
OR2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_504), .Y(n_487) );
OR2x2_ASAP7_75t_L g662 ( .A(n_488), .B(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_489), .B(n_497), .Y(n_488) );
OR2x2_ASAP7_75t_L g537 ( .A(n_489), .B(n_497), .Y(n_537) );
AND2x2_ASAP7_75t_L g580 ( .A(n_489), .B(n_581), .Y(n_580) );
INVx2_ASAP7_75t_SL g588 ( .A(n_489), .Y(n_588) );
BUFx2_ASAP7_75t_L g638 ( .A(n_489), .Y(n_638) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_493), .A2(n_529), .B(n_530), .Y(n_528) );
OAI21x1_ASAP7_75t_L g557 ( .A1(n_493), .A2(n_558), .B(n_559), .Y(n_557) );
INVx1_ASAP7_75t_L g552 ( .A(n_494), .Y(n_552) );
AND2x2_ASAP7_75t_L g583 ( .A(n_497), .B(n_520), .Y(n_583) );
INVx1_ASAP7_75t_L g590 ( .A(n_497), .Y(n_590) );
INVx1_ASAP7_75t_L g595 ( .A(n_497), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_497), .B(n_588), .Y(n_657) );
INVx1_ASAP7_75t_L g678 ( .A(n_497), .Y(n_678) );
NOR2xp33_ASAP7_75t_L g748 ( .A(n_497), .B(n_581), .Y(n_748) );
INVx1_ASAP7_75t_L g641 ( .A(n_504), .Y(n_641) );
OR2x2_ASAP7_75t_L g693 ( .A(n_504), .B(n_657), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_505), .B(n_520), .Y(n_504) );
AND2x2_ASAP7_75t_L g538 ( .A(n_505), .B(n_539), .Y(n_538) );
OR2x2_ASAP7_75t_L g586 ( .A(n_505), .B(n_587), .Y(n_586) );
INVxp67_ASAP7_75t_L g592 ( .A(n_505), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_505), .B(n_535), .Y(n_669) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx2_ASAP7_75t_L g581 ( .A(n_506), .Y(n_581) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_515), .B(n_518), .Y(n_507) );
OAI21xp5_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_511), .B(n_513), .Y(n_508) );
BUFx4f_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_514), .B(n_527), .Y(n_526) );
INVx3_ASAP7_75t_L g535 ( .A(n_520), .Y(n_535) );
INVx1_ASAP7_75t_L g635 ( .A(n_520), .Y(n_635) );
AND2x2_ASAP7_75t_L g637 ( .A(n_520), .B(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g655 ( .A(n_520), .B(n_656), .Y(n_655) );
OR2x2_ASAP7_75t_L g677 ( .A(n_520), .B(n_678), .Y(n_677) );
NAND2x1p5_ASAP7_75t_SL g688 ( .A(n_520), .B(n_664), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_520), .B(n_595), .Y(n_778) );
AND2x4_ASAP7_75t_L g520 ( .A(n_521), .B(n_522), .Y(n_520) );
OAI21xp5_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_528), .B(n_531), .Y(n_522) );
AND2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_538), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g716 ( .A1(n_533), .A2(n_717), .B1(n_718), .B2(n_720), .Y(n_716) );
AND2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_536), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_534), .B(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_534), .B(n_773), .Y(n_772) );
OR2x2_ASAP7_75t_L g795 ( .A(n_534), .B(n_653), .Y(n_795) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AND2x4_ASAP7_75t_L g594 ( .A(n_535), .B(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_535), .B(n_664), .Y(n_663) );
OR2x2_ASAP7_75t_L g683 ( .A(n_535), .B(n_684), .Y(n_683) );
AND2x4_ASAP7_75t_L g634 ( .A(n_536), .B(n_635), .Y(n_634) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx2_ASAP7_75t_L g724 ( .A(n_537), .Y(n_724) );
OR2x2_ASAP7_75t_L g798 ( .A(n_537), .B(n_725), .Y(n_798) );
INVx1_ASAP7_75t_L g629 ( .A(n_538), .Y(n_629) );
INVx3_ASAP7_75t_L g633 ( .A(n_539), .Y(n_633) );
BUFx2_ASAP7_75t_L g644 ( .A(n_539), .Y(n_644) );
BUFx3_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g614 ( .A(n_540), .B(n_565), .Y(n_614) );
INVx2_ASAP7_75t_L g660 ( .A(n_540), .Y(n_660) );
INVx1_ASAP7_75t_L g692 ( .A(n_540), .Y(n_692) );
AND2x2_ASAP7_75t_L g705 ( .A(n_540), .B(n_602), .Y(n_705) );
AND2x2_ASAP7_75t_L g727 ( .A(n_540), .B(n_626), .Y(n_727) );
NAND2x1p5_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
OAI21x1_ASAP7_75t_L g542 ( .A1(n_543), .A2(n_548), .B(n_551), .Y(n_542) );
INVx2_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
HB1xp67_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g718 ( .A(n_554), .B(n_719), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_554), .B(n_727), .Y(n_726) );
AND2x2_ASAP7_75t_L g743 ( .A(n_554), .B(n_611), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_554), .B(n_745), .Y(n_744) );
AND2x4_ASAP7_75t_L g554 ( .A(n_555), .B(n_565), .Y(n_554) );
INVx2_ASAP7_75t_L g600 ( .A(n_555), .Y(n_600) );
AND2x2_ASAP7_75t_L g627 ( .A(n_555), .B(n_628), .Y(n_627) );
AOI21x1_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_560), .B(n_563), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g601 ( .A(n_565), .B(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g620 ( .A(n_565), .Y(n_620) );
INVx2_ASAP7_75t_L g628 ( .A(n_565), .Y(n_628) );
OR2x2_ASAP7_75t_L g648 ( .A(n_565), .B(n_602), .Y(n_648) );
AND2x2_ASAP7_75t_L g659 ( .A(n_565), .B(n_660), .Y(n_659) );
OAI221xp5_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_582), .B1(n_584), .B2(n_589), .C(n_591), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
OAI32xp33_ASAP7_75t_L g689 ( .A1(n_579), .A2(n_593), .A3(n_690), .B1(n_693), .B2(n_694), .Y(n_689) );
HB1xp67_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
INVx1_ASAP7_75t_L g679 ( .A(n_580), .Y(n_679) );
AND2x2_ASAP7_75t_L g715 ( .A(n_580), .B(n_594), .Y(n_715) );
INVx1_ASAP7_75t_L g779 ( .A(n_580), .Y(n_779) );
OR2x2_ASAP7_75t_L g653 ( .A(n_581), .B(n_588), .Y(n_653) );
INVx2_ASAP7_75t_L g664 ( .A(n_581), .Y(n_664) );
BUFx2_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g803 ( .A(n_583), .B(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVxp67_ASAP7_75t_L g790 ( .A(n_586), .Y(n_790) );
INVx1_ASAP7_75t_L g804 ( .A(n_586), .Y(n_804) );
OR2x2_ASAP7_75t_L g684 ( .A(n_587), .B(n_664), .Y(n_684) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
NOR2xp33_ASAP7_75t_L g706 ( .A(n_589), .B(n_684), .Y(n_706) );
INVx1_ASAP7_75t_L g737 ( .A(n_589), .Y(n_737) );
BUFx3_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g771 ( .A(n_590), .Y(n_771) );
OR2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
NAND2x1_ASAP7_75t_L g740 ( .A(n_592), .B(n_741), .Y(n_740) );
OAI21xp5_ASAP7_75t_SL g762 ( .A1(n_593), .A2(n_763), .B(n_768), .Y(n_762) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_SL g596 ( .A(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_598), .B(n_601), .Y(n_597) );
AND2x2_ASAP7_75t_L g672 ( .A(n_598), .B(n_614), .Y(n_672) );
INVxp67_ASAP7_75t_SL g802 ( .A(n_598), .Y(n_802) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g704 ( .A(n_599), .Y(n_704) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g686 ( .A(n_600), .B(n_660), .Y(n_686) );
AND2x2_ASAP7_75t_L g757 ( .A(n_600), .B(n_628), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_601), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g685 ( .A(n_601), .B(n_686), .Y(n_685) );
AND2x2_ASAP7_75t_L g764 ( .A(n_601), .B(n_765), .Y(n_764) );
INVx2_ASAP7_75t_L g613 ( .A(n_602), .Y(n_613) );
INVx2_ASAP7_75t_L g626 ( .A(n_602), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_602), .B(n_617), .Y(n_674) );
AND2x2_ASAP7_75t_L g734 ( .A(n_602), .B(n_628), .Y(n_734) );
NAND2xp33_ASAP7_75t_SL g608 ( .A(n_609), .B(n_615), .Y(n_608) );
INVx2_ASAP7_75t_SL g609 ( .A(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_614), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g709 ( .A(n_612), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_612), .B(n_692), .Y(n_784) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
OR2x2_ASAP7_75t_L g616 ( .A(n_613), .B(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g745 ( .A(n_613), .B(n_660), .Y(n_745) );
OR2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_619), .Y(n_615) );
OR2x2_ASAP7_75t_L g690 ( .A(n_616), .B(n_691), .Y(n_690) );
INVx2_ASAP7_75t_L g647 ( .A(n_617), .Y(n_647) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
OR2x2_ASAP7_75t_L g673 ( .A(n_620), .B(n_674), .Y(n_673) );
AOI22xp5_ASAP7_75t_L g621 ( .A1(n_622), .A2(n_634), .B1(n_636), .B2(n_637), .Y(n_621) );
OAI21xp33_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_629), .B(n_630), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g636 ( .A(n_624), .B(n_633), .Y(n_636) );
BUFx2_ASAP7_75t_L g654 ( .A(n_624), .Y(n_654) );
AND2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_627), .Y(n_624) );
INVx1_ASAP7_75t_L g665 ( .A(n_625), .Y(n_665) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g680 ( .A(n_627), .B(n_644), .Y(n_680) );
INVx2_ASAP7_75t_L g696 ( .A(n_627), .Y(n_696) );
AND2x2_ASAP7_75t_L g738 ( .A(n_627), .B(n_660), .Y(n_738) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g713 ( .A(n_633), .B(n_714), .Y(n_713) );
AND2x2_ASAP7_75t_L g760 ( .A(n_634), .B(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g791 ( .A(n_635), .Y(n_791) );
INVx2_ASAP7_75t_L g730 ( .A(n_638), .Y(n_730) );
NAND4xp25_ASAP7_75t_L g639 ( .A(n_640), .B(n_649), .C(n_666), .D(n_681), .Y(n_639) );
NAND2xp33_ASAP7_75t_SL g640 ( .A(n_641), .B(n_642), .Y(n_640) );
AOI221xp5_ASAP7_75t_L g735 ( .A1(n_642), .A2(n_720), .B1(n_736), .B2(n_738), .C(n_739), .Y(n_735) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
NAND2x1_ASAP7_75t_L g643 ( .A(n_644), .B(n_645), .Y(n_643) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g717 ( .A(n_646), .Y(n_717) );
OR2x2_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
INVx2_ASAP7_75t_L g710 ( .A(n_647), .Y(n_710) );
INVx2_ASAP7_75t_L g782 ( .A(n_648), .Y(n_782) );
AOI222xp33_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_654), .B1(n_655), .B2(n_658), .C1(n_661), .C2(n_665), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g736 ( .A(n_652), .B(n_737), .Y(n_736) );
AOI21xp5_ASAP7_75t_L g763 ( .A1(n_652), .A2(n_764), .B(n_766), .Y(n_763) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
OR2x2_ASAP7_75t_L g775 ( .A(n_653), .B(n_719), .Y(n_775) );
OAI21xp33_ASAP7_75t_SL g749 ( .A1(n_654), .A2(n_675), .B(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
OR2x2_ASAP7_75t_L g668 ( .A(n_657), .B(n_669), .Y(n_668) );
INVxp67_ASAP7_75t_SL g720 ( .A(n_657), .Y(n_720) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
BUFx2_ASAP7_75t_L g719 ( .A(n_660), .Y(n_719) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g725 ( .A(n_664), .Y(n_725) );
AOI22xp33_ASAP7_75t_SL g666 ( .A1(n_667), .A2(n_670), .B1(n_675), .B2(n_680), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_671), .B(n_673), .Y(n_670) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AOI221xp5_ASAP7_75t_L g681 ( .A1(n_672), .A2(n_682), .B1(n_685), .B2(n_687), .C(n_689), .Y(n_681) );
INVx3_ASAP7_75t_R g796 ( .A(n_673), .Y(n_796) );
INVx1_ASAP7_75t_L g714 ( .A(n_674), .Y(n_714) );
INVx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OR2x2_ASAP7_75t_L g676 ( .A(n_677), .B(n_679), .Y(n_676) );
INVxp67_ASAP7_75t_SL g731 ( .A(n_677), .Y(n_731) );
INVx1_ASAP7_75t_L g741 ( .A(n_677), .Y(n_741) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_686), .B(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g759 ( .A(n_686), .Y(n_759) );
AND2x2_ASAP7_75t_L g787 ( .A(n_686), .B(n_734), .Y(n_787) );
INVx2_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
AND2x2_ASAP7_75t_L g781 ( .A(n_691), .B(n_782), .Y(n_781) );
INVx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx3_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
NOR2x1_ASAP7_75t_L g697 ( .A(n_698), .B(n_753), .Y(n_697) );
NAND3xp33_ASAP7_75t_L g698 ( .A(n_699), .B(n_735), .C(n_749), .Y(n_698) );
NOR3xp33_ASAP7_75t_L g699 ( .A(n_700), .B(n_711), .C(n_721), .Y(n_699) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
OAI21xp33_ASAP7_75t_L g712 ( .A1(n_702), .A2(n_713), .B(n_715), .Y(n_712) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_704), .B(n_705), .Y(n_703) );
INVx1_ASAP7_75t_L g752 ( .A(n_704), .Y(n_752) );
AND2x2_ASAP7_75t_L g793 ( .A(n_704), .B(n_782), .Y(n_793) );
NAND2x1_ASAP7_75t_L g751 ( .A(n_705), .B(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
INVx1_ASAP7_75t_L g773 ( .A(n_710), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_712), .B(n_716), .Y(n_711) );
INVx1_ASAP7_75t_L g765 ( .A(n_719), .Y(n_765) );
OAI22xp33_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_726), .B1(n_728), .B2(n_732), .Y(n_721) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .Y(n_723) );
INVx1_ASAP7_75t_L g761 ( .A(n_725), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g767 ( .A(n_727), .B(n_757), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_729), .B(n_731), .Y(n_728) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g800 ( .A(n_733), .Y(n_800) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
OAI22xp33_ASAP7_75t_SL g739 ( .A1(n_740), .A2(n_742), .B1(n_744), .B2(n_746), .Y(n_739) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
HB1xp67_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx2_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_754), .B(n_780), .Y(n_753) );
O2A1O1Ixp33_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_758), .B(n_760), .C(n_762), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
OAI21xp33_ASAP7_75t_L g769 ( .A1(n_756), .A2(n_770), .B(n_772), .Y(n_769) );
INVx2_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
O2A1O1Ixp5_ASAP7_75t_SL g780 ( .A1(n_760), .A2(n_781), .B(n_783), .C(n_785), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_764), .A2(n_769), .B1(n_774), .B2(n_776), .Y(n_768) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
OR2x2_ASAP7_75t_L g777 ( .A(n_778), .B(n_779), .Y(n_777) );
INVx2_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
OAI211xp5_ASAP7_75t_L g785 ( .A1(n_786), .A2(n_788), .B(n_792), .C(n_799), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
INVx2_ASAP7_75t_L g788 ( .A(n_789), .Y(n_788) );
AND2x2_ASAP7_75t_L g789 ( .A(n_790), .B(n_791), .Y(n_789) );
AOI22xp5_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_794), .B1(n_796), .B2(n_797), .Y(n_792) );
INVx2_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
INVx2_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
OAI21xp5_ASAP7_75t_SL g799 ( .A1(n_800), .A2(n_801), .B(n_803), .Y(n_799) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
NOR2x1_ASAP7_75t_R g806 ( .A(n_807), .B(n_813), .Y(n_806) );
NOR2xp67_ASAP7_75t_SL g815 ( .A(n_807), .B(n_816), .Y(n_815) );
INVx5_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
AND2x6_ASAP7_75t_SL g808 ( .A(n_809), .B(n_810), .Y(n_808) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx4_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
CKINVDCx5p33_ASAP7_75t_R g817 ( .A(n_818), .Y(n_817) );
AND2x2_ASAP7_75t_L g826 ( .A(n_818), .B(n_827), .Y(n_826) );
NOR2xp33_ASAP7_75t_L g819 ( .A(n_820), .B(n_821), .Y(n_819) );
BUFx6f_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
INVx2_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
BUFx10_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx5_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
endmodule