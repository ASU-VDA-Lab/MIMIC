module fake_jpeg_22010_n_325 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_325);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_325;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_SL g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx5_ASAP7_75t_SL g28 ( 
.A(n_27),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_28),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_17),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_20),
.Y(n_42)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_34),
.Y(n_43)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

OAI21xp33_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_47),
.B(n_49),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_31),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_46),
.Y(n_73)
);

AND2x2_ASAP7_75t_SL g47 ( 
.A(n_28),
.B(n_27),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_32),
.A2(n_24),
.B1(n_20),
.B2(n_16),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_48),
.A2(n_32),
.B1(n_24),
.B2(n_20),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_28),
.B(n_17),
.Y(n_49)
);

AOI21xp33_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_24),
.B(n_27),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_51),
.Y(n_64)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_54),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_63),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_62),
.A2(n_32),
.B1(n_13),
.B2(n_23),
.Y(n_97)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_68),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_67),
.Y(n_83)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_69),
.B(n_75),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_37),
.Y(n_72)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx3_ASAP7_75t_SL g84 ( 
.A(n_74),
.Y(n_84)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_77),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_47),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_82),
.B(n_87),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_73),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_88),
.Y(n_102)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_93),
.Y(n_108)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_94),
.A2(n_97),
.B1(n_98),
.B2(n_61),
.Y(n_109)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_61),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_56),
.B(n_47),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_82),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_67),
.B(n_51),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_100),
.A2(n_47),
.B(n_52),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_85),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_106),
.Y(n_124)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_103),
.B(n_114),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_105),
.B(n_37),
.Y(n_148)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_80),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_111),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_109),
.A2(n_112),
.B1(n_115),
.B2(n_123),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_110),
.A2(n_121),
.B(n_81),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_80),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_100),
.A2(n_32),
.B1(n_52),
.B2(n_50),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_52),
.C(n_36),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_81),
.C(n_93),
.Y(n_144)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_100),
.A2(n_50),
.B1(n_41),
.B2(n_36),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_97),
.A2(n_86),
.B1(n_96),
.B2(n_36),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_116),
.A2(n_78),
.B1(n_79),
.B2(n_84),
.Y(n_127)
);

FAx1_ASAP7_75t_SL g117 ( 
.A(n_96),
.B(n_49),
.CI(n_27),
.CON(n_117),
.SN(n_117)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_117),
.B(n_14),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_94),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_119),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_89),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_86),
.A2(n_14),
.B(n_46),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_120),
.A2(n_114),
.B(n_103),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_78),
.B(n_27),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_79),
.Y(n_122)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_84),
.A2(n_50),
.B1(n_41),
.B2(n_35),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_132),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_110),
.A2(n_113),
.B(n_104),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_126),
.A2(n_129),
.B(n_131),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_127),
.A2(n_128),
.B1(n_142),
.B2(n_57),
.Y(n_164)
);

AO22x2_ASAP7_75t_SL g128 ( 
.A1(n_112),
.A2(n_40),
.B1(n_16),
.B2(n_26),
.Y(n_128)
);

OA21x2_ASAP7_75t_L g130 ( 
.A1(n_116),
.A2(n_49),
.B(n_26),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_130),
.A2(n_140),
.B(n_141),
.Y(n_150)
);

O2A1O1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_104),
.A2(n_16),
.B(n_26),
.C(n_59),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_135),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_137),
.A2(n_141),
.B(n_129),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_120),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_107),
.A2(n_84),
.B1(n_88),
.B2(n_87),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_143),
.A2(n_149),
.B(n_37),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_121),
.C(n_118),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_101),
.B(n_31),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_145),
.Y(n_156)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_119),
.Y(n_146)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_146),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_117),
.B(n_95),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_147),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_121),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_SL g149 ( 
.A1(n_111),
.A2(n_70),
.B(n_92),
.C(n_83),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_135),
.A2(n_105),
.B1(n_106),
.B2(n_122),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_153),
.A2(n_163),
.B1(n_174),
.B2(n_149),
.Y(n_187)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_117),
.Y(n_154)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_154),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_155),
.B(n_171),
.C(n_172),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_157),
.B(n_175),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_158),
.A2(n_90),
.B1(n_34),
.B2(n_35),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_126),
.B(n_148),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_159),
.B(n_162),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_139),
.A2(n_83),
.B1(n_92),
.B2(n_63),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_160),
.A2(n_167),
.B1(n_173),
.B2(n_176),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_127),
.A2(n_140),
.B1(n_143),
.B2(n_142),
.Y(n_163)
);

OA22x2_ASAP7_75t_L g188 ( 
.A1(n_164),
.A2(n_166),
.B1(n_25),
.B2(n_19),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_133),
.A2(n_14),
.B(n_23),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_128),
.A2(n_92),
.B1(n_83),
.B2(n_98),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_124),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_168),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_128),
.B(n_0),
.Y(n_170)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_170),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_134),
.B(n_35),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_55),
.C(n_53),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_131),
.A2(n_41),
.B1(n_66),
.B2(n_60),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_130),
.A2(n_68),
.B1(n_65),
.B2(n_74),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_136),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_130),
.A2(n_90),
.B1(n_76),
.B2(n_95),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_149),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_177),
.B(n_149),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_181),
.A2(n_203),
.B(n_170),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_132),
.Y(n_184)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_184),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_159),
.B(n_125),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_185),
.B(n_193),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_138),
.Y(n_186)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_186),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_187),
.A2(n_190),
.B1(n_160),
.B2(n_199),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_188),
.B(n_191),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_153),
.B(n_95),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_189),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_177),
.A2(n_90),
.B1(n_53),
.B2(n_55),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_152),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_167),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_192),
.B(n_195),
.Y(n_217)
);

XOR2x1_ASAP7_75t_L g193 ( 
.A(n_157),
.B(n_25),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_194),
.A2(n_174),
.B1(n_53),
.B2(n_35),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_172),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_18),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_196),
.B(n_199),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_165),
.B(n_18),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_163),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_200),
.B(n_201),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_173),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_165),
.B(n_169),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_202),
.Y(n_218)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_158),
.Y(n_203)
);

BUFx12f_ASAP7_75t_SL g205 ( 
.A(n_193),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_205),
.A2(n_226),
.B(n_196),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_155),
.C(n_162),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_206),
.B(n_212),
.C(n_178),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_207),
.A2(n_187),
.B1(n_192),
.B2(n_205),
.Y(n_231)
);

INVxp67_ASAP7_75t_SL g208 ( 
.A(n_189),
.Y(n_208)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_208),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_185),
.B(n_150),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_225),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_154),
.C(n_150),
.Y(n_212)
);

INVx13_ASAP7_75t_L g215 ( 
.A(n_186),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_215),
.B(n_188),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_179),
.B(n_156),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_216),
.B(n_222),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_219),
.A2(n_197),
.B1(n_195),
.B2(n_182),
.Y(n_240)
);

BUFx12f_ASAP7_75t_L g220 ( 
.A(n_184),
.Y(n_220)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_220),
.Y(n_235)
);

HB1xp67_ASAP7_75t_L g221 ( 
.A(n_190),
.Y(n_221)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_221),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_180),
.B(n_166),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_178),
.B(n_154),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_220),
.Y(n_228)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_228),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_19),
.C(n_34),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_212),
.B(n_202),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_230),
.B(n_242),
.Y(n_262)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_231),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_211),
.A2(n_203),
.B1(n_181),
.B2(n_183),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_232),
.B(n_236),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_218),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_233),
.A2(n_240),
.B1(n_247),
.B2(n_34),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_218),
.A2(n_183),
.B1(n_182),
.B2(n_176),
.Y(n_236)
);

HB1xp67_ASAP7_75t_L g238 ( 
.A(n_220),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_238),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_206),
.B(n_217),
.C(n_204),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_245),
.C(n_242),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_223),
.A2(n_188),
.B(n_170),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_243),
.B(n_244),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_209),
.B(n_197),
.C(n_188),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_15),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_13),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_219),
.A2(n_223),
.B1(n_226),
.B2(n_210),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_247),
.A2(n_207),
.B1(n_225),
.B2(n_75),
.Y(n_248)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_248),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_250),
.A2(n_257),
.B1(n_43),
.B2(n_25),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_227),
.B(n_12),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_243),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_255),
.C(n_260),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_43),
.C(n_15),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_245),
.A2(n_31),
.B1(n_34),
.B2(n_13),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_261),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_229),
.B(n_30),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_235),
.B(n_43),
.C(n_33),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_265),
.C(n_266),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_234),
.B(n_10),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_264),
.B(n_0),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_230),
.B(n_43),
.C(n_33),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_237),
.B(n_227),
.C(n_241),
.Y(n_266)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_268),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_30),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_269),
.B(n_277),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_258),
.A2(n_23),
.B1(n_10),
.B2(n_12),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_270),
.B(n_271),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_252),
.A2(n_12),
.B1(n_1),
.B2(n_2),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_281),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_254),
.A2(n_22),
.B1(n_18),
.B2(n_2),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_273),
.B(n_274),
.Y(n_285)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_253),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_249),
.A2(n_30),
.B(n_29),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_30),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_33),
.C(n_22),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_262),
.A2(n_0),
.B(n_1),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_280),
.B(n_3),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_256),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_282),
.B(n_3),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_267),
.A2(n_266),
.B1(n_265),
.B2(n_255),
.Y(n_283)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_283),
.Y(n_300)
);

FAx1_ASAP7_75t_SL g286 ( 
.A(n_268),
.B(n_263),
.CI(n_22),
.CON(n_286),
.SN(n_286)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_286),
.B(n_293),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_29),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_291),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_275),
.A2(n_22),
.B1(n_18),
.B2(n_5),
.Y(n_290)
);

O2A1O1Ixp33_ASAP7_75t_L g296 ( 
.A1(n_290),
.A2(n_269),
.B(n_272),
.C(n_280),
.Y(n_296)
);

OAI22xp33_ASAP7_75t_L g298 ( 
.A1(n_292),
.A2(n_284),
.B1(n_285),
.B2(n_288),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_29),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_279),
.Y(n_299)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_296),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_278),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_297),
.B(n_304),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_299),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_286),
.A2(n_275),
.B1(n_6),
.B2(n_7),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_301),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_SL g302 ( 
.A(n_289),
.B(n_33),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_295),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_294),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_304)
);

AOI211xp5_ASAP7_75t_L g305 ( 
.A1(n_292),
.A2(n_33),
.B(n_7),
.C(n_8),
.Y(n_305)
);

AO21x1_ASAP7_75t_L g308 ( 
.A1(n_305),
.A2(n_4),
.B(n_7),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_308),
.B(n_8),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_311),
.B(n_306),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_300),
.A2(n_4),
.B(n_8),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_312),
.B(n_306),
.C(n_303),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_299),
.Y(n_314)
);

AO21x1_ASAP7_75t_L g318 ( 
.A1(n_314),
.A2(n_315),
.B(n_316),
.Y(n_318)
);

MAJx2_ASAP7_75t_L g319 ( 
.A(n_317),
.B(n_310),
.C(n_307),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_319),
.B(n_314),
.C(n_318),
.Y(n_320)
);

NOR2xp67_ASAP7_75t_L g321 ( 
.A(n_320),
.B(n_309),
.Y(n_321)
);

INVxp33_ASAP7_75t_L g322 ( 
.A(n_321),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_9),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_323),
.B(n_9),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_9),
.B(n_145),
.Y(n_325)
);


endmodule