module fake_jpeg_26544_n_34 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_34);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_34;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_32;
wire n_15;

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_SL g17 ( 
.A(n_3),
.B(n_6),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_15),
.A2(n_7),
.B1(n_10),
.B2(n_9),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_18),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_26)
);

INVx1_ASAP7_75t_SL g19 ( 
.A(n_16),
.Y(n_19)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_17),
.B(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_26),
.A2(n_19),
.B1(n_14),
.B2(n_13),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_28),
.A2(n_26),
.B1(n_23),
.B2(n_25),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_22),
.C(n_12),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_29),
.B(n_30),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_27),
.A2(n_0),
.B(n_1),
.Y(n_30)
);

AOI322xp5_ASAP7_75t_L g33 ( 
.A1(n_32),
.A2(n_2),
.A3(n_4),
.B1(n_5),
.B2(n_8),
.C1(n_31),
.C2(n_26),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_32),
.C(n_2),
.Y(n_34)
);


endmodule