module fake_jpeg_15374_n_158 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_158);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_158;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx11_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx6_ASAP7_75t_SL g28 ( 
.A(n_6),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_6),
.B(n_4),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_4),
.B(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_34),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx5_ASAP7_75t_SL g34 ( 
.A(n_28),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_40),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_14),
.A2(n_1),
.B1(n_2),
.B2(n_5),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_36),
.A2(n_38),
.B1(n_23),
.B2(n_24),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_16),
.A2(n_1),
.B1(n_5),
.B2(n_6),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_39),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_5),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

HAxp5_ASAP7_75t_SL g42 ( 
.A(n_30),
.B(n_7),
.CON(n_42),
.SN(n_42)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_42),
.A2(n_19),
.B(n_18),
.Y(n_64)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_15),
.A2(n_7),
.B1(n_12),
.B2(n_10),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_45),
.A2(n_31),
.B1(n_17),
.B2(n_26),
.Y(n_59)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_47),
.Y(n_57)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_30),
.B(n_20),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_51),
.Y(n_61)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_25),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_25),
.B(n_27),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_21),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_54),
.B(n_58),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_32),
.B(n_31),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_55),
.A2(n_64),
.B(n_69),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_21),
.Y(n_58)
);

OA22x2_ASAP7_75t_L g95 ( 
.A1(n_59),
.A2(n_62),
.B1(n_52),
.B2(n_65),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_26),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_66),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_19),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_13),
.Y(n_67)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_50),
.B(n_13),
.Y(n_68)
);

NOR3xp33_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_70),
.C(n_78),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_39),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_38),
.B(n_18),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_72),
.A2(n_63),
.B1(n_61),
.B2(n_56),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_23),
.Y(n_76)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_24),
.Y(n_77)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_43),
.B(n_27),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_37),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_73),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_70),
.A2(n_33),
.B1(n_34),
.B2(n_66),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_82),
.A2(n_89),
.B1(n_92),
.B2(n_100),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_71),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_90),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_86),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_54),
.B(n_53),
.C(n_58),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_57),
.C(n_78),
.Y(n_105)
);

NOR2x1_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_64),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_88),
.A2(n_101),
.B(n_99),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_75),
.B1(n_53),
.B2(n_65),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_67),
.Y(n_91)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_77),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_93),
.B(n_99),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_95),
.A2(n_98),
.B1(n_94),
.B2(n_96),
.Y(n_110)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_55),
.B(n_69),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_52),
.A2(n_61),
.B1(n_60),
.B2(n_73),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_62),
.A2(n_60),
.B1(n_76),
.B2(n_56),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_98),
.Y(n_102)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_103),
.Y(n_130)
);

OR2x6_ASAP7_75t_L g104 ( 
.A(n_88),
.B(n_69),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_104),
.A2(n_83),
.B(n_116),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_105),
.B(n_82),
.Y(n_123)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_106),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_80),
.C(n_85),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_117),
.C(n_95),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_92),
.B(n_97),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_108),
.B(n_114),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_104),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_96),
.B(n_90),
.Y(n_112)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_112),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_100),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_85),
.C(n_97),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_101),
.B(n_81),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_123),
.B(n_126),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_107),
.B(n_89),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_124),
.B(n_127),
.C(n_117),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_126),
.A2(n_128),
.B1(n_110),
.B2(n_103),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_115),
.A2(n_83),
.B1(n_95),
.B2(n_104),
.Y(n_128)
);

AO22x1_ASAP7_75t_L g138 ( 
.A1(n_131),
.A2(n_115),
.B1(n_129),
.B2(n_123),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_133),
.C(n_134),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_105),
.C(n_113),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_104),
.C(n_109),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_104),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_136),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_139),
.Y(n_146)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_138),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_122),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_131),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_140),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_120),
.C(n_125),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_141),
.Y(n_148)
);

NOR3xp33_ASAP7_75t_SL g144 ( 
.A(n_138),
.B(n_125),
.C(n_140),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_144),
.B(n_136),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_R g153 ( 
.A(n_149),
.B(n_150),
.C(n_151),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_146),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_142),
.A2(n_143),
.B1(n_148),
.B2(n_147),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_151),
.B(n_152),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_145),
.B(n_132),
.C(n_147),
.Y(n_152)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_153),
.Y(n_155)
);

BUFx24_ASAP7_75t_SL g156 ( 
.A(n_154),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_152),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_155),
.Y(n_158)
);


endmodule