module fake_jpeg_20325_n_319 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_319);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_319;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_26),
.B(n_0),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g75 ( 
.A(n_43),
.B(n_45),
.Y(n_75)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_10),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_50),
.Y(n_51)
);

OAI22xp33_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_24),
.B1(n_38),
.B2(n_29),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_52),
.A2(n_57),
.B1(n_65),
.B2(n_69),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_54),
.B(n_64),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_24),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_58),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_50),
.A2(n_24),
.B1(n_17),
.B2(n_29),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_43),
.B(n_17),
.Y(n_58)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_43),
.B(n_29),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_62),
.B(n_74),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_39),
.B(n_19),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_48),
.A2(n_34),
.B1(n_20),
.B2(n_21),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_19),
.Y(n_67)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_67),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_37),
.Y(n_68)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_48),
.A2(n_18),
.B1(n_21),
.B2(n_32),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_46),
.B(n_28),
.Y(n_72)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_47),
.B(n_42),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_28),
.Y(n_76)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

AND2x4_ASAP7_75t_L g77 ( 
.A(n_47),
.B(n_35),
.Y(n_77)
);

OAI21xp33_ASAP7_75t_L g93 ( 
.A1(n_77),
.A2(n_47),
.B(n_36),
.Y(n_93)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_78),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_77),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_81),
.B(n_51),
.Y(n_128)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_82),
.Y(n_137)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_75),
.A2(n_46),
.B1(n_31),
.B2(n_30),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_84),
.A2(n_87),
.B1(n_92),
.B2(n_100),
.Y(n_126)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_75),
.A2(n_31),
.B1(n_30),
.B2(n_22),
.Y(n_87)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_66),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_89),
.B(n_105),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_77),
.A2(n_41),
.B1(n_21),
.B2(n_18),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_91),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_75),
.A2(n_42),
.B1(n_40),
.B2(n_22),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_93),
.B(n_61),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_95),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_52),
.A2(n_41),
.B1(n_18),
.B2(n_32),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_96),
.A2(n_117),
.B1(n_63),
.B2(n_73),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_53),
.Y(n_98)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_98),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_77),
.A2(n_27),
.B1(n_32),
.B2(n_36),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_99),
.A2(n_114),
.B(n_20),
.Y(n_130)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_55),
.A2(n_23),
.B(n_27),
.C(n_34),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g142 ( 
.A1(n_102),
.A2(n_99),
.B(n_85),
.C(n_104),
.Y(n_142)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_109),
.Y(n_134)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_59),
.Y(n_108)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

INVxp33_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_66),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_113),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_58),
.A2(n_47),
.B(n_2),
.Y(n_114)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_51),
.Y(n_115)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_61),
.Y(n_116)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_71),
.A2(n_26),
.B1(n_20),
.B2(n_34),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_62),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_118),
.B(n_149),
.Y(n_156)
);

NAND2xp33_ASAP7_75t_SL g120 ( 
.A(n_109),
.B(n_47),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_120),
.A2(n_130),
.B(n_147),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_78),
.C(n_42),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_124),
.B(n_86),
.C(n_106),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_90),
.B(n_15),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_125),
.B(n_9),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_126),
.B(n_145),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_128),
.B(n_148),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_83),
.A2(n_112),
.B1(n_94),
.B2(n_102),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_131),
.A2(n_133),
.B1(n_139),
.B2(n_150),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_101),
.A2(n_60),
.B1(n_63),
.B2(n_73),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_132),
.A2(n_151),
.B1(n_0),
.B2(n_5),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_94),
.A2(n_63),
.B1(n_73),
.B2(n_59),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_81),
.A2(n_71),
.B1(n_70),
.B2(n_59),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_138),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_97),
.A2(n_70),
.B1(n_12),
.B2(n_4),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_142),
.A2(n_35),
.B(n_5),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_80),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_88),
.Y(n_146)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_146),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_25),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_80),
.B(n_25),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_103),
.A2(n_35),
.B1(n_2),
.B2(n_0),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_115),
.A2(n_11),
.B1(n_5),
.B2(n_6),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_88),
.Y(n_153)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_153),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_135),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_154),
.B(n_163),
.Y(n_195)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

INVx8_ASAP7_75t_L g191 ( 
.A(n_157),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_118),
.B(n_110),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_158),
.B(n_182),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_160),
.A2(n_166),
.B(n_151),
.Y(n_188)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_121),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_161),
.B(n_167),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_127),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_164),
.B(n_128),
.C(n_136),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_143),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_165),
.B(n_168),
.Y(n_209)
);

OA21x2_ASAP7_75t_L g166 ( 
.A1(n_140),
.A2(n_98),
.B(n_82),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_119),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_125),
.B(n_105),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_122),
.A2(n_113),
.B1(n_108),
.B2(n_107),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_170),
.A2(n_172),
.B1(n_179),
.B2(n_183),
.Y(n_214)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_129),
.Y(n_171)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_171),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_133),
.A2(n_152),
.B1(n_122),
.B2(n_140),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_143),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_174),
.B(n_184),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_145),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g210 ( 
.A(n_175),
.B(n_137),
.Y(n_210)
);

FAx1_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_130),
.CI(n_152),
.CON(n_177),
.SN(n_177)
);

MAJIxp5_ASAP7_75t_SL g202 ( 
.A(n_177),
.B(n_120),
.C(n_128),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_147),
.A2(n_106),
.B1(n_116),
.B2(n_8),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_180),
.B(n_126),
.Y(n_199)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_129),
.Y(n_181)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_181),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_124),
.B(n_8),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_147),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_134),
.Y(n_185)
);

INVxp33_ASAP7_75t_L g212 ( 
.A(n_185),
.Y(n_212)
);

NOR2x1_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_142),
.Y(n_187)
);

NAND2xp33_ASAP7_75t_L g216 ( 
.A(n_187),
.B(n_160),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_188),
.A2(n_202),
.B(n_205),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_148),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_189),
.B(n_182),
.Y(n_235)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_167),
.Y(n_190)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_190),
.Y(n_232)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_157),
.Y(n_196)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_196),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_171),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_197),
.B(n_206),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_199),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_156),
.B(n_136),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_200),
.B(n_204),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_164),
.C(n_178),
.Y(n_221)
);

INVx5_ASAP7_75t_SL g203 ( 
.A(n_165),
.Y(n_203)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_203),
.Y(n_217)
);

AO22x1_ASAP7_75t_SL g204 ( 
.A1(n_177),
.A2(n_132),
.B1(n_149),
.B2(n_137),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_172),
.B(n_119),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_156),
.B(n_153),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_181),
.Y(n_207)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_207),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_161),
.Y(n_208)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_208),
.Y(n_228)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_210),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g211 ( 
.A(n_154),
.B(n_9),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_211),
.B(n_215),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_173),
.B(n_123),
.Y(n_213)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_213),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_216),
.B(n_219),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_187),
.B(n_177),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_235),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_225),
.C(n_236),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_205),
.A2(n_186),
.B1(n_169),
.B2(n_180),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_223),
.A2(n_230),
.B1(n_176),
.B2(n_204),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_195),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_224),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_158),
.C(n_186),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_205),
.A2(n_186),
.B1(n_169),
.B2(n_159),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_189),
.B(n_159),
.C(n_179),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_204),
.A2(n_200),
.B1(n_206),
.B2(n_202),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_237),
.A2(n_214),
.B1(n_185),
.B2(n_203),
.Y(n_251)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_208),
.Y(n_238)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_238),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_194),
.B(n_162),
.C(n_155),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_207),
.C(n_198),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_240),
.A2(n_248),
.B1(n_253),
.B2(n_229),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_194),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_235),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_217),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_242),
.B(n_256),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_209),
.Y(n_244)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_244),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_227),
.B(n_197),
.Y(n_246)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_246),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_227),
.A2(n_176),
.B1(n_210),
.B2(n_188),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_249),
.B(n_250),
.C(n_239),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_198),
.C(n_193),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_251),
.A2(n_252),
.B1(n_230),
.B2(n_223),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_237),
.A2(n_193),
.B1(n_191),
.B2(n_192),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_220),
.A2(n_211),
.B1(n_166),
.B2(n_183),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_162),
.Y(n_255)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_255),
.Y(n_267)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_222),
.Y(n_256)
);

AOI221xp5_ASAP7_75t_L g257 ( 
.A1(n_218),
.A2(n_212),
.B1(n_166),
.B2(n_155),
.C(n_123),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_226),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_259),
.B(n_265),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_229),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_261),
.B(n_275),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_245),
.B(n_233),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_262),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_273),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_243),
.B(n_247),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_258),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_266),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_268),
.B(n_271),
.C(n_272),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_270),
.A2(n_240),
.B1(n_244),
.B2(n_248),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_236),
.C(n_228),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_191),
.C(n_232),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_246),
.A2(n_212),
.B(n_238),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_243),
.B(n_226),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_242),
.Y(n_286)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_269),
.Y(n_276)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_276),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_263),
.A2(n_251),
.B1(n_252),
.B2(n_255),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_278),
.A2(n_280),
.B1(n_146),
.B2(n_144),
.Y(n_296)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_266),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_285),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_260),
.B(n_241),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_286),
.B(n_272),
.C(n_274),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_254),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_144),
.C(n_12),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_282),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_279),
.A2(n_267),
.B1(n_273),
.B2(n_268),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_296),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_SL g291 ( 
.A1(n_279),
.A2(n_275),
.B(n_261),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_282),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_288),
.A2(n_265),
.B(n_259),
.Y(n_292)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_292),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_278),
.A2(n_196),
.B1(n_232),
.B2(n_190),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_295),
.A2(n_284),
.B1(n_277),
.B2(n_286),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_297),
.B(n_10),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_283),
.C(n_297),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_300),
.B(n_301),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_277),
.C(n_287),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_302),
.B(n_304),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_294),
.B(n_293),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_305),
.A2(n_295),
.B(n_283),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_306),
.B(n_298),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_303),
.B(n_291),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_308),
.A2(n_310),
.B(n_305),
.Y(n_312)
);

OAI21x1_ASAP7_75t_SL g314 ( 
.A1(n_311),
.A2(n_312),
.B(n_313),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_309),
.B(n_299),
.Y(n_313)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g315 ( 
.A1(n_312),
.A2(n_307),
.B(n_301),
.C(n_15),
.D(n_16),
.Y(n_315)
);

AOI321xp33_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_13),
.A3(n_14),
.B1(n_15),
.B2(n_175),
.C(n_216),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_316),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_314),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_318),
.B(n_13),
.Y(n_319)
);


endmodule