module fake_netlist_1_5250_n_584 (n_117, n_44, n_133, n_149, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_125, n_9, n_161, n_10, n_130, n_103, n_19, n_87, n_137, n_104, n_160, n_98, n_74, n_154, n_7, n_29, n_165, n_146, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_139, n_16, n_13, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_24, n_78, n_6, n_4, n_127, n_40, n_111, n_157, n_79, n_38, n_64, n_142, n_46, n_31, n_58, n_122, n_138, n_126, n_118, n_32, n_0, n_84, n_131, n_112, n_55, n_12, n_86, n_143, n_166, n_162, n_75, n_163, n_105, n_159, n_72, n_136, n_43, n_76, n_89, n_68, n_144, n_27, n_53, n_67, n_77, n_20, n_2, n_147, n_54, n_148, n_123, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_150, n_3, n_18, n_110, n_66, n_134, n_1, n_164, n_82, n_106, n_15, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_96, n_39, n_584);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_125;
input n_9;
input n_161;
input n_10;
input n_130;
input n_103;
input n_19;
input n_87;
input n_137;
input n_104;
input n_160;
input n_98;
input n_74;
input n_154;
input n_7;
input n_29;
input n_165;
input n_146;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_139;
input n_16;
input n_13;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_127;
input n_40;
input n_111;
input n_157;
input n_79;
input n_38;
input n_64;
input n_142;
input n_46;
input n_31;
input n_58;
input n_122;
input n_138;
input n_126;
input n_118;
input n_32;
input n_0;
input n_84;
input n_131;
input n_112;
input n_55;
input n_12;
input n_86;
input n_143;
input n_166;
input n_162;
input n_75;
input n_163;
input n_105;
input n_159;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_68;
input n_144;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_54;
input n_148;
input n_123;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_164;
input n_82;
input n_106;
input n_15;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_96;
input n_39;
output n_584;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_431;
wire n_484;
wire n_496;
wire n_177;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_202;
wire n_386;
wire n_432;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_205;
wire n_330;
wire n_387;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_563;
wire n_517;
wire n_560;
wire n_479;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_533;
wire n_506;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_450;
wire n_579;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_379;
wire n_527;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_574;
wire n_217;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_178;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_295;
wire n_263;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_552;
wire n_344;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_429;
wire n_488;
wire n_233;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_300;
wire n_524;
wire n_497;
wire n_339;
wire n_583;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_198;
wire n_169;
wire n_424;
wire n_569;
wire n_297;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_187;
wire n_375;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_421;
wire n_175;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_137), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_9), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_1), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_126), .Y(n_171) );
OR2x2_ASAP7_75t_L g172 ( .A(n_96), .B(n_68), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_138), .Y(n_173) );
NOR2xp67_ASAP7_75t_L g174 ( .A(n_156), .B(n_143), .Y(n_174) );
CKINVDCx16_ASAP7_75t_R g175 ( .A(n_127), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_120), .Y(n_176) );
BUFx2_ASAP7_75t_L g177 ( .A(n_113), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_18), .Y(n_178) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_148), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_164), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_16), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_132), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_71), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_20), .Y(n_184) );
CKINVDCx5p33_ASAP7_75t_R g185 ( .A(n_112), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_7), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_82), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_50), .Y(n_188) );
CKINVDCx14_ASAP7_75t_R g189 ( .A(n_28), .Y(n_189) );
INVxp67_ASAP7_75t_L g190 ( .A(n_151), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_69), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_79), .Y(n_192) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_130), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_63), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_135), .Y(n_195) );
CKINVDCx5p33_ASAP7_75t_R g196 ( .A(n_118), .Y(n_196) );
BUFx3_ASAP7_75t_L g197 ( .A(n_153), .Y(n_197) );
CKINVDCx16_ASAP7_75t_R g198 ( .A(n_145), .Y(n_198) );
CKINVDCx20_ASAP7_75t_R g199 ( .A(n_75), .Y(n_199) );
CKINVDCx5p33_ASAP7_75t_R g200 ( .A(n_116), .Y(n_200) );
CKINVDCx5p33_ASAP7_75t_R g201 ( .A(n_136), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_150), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_80), .Y(n_203) );
CKINVDCx16_ASAP7_75t_R g204 ( .A(n_2), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_146), .Y(n_205) );
CKINVDCx5p33_ASAP7_75t_R g206 ( .A(n_166), .Y(n_206) );
CKINVDCx5p33_ASAP7_75t_R g207 ( .A(n_161), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_163), .B(n_77), .Y(n_208) );
CKINVDCx5p33_ASAP7_75t_R g209 ( .A(n_123), .Y(n_209) );
CKINVDCx5p33_ASAP7_75t_R g210 ( .A(n_133), .Y(n_210) );
BUFx10_ASAP7_75t_L g211 ( .A(n_155), .Y(n_211) );
CKINVDCx20_ASAP7_75t_R g212 ( .A(n_10), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_103), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_149), .Y(n_214) );
CKINVDCx5p33_ASAP7_75t_R g215 ( .A(n_15), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_42), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_139), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_34), .Y(n_218) );
CKINVDCx5p33_ASAP7_75t_R g219 ( .A(n_97), .Y(n_219) );
CKINVDCx5p33_ASAP7_75t_R g220 ( .A(n_49), .Y(n_220) );
INVx1_ASAP7_75t_SL g221 ( .A(n_124), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_100), .Y(n_222) );
INVxp67_ASAP7_75t_SL g223 ( .A(n_131), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_144), .Y(n_224) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_8), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_33), .Y(n_226) );
INVx2_ASAP7_75t_L g227 ( .A(n_51), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g228 ( .A(n_121), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_115), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_119), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_92), .Y(n_231) );
INVx1_ASAP7_75t_SL g232 ( .A(n_59), .Y(n_232) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_140), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_78), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_95), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_35), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_62), .Y(n_237) );
CKINVDCx5p33_ASAP7_75t_R g238 ( .A(n_159), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_7), .Y(n_239) );
INVx1_ASAP7_75t_SL g240 ( .A(n_110), .Y(n_240) );
CKINVDCx5p33_ASAP7_75t_R g241 ( .A(n_76), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_6), .Y(n_242) );
BUFx2_ASAP7_75t_L g243 ( .A(n_65), .Y(n_243) );
BUFx2_ASAP7_75t_SL g244 ( .A(n_46), .Y(n_244) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_91), .Y(n_245) );
NOR2xp67_ASAP7_75t_L g246 ( .A(n_52), .B(n_23), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_141), .Y(n_247) );
INVxp67_ASAP7_75t_SL g248 ( .A(n_14), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_154), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_142), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_167), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_129), .Y(n_252) );
CKINVDCx20_ASAP7_75t_R g253 ( .A(n_37), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_101), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_36), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_43), .Y(n_256) );
INVxp33_ASAP7_75t_SL g257 ( .A(n_125), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_147), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_39), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_81), .B(n_160), .Y(n_260) );
INVx1_ASAP7_75t_SL g261 ( .A(n_128), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_105), .Y(n_262) );
BUFx10_ASAP7_75t_L g263 ( .A(n_152), .Y(n_263) );
CKINVDCx16_ASAP7_75t_R g264 ( .A(n_88), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_134), .B(n_157), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_122), .Y(n_266) );
CKINVDCx20_ASAP7_75t_R g267 ( .A(n_44), .Y(n_267) );
INVx2_ASAP7_75t_L g268 ( .A(n_45), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_158), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_114), .Y(n_270) );
INVxp67_ASAP7_75t_L g271 ( .A(n_93), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_117), .Y(n_272) );
OAI22xp5_ASAP7_75t_SL g273 ( .A1(n_204), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_177), .B(n_0), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_243), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_199), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_178), .B(n_3), .Y(n_277) );
NOR2x1_ASAP7_75t_L g278 ( .A(n_170), .B(n_11), .Y(n_278) );
OAI22xp5_ASAP7_75t_SL g279 ( .A1(n_186), .A2(n_3), .B1(n_4), .B2(n_5), .Y(n_279) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_239), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_202), .Y(n_281) );
NAND2xp33_ASAP7_75t_L g282 ( .A(n_172), .B(n_165), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_222), .Y(n_283) );
AND2x4_ASAP7_75t_L g284 ( .A(n_242), .B(n_4), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_227), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_234), .B(n_5), .Y(n_286) );
AND2x4_ASAP7_75t_L g287 ( .A(n_237), .B(n_6), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_211), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_252), .Y(n_289) );
AND2x2_ASAP7_75t_SL g290 ( .A(n_175), .B(n_8), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_211), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_263), .Y(n_292) );
BUFx6f_ASAP7_75t_L g293 ( .A(n_225), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_268), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_281), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_275), .B(n_198), .Y(n_296) );
INVx3_ASAP7_75t_L g297 ( .A(n_284), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_283), .Y(n_298) );
NOR2xp33_ASAP7_75t_SL g299 ( .A(n_290), .B(n_264), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_285), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g301 ( .A(n_288), .B(n_190), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_291), .B(n_189), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_292), .B(n_168), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_287), .Y(n_304) );
AND2x6_ASAP7_75t_L g305 ( .A(n_287), .B(n_260), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_289), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g307 ( .A(n_280), .B(n_294), .Y(n_307) );
CKINVDCx20_ASAP7_75t_R g308 ( .A(n_276), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_284), .Y(n_309) );
AOI22xp5_ASAP7_75t_L g310 ( .A1(n_299), .A2(n_274), .B1(n_282), .B2(n_273), .Y(n_310) );
INVx2_ASAP7_75t_SL g311 ( .A(n_297), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_296), .B(n_263), .Y(n_312) );
OR2x6_ASAP7_75t_L g313 ( .A(n_309), .B(n_279), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g314 ( .A1(n_304), .A2(n_228), .B1(n_253), .B2(n_212), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_295), .Y(n_315) );
AOI21xp5_ASAP7_75t_L g316 ( .A1(n_302), .A2(n_286), .B(n_277), .Y(n_316) );
OAI22xp5_ASAP7_75t_L g317 ( .A1(n_307), .A2(n_267), .B1(n_257), .B2(n_271), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_305), .B(n_179), .Y(n_318) );
INVx8_ASAP7_75t_L g319 ( .A(n_305), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_298), .Y(n_320) );
AND2x4_ASAP7_75t_L g321 ( .A(n_303), .B(n_278), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_305), .B(n_301), .Y(n_322) );
INVx2_ASAP7_75t_SL g323 ( .A(n_300), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g324 ( .A1(n_306), .A2(n_225), .B1(n_244), .B2(n_169), .Y(n_324) );
AOI21xp5_ASAP7_75t_L g325 ( .A1(n_316), .A2(n_265), .B(n_248), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_312), .B(n_221), .Y(n_326) );
NAND2x1p5_ASAP7_75t_L g327 ( .A(n_323), .B(n_225), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g328 ( .A1(n_321), .A2(n_173), .B1(n_176), .B2(n_171), .Y(n_328) );
INVxp67_ASAP7_75t_L g329 ( .A(n_314), .Y(n_329) );
BUFx2_ASAP7_75t_L g330 ( .A(n_319), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_322), .B(n_232), .Y(n_331) );
A2O1A1Ixp33_ASAP7_75t_L g332 ( .A1(n_321), .A2(n_180), .B(n_182), .C(n_181), .Y(n_332) );
OR2x6_ASAP7_75t_SL g333 ( .A(n_317), .B(n_308), .Y(n_333) );
OR2x6_ASAP7_75t_SL g334 ( .A(n_319), .B(n_185), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_310), .B(n_261), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_313), .B(n_261), .Y(n_336) );
O2A1O1Ixp33_ASAP7_75t_L g337 ( .A1(n_313), .A2(n_183), .B(n_187), .C(n_184), .Y(n_337) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_320), .B(n_223), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_311), .B(n_240), .Y(n_339) );
O2A1O1Ixp5_ASAP7_75t_L g340 ( .A1(n_318), .A2(n_188), .B(n_192), .C(n_191), .Y(n_340) );
INVx6_ASAP7_75t_L g341 ( .A(n_336), .Y(n_341) );
OAI21x1_ASAP7_75t_SL g342 ( .A1(n_325), .A2(n_324), .B(n_195), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_338), .Y(n_343) );
OAI22xp5_ASAP7_75t_L g344 ( .A1(n_328), .A2(n_315), .B1(n_193), .B2(n_200), .Y(n_344) );
AOI21x1_ASAP7_75t_L g345 ( .A1(n_331), .A2(n_246), .B(n_174), .Y(n_345) );
CKINVDCx5p33_ASAP7_75t_R g346 ( .A(n_334), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_335), .B(n_194), .Y(n_347) );
OAI21x1_ASAP7_75t_L g348 ( .A1(n_327), .A2(n_205), .B(n_203), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_326), .Y(n_349) );
INVx2_ASAP7_75t_SL g350 ( .A(n_330), .Y(n_350) );
A2O1A1Ixp33_ASAP7_75t_L g351 ( .A1(n_340), .A2(n_249), .B(n_272), .C(n_270), .Y(n_351) );
INVx3_ASAP7_75t_L g352 ( .A(n_327), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_332), .Y(n_353) );
AO21x1_ASAP7_75t_L g354 ( .A1(n_337), .A2(n_214), .B(n_213), .Y(n_354) );
AO31x2_ASAP7_75t_L g355 ( .A1(n_339), .A2(n_247), .A3(n_269), .B(n_266), .Y(n_355) );
OA21x2_ASAP7_75t_L g356 ( .A1(n_329), .A2(n_217), .B(n_216), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_333), .B(n_218), .Y(n_357) );
INVx3_ASAP7_75t_SL g358 ( .A(n_336), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_327), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_329), .B(n_196), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_335), .B(n_226), .Y(n_361) );
AO31x2_ASAP7_75t_L g362 ( .A1(n_351), .A2(n_250), .A3(n_262), .B(n_259), .Y(n_362) );
INVx3_ASAP7_75t_L g363 ( .A(n_352), .Y(n_363) );
OAI21x1_ASAP7_75t_L g364 ( .A1(n_359), .A2(n_230), .B(n_229), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_343), .Y(n_365) );
AND2x4_ASAP7_75t_L g366 ( .A(n_349), .B(n_235), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_353), .B(n_236), .Y(n_367) );
INVx2_ASAP7_75t_L g368 ( .A(n_348), .Y(n_368) );
INVx2_ASAP7_75t_SL g369 ( .A(n_350), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_342), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_347), .B(n_251), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_361), .B(n_254), .Y(n_372) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_341), .Y(n_373) );
OAI21x1_ASAP7_75t_L g374 ( .A1(n_345), .A2(n_256), .B(n_255), .Y(n_374) );
OA21x2_ASAP7_75t_L g375 ( .A1(n_354), .A2(n_258), .B(n_208), .Y(n_375) );
OA21x2_ASAP7_75t_L g376 ( .A1(n_357), .A2(n_206), .B(n_201), .Y(n_376) );
NOR2xp33_ASAP7_75t_SL g377 ( .A(n_346), .B(n_197), .Y(n_377) );
OAI21x1_ASAP7_75t_L g378 ( .A1(n_356), .A2(n_12), .B(n_13), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_356), .Y(n_379) );
OA21x2_ASAP7_75t_L g380 ( .A1(n_360), .A2(n_209), .B(n_207), .Y(n_380) );
INVx2_ASAP7_75t_L g381 ( .A(n_355), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_355), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_344), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_353), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_358), .B(n_210), .Y(n_385) );
BUFx12f_ASAP7_75t_L g386 ( .A(n_346), .Y(n_386) );
AND2x4_ASAP7_75t_L g387 ( .A(n_352), .B(n_17), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_343), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_353), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_353), .Y(n_390) );
OAI21xp5_ASAP7_75t_L g391 ( .A1(n_353), .A2(n_219), .B(n_215), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_358), .B(n_220), .Y(n_392) );
OAI21x1_ASAP7_75t_L g393 ( .A1(n_359), .A2(n_19), .B(n_21), .Y(n_393) );
OAI21x1_ASAP7_75t_L g394 ( .A1(n_359), .A2(n_22), .B(n_24), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_343), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_384), .Y(n_396) );
INVx3_ASAP7_75t_L g397 ( .A(n_387), .Y(n_397) );
INVx4_ASAP7_75t_L g398 ( .A(n_387), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_389), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_389), .Y(n_400) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_388), .Y(n_401) );
BUFx2_ASAP7_75t_L g402 ( .A(n_369), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_395), .B(n_224), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_381), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_382), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_366), .B(n_293), .Y(n_406) );
AO21x2_ASAP7_75t_L g407 ( .A1(n_379), .A2(n_293), .B(n_231), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_390), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_390), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_367), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_363), .Y(n_411) );
HB1xp67_ASAP7_75t_L g412 ( .A(n_373), .Y(n_412) );
BUFx2_ASAP7_75t_L g413 ( .A(n_363), .Y(n_413) );
BUFx2_ASAP7_75t_L g414 ( .A(n_385), .Y(n_414) );
AND2x4_ASAP7_75t_L g415 ( .A(n_383), .B(n_25), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_370), .Y(n_416) );
BUFx2_ASAP7_75t_L g417 ( .A(n_376), .Y(n_417) );
AOI21xp5_ASAP7_75t_L g418 ( .A1(n_368), .A2(n_245), .B(n_241), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_372), .B(n_233), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_378), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_383), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_372), .B(n_371), .Y(n_422) );
OR2x6_ASAP7_75t_L g423 ( .A(n_392), .B(n_26), .Y(n_423) );
OR2x6_ASAP7_75t_L g424 ( .A(n_391), .B(n_27), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_374), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_364), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_375), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_380), .B(n_238), .Y(n_428) );
AND2x4_ASAP7_75t_L g429 ( .A(n_362), .B(n_29), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_362), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_362), .Y(n_431) );
OA21x2_ASAP7_75t_L g432 ( .A1(n_393), .A2(n_30), .B(n_31), .Y(n_432) );
AND2x4_ASAP7_75t_L g433 ( .A(n_394), .B(n_32), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_377), .B(n_38), .Y(n_434) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_377), .B(n_40), .Y(n_435) );
OR2x6_ASAP7_75t_L g436 ( .A(n_386), .B(n_41), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_365), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_365), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_365), .B(n_162), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_365), .Y(n_440) );
HB1xp67_ASAP7_75t_L g441 ( .A(n_365), .Y(n_441) );
INVx1_ASAP7_75t_SL g442 ( .A(n_413), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_401), .B(n_47), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_440), .B(n_48), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_441), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_437), .Y(n_446) );
BUFx3_ASAP7_75t_L g447 ( .A(n_402), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_421), .B(n_53), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_421), .B(n_54), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_404), .Y(n_450) );
BUFx6f_ASAP7_75t_L g451 ( .A(n_398), .Y(n_451) );
BUFx2_ASAP7_75t_L g452 ( .A(n_398), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_438), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_396), .Y(n_454) );
INVx3_ASAP7_75t_L g455 ( .A(n_397), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_408), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_414), .B(n_55), .Y(n_457) );
AND2x4_ASAP7_75t_L g458 ( .A(n_397), .B(n_56), .Y(n_458) );
INVx3_ASAP7_75t_L g459 ( .A(n_415), .Y(n_459) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_406), .Y(n_460) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_405), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_403), .B(n_57), .Y(n_462) );
INVx5_ASAP7_75t_SL g463 ( .A(n_436), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_412), .B(n_58), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_422), .A2(n_60), .B1(n_61), .B2(n_64), .Y(n_465) );
BUFx2_ASAP7_75t_L g466 ( .A(n_423), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_399), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_400), .B(n_66), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_400), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_410), .B(n_67), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_409), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_411), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_423), .B(n_70), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_416), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_428), .B(n_72), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_416), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_430), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_431), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_425), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_427), .Y(n_480) );
INVxp67_ASAP7_75t_SL g481 ( .A(n_415), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_434), .B(n_73), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_426), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_439), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_429), .Y(n_485) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_429), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_417), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_424), .Y(n_488) );
BUFx3_ASAP7_75t_L g489 ( .A(n_424), .Y(n_489) );
INVx3_ASAP7_75t_L g490 ( .A(n_433), .Y(n_490) );
INVxp67_ASAP7_75t_L g491 ( .A(n_407), .Y(n_491) );
INVx3_ASAP7_75t_L g492 ( .A(n_433), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_435), .B(n_74), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_467), .Y(n_494) );
INVx1_ASAP7_75t_L g495 ( .A(n_467), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_445), .B(n_420), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_446), .B(n_419), .Y(n_497) );
BUFx2_ASAP7_75t_L g498 ( .A(n_447), .Y(n_498) );
BUFx6f_ASAP7_75t_L g499 ( .A(n_451), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_471), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_453), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_454), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_456), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_442), .B(n_418), .Y(n_504) );
INVxp67_ASAP7_75t_L g505 ( .A(n_447), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_461), .B(n_432), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_469), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_469), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_472), .B(n_83), .Y(n_509) );
BUFx2_ASAP7_75t_L g510 ( .A(n_452), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_474), .B(n_84), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_488), .B(n_85), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_489), .B(n_86), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_476), .B(n_87), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_477), .Y(n_515) );
HB1xp67_ASAP7_75t_L g516 ( .A(n_466), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_460), .B(n_481), .Y(n_517) );
AND2x4_ASAP7_75t_L g518 ( .A(n_481), .B(n_89), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_450), .Y(n_519) );
OR2x2_ASAP7_75t_L g520 ( .A(n_450), .B(n_90), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_480), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_478), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_479), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_483), .Y(n_524) );
INVxp67_ASAP7_75t_SL g525 ( .A(n_510), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_498), .B(n_486), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_500), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_515), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_496), .B(n_459), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_517), .B(n_490), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_502), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_522), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_516), .B(n_492), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_522), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_523), .B(n_487), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_505), .B(n_492), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g537 ( .A(n_499), .B(n_463), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_503), .B(n_501), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_521), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_523), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_494), .B(n_485), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_508), .B(n_455), .Y(n_542) );
NOR4xp25_ASAP7_75t_L g543 ( .A(n_497), .B(n_473), .C(n_468), .D(n_457), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_507), .B(n_455), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_538), .B(n_524), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_530), .B(n_495), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_532), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_533), .B(n_519), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_525), .B(n_524), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_526), .B(n_506), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_529), .B(n_504), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_536), .B(n_513), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_527), .B(n_491), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_543), .B(n_518), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_534), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_539), .Y(n_556) );
OAI21xp5_ASAP7_75t_L g557 ( .A1(n_554), .A2(n_543), .B(n_537), .Y(n_557) );
INVx2_ASAP7_75t_SL g558 ( .A(n_546), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_549), .B(n_528), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_551), .A2(n_518), .B1(n_475), .B2(n_512), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_545), .B(n_531), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_552), .A2(n_542), .B1(n_535), .B2(n_540), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_547), .Y(n_563) );
AOI22xp5_ASAP7_75t_L g564 ( .A1(n_557), .A2(n_550), .B1(n_548), .B2(n_553), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_558), .A2(n_556), .B1(n_555), .B2(n_541), .Y(n_565) );
OAI22xp33_ASAP7_75t_SL g566 ( .A1(n_559), .A2(n_514), .B1(n_511), .B2(n_520), .Y(n_566) );
NAND3xp33_ASAP7_75t_L g567 ( .A(n_563), .B(n_465), .C(n_544), .Y(n_567) );
OAI21xp5_ASAP7_75t_L g568 ( .A1(n_560), .A2(n_458), .B(n_482), .Y(n_568) );
AOI32xp33_ASAP7_75t_L g569 ( .A1(n_561), .A2(n_464), .A3(n_443), .B1(n_444), .B2(n_509), .Y(n_569) );
AOI322xp5_ASAP7_75t_L g570 ( .A1(n_562), .A2(n_448), .A3(n_449), .B1(n_470), .B2(n_462), .C1(n_484), .C2(n_493), .Y(n_570) );
NAND4xp25_ASAP7_75t_L g571 ( .A(n_564), .B(n_570), .C(n_569), .D(n_568), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_565), .Y(n_572) );
NAND4xp25_ASAP7_75t_L g573 ( .A(n_571), .B(n_567), .C(n_566), .D(n_98), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_572), .Y(n_574) );
INVx1_ASAP7_75t_SL g575 ( .A(n_574), .Y(n_575) );
AND2x4_ASAP7_75t_L g576 ( .A(n_573), .B(n_94), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_575), .Y(n_577) );
INVx3_ASAP7_75t_L g578 ( .A(n_576), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_577), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_579), .A2(n_578), .B1(n_99), .B2(n_102), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_580), .Y(n_581) );
NOR2x1_ASAP7_75t_R g582 ( .A(n_581), .B(n_104), .Y(n_582) );
AO21x2_ASAP7_75t_L g583 ( .A1(n_582), .A2(n_106), .B(n_107), .Y(n_583) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_583), .A2(n_108), .B1(n_109), .B2(n_111), .Y(n_584) );
endmodule