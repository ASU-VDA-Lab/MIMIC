module fake_jpeg_1581_n_219 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_219);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_219;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_140;
wire n_82;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_9),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_16),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_26),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_27),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_35),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_23),
.Y(n_65)
);

BUFx16f_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_7),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_30),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_13),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_4),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_12),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_11),
.Y(n_73)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_74),
.Y(n_76)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_0),
.Y(n_77)
);

NAND3xp33_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_63),
.C(n_70),
.Y(n_86)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_66),
.Y(n_78)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_61),
.Y(n_82)
);

NAND2xp33_ASAP7_75t_SL g96 ( 
.A(n_82),
.B(n_83),
.Y(n_96)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx13_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_84),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_71),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_86),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_62),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_87),
.B(n_89),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_79),
.B(n_73),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_76),
.A2(n_72),
.B1(n_55),
.B2(n_73),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_92),
.A2(n_53),
.B1(n_58),
.B2(n_57),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_81),
.B(n_51),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_65),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_78),
.A2(n_68),
.B1(n_72),
.B2(n_55),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_94),
.A2(n_74),
.B1(n_68),
.B2(n_63),
.Y(n_104)
);

O2A1O1Ixp33_ASAP7_75t_SL g98 ( 
.A1(n_96),
.A2(n_57),
.B(n_58),
.C(n_51),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_98),
.A2(n_105),
.B1(n_116),
.B2(n_90),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_61),
.C(n_75),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_100),
.B(n_102),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_93),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_101),
.B(n_107),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_52),
.C(n_67),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_104),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_52),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_109),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_95),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_67),
.Y(n_109)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_113),
.B(n_90),
.Y(n_121)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_114),
.Y(n_128)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

OAI22xp33_ASAP7_75t_L g116 ( 
.A1(n_92),
.A2(n_60),
.B1(n_59),
.B2(n_56),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_64),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_131),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_112),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_120),
.B(n_122),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_121),
.B(n_130),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_103),
.B(n_0),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_99),
.B(n_1),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_123),
.B(n_2),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_124),
.A2(n_125),
.B(n_119),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_95),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_53),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_84),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_134),
.B(n_84),
.C(n_58),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_110),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_18),
.Y(n_152)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_136),
.Y(n_144)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_137),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_117),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_146),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_124),
.A2(n_98),
.B1(n_108),
.B2(n_88),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_140),
.A2(n_148),
.B1(n_6),
.B2(n_7),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_37),
.C(n_36),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_143),
.A2(n_160),
.B(n_3),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_126),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_1),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_147),
.B(n_155),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_134),
.A2(n_57),
.B1(n_19),
.B2(n_22),
.Y(n_148)
);

AND2x6_ASAP7_75t_L g150 ( 
.A(n_118),
.B(n_132),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_151),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_127),
.Y(n_151)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_152),
.Y(n_162)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_153),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_125),
.A2(n_17),
.B1(n_46),
.B2(n_45),
.Y(n_154)
);

BUFx8_ASAP7_75t_L g173 ( 
.A(n_154),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_128),
.B(n_2),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_156),
.B(n_159),
.Y(n_175)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_129),
.Y(n_157)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_157),
.Y(n_165)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_133),
.Y(n_158)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

AO22x1_ASAP7_75t_L g159 ( 
.A1(n_126),
.A2(n_50),
.B1(n_44),
.B2(n_41),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_117),
.A2(n_3),
.B(n_4),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_117),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_5),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_163),
.A2(n_177),
.B(n_179),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_145),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_170),
.Y(n_187)
);

MAJx2_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_40),
.C(n_38),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_169),
.B(n_180),
.Y(n_186)
);

NOR2xp67_ASAP7_75t_R g172 ( 
.A(n_139),
.B(n_5),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_172),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_179),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_176),
.A2(n_149),
.B1(n_151),
.B2(n_153),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_160),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_178),
.B(n_141),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_142),
.B(n_33),
.C(n_32),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_148),
.B(n_31),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_144),
.Y(n_181)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_181),
.Y(n_184)
);

OA21x2_ASAP7_75t_SL g198 ( 
.A1(n_182),
.A2(n_180),
.B(n_8),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_171),
.A2(n_140),
.B(n_154),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g195 ( 
.A1(n_185),
.A2(n_173),
.B(n_176),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_188),
.A2(n_189),
.B1(n_192),
.B2(n_174),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_175),
.A2(n_159),
.B1(n_8),
.B2(n_9),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_165),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_191),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_167),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_184),
.A2(n_168),
.B1(n_173),
.B2(n_164),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_194),
.A2(n_196),
.B1(n_202),
.B2(n_186),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_195),
.B(n_197),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_187),
.A2(n_173),
.B1(n_169),
.B2(n_162),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_198),
.B(n_199),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_193),
.B(n_6),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_183),
.B(n_28),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_201),
.B(n_183),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_193),
.A2(n_24),
.B(n_11),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_200),
.Y(n_203)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_203),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_194),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_204),
.B(n_206),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_207),
.B(n_186),
.C(n_196),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_211),
.B(n_201),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_212),
.B(n_213),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_209),
.B(n_205),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_214),
.A2(n_208),
.B(n_210),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_215),
.B(n_204),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_10),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_217),
.B(n_14),
.C(n_12),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_10),
.Y(n_219)
);


endmodule