module fake_jpeg_16995_n_184 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_184);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_184;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx2_ASAP7_75t_SL g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_5),
.B(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_34),
.Y(n_52)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_30),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_35),
.B(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

CKINVDCx9p33_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_38),
.B(n_49),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_23),
.B(n_1),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_17),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_47),
.A2(n_20),
.B1(n_24),
.B2(n_28),
.Y(n_63)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_48),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_26),
.B(n_1),
.Y(n_49)
);

BUFx8_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_50),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_26),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_55),
.B(n_56),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_15),
.Y(n_56)
);

OA22x2_ASAP7_75t_SL g57 ( 
.A1(n_42),
.A2(n_43),
.B1(n_40),
.B2(n_41),
.Y(n_57)
);

AO22x1_ASAP7_75t_SL g99 ( 
.A1(n_57),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_33),
.B(n_15),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_67),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_46),
.A2(n_18),
.B1(n_31),
.B2(n_21),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_60),
.A2(n_68),
.B1(n_69),
.B2(n_61),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_63),
.A2(n_25),
.B1(n_32),
.B2(n_11),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_36),
.B(n_21),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_70),
.Y(n_83)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_48),
.A2(n_16),
.B1(n_31),
.B2(n_22),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_34),
.A2(n_16),
.B1(n_22),
.B2(n_27),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_36),
.B(n_18),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_39),
.B(n_27),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_72),
.B(n_76),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_45),
.B(n_28),
.Y(n_76)
);

AND2x6_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_2),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_77),
.A2(n_81),
.B1(n_91),
.B2(n_92),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_78),
.Y(n_116)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_44),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_80),
.B(n_86),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_62),
.A2(n_24),
.B1(n_20),
.B2(n_25),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_44),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_98),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_64),
.B(n_3),
.Y(n_86)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_87),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_54),
.B(n_32),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_90),
.Y(n_102)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_57),
.A2(n_25),
.B1(n_6),
.B2(n_7),
.Y(n_91)
);

AND2x6_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_4),
.Y(n_92)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_94),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_95),
.B(n_97),
.Y(n_114)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_101),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_66),
.A2(n_32),
.B1(n_8),
.B2(n_11),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_4),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_99),
.B(n_100),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_52),
.B(n_8),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_66),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_80),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_103),
.B(n_110),
.Y(n_124)
);

NOR2x1_ASAP7_75t_L g105 ( 
.A(n_99),
.B(n_50),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_105),
.B(n_113),
.Y(n_138)
);

NAND3xp33_ASAP7_75t_L g110 ( 
.A(n_84),
.B(n_71),
.C(n_13),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_93),
.B(n_13),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_73),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_119),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_93),
.B(n_12),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_118),
.B(n_81),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_51),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_82),
.B(n_58),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_120),
.A2(n_90),
.B1(n_87),
.B2(n_94),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_79),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_121),
.B(n_67),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_116),
.A2(n_83),
.B1(n_96),
.B2(n_77),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_122),
.A2(n_126),
.B1(n_112),
.B2(n_114),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_123),
.B(n_127),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_116),
.A2(n_111),
.B1(n_105),
.B2(n_91),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_125),
.A2(n_131),
.B1(n_120),
.B2(n_102),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_111),
.A2(n_78),
.B1(n_92),
.B2(n_99),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_104),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_104),
.Y(n_145)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_129),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_105),
.A2(n_85),
.B1(n_98),
.B2(n_86),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_134),
.Y(n_148)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_133),
.Y(n_142)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_115),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_107),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_107),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_117),
.B(n_100),
.C(n_80),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_137),
.C(n_109),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_58),
.C(n_51),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g139 ( 
.A(n_130),
.B(n_103),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_139),
.B(n_144),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_140),
.B(n_145),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_122),
.A2(n_112),
.B1(n_119),
.B2(n_114),
.Y(n_141)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_141),
.Y(n_153)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_143),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_130),
.B(n_106),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_147),
.B(n_136),
.C(n_128),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_149),
.B(n_151),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_120),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_156),
.C(n_159),
.Y(n_166)
);

INVx2_ASAP7_75t_SL g155 ( 
.A(n_143),
.Y(n_155)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_155),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_147),
.B(n_126),
.C(n_134),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_145),
.B(n_151),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_144),
.B(n_149),
.C(n_140),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_161),
.Y(n_163)
);

AOI321xp33_ASAP7_75t_L g164 ( 
.A1(n_159),
.A2(n_139),
.A3(n_141),
.B1(n_148),
.B2(n_138),
.C(n_109),
.Y(n_164)
);

AOI21xp33_ASAP7_75t_L g173 ( 
.A1(n_164),
.A2(n_167),
.B(n_133),
.Y(n_173)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_155),
.Y(n_165)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_165),
.Y(n_171)
);

AOI322xp5_ASAP7_75t_L g167 ( 
.A1(n_158),
.A2(n_153),
.A3(n_156),
.B1(n_161),
.B2(n_154),
.C1(n_157),
.C2(n_138),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_160),
.A2(n_142),
.B1(n_150),
.B2(n_146),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_168),
.A2(n_152),
.B1(n_118),
.B2(n_139),
.Y(n_172)
);

NOR3xp33_ASAP7_75t_L g169 ( 
.A(n_164),
.B(n_124),
.C(n_113),
.Y(n_169)
);

AO21x1_ASAP7_75t_L g174 ( 
.A1(n_169),
.A2(n_173),
.B(n_163),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_162),
.A2(n_142),
.B(n_154),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_170),
.A2(n_168),
.B(n_129),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_172),
.A2(n_166),
.B1(n_135),
.B2(n_115),
.Y(n_177)
);

OAI21x1_ASAP7_75t_L g180 ( 
.A1(n_174),
.A2(n_175),
.B(n_12),
.Y(n_180)
);

XNOR2x1_ASAP7_75t_L g175 ( 
.A(n_170),
.B(n_166),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_176),
.B(n_177),
.C(n_53),
.Y(n_179)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_177),
.B(n_171),
.Y(n_178)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_178),
.Y(n_182)
);

MAJx2_ASAP7_75t_L g181 ( 
.A(n_179),
.B(n_180),
.C(n_53),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_181),
.B(n_182),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_183),
.B(n_89),
.C(n_50),
.Y(n_184)
);


endmodule