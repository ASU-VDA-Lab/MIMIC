module fake_jpeg_2432_n_556 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_556);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_556;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_18),
.B(n_4),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_8),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_SL g39 ( 
.A(n_13),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_11),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_12),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_55),
.Y(n_128)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_56),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_29),
.B(n_18),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_57),
.B(n_63),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_58),
.Y(n_119)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_23),
.Y(n_59)
);

INVx3_ASAP7_75t_SL g160 ( 
.A(n_59),
.Y(n_160)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_60),
.Y(n_117)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_62),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_29),
.B(n_18),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_35),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_64),
.B(n_69),
.Y(n_147)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_65),
.Y(n_145)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_49),
.Y(n_66)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_66),
.Y(n_126)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_67),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_35),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_70),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_35),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_71),
.B(n_75),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

INVxp67_ASAP7_75t_SL g74 ( 
.A(n_30),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_74),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_48),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_19),
.B(n_0),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_76),
.B(n_39),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_19),
.B(n_0),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_77),
.B(n_81),
.Y(n_120)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_78),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_37),
.B(n_0),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_80),
.B(n_2),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_21),
.B(n_1),
.Y(n_81)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_32),
.Y(n_82)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_82),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_48),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_83),
.B(n_84),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_48),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_21),
.Y(n_85)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_85),
.Y(n_131)
);

INVx4_ASAP7_75t_SL g86 ( 
.A(n_32),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g163 ( 
.A(n_86),
.B(n_106),
.Y(n_163)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_87),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_39),
.B(n_1),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_88),
.B(n_94),
.Y(n_143)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_34),
.Y(n_89)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_89),
.Y(n_137)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_90),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_33),
.Y(n_92)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_92),
.Y(n_164)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_34),
.Y(n_93)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_93),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_25),
.Y(n_94)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_30),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_95),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_52),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_96),
.B(n_102),
.Y(n_108)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_97),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_25),
.Y(n_98)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_22),
.Y(n_99)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_99),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_24),
.Y(n_100)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_100),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g101 ( 
.A(n_33),
.Y(n_101)
);

AOI21xp33_ASAP7_75t_SL g159 ( 
.A1(n_101),
.A2(n_33),
.B(n_52),
.Y(n_159)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_32),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_27),
.B(n_1),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_103),
.B(n_28),
.Y(n_146)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_27),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_105),
.Y(n_127)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_44),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_52),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_92),
.A2(n_39),
.B1(n_49),
.B2(n_45),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_107),
.A2(n_129),
.B1(n_135),
.B2(n_144),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_110),
.B(n_122),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_80),
.B(n_31),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_123),
.B(n_130),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_97),
.A2(n_44),
.B1(n_47),
.B2(n_31),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_124),
.A2(n_78),
.B(n_26),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_92),
.A2(n_86),
.B1(n_106),
.B2(n_96),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_88),
.B(n_51),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_64),
.A2(n_45),
.B1(n_41),
.B2(n_51),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_61),
.B(n_67),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_150),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_69),
.A2(n_45),
.B1(n_43),
.B2(n_46),
.Y(n_144)
);

OAI21xp33_ASAP7_75t_L g203 ( 
.A1(n_146),
.A2(n_159),
.B(n_2),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_71),
.A2(n_28),
.B1(n_36),
.B2(n_50),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_148),
.A2(n_124),
.B1(n_142),
.B2(n_138),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_89),
.B(n_46),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_75),
.A2(n_45),
.B1(n_43),
.B2(n_41),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_151),
.A2(n_155),
.B1(n_158),
.B2(n_55),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_84),
.A2(n_47),
.B1(n_44),
.B2(n_50),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_153),
.A2(n_54),
.B1(n_98),
.B2(n_73),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_66),
.A2(n_45),
.B1(n_40),
.B2(n_36),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_90),
.A2(n_40),
.B1(n_47),
.B2(n_44),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_85),
.B(n_47),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_162),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_87),
.B(n_2),
.Y(n_162)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_111),
.Y(n_167)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_167),
.Y(n_268)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_119),
.Y(n_168)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_168),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_123),
.A2(n_93),
.B1(n_105),
.B2(n_59),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_170),
.A2(n_177),
.B1(n_216),
.B2(n_156),
.Y(n_253)
);

INVx4_ASAP7_75t_SL g171 ( 
.A(n_163),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_171),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_109),
.B(n_104),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_172),
.B(n_173),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_120),
.B(n_99),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_56),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_174),
.B(n_191),
.Y(n_233)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_111),
.Y(n_175)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_175),
.Y(n_232)
);

A2O1A1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_130),
.A2(n_65),
.B(n_101),
.C(n_91),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_176),
.B(n_181),
.Y(n_256)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_114),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_180),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_110),
.B(n_79),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_122),
.B(n_102),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_183),
.B(n_211),
.Y(n_231)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_164),
.Y(n_184)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_184),
.Y(n_252)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_136),
.Y(n_185)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_185),
.Y(n_276)
);

BUFx2_ASAP7_75t_L g186 ( 
.A(n_164),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_186),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_150),
.A2(n_62),
.B1(n_68),
.B2(n_72),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_187),
.A2(n_217),
.B1(n_160),
.B2(n_116),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_163),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_188),
.B(n_203),
.Y(n_248)
);

INVx4_ASAP7_75t_SL g189 ( 
.A(n_117),
.Y(n_189)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_189),
.Y(n_255)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_112),
.Y(n_190)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_190),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_125),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_131),
.B(n_58),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_192),
.B(n_193),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_131),
.B(n_58),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_132),
.B(n_95),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_194),
.B(n_196),
.Y(n_254)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_119),
.Y(n_195)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_195),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_132),
.B(n_55),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_197),
.Y(n_242)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_112),
.Y(n_198)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_198),
.Y(n_266)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_115),
.Y(n_199)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_199),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_200),
.Y(n_257)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_136),
.Y(n_201)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_201),
.Y(n_271)
);

OAI32xp33_ASAP7_75t_L g202 ( 
.A1(n_140),
.A2(n_100),
.A3(n_70),
.B1(n_82),
.B2(n_60),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_202),
.A2(n_128),
.B(n_154),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_147),
.A2(n_100),
.B1(n_70),
.B2(n_53),
.Y(n_204)
);

OAI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_204),
.A2(n_20),
.B1(n_128),
.B2(n_117),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_113),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_205),
.B(n_212),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_108),
.B(n_4),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_206),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_127),
.A2(n_53),
.B1(n_38),
.B2(n_26),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_207),
.A2(n_7),
.B(n_9),
.Y(n_263)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_117),
.Y(n_208)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_208),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_108),
.A2(n_38),
.B1(n_26),
.B2(n_20),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_209),
.A2(n_221),
.B1(n_223),
.B2(n_145),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_126),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_210),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_142),
.B(n_4),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_108),
.B(n_6),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_157),
.B(n_6),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_213),
.B(n_219),
.Y(n_246)
);

OR2x2_ASAP7_75t_SL g214 ( 
.A(n_134),
.B(n_53),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_214),
.B(n_225),
.C(n_152),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_127),
.A2(n_138),
.B1(n_137),
.B2(n_118),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_127),
.Y(n_218)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_218),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_137),
.B(n_6),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_114),
.Y(n_220)
);

INVx6_ASAP7_75t_L g238 ( 
.A(n_220),
.Y(n_238)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_115),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_165),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_222),
.B(n_224),
.Y(n_264)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_116),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_157),
.B(n_6),
.Y(n_224)
);

AND2x2_ASAP7_75t_SL g225 ( 
.A(n_165),
.B(n_38),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_227),
.A2(n_234),
.B1(n_235),
.B2(n_237),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_230),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_179),
.A2(n_139),
.B1(n_118),
.B2(n_121),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_179),
.A2(n_139),
.B1(n_160),
.B2(n_121),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_187),
.A2(n_160),
.B1(n_134),
.B2(n_126),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_171),
.A2(n_145),
.B1(n_133),
.B2(n_166),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_239),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_176),
.A2(n_133),
.B(n_149),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_240),
.A2(n_243),
.B(n_208),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_194),
.A2(n_149),
.B(n_152),
.Y(n_243)
);

AO22x1_ASAP7_75t_SL g247 ( 
.A1(n_218),
.A2(n_141),
.B1(n_156),
.B2(n_117),
.Y(n_247)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_247),
.B(n_250),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_178),
.B(n_154),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_225),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_253),
.A2(n_261),
.B1(n_265),
.B2(n_220),
.Y(n_320)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_258),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g289 ( 
.A1(n_259),
.A2(n_171),
.B1(n_189),
.B2(n_214),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_183),
.A2(n_20),
.B1(n_9),
.B2(n_10),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_170),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_262),
.A2(n_211),
.B1(n_182),
.B2(n_186),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_263),
.B(n_188),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_177),
.A2(n_17),
.B1(n_11),
.B2(n_12),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_178),
.B(n_10),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_219),
.Y(n_282)
);

AND2x4_ASAP7_75t_SL g273 ( 
.A(n_184),
.B(n_12),
.Y(n_273)
);

INVx2_ASAP7_75t_SL g313 ( 
.A(n_273),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_233),
.B(n_205),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g337 ( 
.A(n_277),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_278),
.B(n_258),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_280),
.B(n_301),
.Y(n_354)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_252),
.Y(n_281)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_281),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_282),
.B(n_288),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_226),
.B(n_191),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_283),
.B(n_284),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_244),
.B(n_169),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_251),
.B(n_215),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_285),
.B(n_286),
.C(n_302),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_231),
.B(n_181),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_287),
.A2(n_290),
.B1(n_298),
.B2(n_309),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_231),
.B(n_225),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_289),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_250),
.A2(n_202),
.B1(n_207),
.B2(n_200),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_252),
.Y(n_291)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_291),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_269),
.B(n_196),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_293),
.B(n_295),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_267),
.B(n_206),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_294),
.B(n_304),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_254),
.B(n_186),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_228),
.Y(n_296)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_296),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_264),
.B(n_195),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_297),
.B(n_299),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_256),
.A2(n_206),
.B1(n_180),
.B2(n_223),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_264),
.B(n_168),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_228),
.Y(n_300)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_300),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_246),
.B(n_212),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_275),
.B(n_217),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_232),
.Y(n_303)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_303),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_246),
.B(n_190),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_275),
.B(n_249),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_305),
.B(n_268),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_274),
.B(n_167),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_307),
.B(n_314),
.Y(n_349)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_232),
.Y(n_308)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_308),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_257),
.A2(n_221),
.B1(n_199),
.B2(n_220),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_260),
.Y(n_310)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_310),
.Y(n_335)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_255),
.Y(n_312)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_312),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_274),
.B(n_198),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g347 ( 
.A(n_315),
.Y(n_347)
);

AOI22x1_ASAP7_75t_L g316 ( 
.A1(n_257),
.A2(n_222),
.B1(n_189),
.B2(n_175),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_316),
.A2(n_229),
.B1(n_240),
.B2(n_247),
.Y(n_334)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_260),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_318),
.Y(n_355)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_266),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_319),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_320),
.A2(n_227),
.B1(n_253),
.B2(n_235),
.Y(n_326)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_266),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_321),
.B(n_323),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_241),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_322),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_229),
.B(n_185),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_326),
.A2(n_334),
.B1(n_341),
.B2(n_351),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_312),
.Y(n_330)
);

CKINVDCx14_ASAP7_75t_R g368 ( 
.A(n_330),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_279),
.B(n_285),
.C(n_278),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_332),
.B(n_339),
.C(n_357),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_333),
.B(n_294),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_286),
.B(n_248),
.C(n_243),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_287),
.A2(n_242),
.B1(n_237),
.B2(n_265),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g403 ( 
.A1(n_340),
.A2(n_353),
.B1(n_359),
.B2(n_361),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_292),
.A2(n_242),
.B1(n_262),
.B2(n_248),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_315),
.A2(n_248),
.B(n_263),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_344),
.Y(n_378)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_313),
.A2(n_255),
.B(n_273),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g374 ( 
.A(n_346),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_292),
.A2(n_247),
.B1(n_261),
.B2(n_234),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_292),
.A2(n_273),
.B1(n_249),
.B2(n_245),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_282),
.B(n_273),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_356),
.B(n_360),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_288),
.B(n_304),
.C(n_302),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_290),
.A2(n_245),
.B1(n_241),
.B2(n_272),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_312),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_320),
.A2(n_238),
.B1(n_245),
.B2(n_270),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_317),
.A2(n_238),
.B1(n_270),
.B2(n_268),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_363),
.A2(n_317),
.B1(n_291),
.B2(n_281),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_365),
.B(n_296),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_337),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_367),
.B(n_381),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_338),
.Y(n_369)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_369),
.Y(n_420)
);

AND2x2_ASAP7_75t_SL g371 ( 
.A(n_347),
.B(n_313),
.Y(n_371)
);

INVx1_ASAP7_75t_SL g423 ( 
.A(n_371),
.Y(n_423)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_372),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_325),
.B(n_301),
.Y(n_373)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_373),
.Y(n_429)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_335),
.Y(n_375)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_375),
.Y(n_406)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_335),
.Y(n_376)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_376),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_328),
.B(n_325),
.Y(n_377)
);

XNOR2x1_ASAP7_75t_L g428 ( 
.A(n_377),
.B(n_308),
.Y(n_428)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_352),
.Y(n_379)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_379),
.Y(n_436)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_352),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_327),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_382),
.B(n_383),
.Y(n_417)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_327),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_384),
.A2(n_363),
.B1(n_326),
.B2(n_334),
.Y(n_410)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_331),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_385),
.B(n_386),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_350),
.B(n_272),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_324),
.A2(n_298),
.B1(n_306),
.B2(n_313),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_388),
.A2(n_394),
.B1(n_395),
.B2(n_401),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_355),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_389),
.B(n_391),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_349),
.B(n_307),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_390),
.Y(n_404)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_331),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_392),
.B(n_328),
.C(n_332),
.Y(n_405)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_345),
.Y(n_393)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_393),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_324),
.A2(n_306),
.B1(n_311),
.B2(n_309),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_351),
.A2(n_311),
.B1(n_314),
.B2(n_323),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_358),
.B(n_236),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g435 ( 
.A(n_396),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_364),
.B(n_236),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_397),
.A2(n_402),
.B1(n_338),
.B2(n_342),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_355),
.Y(n_398)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_398),
.A2(n_330),
.B(n_360),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_349),
.B(n_303),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_399),
.B(n_400),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_336),
.B(n_321),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_340),
.A2(n_316),
.B1(n_318),
.B2(n_310),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_354),
.B(n_271),
.Y(n_402)
);

MAJx2_ASAP7_75t_L g448 ( 
.A(n_405),
.B(n_413),
.C(n_428),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g407 ( 
.A1(n_378),
.A2(n_347),
.B(n_353),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_407),
.A2(n_419),
.B(n_433),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_410),
.A2(n_414),
.B1(n_415),
.B2(n_421),
.Y(n_455)
);

INVxp67_ASAP7_75t_SL g437 ( 
.A(n_412),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_380),
.B(n_333),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_370),
.A2(n_359),
.B1(n_329),
.B2(n_336),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_370),
.A2(n_329),
.B1(n_344),
.B2(n_356),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_380),
.B(n_357),
.C(n_339),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g438 ( 
.A(n_416),
.B(n_422),
.C(n_426),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_403),
.A2(n_361),
.B1(n_341),
.B2(n_342),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_392),
.B(n_346),
.C(n_348),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_377),
.B(n_348),
.C(n_345),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_374),
.B(n_362),
.C(n_316),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_427),
.B(n_432),
.C(n_422),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_374),
.B(n_362),
.C(n_300),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_378),
.A2(n_343),
.B(n_322),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_403),
.A2(n_343),
.B1(n_366),
.B2(n_319),
.Y(n_434)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_434),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_413),
.B(n_387),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_439),
.B(n_440),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_405),
.B(n_416),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_408),
.Y(n_441)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_441),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_435),
.B(n_367),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_SL g468 ( 
.A(n_442),
.B(n_453),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_426),
.B(n_387),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_443),
.B(n_393),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_428),
.B(n_379),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_444),
.B(n_450),
.Y(n_470)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_408),
.Y(n_445)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_445),
.Y(n_477)
);

AOI22xp33_ASAP7_75t_SL g446 ( 
.A1(n_423),
.A2(n_389),
.B1(n_398),
.B2(n_385),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_446),
.A2(n_460),
.B1(n_433),
.B2(n_419),
.Y(n_472)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_430),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_447),
.B(n_449),
.Y(n_479)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_417),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_432),
.B(n_381),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_451),
.B(n_452),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_415),
.B(n_373),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_411),
.B(n_271),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_SL g454 ( 
.A(n_429),
.B(n_400),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_454),
.B(n_461),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_424),
.B(n_399),
.Y(n_456)
);

CKINVDCx14_ASAP7_75t_R g465 ( 
.A(n_456),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_436),
.B(n_371),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_458),
.B(n_464),
.Y(n_486)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_417),
.Y(n_459)
);

BUFx2_ASAP7_75t_L g487 ( 
.A(n_459),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_407),
.A2(n_401),
.B(n_395),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_460),
.A2(n_391),
.B(n_383),
.Y(n_485)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_425),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_436),
.B(n_371),
.C(n_388),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_462),
.B(n_406),
.C(n_431),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_424),
.B(n_390),
.Y(n_464)
);

BUFx12_ASAP7_75t_L g466 ( 
.A(n_463),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_466),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_455),
.A2(n_421),
.B1(n_410),
.B2(n_404),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_467),
.A2(n_476),
.B1(n_457),
.B2(n_444),
.Y(n_491)
);

NAND4xp25_ASAP7_75t_SL g469 ( 
.A(n_456),
.B(n_394),
.C(n_412),
.D(n_384),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_469),
.B(n_448),
.Y(n_499)
);

A2O1A1O1Ixp25_ASAP7_75t_L g471 ( 
.A1(n_437),
.A2(n_427),
.B(n_423),
.C(n_409),
.D(n_414),
.Y(n_471)
);

AOI21xp33_ASAP7_75t_L g494 ( 
.A1(n_471),
.A2(n_443),
.B(n_439),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_472),
.A2(n_420),
.B1(n_369),
.B2(n_382),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_473),
.B(n_482),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_463),
.A2(n_458),
.B(n_462),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_474),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_455),
.A2(n_434),
.B1(n_409),
.B2(n_431),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_440),
.B(n_406),
.C(n_368),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_480),
.B(n_483),
.C(n_438),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_438),
.B(n_375),
.C(n_376),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_485),
.Y(n_498)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_484),
.Y(n_488)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_488),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_485),
.A2(n_457),
.B1(n_452),
.B2(n_464),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_489),
.A2(n_495),
.B1(n_481),
.B2(n_486),
.Y(n_513)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_479),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_490),
.B(n_499),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_491),
.A2(n_496),
.B1(n_487),
.B2(n_477),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_492),
.B(n_470),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g507 ( 
.A1(n_494),
.A2(n_480),
.B(n_482),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_465),
.A2(n_418),
.B1(n_450),
.B2(n_451),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_475),
.A2(n_369),
.B1(n_420),
.B2(n_448),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_497),
.B(n_504),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_483),
.B(n_276),
.C(n_201),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_502),
.B(n_503),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_468),
.B(n_276),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_478),
.B(n_13),
.C(n_15),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_487),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_505),
.B(n_473),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_SL g506 ( 
.A1(n_493),
.A2(n_474),
.B(n_471),
.Y(n_506)
);

OAI21xp5_ASAP7_75t_L g533 ( 
.A1(n_506),
.A2(n_507),
.B(n_513),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_509),
.A2(n_466),
.B1(n_469),
.B2(n_16),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_492),
.B(n_478),
.C(n_501),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_510),
.B(n_511),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g511 ( 
.A(n_500),
.Y(n_511)
);

HB1xp67_ASAP7_75t_L g514 ( 
.A(n_501),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_514),
.B(n_517),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_495),
.B(n_481),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_516),
.B(n_521),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_493),
.B(n_470),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_518),
.B(n_519),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_502),
.B(n_486),
.C(n_476),
.Y(n_521)
);

INVxp67_ASAP7_75t_L g522 ( 
.A(n_512),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_522),
.B(n_530),
.Y(n_543)
);

OR2x2_ASAP7_75t_L g523 ( 
.A(n_509),
.B(n_489),
.Y(n_523)
);

OAI21x1_ASAP7_75t_L g539 ( 
.A1(n_523),
.A2(n_516),
.B(n_521),
.Y(n_539)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_515),
.A2(n_467),
.B1(n_498),
.B2(n_491),
.Y(n_525)
);

OR2x2_ASAP7_75t_L g537 ( 
.A(n_525),
.B(n_527),
.Y(n_537)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_508),
.A2(n_498),
.B1(n_504),
.B2(n_496),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_510),
.B(n_466),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_529),
.B(n_532),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_507),
.B(n_13),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_531),
.B(n_17),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_519),
.B(n_13),
.C(n_15),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_524),
.B(n_511),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_536),
.B(n_539),
.Y(n_546)
);

NAND3xp33_ASAP7_75t_SL g538 ( 
.A(n_533),
.B(n_520),
.C(n_513),
.Y(n_538)
);

CKINVDCx14_ASAP7_75t_R g544 ( 
.A(n_538),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_522),
.B(n_15),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_540),
.B(n_541),
.C(n_531),
.Y(n_545)
);

NOR2xp67_ASAP7_75t_L g541 ( 
.A(n_534),
.B(n_16),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g548 ( 
.A(n_542),
.B(n_532),
.C(n_523),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_545),
.B(n_547),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_537),
.B(n_526),
.C(n_528),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_548),
.B(n_535),
.Y(n_550)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_550),
.Y(n_553)
);

AOI21xp5_ASAP7_75t_L g551 ( 
.A1(n_546),
.A2(n_544),
.B(n_543),
.Y(n_551)
);

OAI21xp5_ASAP7_75t_L g552 ( 
.A1(n_551),
.A2(n_543),
.B(n_530),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_552),
.B(n_549),
.Y(n_554)
);

XOR2xp5_ASAP7_75t_L g555 ( 
.A(n_554),
.B(n_553),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_SL g556 ( 
.A(n_555),
.B(n_17),
.Y(n_556)
);


endmodule