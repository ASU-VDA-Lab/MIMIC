module fake_jpeg_29700_n_390 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_390);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_390;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx24_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx16f_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_16),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_46),
.B(n_47),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_23),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_53),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_54),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_15),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_62),
.Y(n_94)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_61),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_25),
.B(n_15),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_63),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_25),
.B(n_14),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_82),
.Y(n_95)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_26),
.B(n_14),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_66),
.B(n_67),
.Y(n_111)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_45),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

INVx8_ASAP7_75t_L g115 ( 
.A(n_68),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_17),
.Y(n_69)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_71),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_26),
.B(n_1),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_72),
.B(n_76),
.Y(n_104)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_73),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_75),
.B(n_77),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_28),
.B(n_30),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_17),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_78),
.B(n_20),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_28),
.B(n_1),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_79),
.B(n_1),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_80),
.B(n_81),
.Y(n_128)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_17),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_51),
.A2(n_56),
.B1(n_80),
.B2(n_75),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_84),
.A2(n_87),
.B1(n_99),
.B2(n_102),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_52),
.A2(n_33),
.B1(n_40),
.B2(n_32),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_85),
.A2(n_89),
.B1(n_97),
.B2(n_106),
.Y(n_156)
);

A2O1A1Ixp33_ASAP7_75t_L g86 ( 
.A1(n_67),
.A2(n_23),
.B(n_32),
.C(n_41),
.Y(n_86)
);

OAI32xp33_ASAP7_75t_L g150 ( 
.A1(n_86),
.A2(n_120),
.A3(n_39),
.B1(n_29),
.B2(n_74),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_48),
.A2(n_36),
.B1(n_38),
.B2(n_43),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_53),
.A2(n_33),
.B1(n_40),
.B2(n_32),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_54),
.B(n_41),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_92),
.B(n_113),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_68),
.A2(n_33),
.B1(n_40),
.B2(n_32),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_70),
.A2(n_33),
.B1(n_40),
.B2(n_30),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_50),
.A2(n_36),
.B1(n_43),
.B2(n_42),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_59),
.A2(n_36),
.B1(n_43),
.B2(n_42),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_103),
.A2(n_121),
.B1(n_2),
.B2(n_3),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_82),
.A2(n_32),
.B1(n_36),
.B2(n_43),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_130),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_61),
.B(n_31),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_63),
.B(n_31),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_117),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_77),
.B(n_44),
.Y(n_117)
);

AO22x1_ASAP7_75t_L g120 ( 
.A1(n_65),
.A2(n_39),
.B1(n_23),
.B2(n_45),
.Y(n_120)
);

OAI22xp33_ASAP7_75t_L g121 ( 
.A1(n_49),
.A2(n_42),
.B1(n_38),
.B2(n_24),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_81),
.B(n_44),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_124),
.B(n_125),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_71),
.B(n_22),
.Y(n_125)
);

OA22x2_ASAP7_75t_L g126 ( 
.A1(n_57),
.A2(n_39),
.B1(n_22),
.B2(n_29),
.Y(n_126)
);

AO22x2_ASAP7_75t_L g161 ( 
.A1(n_126),
.A2(n_39),
.B1(n_29),
.B2(n_37),
.Y(n_161)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_98),
.Y(n_132)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_132),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_133),
.Y(n_178)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_134),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_83),
.Y(n_135)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_135),
.Y(n_196)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_139),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_120),
.A2(n_38),
.B1(n_42),
.B2(n_29),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_L g185 ( 
.A1(n_140),
.A2(n_171),
.B1(n_176),
.B2(n_129),
.Y(n_185)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_98),
.Y(n_141)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_141),
.Y(n_194)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_142),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_95),
.B(n_69),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_143),
.B(n_148),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_104),
.B(n_60),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_145),
.B(n_147),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_60),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_146),
.B(n_155),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_90),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_73),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_105),
.Y(n_149)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_149),
.Y(n_202)
);

AO22x2_ASAP7_75t_L g184 ( 
.A1(n_150),
.A2(n_161),
.B1(n_91),
.B2(n_93),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_92),
.B(n_55),
.C(n_38),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_151),
.B(n_162),
.C(n_163),
.Y(n_199)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_110),
.Y(n_152)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_152),
.Y(n_195)
);

INVx4_ASAP7_75t_SL g153 ( 
.A(n_100),
.Y(n_153)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_153),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_108),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_154),
.B(n_158),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_94),
.Y(n_155)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_131),
.Y(n_157)
);

INVx8_ASAP7_75t_L g186 ( 
.A(n_157),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_118),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_108),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_159),
.B(n_167),
.Y(n_204)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_110),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_160),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_29),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_118),
.B(n_37),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_118),
.B(n_1),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_164),
.B(n_144),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_112),
.Y(n_165)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_165),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_128),
.Y(n_167)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_131),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_168),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_86),
.B(n_37),
.C(n_24),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_169),
.A2(n_93),
.B(n_91),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_170),
.A2(n_166),
.B1(n_156),
.B2(n_148),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_122),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_83),
.B(n_2),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_172),
.B(n_173),
.Y(n_215)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_119),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_128),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_174),
.B(n_175),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_101),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_122),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_138),
.B(n_101),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_177),
.B(n_200),
.Y(n_224)
);

OAI32xp33_ASAP7_75t_L g180 ( 
.A1(n_136),
.A2(n_121),
.A3(n_128),
.B1(n_88),
.B2(n_107),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_180),
.B(n_181),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_133),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_184),
.B(n_10),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_185),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_189),
.A2(n_190),
.B1(n_192),
.B2(n_214),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_162),
.A2(n_148),
.B1(n_156),
.B2(n_143),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_162),
.A2(n_129),
.B1(n_112),
.B2(n_115),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_198),
.B(n_210),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_144),
.B(n_96),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_157),
.Y(n_203)
);

INVxp67_ASAP7_75t_SL g223 ( 
.A(n_203),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_136),
.B(n_107),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_207),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_137),
.B(n_123),
.Y(n_207)
);

O2A1O1Ixp33_ASAP7_75t_L g210 ( 
.A1(n_155),
.A2(n_127),
.B(n_106),
.C(n_85),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_168),
.Y(n_211)
);

INVxp67_ASAP7_75t_SL g227 ( 
.A(n_211),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_212),
.A2(n_9),
.B(n_10),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_169),
.A2(n_127),
.B(n_5),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_213),
.A2(n_4),
.B(n_5),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_143),
.A2(n_123),
.B1(n_115),
.B2(n_96),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_182),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_217),
.B(n_208),
.Y(n_256)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_191),
.Y(n_218)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_218),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_179),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_221),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_188),
.B(n_137),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_222),
.B(n_236),
.Y(n_252)
);

AOI22x1_ASAP7_75t_L g225 ( 
.A1(n_184),
.A2(n_150),
.B1(n_161),
.B2(n_163),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_225),
.B(n_229),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_199),
.B(n_151),
.C(n_146),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_226),
.B(n_233),
.C(n_197),
.Y(n_267)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_191),
.Y(n_228)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_228),
.Y(n_255)
);

AND2x4_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_161),
.Y(n_229)
);

AOI221xp5_ASAP7_75t_SL g230 ( 
.A1(n_188),
.A2(n_161),
.B1(n_164),
.B2(n_163),
.C(n_149),
.Y(n_230)
);

NOR2x1_ASAP7_75t_R g266 ( 
.A(n_230),
.B(n_184),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_198),
.B(n_132),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_231),
.B(n_234),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_232),
.A2(n_192),
.B(n_211),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_199),
.B(n_142),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_200),
.B(n_160),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_216),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_235),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_204),
.B(n_175),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_189),
.A2(n_161),
.B1(n_165),
.B2(n_153),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_237),
.A2(n_242),
.B1(n_248),
.B2(n_213),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_207),
.B(n_152),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_241),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_177),
.B(n_159),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g242 ( 
.A1(n_210),
.A2(n_173),
.B1(n_134),
.B2(n_154),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_243),
.A2(n_251),
.B1(n_209),
.B2(n_203),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_183),
.B(n_6),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_244),
.B(n_245),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_183),
.B(n_8),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_215),
.B(n_9),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_246),
.B(n_250),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_247),
.B(n_214),
.Y(n_261)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_195),
.Y(n_249)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_249),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_201),
.B(n_11),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_184),
.A2(n_11),
.B1(n_12),
.B2(n_212),
.Y(n_251)
);

OAI22x1_ASAP7_75t_L g253 ( 
.A1(n_230),
.A2(n_184),
.B1(n_180),
.B2(n_190),
.Y(n_253)
);

OA22x2_ASAP7_75t_L g284 ( 
.A1(n_253),
.A2(n_260),
.B1(n_266),
.B2(n_251),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_256),
.B(n_258),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_201),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_261),
.B(n_248),
.Y(n_286)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_218),
.Y(n_265)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_265),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_267),
.B(n_268),
.C(n_275),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_233),
.B(n_202),
.C(n_197),
.Y(n_268)
);

NOR3xp33_ASAP7_75t_L g269 ( 
.A(n_235),
.B(n_208),
.C(n_181),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_269),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_270),
.A2(n_247),
.B(n_248),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_226),
.B(n_202),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_271),
.B(n_178),
.C(n_223),
.Y(n_305)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_228),
.Y(n_273)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_273),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_221),
.B(n_196),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_274),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_222),
.B(n_194),
.C(n_196),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_276),
.A2(n_219),
.B1(n_238),
.B2(n_234),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_237),
.A2(n_194),
.B1(n_187),
.B2(n_209),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_277),
.A2(n_242),
.B1(n_243),
.B2(n_229),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_220),
.B(n_206),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_244),
.C(n_245),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_220),
.B(n_187),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_281),
.B(n_195),
.Y(n_303)
);

AOI322xp5_ASAP7_75t_L g283 ( 
.A1(n_253),
.A2(n_238),
.A3(n_219),
.B1(n_239),
.B2(n_224),
.C1(n_248),
.C2(n_225),
.Y(n_283)
);

NAND3xp33_ASAP7_75t_L g314 ( 
.A(n_283),
.B(n_252),
.C(n_280),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_284),
.B(n_285),
.Y(n_307)
);

XNOR2x1_ASAP7_75t_L g317 ( 
.A(n_286),
.B(n_295),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_288),
.A2(n_299),
.B(n_262),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_266),
.A2(n_239),
.B1(n_240),
.B2(n_224),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_289),
.B(n_293),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_290),
.A2(n_297),
.B1(n_302),
.B2(n_280),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_257),
.A2(n_229),
.B1(n_225),
.B2(n_231),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_257),
.A2(n_229),
.B1(n_225),
.B2(n_246),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_294),
.B(n_303),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_267),
.B(n_236),
.C(n_229),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_296),
.B(n_300),
.C(n_305),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_260),
.A2(n_232),
.B1(n_250),
.B2(n_186),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_257),
.A2(n_227),
.B(n_223),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_271),
.B(n_193),
.C(n_186),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_277),
.A2(n_186),
.B1(n_193),
.B2(n_249),
.Y(n_302)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_254),
.Y(n_304)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_304),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_268),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_306),
.B(n_305),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_298),
.B(n_272),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_309),
.B(n_314),
.Y(n_330)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_287),
.Y(n_310)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_310),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_311),
.B(n_325),
.Y(n_326)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_287),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_313),
.B(n_321),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_291),
.B(n_278),
.C(n_275),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_316),
.B(n_320),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_318),
.A2(n_324),
.B1(n_285),
.B2(n_294),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_300),
.B(n_281),
.C(n_252),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_292),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_296),
.B(n_262),
.C(n_261),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_322),
.B(n_301),
.Y(n_336)
);

NOR3xp33_ASAP7_75t_L g323 ( 
.A(n_282),
.B(n_272),
.C(n_259),
.Y(n_323)
);

NOR3xp33_ASAP7_75t_L g331 ( 
.A(n_323),
.B(n_310),
.C(n_321),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_297),
.A2(n_259),
.B1(n_270),
.B2(n_273),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_299),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_327),
.B(n_329),
.Y(n_355)
);

NAND4xp25_ASAP7_75t_L g328 ( 
.A(n_324),
.B(n_282),
.C(n_293),
.D(n_298),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_328),
.A2(n_331),
.B(n_312),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g333 ( 
.A1(n_308),
.A2(n_288),
.B(n_284),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_333),
.A2(n_334),
.B(n_337),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_312),
.B(n_303),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_318),
.A2(n_290),
.B1(n_302),
.B2(n_286),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_335),
.A2(n_338),
.B1(n_320),
.B2(n_279),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_336),
.B(n_339),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_313),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_307),
.A2(n_289),
.B1(n_284),
.B2(n_301),
.Y(n_338)
);

XNOR2x1_ASAP7_75t_L g339 ( 
.A(n_322),
.B(n_284),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_308),
.A2(n_292),
.B(n_304),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_341),
.A2(n_255),
.B(n_265),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_343),
.A2(n_341),
.B(n_338),
.Y(n_357)
);

A2O1A1O1Ixp25_ASAP7_75t_L g344 ( 
.A1(n_326),
.A2(n_307),
.B(n_311),
.C(n_317),
.D(n_325),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_344),
.B(n_353),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_329),
.B(n_316),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_347),
.B(n_348),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_339),
.B(n_315),
.Y(n_348)
);

AOI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_328),
.A2(n_319),
.B(n_279),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_349),
.B(n_351),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_332),
.B(n_315),
.C(n_306),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_350),
.B(n_327),
.C(n_295),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g352 ( 
.A(n_330),
.B(n_263),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_352),
.B(n_354),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_333),
.B(n_317),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_349),
.A2(n_335),
.B1(n_326),
.B2(n_334),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_356),
.B(n_358),
.Y(n_371)
);

OAI21xp33_ASAP7_75t_SL g370 ( 
.A1(n_357),
.A2(n_346),
.B(n_355),
.Y(n_370)
);

INVx11_ASAP7_75t_L g358 ( 
.A(n_345),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_360),
.B(n_364),
.C(n_365),
.Y(n_368)
);

OR2x2_ASAP7_75t_L g361 ( 
.A(n_351),
.B(n_337),
.Y(n_361)
);

AOI31xp33_ASAP7_75t_L g369 ( 
.A1(n_361),
.A2(n_358),
.A3(n_344),
.B(n_357),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_350),
.B(n_342),
.C(n_340),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_347),
.B(n_342),
.C(n_340),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_363),
.A2(n_346),
.B(n_353),
.Y(n_367)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_367),
.A2(n_373),
.B(n_361),
.Y(n_378)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_369),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_370),
.A2(n_374),
.B(n_366),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_360),
.B(n_355),
.C(n_348),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g379 ( 
.A(n_372),
.B(n_375),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_362),
.A2(n_254),
.B(n_255),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_364),
.A2(n_264),
.B(n_263),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_359),
.B(n_264),
.C(n_178),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_368),
.B(n_365),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_376),
.B(n_380),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_378),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_369),
.A2(n_366),
.B1(n_356),
.B2(n_359),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_381),
.A2(n_382),
.B(n_12),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_371),
.B(n_227),
.C(n_11),
.Y(n_382)
);

OAI21x1_ASAP7_75t_L g388 ( 
.A1(n_383),
.A2(n_386),
.B(n_377),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_377),
.A2(n_379),
.B(n_382),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_385),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_387),
.B(n_388),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_389),
.B(n_384),
.Y(n_390)
);


endmodule