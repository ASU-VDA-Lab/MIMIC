module fake_netlist_5_2002_n_1840 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1840);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1840;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_1809;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_604;
wire n_314;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1406;
wire n_1279;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_681;
wire n_584;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_990;
wire n_836;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1747;
wire n_714;
wire n_1817;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_174),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_33),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_49),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_87),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_100),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_28),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_170),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_150),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_19),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_59),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_103),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_161),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_99),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_133),
.Y(n_198)
);

BUFx10_ASAP7_75t_L g199 ( 
.A(n_33),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_173),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_121),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_83),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_85),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_111),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_71),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_15),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_10),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_153),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_182),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_152),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_167),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_106),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_21),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_125),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_180),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_9),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_34),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_30),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_25),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_9),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g221 ( 
.A(n_155),
.Y(n_221)
);

BUFx5_ASAP7_75t_L g222 ( 
.A(n_61),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_77),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_39),
.Y(n_224)
);

BUFx10_ASAP7_75t_L g225 ( 
.A(n_38),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_26),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_63),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_101),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_7),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_151),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_122),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_139),
.Y(n_232)
);

INVx2_ASAP7_75t_SL g233 ( 
.A(n_114),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_41),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_81),
.Y(n_235)
);

BUFx5_ASAP7_75t_L g236 ( 
.A(n_34),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_118),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_175),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_50),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_128),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_94),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_22),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_115),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_145),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_18),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_110),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_72),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_76),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_109),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_63),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_65),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_93),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_119),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_15),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_66),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_95),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_46),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_79),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_51),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_31),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_19),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_52),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_104),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_64),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_0),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_22),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_3),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_75),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_140),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_56),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_162),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_141),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_96),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_57),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_5),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_2),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_159),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_172),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_129),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_32),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_144),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_17),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_98),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_88),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_73),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_3),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_91),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_32),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_23),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_28),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_179),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_38),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_21),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_135),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_1),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_183),
.Y(n_296)
);

INVx2_ASAP7_75t_SL g297 ( 
.A(n_105),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_74),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_160),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_39),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_120),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_146),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_132),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_130),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_149),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_36),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_57),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_45),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_30),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_84),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_70),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_126),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_134),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_127),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_78),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_64),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_143),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_181),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_178),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_42),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_52),
.Y(n_321)
);

BUFx5_ASAP7_75t_L g322 ( 
.A(n_13),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_29),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_171),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_80),
.Y(n_325)
);

INVx2_ASAP7_75t_SL g326 ( 
.A(n_92),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_40),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_13),
.Y(n_328)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_6),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_50),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_24),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_86),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_46),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_26),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_89),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_69),
.Y(n_336)
);

BUFx10_ASAP7_75t_L g337 ( 
.A(n_102),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_117),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_147),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_20),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_1),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_123),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_62),
.Y(n_343)
);

BUFx10_ASAP7_75t_L g344 ( 
.A(n_44),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_158),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_7),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_107),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_55),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_20),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_24),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_113),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_2),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_53),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_154),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_56),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_67),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_131),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_43),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_29),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_49),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_25),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_60),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_163),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_202),
.Y(n_364)
);

INVxp67_ASAP7_75t_SL g365 ( 
.A(n_221),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_267),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_222),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_222),
.Y(n_368)
);

BUFx10_ASAP7_75t_L g369 ( 
.A(n_334),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_222),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_222),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_222),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_222),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_202),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_222),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_236),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_236),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_236),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_227),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_236),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g381 ( 
.A(n_186),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_307),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_199),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_237),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_236),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_236),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_236),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_322),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_322),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_187),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_322),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_322),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_322),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_322),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_322),
.Y(n_395)
);

INVxp67_ASAP7_75t_SL g396 ( 
.A(n_269),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_190),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_190),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_237),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_190),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_194),
.Y(n_401)
);

INVx1_ASAP7_75t_SL g402 ( 
.A(n_199),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_216),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_225),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_190),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_234),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_234),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_234),
.Y(n_408)
);

INVxp67_ASAP7_75t_SL g409 ( 
.A(n_311),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_234),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_343),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_343),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_217),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_343),
.Y(n_414)
);

INVxp67_ASAP7_75t_SL g415 ( 
.A(n_343),
.Y(n_415)
);

INVxp67_ASAP7_75t_SL g416 ( 
.A(n_350),
.Y(n_416)
);

INVxp33_ASAP7_75t_SL g417 ( 
.A(n_186),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_350),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_350),
.Y(n_419)
);

INVx3_ASAP7_75t_L g420 ( 
.A(n_350),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_193),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_225),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_213),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_218),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_247),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_224),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_247),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_250),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_219),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_257),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_225),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_344),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_262),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_273),
.Y(n_434)
);

INVxp67_ASAP7_75t_SL g435 ( 
.A(n_192),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_264),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_275),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_280),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_206),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_220),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_286),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_344),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_273),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_293),
.Y(n_444)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_203),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_295),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_300),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_226),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_306),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_316),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_260),
.Y(n_451)
);

CKINVDCx16_ASAP7_75t_R g452 ( 
.A(n_287),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_301),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_260),
.Y(n_454)
);

INVxp33_ASAP7_75t_L g455 ( 
.A(n_320),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_321),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_301),
.Y(n_457)
);

INVxp67_ASAP7_75t_SL g458 ( 
.A(n_195),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_327),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_330),
.Y(n_460)
);

INVx1_ASAP7_75t_SL g461 ( 
.A(n_344),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_206),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_346),
.Y(n_463)
);

INVxp33_ASAP7_75t_SL g464 ( 
.A(n_207),
.Y(n_464)
);

BUFx2_ASAP7_75t_L g465 ( 
.A(n_207),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_229),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_189),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_367),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_368),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_397),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_373),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_397),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_435),
.B(n_208),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_373),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_370),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_366),
.B(n_337),
.Y(n_476)
);

INVxp33_ASAP7_75t_SL g477 ( 
.A(n_379),
.Y(n_477)
);

BUFx8_ASAP7_75t_L g478 ( 
.A(n_381),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_415),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_371),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_467),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_375),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_416),
.Y(n_483)
);

INVx5_ASAP7_75t_L g484 ( 
.A(n_420),
.Y(n_484)
);

AND2x2_ASAP7_75t_SL g485 ( 
.A(n_445),
.B(n_191),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_364),
.A2(n_276),
.B1(n_288),
.B2(n_270),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_420),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_372),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g489 ( 
.A(n_439),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_390),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_398),
.Y(n_491)
);

CKINVDCx8_ASAP7_75t_R g492 ( 
.A(n_379),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_390),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_458),
.B(n_208),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_375),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_400),
.Y(n_496)
);

BUFx8_ASAP7_75t_L g497 ( 
.A(n_381),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_405),
.B(n_233),
.Y(n_498)
);

AND2x2_ASAP7_75t_SL g499 ( 
.A(n_452),
.B(n_191),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_406),
.B(n_233),
.Y(n_500)
);

OAI21x1_ASAP7_75t_L g501 ( 
.A1(n_376),
.A2(n_315),
.B(n_249),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_407),
.B(n_297),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_408),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_376),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_401),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_377),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_377),
.B(n_297),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_410),
.B(n_411),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_378),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_412),
.B(n_326),
.Y(n_510)
);

HB1xp67_ASAP7_75t_L g511 ( 
.A(n_462),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_378),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_414),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_418),
.Y(n_514)
);

AND2x4_ASAP7_75t_L g515 ( 
.A(n_380),
.B(n_326),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_419),
.B(n_249),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_380),
.B(n_185),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_385),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_385),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_386),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_386),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_387),
.B(n_315),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_387),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_388),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_388),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_403),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_389),
.B(n_185),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_389),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_391),
.Y(n_529)
);

AND2x4_ASAP7_75t_L g530 ( 
.A(n_391),
.B(n_198),
.Y(n_530)
);

BUFx3_ASAP7_75t_L g531 ( 
.A(n_392),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_392),
.B(n_200),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_393),
.B(n_201),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_394),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_394),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_395),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_395),
.B(n_204),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_451),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_451),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_454),
.Y(n_540)
);

INVxp33_ASAP7_75t_SL g541 ( 
.A(n_382),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_454),
.Y(n_542)
);

OA21x2_ASAP7_75t_L g543 ( 
.A1(n_421),
.A2(n_362),
.B(n_360),
.Y(n_543)
);

CKINVDCx16_ASAP7_75t_R g544 ( 
.A(n_374),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_423),
.B(n_200),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_L g546 ( 
.A1(n_499),
.A2(n_396),
.B1(n_409),
.B2(n_365),
.Y(n_546)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_474),
.Y(n_547)
);

NAND3xp33_ASAP7_75t_L g548 ( 
.A(n_545),
.B(n_424),
.C(n_413),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_508),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_499),
.B(n_413),
.Y(n_550)
);

INVx2_ASAP7_75t_SL g551 ( 
.A(n_485),
.Y(n_551)
);

INVx4_ASAP7_75t_L g552 ( 
.A(n_474),
.Y(n_552)
);

BUFx4f_ASAP7_75t_L g553 ( 
.A(n_543),
.Y(n_553)
);

AND3x4_ASAP7_75t_L g554 ( 
.A(n_486),
.B(n_399),
.C(n_384),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_473),
.B(n_424),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_479),
.B(n_417),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_479),
.B(n_417),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_474),
.Y(n_558)
);

BUFx6f_ASAP7_75t_L g559 ( 
.A(n_474),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_495),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_485),
.B(n_429),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_485),
.Y(n_562)
);

BUFx4f_ASAP7_75t_L g563 ( 
.A(n_543),
.Y(n_563)
);

INVxp33_ASAP7_75t_SL g564 ( 
.A(n_490),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_473),
.B(n_483),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_508),
.Y(n_566)
);

AND2x2_ASAP7_75t_SL g567 ( 
.A(n_543),
.B(n_188),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_495),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_508),
.Y(n_569)
);

NAND2xp33_ASAP7_75t_L g570 ( 
.A(n_517),
.B(n_188),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_531),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_474),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_473),
.B(n_429),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_483),
.B(n_464),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_495),
.Y(n_575)
);

AO21x2_ASAP7_75t_L g576 ( 
.A1(n_517),
.A2(n_211),
.B(n_209),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_506),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_531),
.B(n_440),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_489),
.B(n_464),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_518),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_527),
.B(n_440),
.Y(n_581)
);

INVx4_ASAP7_75t_L g582 ( 
.A(n_474),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_518),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_474),
.Y(n_584)
);

AO21x2_ASAP7_75t_L g585 ( 
.A1(n_527),
.A2(n_532),
.B(n_501),
.Y(n_585)
);

INVx4_ASAP7_75t_L g586 ( 
.A(n_504),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_506),
.Y(n_587)
);

BUFx10_ASAP7_75t_L g588 ( 
.A(n_493),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_489),
.B(n_448),
.Y(n_589)
);

OR2x2_ASAP7_75t_L g590 ( 
.A(n_532),
.B(n_465),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_519),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_506),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_519),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_520),
.B(n_448),
.Y(n_594)
);

OR2x2_ASAP7_75t_L g595 ( 
.A(n_511),
.B(n_465),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_520),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_512),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_523),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_523),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_481),
.Y(n_600)
);

BUFx10_ASAP7_75t_L g601 ( 
.A(n_505),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_512),
.Y(n_602)
);

INVx2_ASAP7_75t_SL g603 ( 
.A(n_511),
.Y(n_603)
);

INVx5_ASAP7_75t_L g604 ( 
.A(n_504),
.Y(n_604)
);

BUFx2_ASAP7_75t_L g605 ( 
.A(n_478),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_512),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_521),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_525),
.Y(n_608)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_476),
.B(n_466),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_525),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_529),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_521),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_529),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_521),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_544),
.Y(n_615)
);

INVxp67_ASAP7_75t_SL g616 ( 
.A(n_471),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_494),
.B(n_382),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_494),
.B(n_402),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_477),
.B(n_431),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_504),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_534),
.Y(n_621)
);

BUFx6f_ASAP7_75t_SL g622 ( 
.A(n_507),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_534),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_504),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_536),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_536),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_507),
.B(n_251),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_541),
.B(n_461),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_524),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_530),
.A2(n_426),
.B1(n_430),
.B2(n_428),
.Y(n_630)
);

BUFx3_ASAP7_75t_L g631 ( 
.A(n_530),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_526),
.B(n_369),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_507),
.B(n_515),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_471),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_524),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_471),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_530),
.B(n_433),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_530),
.B(n_436),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_504),
.Y(n_639)
);

INVx4_ASAP7_75t_L g640 ( 
.A(n_504),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_524),
.Y(n_641)
);

NAND3xp33_ASAP7_75t_L g642 ( 
.A(n_545),
.B(n_404),
.C(n_383),
.Y(n_642)
);

AOI21x1_ASAP7_75t_L g643 ( 
.A1(n_522),
.A2(n_215),
.B(n_212),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_535),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_535),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_504),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_535),
.Y(n_647)
);

BUFx6f_ASAP7_75t_L g648 ( 
.A(n_509),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_507),
.B(n_336),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_507),
.B(n_196),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_491),
.B(n_422),
.Y(n_651)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_509),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_515),
.B(n_197),
.Y(n_653)
);

NOR2x1p5_ASAP7_75t_L g654 ( 
.A(n_500),
.B(n_355),
.Y(n_654)
);

INVx4_ASAP7_75t_L g655 ( 
.A(n_509),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_492),
.B(n_369),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_468),
.Y(n_657)
);

INVx6_ASAP7_75t_L g658 ( 
.A(n_484),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_492),
.B(n_432),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_491),
.B(n_442),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_468),
.Y(n_661)
);

INVx5_ASAP7_75t_L g662 ( 
.A(n_509),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_537),
.A2(n_437),
.B1(n_441),
.B2(n_438),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_482),
.Y(n_664)
);

NAND3xp33_ASAP7_75t_SL g665 ( 
.A(n_500),
.B(n_276),
.C(n_270),
.Y(n_665)
);

AOI22xp33_ASAP7_75t_L g666 ( 
.A1(n_537),
.A2(n_463),
.B1(n_460),
.B2(n_459),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_537),
.A2(n_449),
.B1(n_456),
.B2(n_446),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_509),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_498),
.B(n_444),
.Y(n_669)
);

INVxp33_ASAP7_75t_L g670 ( 
.A(n_486),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_482),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_468),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_469),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_482),
.Y(n_674)
);

BUFx3_ASAP7_75t_L g675 ( 
.A(n_533),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_469),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_482),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_509),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_498),
.B(n_447),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_469),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_496),
.B(n_455),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_475),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_503),
.B(n_425),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_475),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_475),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_631),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_618),
.B(n_515),
.Y(n_687)
);

AND2x4_ASAP7_75t_L g688 ( 
.A(n_637),
.B(n_638),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_560),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_631),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_580),
.B(n_533),
.Y(n_691)
);

HB1xp67_ASAP7_75t_L g692 ( 
.A(n_603),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_603),
.B(n_556),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_580),
.B(n_533),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_583),
.B(n_533),
.Y(n_695)
);

BUFx5_ASAP7_75t_L g696 ( 
.A(n_567),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_675),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_553),
.B(n_563),
.Y(n_698)
);

NAND2x1_ASAP7_75t_L g699 ( 
.A(n_658),
.B(n_533),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_669),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_553),
.B(n_509),
.Y(n_701)
);

NAND2xp33_ASAP7_75t_L g702 ( 
.A(n_551),
.B(n_228),
.Y(n_702)
);

OAI22xp5_ASAP7_75t_SL g703 ( 
.A1(n_554),
.A2(n_434),
.B1(n_443),
.B2(n_427),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_583),
.B(n_522),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_675),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_611),
.B(n_522),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_560),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_553),
.B(n_528),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_611),
.B(n_543),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_563),
.B(n_528),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_613),
.B(n_543),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_581),
.B(n_551),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_600),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_568),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_591),
.B(n_528),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_593),
.B(n_528),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_571),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_596),
.B(n_528),
.Y(n_718)
);

O2A1O1Ixp33_ASAP7_75t_L g719 ( 
.A1(n_562),
.A2(n_565),
.B(n_573),
.C(n_555),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_568),
.Y(n_720)
);

INVx1_ASAP7_75t_SL g721 ( 
.A(n_595),
.Y(n_721)
);

OR2x6_ASAP7_75t_L g722 ( 
.A(n_605),
.B(n_450),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_575),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_598),
.B(n_528),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_562),
.B(n_617),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_575),
.Y(n_726)
);

OR2x2_ASAP7_75t_L g727 ( 
.A(n_595),
.B(n_544),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_577),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_599),
.B(n_480),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_549),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_590),
.B(n_254),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_608),
.B(n_480),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_610),
.B(n_480),
.Y(n_733)
);

AOI22xp5_ASAP7_75t_L g734 ( 
.A1(n_550),
.A2(n_453),
.B1(n_457),
.B2(n_271),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_561),
.A2(n_305),
.B1(n_291),
.B2(n_258),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_577),
.Y(n_736)
);

NOR3xp33_ASAP7_75t_L g737 ( 
.A(n_619),
.B(n_290),
.C(n_265),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_563),
.B(n_188),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_567),
.B(n_188),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_621),
.B(n_488),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_594),
.B(n_309),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_566),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_569),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_633),
.B(n_497),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_623),
.B(n_516),
.Y(n_745)
);

OAI22xp5_ASAP7_75t_L g746 ( 
.A1(n_627),
.A2(n_277),
.B1(n_304),
.B2(n_303),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_625),
.B(n_516),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_557),
.B(n_329),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_626),
.B(n_516),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_637),
.Y(n_750)
);

INVx8_ASAP7_75t_L g751 ( 
.A(n_622),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_616),
.B(n_637),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_600),
.Y(n_753)
);

INVxp67_ASAP7_75t_L g754 ( 
.A(n_579),
.Y(n_754)
);

O2A1O1Ixp5_ASAP7_75t_L g755 ( 
.A1(n_634),
.A2(n_510),
.B(n_498),
.C(n_502),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_587),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_638),
.B(n_502),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_638),
.B(n_649),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_574),
.B(n_205),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_578),
.B(n_497),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_L g761 ( 
.A1(n_609),
.A2(n_248),
.B1(n_243),
.B2(n_241),
.Y(n_761)
);

NAND2xp33_ASAP7_75t_L g762 ( 
.A(n_650),
.B(n_231),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_592),
.Y(n_763)
);

INVxp67_ASAP7_75t_L g764 ( 
.A(n_628),
.Y(n_764)
);

INVx2_ASAP7_75t_SL g765 ( 
.A(n_669),
.Y(n_765)
);

INVx2_ASAP7_75t_L g766 ( 
.A(n_592),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_589),
.B(n_223),
.Y(n_767)
);

BUFx3_ASAP7_75t_L g768 ( 
.A(n_588),
.Y(n_768)
);

NOR3xp33_ASAP7_75t_L g769 ( 
.A(n_665),
.B(n_242),
.C(n_239),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_681),
.B(n_502),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_548),
.B(n_546),
.Y(n_771)
);

INVx2_ASAP7_75t_SL g772 ( 
.A(n_679),
.Y(n_772)
);

AOI22xp33_ASAP7_75t_L g773 ( 
.A1(n_576),
.A2(n_501),
.B1(n_348),
.B2(n_288),
.Y(n_773)
);

INVx2_ASAP7_75t_SL g774 ( 
.A(n_679),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_642),
.B(n_205),
.Y(n_775)
);

AOI22xp33_ASAP7_75t_L g776 ( 
.A1(n_576),
.A2(n_501),
.B1(n_348),
.B2(n_353),
.Y(n_776)
);

BUFx12f_ASAP7_75t_L g777 ( 
.A(n_588),
.Y(n_777)
);

INVx3_ASAP7_75t_L g778 ( 
.A(n_622),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_636),
.B(n_664),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_671),
.B(n_674),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_597),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_659),
.B(n_210),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_564),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_683),
.B(n_210),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_677),
.B(n_653),
.Y(n_785)
);

OAI22xp5_ASAP7_75t_L g786 ( 
.A1(n_622),
.A2(n_299),
.B1(n_294),
.B2(n_279),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_651),
.B(n_214),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_657),
.B(n_230),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_576),
.B(n_487),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_660),
.B(n_214),
.Y(n_790)
);

INVx2_ASAP7_75t_SL g791 ( 
.A(n_654),
.Y(n_791)
);

INVxp67_ASAP7_75t_L g792 ( 
.A(n_632),
.Y(n_792)
);

BUFx3_ASAP7_75t_L g793 ( 
.A(n_588),
.Y(n_793)
);

OAI22xp5_ASAP7_75t_L g794 ( 
.A1(n_630),
.A2(n_272),
.B1(n_268),
.B2(n_263),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_602),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_558),
.B(n_572),
.Y(n_796)
);

BUFx6f_ASAP7_75t_L g797 ( 
.A(n_547),
.Y(n_797)
);

A2O1A1Ixp33_ASAP7_75t_L g798 ( 
.A1(n_645),
.A2(n_325),
.B(n_232),
.C(n_246),
.Y(n_798)
);

INVx2_ASAP7_75t_SL g799 ( 
.A(n_601),
.Y(n_799)
);

AND2x4_ASAP7_75t_L g800 ( 
.A(n_663),
.B(n_666),
.Y(n_800)
);

NAND2x1p5_ASAP7_75t_L g801 ( 
.A(n_558),
.B(n_244),
.Y(n_801)
);

INVx2_ASAP7_75t_SL g802 ( 
.A(n_601),
.Y(n_802)
);

INVx2_ASAP7_75t_SL g803 ( 
.A(n_601),
.Y(n_803)
);

BUFx8_ASAP7_75t_L g804 ( 
.A(n_605),
.Y(n_804)
);

NOR2x1p5_ASAP7_75t_L g805 ( 
.A(n_615),
.B(n_358),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_685),
.Y(n_806)
);

INVx2_ASAP7_75t_SL g807 ( 
.A(n_615),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_564),
.B(n_356),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_602),
.Y(n_809)
);

INVxp67_ASAP7_75t_SL g810 ( 
.A(n_547),
.Y(n_810)
);

OAI22xp5_ASAP7_75t_SL g811 ( 
.A1(n_554),
.A2(n_323),
.B1(n_353),
.B2(n_361),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_645),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_606),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_656),
.B(n_356),
.Y(n_814)
);

AOI22xp33_ASAP7_75t_L g815 ( 
.A1(n_585),
.A2(n_323),
.B1(n_361),
.B2(n_339),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_657),
.B(n_252),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_620),
.B(n_470),
.Y(n_817)
);

NOR2x1p5_ASAP7_75t_L g818 ( 
.A(n_643),
.B(n_359),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_647),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_585),
.B(n_647),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_661),
.B(n_253),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_684),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_585),
.B(n_363),
.Y(n_823)
);

INVxp67_ASAP7_75t_L g824 ( 
.A(n_667),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_661),
.B(n_312),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_620),
.B(n_470),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_620),
.B(n_624),
.Y(n_827)
);

NAND2xp33_ASAP7_75t_L g828 ( 
.A(n_547),
.B(n_235),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_672),
.B(n_313),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_624),
.B(n_472),
.Y(n_830)
);

INVx8_ASAP7_75t_L g831 ( 
.A(n_547),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_672),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_673),
.B(n_318),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_L g834 ( 
.A(n_764),
.B(n_754),
.Y(n_834)
);

CKINVDCx20_ASAP7_75t_R g835 ( 
.A(n_713),
.Y(n_835)
);

NOR2x1p5_ASAP7_75t_L g836 ( 
.A(n_768),
.B(n_245),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_717),
.Y(n_837)
);

INVx6_ASAP7_75t_L g838 ( 
.A(n_804),
.Y(n_838)
);

BUFx4f_ASAP7_75t_L g839 ( 
.A(n_751),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_712),
.B(n_607),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_696),
.B(n_363),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_806),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_696),
.B(n_607),
.Y(n_843)
);

OAI22xp5_ASAP7_75t_L g844 ( 
.A1(n_815),
.A2(n_670),
.B1(n_259),
.B2(n_341),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_696),
.B(n_612),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_696),
.B(n_612),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_696),
.B(n_614),
.Y(n_847)
);

HB1xp67_ASAP7_75t_L g848 ( 
.A(n_692),
.Y(n_848)
);

OAI21xp5_ASAP7_75t_L g849 ( 
.A1(n_820),
.A2(n_643),
.B(n_629),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_812),
.Y(n_850)
);

OR2x2_ASAP7_75t_L g851 ( 
.A(n_721),
.B(n_670),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_696),
.B(n_614),
.Y(n_852)
);

INVx3_ASAP7_75t_L g853 ( 
.A(n_688),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_819),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_701),
.A2(n_582),
.B(n_552),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_687),
.B(n_635),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_730),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_742),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_770),
.B(n_635),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_693),
.B(n_539),
.Y(n_860)
);

OAI22xp5_ASAP7_75t_L g861 ( 
.A1(n_815),
.A2(n_261),
.B1(n_266),
.B2(n_274),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_689),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_743),
.Y(n_863)
);

AND3x1_ASAP7_75t_L g864 ( 
.A(n_769),
.B(n_324),
.C(n_319),
.Y(n_864)
);

AND2x2_ASAP7_75t_SL g865 ( 
.A(n_784),
.B(n_570),
.Y(n_865)
);

BUFx5_ASAP7_75t_L g866 ( 
.A(n_697),
.Y(n_866)
);

AND2x6_ASAP7_75t_L g867 ( 
.A(n_820),
.B(n_624),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_705),
.Y(n_868)
);

HB1xp67_ASAP7_75t_L g869 ( 
.A(n_692),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_759),
.B(n_641),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_784),
.B(n_582),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_686),
.Y(n_872)
);

BUFx8_ASAP7_75t_L g873 ( 
.A(n_777),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_719),
.B(n_641),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_704),
.B(n_644),
.Y(n_875)
);

BUFx2_ASAP7_75t_L g876 ( 
.A(n_727),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_731),
.B(n_539),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_707),
.Y(n_878)
);

AND2x4_ASAP7_75t_L g879 ( 
.A(n_688),
.B(n_542),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_714),
.Y(n_880)
);

BUFx6f_ASAP7_75t_L g881 ( 
.A(n_751),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_690),
.Y(n_882)
);

AND2x4_ASAP7_75t_L g883 ( 
.A(n_750),
.B(n_542),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_706),
.B(n_644),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_700),
.B(n_559),
.Y(n_885)
);

AND2x4_ASAP7_75t_L g886 ( 
.A(n_765),
.B(n_513),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_731),
.B(n_282),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_758),
.B(n_673),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_822),
.Y(n_889)
);

NAND2x1_ASAP7_75t_L g890 ( 
.A(n_797),
.B(n_652),
.Y(n_890)
);

BUFx2_ASAP7_75t_L g891 ( 
.A(n_753),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_725),
.B(n_676),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_SL g893 ( 
.A(n_772),
.B(n_559),
.Y(n_893)
);

NAND3xp33_ASAP7_75t_L g894 ( 
.A(n_759),
.B(n_570),
.C(n_292),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_771),
.A2(n_652),
.B1(n_668),
.B2(n_678),
.Y(n_895)
);

INVx2_ASAP7_75t_SL g896 ( 
.A(n_791),
.Y(n_896)
);

INVx1_ASAP7_75t_SL g897 ( 
.A(n_774),
.Y(n_897)
);

OAI22xp5_ASAP7_75t_L g898 ( 
.A1(n_773),
.A2(n_776),
.B1(n_771),
.B2(n_824),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_720),
.Y(n_899)
);

INVx3_ASAP7_75t_L g900 ( 
.A(n_797),
.Y(n_900)
);

XOR2x2_ASAP7_75t_L g901 ( 
.A(n_811),
.B(n_0),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_741),
.B(n_582),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_832),
.Y(n_903)
);

NAND2x1p5_ASAP7_75t_L g904 ( 
.A(n_778),
.B(n_586),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_741),
.B(n_586),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_752),
.B(n_676),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_709),
.B(n_680),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_723),
.Y(n_908)
);

INVx3_ASAP7_75t_L g909 ( 
.A(n_831),
.Y(n_909)
);

AOI22xp33_ASAP7_75t_L g910 ( 
.A1(n_823),
.A2(n_682),
.B1(n_680),
.B2(n_335),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_729),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_711),
.B(n_682),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_783),
.Y(n_913)
);

AND2x4_ASAP7_75t_L g914 ( 
.A(n_778),
.B(n_514),
.Y(n_914)
);

BUFx3_ASAP7_75t_L g915 ( 
.A(n_793),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_787),
.B(n_289),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_800),
.B(n_559),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_726),
.Y(n_918)
);

AND2x6_ASAP7_75t_L g919 ( 
.A(n_800),
.B(n_652),
.Y(n_919)
);

AOI22xp5_ASAP7_75t_L g920 ( 
.A1(n_823),
.A2(n_678),
.B1(n_668),
.B2(n_655),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_732),
.Y(n_921)
);

BUFx2_ASAP7_75t_L g922 ( 
.A(n_722),
.Y(n_922)
);

HB1xp67_ASAP7_75t_L g923 ( 
.A(n_722),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_691),
.B(n_694),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_814),
.B(n_559),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_733),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_695),
.B(n_678),
.Y(n_927)
);

OR2x6_ASAP7_75t_L g928 ( 
.A(n_751),
.B(n_354),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_698),
.A2(n_668),
.B(n_586),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_728),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_814),
.B(n_559),
.Y(n_931)
);

BUFx6f_ASAP7_75t_L g932 ( 
.A(n_831),
.Y(n_932)
);

BUFx2_ASAP7_75t_L g933 ( 
.A(n_722),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_787),
.B(n_640),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_790),
.B(n_640),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_757),
.B(n_584),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_790),
.B(n_640),
.Y(n_937)
);

NOR2xp33_ASAP7_75t_L g938 ( 
.A(n_792),
.B(n_655),
.Y(n_938)
);

AND2x4_ASAP7_75t_L g939 ( 
.A(n_799),
.B(n_357),
.Y(n_939)
);

AOI22xp5_ASAP7_75t_L g940 ( 
.A1(n_785),
.A2(n_655),
.B1(n_238),
.B2(n_240),
.Y(n_940)
);

AOI22xp5_ASAP7_75t_L g941 ( 
.A1(n_785),
.A2(n_255),
.B1(n_256),
.B2(n_278),
.Y(n_941)
);

NOR2xp33_ASAP7_75t_L g942 ( 
.A(n_782),
.B(n_308),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_773),
.B(n_584),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_831),
.Y(n_944)
);

INVx2_ASAP7_75t_L g945 ( 
.A(n_736),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_SL g946 ( 
.A(n_802),
.B(n_337),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_756),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_782),
.B(n_584),
.Y(n_948)
);

AOI22xp33_ASAP7_75t_L g949 ( 
.A1(n_776),
.A2(n_648),
.B1(n_646),
.B2(n_639),
.Y(n_949)
);

AND2x6_ASAP7_75t_L g950 ( 
.A(n_789),
.B(n_584),
.Y(n_950)
);

INVx4_ASAP7_75t_L g951 ( 
.A(n_803),
.Y(n_951)
);

BUFx6f_ASAP7_75t_L g952 ( 
.A(n_699),
.Y(n_952)
);

INVx2_ASAP7_75t_SL g953 ( 
.A(n_805),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_740),
.Y(n_954)
);

INVx2_ASAP7_75t_SL g955 ( 
.A(n_807),
.Y(n_955)
);

BUFx12f_ASAP7_75t_SL g956 ( 
.A(n_804),
.Y(n_956)
);

HB1xp67_ASAP7_75t_L g957 ( 
.A(n_745),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_763),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_766),
.Y(n_959)
);

NOR2xp67_ASAP7_75t_L g960 ( 
.A(n_734),
.B(n_281),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_760),
.B(n_744),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_781),
.Y(n_962)
);

AOI22xp33_ASAP7_75t_L g963 ( 
.A1(n_818),
.A2(n_648),
.B1(n_646),
.B2(n_639),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_747),
.B(n_639),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_795),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_703),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_735),
.B(n_639),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_809),
.Y(n_968)
);

HB1xp67_ASAP7_75t_L g969 ( 
.A(n_749),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_813),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_779),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_779),
.Y(n_972)
);

A2O1A1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_775),
.A2(n_472),
.B(n_284),
.C(n_285),
.Y(n_973)
);

INVx5_ASAP7_75t_L g974 ( 
.A(n_698),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_780),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_796),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_780),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_817),
.Y(n_978)
);

INVxp67_ASAP7_75t_L g979 ( 
.A(n_775),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_826),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_738),
.B(n_639),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_830),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_761),
.B(n_646),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_827),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_738),
.B(n_646),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_739),
.B(n_715),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_739),
.B(n_646),
.Y(n_987)
);

AND2x6_ASAP7_75t_L g988 ( 
.A(n_716),
.B(n_648),
.Y(n_988)
);

AND2x4_ASAP7_75t_L g989 ( 
.A(n_760),
.B(n_538),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_718),
.B(n_724),
.Y(n_990)
);

INVx3_ASAP7_75t_L g991 ( 
.A(n_801),
.Y(n_991)
);

A2O1A1Ixp33_ASAP7_75t_L g992 ( 
.A1(n_755),
.A2(n_283),
.B(n_296),
.C(n_298),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_701),
.B(n_648),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_708),
.B(n_648),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_708),
.B(n_604),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_788),
.Y(n_996)
);

BUFx3_ASAP7_75t_L g997 ( 
.A(n_794),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_710),
.B(n_604),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_834),
.B(n_767),
.Y(n_999)
);

BUFx8_ASAP7_75t_SL g1000 ( 
.A(n_835),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_957),
.B(n_767),
.Y(n_1001)
);

O2A1O1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_898),
.A2(n_746),
.B(n_798),
.C(n_833),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_924),
.A2(n_710),
.B(n_810),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_L g1004 ( 
.A(n_979),
.B(n_808),
.Y(n_1004)
);

O2A1O1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_898),
.A2(n_833),
.B(n_829),
.C(n_788),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_924),
.A2(n_702),
.B(n_828),
.Y(n_1006)
);

AND2x2_ASAP7_75t_L g1007 ( 
.A(n_887),
.B(n_737),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_856),
.A2(n_801),
.B(n_662),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_857),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_851),
.B(n_786),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_858),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_877),
.B(n_302),
.Y(n_1012)
);

OAI21xp33_ASAP7_75t_SL g1013 ( 
.A1(n_949),
.A2(n_865),
.B(n_917),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_969),
.B(n_762),
.Y(n_1014)
);

BUFx6f_ASAP7_75t_L g1015 ( 
.A(n_932),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_881),
.B(n_816),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_942),
.B(n_829),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_856),
.A2(n_662),
.B(n_604),
.Y(n_1018)
);

NOR2xp67_ASAP7_75t_L g1019 ( 
.A(n_913),
.B(n_816),
.Y(n_1019)
);

NAND2xp33_ASAP7_75t_R g1020 ( 
.A(n_876),
.B(n_310),
.Y(n_1020)
);

AO32x1_ASAP7_75t_L g1021 ( 
.A1(n_861),
.A2(n_540),
.A3(n_538),
.B1(n_825),
.B2(n_821),
.Y(n_1021)
);

CKINVDCx6p67_ASAP7_75t_R g1022 ( 
.A(n_915),
.Y(n_1022)
);

A2O1A1Ixp33_ASAP7_75t_L g1023 ( 
.A1(n_916),
.A2(n_345),
.B(n_314),
.C(n_317),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_932),
.Y(n_1024)
);

NOR2xp33_ASAP7_75t_L g1025 ( 
.A(n_897),
.B(n_328),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_956),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_863),
.Y(n_1027)
);

O2A1O1Ixp5_ASAP7_75t_SL g1028 ( 
.A1(n_925),
.A2(n_352),
.B(n_349),
.C(n_340),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_860),
.B(n_538),
.Y(n_1029)
);

BUFx2_ASAP7_75t_L g1030 ( 
.A(n_891),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_888),
.A2(n_662),
.B(n_604),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_848),
.B(n_331),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_911),
.B(n_540),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_873),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_888),
.A2(n_662),
.B(n_604),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_869),
.B(n_333),
.Y(n_1036)
);

OAI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_986),
.A2(n_662),
.B(n_540),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_837),
.Y(n_1038)
);

INVx2_ASAP7_75t_SL g1039 ( 
.A(n_955),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_990),
.A2(n_484),
.B(n_347),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_921),
.B(n_332),
.Y(n_1041)
);

AO21x2_ASAP7_75t_L g1042 ( 
.A1(n_849),
.A2(n_338),
.B(n_351),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_997),
.B(n_342),
.Y(n_1043)
);

HB1xp67_ASAP7_75t_L g1044 ( 
.A(n_923),
.Y(n_1044)
);

AOI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_961),
.A2(n_853),
.B1(n_919),
.B2(n_905),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_844),
.B(n_926),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_862),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_878),
.Y(n_1048)
);

OAI21x1_ASAP7_75t_L g1049 ( 
.A1(n_855),
.A2(n_68),
.B(n_184),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_880),
.Y(n_1050)
);

BUFx12f_ASAP7_75t_L g1051 ( 
.A(n_873),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_844),
.B(n_4),
.Y(n_1052)
);

BUFx2_ASAP7_75t_L g1053 ( 
.A(n_922),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_899),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_L g1055 ( 
.A(n_954),
.B(n_8),
.Y(n_1055)
);

BUFx3_ASAP7_75t_L g1056 ( 
.A(n_881),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_908),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_902),
.B(n_8),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_871),
.B(n_11),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_934),
.B(n_11),
.Y(n_1060)
);

BUFx6f_ASAP7_75t_L g1061 ( 
.A(n_881),
.Y(n_1061)
);

HB1xp67_ASAP7_75t_L g1062 ( 
.A(n_879),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_918),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_935),
.B(n_12),
.Y(n_1064)
);

O2A1O1Ixp5_ASAP7_75t_SL g1065 ( 
.A1(n_931),
.A2(n_14),
.B(n_16),
.C(n_18),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_868),
.B(n_16),
.Y(n_1066)
);

INVx1_ASAP7_75t_SL g1067 ( 
.A(n_933),
.Y(n_1067)
);

HB1xp67_ASAP7_75t_L g1068 ( 
.A(n_879),
.Y(n_1068)
);

OAI21xp33_ASAP7_75t_L g1069 ( 
.A1(n_946),
.A2(n_23),
.B(n_27),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_906),
.A2(n_484),
.B(n_658),
.Y(n_1070)
);

BUFx4f_ASAP7_75t_SL g1071 ( 
.A(n_953),
.Y(n_1071)
);

BUFx2_ASAP7_75t_L g1072 ( 
.A(n_914),
.Y(n_1072)
);

A2O1A1Ixp33_ASAP7_75t_L g1073 ( 
.A1(n_937),
.A2(n_27),
.B(n_35),
.C(n_36),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_946),
.B(n_90),
.Y(n_1074)
);

INVx5_ASAP7_75t_L g1075 ( 
.A(n_867),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_930),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_842),
.Y(n_1077)
);

INVx4_ASAP7_75t_L g1078 ( 
.A(n_909),
.Y(n_1078)
);

O2A1O1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_859),
.A2(n_35),
.B(n_37),
.C(n_40),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_850),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_978),
.B(n_37),
.Y(n_1081)
);

A2O1A1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_972),
.A2(n_41),
.B(n_42),
.C(n_43),
.Y(n_1082)
);

INVx2_ASAP7_75t_L g1083 ( 
.A(n_945),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_906),
.A2(n_658),
.B(n_116),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_907),
.A2(n_112),
.B(n_176),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_854),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_889),
.Y(n_1087)
);

BUFx3_ASAP7_75t_L g1088 ( 
.A(n_838),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_886),
.B(n_44),
.Y(n_1089)
);

HB1xp67_ASAP7_75t_L g1090 ( 
.A(n_984),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_886),
.B(n_45),
.Y(n_1091)
);

NOR3xp33_ASAP7_75t_L g1092 ( 
.A(n_861),
.B(n_47),
.C(n_48),
.Y(n_1092)
);

NAND2x1p5_ASAP7_75t_L g1093 ( 
.A(n_944),
.B(n_124),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_SL g1094 ( 
.A(n_839),
.B(n_108),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_980),
.B(n_47),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_907),
.A2(n_136),
.B(n_169),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_912),
.A2(n_97),
.B(n_168),
.Y(n_1097)
);

A2O1A1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_975),
.A2(n_48),
.B(n_53),
.C(n_54),
.Y(n_1098)
);

INVxp67_ASAP7_75t_L g1099 ( 
.A(n_872),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_912),
.A2(n_138),
.B(n_166),
.Y(n_1100)
);

OR2x2_ASAP7_75t_L g1101 ( 
.A(n_882),
.B(n_55),
.Y(n_1101)
);

AOI22xp33_ASAP7_75t_L g1102 ( 
.A1(n_919),
.A2(n_58),
.B1(n_61),
.B2(n_62),
.Y(n_1102)
);

INVx3_ASAP7_75t_L g1103 ( 
.A(n_952),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_982),
.B(n_58),
.Y(n_1104)
);

BUFx2_ASAP7_75t_L g1105 ( 
.A(n_914),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_927),
.A2(n_82),
.B(n_137),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_947),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_958),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_939),
.B(n_142),
.Y(n_1109)
);

OR2x6_ASAP7_75t_SL g1110 ( 
.A(n_966),
.B(n_148),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_959),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_927),
.A2(n_156),
.B(n_157),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_843),
.A2(n_164),
.B(n_165),
.Y(n_1113)
);

AND2x2_ASAP7_75t_L g1114 ( 
.A(n_939),
.B(n_177),
.Y(n_1114)
);

INVx6_ASAP7_75t_L g1115 ( 
.A(n_951),
.Y(n_1115)
);

BUFx6f_ASAP7_75t_L g1116 ( 
.A(n_944),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_843),
.A2(n_852),
.B(n_847),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_845),
.A2(n_852),
.B(n_847),
.Y(n_1118)
);

OAI21x1_ASAP7_75t_L g1119 ( 
.A1(n_993),
.A2(n_994),
.B(n_846),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_845),
.A2(n_846),
.B(n_981),
.Y(n_1120)
);

INVx1_ASAP7_75t_SL g1121 ( 
.A(n_896),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_900),
.Y(n_1122)
);

NOR2xp33_ASAP7_75t_L g1123 ( 
.A(n_977),
.B(n_971),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_981),
.A2(n_985),
.B(n_964),
.Y(n_1124)
);

BUFx2_ASAP7_75t_L g1125 ( 
.A(n_989),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_985),
.A2(n_875),
.B(n_884),
.Y(n_1126)
);

AOI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_919),
.A2(n_960),
.B1(n_989),
.B2(n_938),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_883),
.B(n_836),
.Y(n_1128)
);

INVx3_ASAP7_75t_L g1129 ( 
.A(n_952),
.Y(n_1129)
);

BUFx2_ASAP7_75t_L g1130 ( 
.A(n_864),
.Y(n_1130)
);

NOR3xp33_ASAP7_75t_L g1131 ( 
.A(n_973),
.B(n_894),
.C(n_841),
.Y(n_1131)
);

NOR2xp33_ASAP7_75t_L g1132 ( 
.A(n_870),
.B(n_883),
.Y(n_1132)
);

A2O1A1Ixp33_ASAP7_75t_SL g1133 ( 
.A1(n_849),
.A2(n_929),
.B(n_910),
.C(n_991),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_1006),
.A2(n_983),
.B(n_967),
.Y(n_1134)
);

BUFx6f_ASAP7_75t_L g1135 ( 
.A(n_1061),
.Y(n_1135)
);

BUFx3_ASAP7_75t_L g1136 ( 
.A(n_1030),
.Y(n_1136)
);

OAI21x1_ASAP7_75t_L g1137 ( 
.A1(n_1119),
.A2(n_929),
.B(n_874),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1003),
.A2(n_986),
.B(n_840),
.Y(n_1138)
);

NOR2xp67_ASAP7_75t_L g1139 ( 
.A(n_1039),
.B(n_951),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_999),
.B(n_884),
.Y(n_1140)
);

AO22x2_ASAP7_75t_L g1141 ( 
.A1(n_1092),
.A2(n_901),
.B1(n_943),
.B2(n_874),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_1120),
.A2(n_993),
.B(n_994),
.Y(n_1142)
);

AND2x4_ASAP7_75t_L g1143 ( 
.A(n_1128),
.B(n_903),
.Y(n_1143)
);

OA21x2_ASAP7_75t_L g1144 ( 
.A1(n_1037),
.A2(n_992),
.B(n_948),
.Y(n_1144)
);

NOR4xp25_ASAP7_75t_L g1145 ( 
.A(n_1069),
.B(n_1052),
.C(n_1073),
.D(n_1079),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1046),
.B(n_1132),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1126),
.A2(n_974),
.B(n_943),
.Y(n_1147)
);

NAND3xp33_ASAP7_75t_L g1148 ( 
.A(n_1017),
.B(n_941),
.C(n_940),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1046),
.B(n_919),
.Y(n_1149)
);

OAI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1017),
.A2(n_895),
.B(n_892),
.Y(n_1150)
);

INVx3_ASAP7_75t_L g1151 ( 
.A(n_1116),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1033),
.Y(n_1152)
);

INVxp67_ASAP7_75t_L g1153 ( 
.A(n_1044),
.Y(n_1153)
);

OAI22x1_ASAP7_75t_L g1154 ( 
.A1(n_1052),
.A2(n_974),
.B1(n_996),
.B2(n_893),
.Y(n_1154)
);

AO31x2_ASAP7_75t_L g1155 ( 
.A1(n_1124),
.A2(n_987),
.A3(n_998),
.B(n_995),
.Y(n_1155)
);

AO31x2_ASAP7_75t_L g1156 ( 
.A1(n_1117),
.A2(n_1118),
.A3(n_1008),
.B(n_1058),
.Y(n_1156)
);

CKINVDCx16_ASAP7_75t_R g1157 ( 
.A(n_1051),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_1009),
.Y(n_1158)
);

NAND3x1_ASAP7_75t_L g1159 ( 
.A(n_1092),
.B(n_838),
.C(n_839),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1049),
.A2(n_998),
.B(n_995),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_1018),
.A2(n_1035),
.B(n_1031),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1084),
.A2(n_936),
.B(n_920),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1038),
.Y(n_1163)
);

BUFx3_ASAP7_75t_L g1164 ( 
.A(n_1022),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_1004),
.B(n_1043),
.Y(n_1165)
);

AO32x2_ASAP7_75t_L g1166 ( 
.A1(n_1021),
.A2(n_867),
.A3(n_950),
.B1(n_866),
.B2(n_963),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1090),
.B(n_976),
.Y(n_1167)
);

O2A1O1Ixp33_ASAP7_75t_SL g1168 ( 
.A1(n_1133),
.A2(n_885),
.B(n_890),
.C(n_962),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_1000),
.Y(n_1169)
);

AO31x2_ASAP7_75t_L g1170 ( 
.A1(n_1059),
.A2(n_970),
.A3(n_968),
.B(n_965),
.Y(n_1170)
);

O2A1O1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_1007),
.A2(n_928),
.B(n_904),
.C(n_867),
.Y(n_1171)
);

AO21x1_ASAP7_75t_L g1172 ( 
.A1(n_1060),
.A2(n_904),
.B(n_950),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_SL g1173 ( 
.A(n_1043),
.B(n_1004),
.Y(n_1173)
);

NAND3xp33_ASAP7_75t_SL g1174 ( 
.A(n_1130),
.B(n_928),
.C(n_866),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_L g1175 ( 
.A1(n_1005),
.A2(n_866),
.B(n_950),
.Y(n_1175)
);

AOI21x1_ASAP7_75t_L g1176 ( 
.A1(n_1064),
.A2(n_950),
.B(n_928),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1075),
.A2(n_1029),
.B(n_1131),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1010),
.B(n_988),
.Y(n_1178)
);

OAI21x1_ASAP7_75t_SL g1179 ( 
.A1(n_1085),
.A2(n_988),
.B(n_1096),
.Y(n_1179)
);

NOR2xp33_ASAP7_75t_SL g1180 ( 
.A(n_1034),
.B(n_988),
.Y(n_1180)
);

OAI21x1_ASAP7_75t_L g1181 ( 
.A1(n_1070),
.A2(n_988),
.B(n_1028),
.Y(n_1181)
);

OR2x2_ASAP7_75t_L g1182 ( 
.A(n_1001),
.B(n_1067),
.Y(n_1182)
);

AOI21xp33_ASAP7_75t_L g1183 ( 
.A1(n_1010),
.A2(n_1025),
.B(n_1020),
.Y(n_1183)
);

HB1xp67_ASAP7_75t_L g1184 ( 
.A(n_1044),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1097),
.A2(n_1100),
.B(n_1113),
.Y(n_1185)
);

BUFx12f_ASAP7_75t_L g1186 ( 
.A(n_1026),
.Y(n_1186)
);

OAI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1106),
.A2(n_1112),
.B(n_1002),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_SL g1188 ( 
.A(n_1088),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1077),
.Y(n_1189)
);

AO31x2_ASAP7_75t_L g1190 ( 
.A1(n_1123),
.A2(n_1021),
.A3(n_1082),
.B(n_1098),
.Y(n_1190)
);

OAI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1123),
.A2(n_1045),
.B(n_1131),
.Y(n_1191)
);

NAND3x1_ASAP7_75t_L g1192 ( 
.A(n_1089),
.B(n_1091),
.C(n_1066),
.Y(n_1192)
);

BUFx10_ASAP7_75t_L g1193 ( 
.A(n_1032),
.Y(n_1193)
);

AO31x2_ASAP7_75t_L g1194 ( 
.A1(n_1021),
.A2(n_1055),
.A3(n_1104),
.B(n_1081),
.Y(n_1194)
);

OAI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1127),
.A2(n_1041),
.B(n_1040),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1055),
.B(n_1011),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1080),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_1019),
.B(n_1072),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1027),
.B(n_1086),
.Y(n_1199)
);

NOR2xp33_ASAP7_75t_L g1200 ( 
.A(n_1025),
.B(n_1014),
.Y(n_1200)
);

O2A1O1Ixp5_ASAP7_75t_L g1201 ( 
.A1(n_1095),
.A2(n_1074),
.B(n_1012),
.C(n_1023),
.Y(n_1201)
);

INVx4_ASAP7_75t_L g1202 ( 
.A(n_1015),
.Y(n_1202)
);

AO32x2_ASAP7_75t_L g1203 ( 
.A1(n_1065),
.A2(n_1042),
.A3(n_1078),
.B1(n_1079),
.B2(n_1102),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1075),
.A2(n_1042),
.B(n_1129),
.Y(n_1204)
);

BUFx3_ASAP7_75t_L g1205 ( 
.A(n_1056),
.Y(n_1205)
);

AOI21xp33_ASAP7_75t_L g1206 ( 
.A1(n_1020),
.A2(n_1032),
.B(n_1036),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1075),
.A2(n_1129),
.B(n_1103),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1099),
.B(n_1125),
.Y(n_1208)
);

AO32x2_ASAP7_75t_L g1209 ( 
.A1(n_1102),
.A2(n_1099),
.A3(n_1101),
.B1(n_1087),
.B2(n_1093),
.Y(n_1209)
);

BUFx6f_ASAP7_75t_L g1210 ( 
.A(n_1061),
.Y(n_1210)
);

INVx6_ASAP7_75t_L g1211 ( 
.A(n_1061),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1047),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1062),
.B(n_1068),
.Y(n_1213)
);

BUFx12f_ASAP7_75t_L g1214 ( 
.A(n_1053),
.Y(n_1214)
);

INVx2_ASAP7_75t_SL g1215 ( 
.A(n_1121),
.Y(n_1215)
);

INVx2_ASAP7_75t_SL g1216 ( 
.A(n_1071),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1048),
.Y(n_1217)
);

AND2x4_ASAP7_75t_L g1218 ( 
.A(n_1062),
.B(n_1068),
.Y(n_1218)
);

AOI221xp5_ASAP7_75t_L g1219 ( 
.A1(n_1105),
.A2(n_1109),
.B1(n_1114),
.B2(n_1083),
.C(n_1063),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1050),
.B(n_1076),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1054),
.Y(n_1221)
);

AND2x4_ASAP7_75t_L g1222 ( 
.A(n_1016),
.B(n_1024),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1057),
.A2(n_1107),
.B(n_1111),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1108),
.Y(n_1224)
);

INVx2_ASAP7_75t_SL g1225 ( 
.A(n_1071),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_SL g1226 ( 
.A(n_1094),
.B(n_1015),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1016),
.A2(n_1116),
.B(n_1122),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1122),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1122),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1122),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1115),
.B(n_1116),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1115),
.A2(n_1006),
.B(n_924),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_SL g1233 ( 
.A(n_1115),
.B(n_1110),
.Y(n_1233)
);

OR2x2_ASAP7_75t_L g1234 ( 
.A(n_1001),
.B(n_721),
.Y(n_1234)
);

OAI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1017),
.A2(n_898),
.B(n_1013),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_999),
.B(n_877),
.Y(n_1236)
);

INVx3_ASAP7_75t_L g1237 ( 
.A(n_1116),
.Y(n_1237)
);

AOI221x1_ASAP7_75t_L g1238 ( 
.A1(n_1092),
.A2(n_898),
.B1(n_1052),
.B2(n_1131),
.C(n_1060),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_999),
.B(n_877),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1006),
.A2(n_924),
.B(n_1003),
.Y(n_1240)
);

OAI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1017),
.A2(n_898),
.B1(n_999),
.B2(n_1046),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_999),
.B(n_877),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1006),
.A2(n_924),
.B(n_1003),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1007),
.B(n_693),
.Y(n_1244)
);

NOR2xp67_ASAP7_75t_SL g1245 ( 
.A(n_1075),
.B(n_777),
.Y(n_1245)
);

INVx4_ASAP7_75t_L g1246 ( 
.A(n_1015),
.Y(n_1246)
);

AO32x2_ASAP7_75t_L g1247 ( 
.A1(n_1021),
.A2(n_898),
.A3(n_844),
.B1(n_861),
.B2(n_551),
.Y(n_1247)
);

O2A1O1Ixp33_ASAP7_75t_SL g1248 ( 
.A1(n_1133),
.A2(n_898),
.B(n_1073),
.C(n_1017),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1007),
.B(n_693),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1017),
.A2(n_898),
.B1(n_999),
.B2(n_1046),
.Y(n_1250)
);

AO32x2_ASAP7_75t_L g1251 ( 
.A1(n_1021),
.A2(n_898),
.A3(n_844),
.B1(n_861),
.B2(n_551),
.Y(n_1251)
);

BUFx3_ASAP7_75t_L g1252 ( 
.A(n_1030),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1006),
.A2(n_924),
.B(n_1003),
.Y(n_1253)
);

NAND3x1_ASAP7_75t_L g1254 ( 
.A(n_1052),
.B(n_1092),
.C(n_748),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1006),
.A2(n_924),
.B(n_1003),
.Y(n_1255)
);

BUFx2_ASAP7_75t_SL g1256 ( 
.A(n_1056),
.Y(n_1256)
);

AOI21xp33_ASAP7_75t_L g1257 ( 
.A1(n_1017),
.A2(n_942),
.B(n_748),
.Y(n_1257)
);

AND2x2_ASAP7_75t_SL g1258 ( 
.A(n_1052),
.B(n_815),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_1061),
.Y(n_1259)
);

NOR4xp25_ASAP7_75t_L g1260 ( 
.A(n_1069),
.B(n_1052),
.C(n_942),
.D(n_1073),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1119),
.A2(n_1120),
.B(n_1124),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1119),
.A2(n_1120),
.B(n_1124),
.Y(n_1262)
);

A2O1A1Ixp33_ASAP7_75t_L g1263 ( 
.A1(n_1017),
.A2(n_771),
.B(n_942),
.C(n_999),
.Y(n_1263)
);

OAI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1017),
.A2(n_898),
.B(n_1013),
.Y(n_1264)
);

OAI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1017),
.A2(n_898),
.B(n_1013),
.Y(n_1265)
);

A2O1A1Ixp33_ASAP7_75t_L g1266 ( 
.A1(n_1017),
.A2(n_771),
.B(n_942),
.C(n_999),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1090),
.Y(n_1267)
);

O2A1O1Ixp5_ASAP7_75t_L g1268 ( 
.A1(n_1017),
.A2(n_942),
.B(n_1060),
.C(n_1059),
.Y(n_1268)
);

O2A1O1Ixp33_ASAP7_75t_L g1269 ( 
.A1(n_999),
.A2(n_942),
.B(n_748),
.C(n_764),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1119),
.A2(n_1120),
.B(n_1124),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1033),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_1000),
.Y(n_1272)
);

O2A1O1Ixp33_ASAP7_75t_L g1273 ( 
.A1(n_999),
.A2(n_942),
.B(n_748),
.C(n_764),
.Y(n_1273)
);

AO31x2_ASAP7_75t_L g1274 ( 
.A1(n_1006),
.A2(n_992),
.A3(n_820),
.B(n_898),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_SL g1275 ( 
.A1(n_1017),
.A2(n_898),
.B(n_924),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_999),
.B(n_877),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1006),
.A2(n_924),
.B(n_1003),
.Y(n_1277)
);

NAND3xp33_ASAP7_75t_SL g1278 ( 
.A(n_1017),
.B(n_942),
.C(n_748),
.Y(n_1278)
);

INVxp67_ASAP7_75t_L g1279 ( 
.A(n_1184),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1244),
.B(n_1249),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1199),
.Y(n_1281)
);

BUFx12f_ASAP7_75t_L g1282 ( 
.A(n_1169),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1161),
.A2(n_1262),
.B(n_1261),
.Y(n_1283)
);

OAI222xp33_ASAP7_75t_L g1284 ( 
.A1(n_1241),
.A2(n_1250),
.B1(n_1269),
.B2(n_1273),
.C1(n_1165),
.C2(n_1173),
.Y(n_1284)
);

AOI211xp5_ASAP7_75t_L g1285 ( 
.A1(n_1257),
.A2(n_1278),
.B(n_1183),
.C(n_1263),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1258),
.A2(n_1141),
.B1(n_1264),
.B2(n_1265),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1270),
.A2(n_1160),
.B(n_1147),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1266),
.A2(n_1254),
.B1(n_1200),
.B2(n_1276),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_L g1289 ( 
.A1(n_1232),
.A2(n_1243),
.B(n_1240),
.Y(n_1289)
);

OR2x6_ASAP7_75t_L g1290 ( 
.A(n_1171),
.B(n_1275),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1242),
.B(n_1146),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1253),
.A2(n_1277),
.B(n_1255),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1141),
.A2(n_1235),
.B1(n_1148),
.B2(n_1206),
.Y(n_1293)
);

NOR2xp33_ASAP7_75t_L g1294 ( 
.A(n_1196),
.B(n_1140),
.Y(n_1294)
);

BUFx2_ASAP7_75t_L g1295 ( 
.A(n_1136),
.Y(n_1295)
);

INVx2_ASAP7_75t_SL g1296 ( 
.A(n_1205),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1137),
.A2(n_1162),
.B(n_1134),
.Y(n_1297)
);

HB1xp67_ASAP7_75t_L g1298 ( 
.A(n_1215),
.Y(n_1298)
);

OR2x2_ASAP7_75t_L g1299 ( 
.A(n_1182),
.B(n_1234),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1175),
.A2(n_1185),
.B(n_1142),
.Y(n_1300)
);

OAI21x1_ASAP7_75t_L g1301 ( 
.A1(n_1138),
.A2(n_1187),
.B(n_1181),
.Y(n_1301)
);

OAI222xp33_ASAP7_75t_L g1302 ( 
.A1(n_1149),
.A2(n_1178),
.B1(n_1208),
.B2(n_1153),
.C1(n_1198),
.C2(n_1167),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1191),
.A2(n_1150),
.B1(n_1233),
.B2(n_1193),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1193),
.A2(n_1219),
.B1(n_1174),
.B2(n_1271),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1189),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1204),
.A2(n_1179),
.B(n_1177),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_SL g1307 ( 
.A1(n_1226),
.A2(n_1192),
.B1(n_1180),
.B2(n_1195),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_L g1308 ( 
.A(n_1213),
.B(n_1218),
.Y(n_1308)
);

OA21x2_ASAP7_75t_L g1309 ( 
.A1(n_1238),
.A2(n_1268),
.B(n_1172),
.Y(n_1309)
);

BUFx6f_ASAP7_75t_L g1310 ( 
.A(n_1135),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1218),
.B(n_1267),
.Y(n_1311)
);

OAI22xp5_ASAP7_75t_L g1312 ( 
.A1(n_1143),
.A2(n_1159),
.B1(n_1139),
.B2(n_1158),
.Y(n_1312)
);

O2A1O1Ixp33_ASAP7_75t_SL g1313 ( 
.A1(n_1152),
.A2(n_1228),
.B(n_1229),
.C(n_1230),
.Y(n_1313)
);

OAI211xp5_ASAP7_75t_L g1314 ( 
.A1(n_1260),
.A2(n_1145),
.B(n_1248),
.C(n_1197),
.Y(n_1314)
);

OAI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1143),
.A2(n_1252),
.B1(n_1197),
.B2(n_1222),
.Y(n_1315)
);

AND2x4_ASAP7_75t_L g1316 ( 
.A(n_1222),
.B(n_1227),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1224),
.Y(n_1317)
);

AO31x2_ASAP7_75t_L g1318 ( 
.A1(n_1154),
.A2(n_1247),
.A3(n_1251),
.B(n_1166),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1223),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1224),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1144),
.A2(n_1207),
.B(n_1201),
.Y(n_1321)
);

OAI21x1_ASAP7_75t_L g1322 ( 
.A1(n_1220),
.A2(n_1237),
.B(n_1151),
.Y(n_1322)
);

AO31x2_ASAP7_75t_L g1323 ( 
.A1(n_1247),
.A2(n_1251),
.A3(n_1166),
.B(n_1156),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1151),
.A2(n_1237),
.B(n_1217),
.Y(n_1324)
);

OAI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1168),
.A2(n_1221),
.B(n_1212),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_SL g1326 ( 
.A1(n_1231),
.A2(n_1202),
.B(n_1246),
.Y(n_1326)
);

BUFx2_ASAP7_75t_L g1327 ( 
.A(n_1214),
.Y(n_1327)
);

OA21x2_ASAP7_75t_L g1328 ( 
.A1(n_1166),
.A2(n_1156),
.B(n_1247),
.Y(n_1328)
);

OA21x2_ASAP7_75t_L g1329 ( 
.A1(n_1251),
.A2(n_1194),
.B(n_1274),
.Y(n_1329)
);

AOI221x1_ASAP7_75t_L g1330 ( 
.A1(n_1203),
.A2(n_1209),
.B1(n_1194),
.B2(n_1190),
.C(n_1246),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1155),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1245),
.A2(n_1188),
.B1(n_1186),
.B2(n_1164),
.Y(n_1332)
);

NAND3xp33_ASAP7_75t_L g1333 ( 
.A(n_1272),
.B(n_1225),
.C(n_1216),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1170),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1190),
.Y(n_1335)
);

OAI21xp5_ASAP7_75t_SL g1336 ( 
.A1(n_1209),
.A2(n_1157),
.B(n_1203),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1188),
.A2(n_1210),
.B1(n_1259),
.B2(n_1211),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1190),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1209),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1274),
.Y(n_1340)
);

OAI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1203),
.A2(n_1194),
.B(n_1211),
.Y(n_1341)
);

INVx5_ASAP7_75t_L g1342 ( 
.A(n_1135),
.Y(n_1342)
);

INVx6_ASAP7_75t_L g1343 ( 
.A(n_1214),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1244),
.B(n_1249),
.Y(n_1344)
);

OAI221xp5_ASAP7_75t_L g1345 ( 
.A1(n_1257),
.A2(n_1263),
.B1(n_1266),
.B2(n_1165),
.C(n_1278),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1199),
.Y(n_1346)
);

AO21x2_ASAP7_75t_L g1347 ( 
.A1(n_1134),
.A2(n_1243),
.B(n_1240),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1161),
.A2(n_1262),
.B(n_1261),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1163),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_L g1350 ( 
.A1(n_1161),
.A2(n_1262),
.B(n_1261),
.Y(n_1350)
);

OAI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1257),
.A2(n_1266),
.B(n_1263),
.Y(n_1351)
);

OR2x2_ASAP7_75t_L g1352 ( 
.A(n_1182),
.B(n_1234),
.Y(n_1352)
);

INVx4_ASAP7_75t_L g1353 ( 
.A(n_1135),
.Y(n_1353)
);

INVx1_ASAP7_75t_SL g1354 ( 
.A(n_1136),
.Y(n_1354)
);

AOI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1258),
.A2(n_1278),
.B1(n_1257),
.B2(n_1241),
.Y(n_1355)
);

AO21x2_ASAP7_75t_L g1356 ( 
.A1(n_1134),
.A2(n_1243),
.B(n_1240),
.Y(n_1356)
);

INVx2_ASAP7_75t_SL g1357 ( 
.A(n_1205),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1163),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1258),
.A2(n_1278),
.B1(n_1257),
.B2(n_1241),
.Y(n_1359)
);

AO32x2_ASAP7_75t_L g1360 ( 
.A1(n_1241),
.A2(n_1250),
.A3(n_898),
.B1(n_1251),
.B2(n_1247),
.Y(n_1360)
);

OAI21xp5_ASAP7_75t_L g1361 ( 
.A1(n_1257),
.A2(n_1266),
.B(n_1263),
.Y(n_1361)
);

OAI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1257),
.A2(n_1266),
.B(n_1263),
.Y(n_1362)
);

OAI21xp5_ASAP7_75t_L g1363 ( 
.A1(n_1257),
.A2(n_1266),
.B(n_1263),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1161),
.A2(n_1262),
.B(n_1261),
.Y(n_1364)
);

OA21x2_ASAP7_75t_L g1365 ( 
.A1(n_1240),
.A2(n_1253),
.B(n_1243),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1161),
.A2(n_1262),
.B(n_1261),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1163),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1161),
.A2(n_1262),
.B(n_1261),
.Y(n_1368)
);

OAI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1257),
.A2(n_1266),
.B(n_1263),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1161),
.A2(n_1262),
.B(n_1261),
.Y(n_1370)
);

NOR2xp33_ASAP7_75t_L g1371 ( 
.A(n_1257),
.B(n_1278),
.Y(n_1371)
);

OAI21xp5_ASAP7_75t_L g1372 ( 
.A1(n_1257),
.A2(n_1266),
.B(n_1263),
.Y(n_1372)
);

AND2x4_ASAP7_75t_L g1373 ( 
.A(n_1222),
.B(n_1218),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_SL g1374 ( 
.A1(n_1258),
.A2(n_1165),
.B1(n_374),
.B2(n_384),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1199),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1258),
.A2(n_1278),
.B1(n_1257),
.B2(n_1241),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_L g1377 ( 
.A(n_1257),
.B(n_1278),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1161),
.A2(n_1262),
.B(n_1261),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1163),
.Y(n_1379)
);

NAND3xp33_ASAP7_75t_L g1380 ( 
.A(n_1257),
.B(n_1266),
.C(n_1263),
.Y(n_1380)
);

AOI21x1_ASAP7_75t_L g1381 ( 
.A1(n_1176),
.A2(n_1204),
.B(n_1177),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1236),
.B(n_1239),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1258),
.A2(n_1278),
.B1(n_1257),
.B2(n_1241),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_1169),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1161),
.A2(n_1262),
.B(n_1261),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1236),
.B(n_1239),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1161),
.A2(n_1262),
.B(n_1261),
.Y(n_1387)
);

OAI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1257),
.A2(n_1266),
.B(n_1263),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1236),
.B(n_1239),
.Y(n_1389)
);

OAI21x1_ASAP7_75t_L g1390 ( 
.A1(n_1161),
.A2(n_1262),
.B(n_1261),
.Y(n_1390)
);

INVx6_ASAP7_75t_L g1391 ( 
.A(n_1214),
.Y(n_1391)
);

OAI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1263),
.A2(n_1266),
.B1(n_1165),
.B2(n_1258),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_L g1393 ( 
.A(n_1257),
.B(n_1278),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1161),
.A2(n_1262),
.B(n_1261),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1161),
.A2(n_1262),
.B(n_1261),
.Y(n_1395)
);

CKINVDCx8_ASAP7_75t_R g1396 ( 
.A(n_1256),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1199),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_1169),
.Y(n_1398)
);

NOR2xp67_ASAP7_75t_L g1399 ( 
.A(n_1215),
.B(n_913),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1161),
.A2(n_1262),
.B(n_1261),
.Y(n_1400)
);

INVx2_ASAP7_75t_SL g1401 ( 
.A(n_1205),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1199),
.Y(n_1402)
);

OAI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1257),
.A2(n_1266),
.B(n_1263),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1236),
.B(n_1239),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1161),
.A2(n_1262),
.B(n_1261),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1199),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1258),
.A2(n_1278),
.B1(n_1257),
.B2(n_1241),
.Y(n_1407)
);

OA21x2_ASAP7_75t_L g1408 ( 
.A1(n_1330),
.A2(n_1301),
.B(n_1292),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_SL g1409 ( 
.A1(n_1345),
.A2(n_1377),
.B(n_1371),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1294),
.B(n_1291),
.Y(n_1410)
);

OR2x2_ASAP7_75t_L g1411 ( 
.A(n_1299),
.B(n_1352),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1382),
.B(n_1386),
.Y(n_1412)
);

A2O1A1Ixp33_ASAP7_75t_L g1413 ( 
.A1(n_1371),
.A2(n_1393),
.B(n_1377),
.C(n_1286),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1389),
.B(n_1404),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_1384),
.Y(n_1415)
);

AND2x4_ASAP7_75t_L g1416 ( 
.A(n_1373),
.B(n_1316),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1303),
.A2(n_1407),
.B1(n_1383),
.B2(n_1376),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1280),
.B(n_1344),
.Y(n_1418)
);

OR2x2_ASAP7_75t_L g1419 ( 
.A(n_1293),
.B(n_1392),
.Y(n_1419)
);

INVx5_ASAP7_75t_L g1420 ( 
.A(n_1290),
.Y(n_1420)
);

NAND2x1p5_ASAP7_75t_L g1421 ( 
.A(n_1316),
.B(n_1324),
.Y(n_1421)
);

O2A1O1Ixp33_ASAP7_75t_L g1422 ( 
.A1(n_1284),
.A2(n_1393),
.B(n_1288),
.C(n_1361),
.Y(n_1422)
);

INVx2_ASAP7_75t_SL g1423 ( 
.A(n_1343),
.Y(n_1423)
);

A2O1A1Ixp33_ASAP7_75t_L g1424 ( 
.A1(n_1380),
.A2(n_1285),
.B(n_1351),
.C(n_1388),
.Y(n_1424)
);

INVx2_ASAP7_75t_SL g1425 ( 
.A(n_1343),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1308),
.B(n_1311),
.Y(n_1426)
);

O2A1O1Ixp33_ASAP7_75t_L g1427 ( 
.A1(n_1362),
.A2(n_1363),
.B(n_1369),
.C(n_1372),
.Y(n_1427)
);

O2A1O1Ixp33_ASAP7_75t_L g1428 ( 
.A1(n_1403),
.A2(n_1407),
.B(n_1355),
.C(n_1359),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_L g1429 ( 
.A(n_1281),
.B(n_1346),
.Y(n_1429)
);

INVx1_ASAP7_75t_SL g1430 ( 
.A(n_1354),
.Y(n_1430)
);

NOR2xp67_ASAP7_75t_L g1431 ( 
.A(n_1333),
.B(n_1298),
.Y(n_1431)
);

OR2x2_ASAP7_75t_L g1432 ( 
.A(n_1293),
.B(n_1308),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1355),
.B(n_1383),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1307),
.A2(n_1304),
.B1(n_1312),
.B2(n_1396),
.Y(n_1434)
);

NAND2x1p5_ASAP7_75t_L g1435 ( 
.A(n_1324),
.B(n_1342),
.Y(n_1435)
);

OAI22xp5_ASAP7_75t_L g1436 ( 
.A1(n_1304),
.A2(n_1315),
.B1(n_1337),
.B2(n_1332),
.Y(n_1436)
);

OAI22xp5_ASAP7_75t_L g1437 ( 
.A1(n_1337),
.A2(n_1332),
.B1(n_1402),
.B2(n_1397),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1375),
.B(n_1406),
.Y(n_1438)
);

O2A1O1Ixp5_ASAP7_75t_L g1439 ( 
.A1(n_1314),
.A2(n_1381),
.B(n_1302),
.C(n_1331),
.Y(n_1439)
);

CKINVDCx5p33_ASAP7_75t_R g1440 ( 
.A(n_1384),
.Y(n_1440)
);

OAI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1399),
.A2(n_1279),
.B1(n_1290),
.B2(n_1295),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1317),
.B(n_1320),
.Y(n_1442)
);

OA21x2_ASAP7_75t_L g1443 ( 
.A1(n_1321),
.A2(n_1289),
.B(n_1292),
.Y(n_1443)
);

OA21x2_ASAP7_75t_L g1444 ( 
.A1(n_1300),
.A2(n_1297),
.B(n_1341),
.Y(n_1444)
);

O2A1O1Ixp33_ASAP7_75t_L g1445 ( 
.A1(n_1336),
.A2(n_1313),
.B(n_1325),
.C(n_1305),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1349),
.B(n_1358),
.Y(n_1446)
);

NOR2x1_ASAP7_75t_SL g1447 ( 
.A(n_1367),
.B(n_1379),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1334),
.Y(n_1448)
);

A2O1A1Ixp33_ASAP7_75t_L g1449 ( 
.A1(n_1341),
.A2(n_1306),
.B(n_1360),
.C(n_1340),
.Y(n_1449)
);

AOI21xp5_ASAP7_75t_SL g1450 ( 
.A1(n_1296),
.A2(n_1401),
.B(n_1357),
.Y(n_1450)
);

AOI21xp5_ASAP7_75t_SL g1451 ( 
.A1(n_1365),
.A2(n_1398),
.B(n_1353),
.Y(n_1451)
);

NOR2xp67_ASAP7_75t_L g1452 ( 
.A(n_1398),
.B(n_1282),
.Y(n_1452)
);

OR2x2_ASAP7_75t_L g1453 ( 
.A(n_1309),
.B(n_1340),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1309),
.B(n_1327),
.Y(n_1454)
);

OAI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1343),
.A2(n_1391),
.B1(n_1342),
.B2(n_1353),
.Y(n_1455)
);

INVxp67_ASAP7_75t_L g1456 ( 
.A(n_1322),
.Y(n_1456)
);

OA21x2_ASAP7_75t_L g1457 ( 
.A1(n_1287),
.A2(n_1297),
.B(n_1300),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1310),
.B(n_1322),
.Y(n_1458)
);

AND2x4_ASAP7_75t_SL g1459 ( 
.A(n_1319),
.B(n_1331),
.Y(n_1459)
);

NOR2xp67_ASAP7_75t_L g1460 ( 
.A(n_1282),
.B(n_1319),
.Y(n_1460)
);

OAI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1391),
.A2(n_1338),
.B1(n_1335),
.B2(n_1339),
.Y(n_1461)
);

HB1xp67_ASAP7_75t_L g1462 ( 
.A(n_1347),
.Y(n_1462)
);

OR2x2_ASAP7_75t_L g1463 ( 
.A(n_1318),
.B(n_1329),
.Y(n_1463)
);

AOI221x1_ASAP7_75t_SL g1464 ( 
.A1(n_1360),
.A2(n_1318),
.B1(n_1391),
.B2(n_1323),
.C(n_1328),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1326),
.B(n_1318),
.Y(n_1465)
);

AND2x2_ASAP7_75t_L g1466 ( 
.A(n_1329),
.B(n_1318),
.Y(n_1466)
);

INVx1_ASAP7_75t_SL g1467 ( 
.A(n_1356),
.Y(n_1467)
);

INVx2_ASAP7_75t_SL g1468 ( 
.A(n_1283),
.Y(n_1468)
);

OA21x2_ASAP7_75t_L g1469 ( 
.A1(n_1283),
.A2(n_1378),
.B(n_1400),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1323),
.B(n_1405),
.Y(n_1470)
);

AND2x4_ASAP7_75t_L g1471 ( 
.A(n_1348),
.B(n_1350),
.Y(n_1471)
);

OR2x2_ASAP7_75t_L g1472 ( 
.A(n_1364),
.B(n_1366),
.Y(n_1472)
);

BUFx12f_ASAP7_75t_L g1473 ( 
.A(n_1366),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1368),
.B(n_1405),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1400),
.B(n_1370),
.Y(n_1475)
);

AOI21xp5_ASAP7_75t_SL g1476 ( 
.A1(n_1385),
.A2(n_1387),
.B(n_1390),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1387),
.B(n_1390),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1394),
.B(n_1395),
.Y(n_1478)
);

BUFx12f_ASAP7_75t_L g1479 ( 
.A(n_1395),
.Y(n_1479)
);

OR2x2_ASAP7_75t_L g1480 ( 
.A(n_1299),
.B(n_1352),
.Y(n_1480)
);

AOI21xp5_ASAP7_75t_SL g1481 ( 
.A1(n_1345),
.A2(n_1266),
.B(n_1263),
.Y(n_1481)
);

BUFx3_ASAP7_75t_L g1482 ( 
.A(n_1295),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1294),
.B(n_1291),
.Y(n_1483)
);

OAI21xp5_ASAP7_75t_SL g1484 ( 
.A1(n_1286),
.A2(n_1257),
.B(n_1278),
.Y(n_1484)
);

A2O1A1Ixp33_ASAP7_75t_L g1485 ( 
.A1(n_1371),
.A2(n_1266),
.B(n_1263),
.C(n_1257),
.Y(n_1485)
);

AOI21xp5_ASAP7_75t_SL g1486 ( 
.A1(n_1345),
.A2(n_1266),
.B(n_1263),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1280),
.B(n_1344),
.Y(n_1487)
);

OA21x2_ASAP7_75t_L g1488 ( 
.A1(n_1330),
.A2(n_1301),
.B(n_1292),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1280),
.B(n_1344),
.Y(n_1489)
);

CKINVDCx5p33_ASAP7_75t_R g1490 ( 
.A(n_1384),
.Y(n_1490)
);

OAI22xp5_ASAP7_75t_L g1491 ( 
.A1(n_1374),
.A2(n_1165),
.B1(n_1266),
.B2(n_1263),
.Y(n_1491)
);

OR2x2_ASAP7_75t_L g1492 ( 
.A(n_1299),
.B(n_1352),
.Y(n_1492)
);

O2A1O1Ixp5_ASAP7_75t_L g1493 ( 
.A1(n_1351),
.A2(n_1257),
.B(n_1266),
.C(n_1263),
.Y(n_1493)
);

O2A1O1Ixp33_ASAP7_75t_L g1494 ( 
.A1(n_1284),
.A2(n_1257),
.B(n_1266),
.C(n_1263),
.Y(n_1494)
);

INVxp33_ASAP7_75t_L g1495 ( 
.A(n_1308),
.Y(n_1495)
);

OR2x2_ASAP7_75t_L g1496 ( 
.A(n_1299),
.B(n_1352),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1280),
.B(n_1344),
.Y(n_1497)
);

AND2x4_ASAP7_75t_L g1498 ( 
.A(n_1373),
.B(n_1316),
.Y(n_1498)
);

OAI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1374),
.A2(n_1165),
.B1(n_1266),
.B2(n_1263),
.Y(n_1499)
);

INVx1_ASAP7_75t_SL g1500 ( 
.A(n_1299),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1299),
.B(n_1352),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1280),
.B(n_1344),
.Y(n_1502)
);

OAI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1374),
.A2(n_1165),
.B1(n_1266),
.B2(n_1263),
.Y(n_1503)
);

AND2x4_ASAP7_75t_L g1504 ( 
.A(n_1373),
.B(n_1316),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1294),
.B(n_1291),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_1470),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1448),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1466),
.B(n_1449),
.Y(n_1508)
);

CKINVDCx20_ASAP7_75t_R g1509 ( 
.A(n_1415),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1463),
.B(n_1453),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1413),
.B(n_1427),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1456),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1408),
.B(n_1488),
.Y(n_1513)
);

HB1xp67_ASAP7_75t_L g1514 ( 
.A(n_1465),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1444),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1458),
.B(n_1462),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1444),
.Y(n_1517)
);

OAI21xp5_ASAP7_75t_L g1518 ( 
.A1(n_1493),
.A2(n_1494),
.B(n_1485),
.Y(n_1518)
);

INVxp67_ASAP7_75t_SL g1519 ( 
.A(n_1427),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1408),
.B(n_1488),
.Y(n_1520)
);

OA21x2_ASAP7_75t_L g1521 ( 
.A1(n_1439),
.A2(n_1493),
.B(n_1467),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1413),
.B(n_1424),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1469),
.Y(n_1523)
);

OR2x6_ASAP7_75t_L g1524 ( 
.A(n_1451),
.B(n_1421),
.Y(n_1524)
);

BUFx3_ASAP7_75t_L g1525 ( 
.A(n_1421),
.Y(n_1525)
);

AO21x2_ASAP7_75t_L g1526 ( 
.A1(n_1476),
.A2(n_1424),
.B(n_1486),
.Y(n_1526)
);

AO21x2_ASAP7_75t_L g1527 ( 
.A1(n_1481),
.A2(n_1454),
.B(n_1484),
.Y(n_1527)
);

OA21x2_ASAP7_75t_L g1528 ( 
.A1(n_1474),
.A2(n_1475),
.B(n_1477),
.Y(n_1528)
);

HB1xp67_ASAP7_75t_L g1529 ( 
.A(n_1461),
.Y(n_1529)
);

AOI21x1_ASAP7_75t_L g1530 ( 
.A1(n_1417),
.A2(n_1478),
.B(n_1471),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1447),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1472),
.Y(n_1532)
);

BUFx2_ASAP7_75t_L g1533 ( 
.A(n_1473),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1410),
.B(n_1483),
.Y(n_1534)
);

BUFx2_ASAP7_75t_L g1535 ( 
.A(n_1479),
.Y(n_1535)
);

AO21x2_ASAP7_75t_L g1536 ( 
.A1(n_1445),
.A2(n_1494),
.B(n_1428),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1457),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1505),
.B(n_1412),
.Y(n_1538)
);

INVxp67_ASAP7_75t_SL g1539 ( 
.A(n_1445),
.Y(n_1539)
);

OA21x2_ASAP7_75t_L g1540 ( 
.A1(n_1468),
.A2(n_1433),
.B(n_1442),
.Y(n_1540)
);

INVx3_ASAP7_75t_L g1541 ( 
.A(n_1457),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1446),
.B(n_1443),
.Y(n_1542)
);

AO21x2_ASAP7_75t_L g1543 ( 
.A1(n_1428),
.A2(n_1422),
.B(n_1409),
.Y(n_1543)
);

NAND2xp5_ASAP7_75t_SL g1544 ( 
.A(n_1422),
.B(n_1491),
.Y(n_1544)
);

AO21x2_ASAP7_75t_L g1545 ( 
.A1(n_1499),
.A2(n_1503),
.B(n_1419),
.Y(n_1545)
);

BUFx2_ASAP7_75t_L g1546 ( 
.A(n_1435),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1464),
.Y(n_1547)
);

AOI21xp5_ASAP7_75t_L g1548 ( 
.A1(n_1544),
.A2(n_1420),
.B(n_1414),
.Y(n_1548)
);

CKINVDCx20_ASAP7_75t_R g1549 ( 
.A(n_1509),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1516),
.B(n_1489),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1538),
.B(n_1500),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1507),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1510),
.B(n_1480),
.Y(n_1553)
);

OR2x2_ASAP7_75t_L g1554 ( 
.A(n_1510),
.B(n_1492),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1516),
.B(n_1487),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1507),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1514),
.Y(n_1557)
);

OR2x2_ASAP7_75t_L g1558 ( 
.A(n_1506),
.B(n_1501),
.Y(n_1558)
);

BUFx3_ASAP7_75t_L g1559 ( 
.A(n_1533),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1506),
.B(n_1411),
.Y(n_1560)
);

INVxp67_ASAP7_75t_L g1561 ( 
.A(n_1538),
.Y(n_1561)
);

AO21x2_ASAP7_75t_L g1562 ( 
.A1(n_1515),
.A2(n_1441),
.B(n_1436),
.Y(n_1562)
);

NOR2x1_ASAP7_75t_L g1563 ( 
.A(n_1526),
.B(n_1460),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1523),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1516),
.B(n_1508),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_SL g1566 ( 
.A1(n_1543),
.A2(n_1434),
.B1(n_1432),
.B2(n_1437),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_SL g1567 ( 
.A1(n_1543),
.A2(n_1504),
.B1(n_1498),
.B2(n_1416),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1506),
.B(n_1496),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1508),
.B(n_1502),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1542),
.B(n_1528),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1542),
.B(n_1497),
.Y(n_1571)
);

INVxp67_ASAP7_75t_L g1572 ( 
.A(n_1534),
.Y(n_1572)
);

AND2x4_ASAP7_75t_L g1573 ( 
.A(n_1525),
.B(n_1459),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1540),
.B(n_1426),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1542),
.B(n_1418),
.Y(n_1575)
);

HB1xp67_ASAP7_75t_L g1576 ( 
.A(n_1514),
.Y(n_1576)
);

BUFx2_ASAP7_75t_L g1577 ( 
.A(n_1525),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1534),
.B(n_1438),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1528),
.B(n_1495),
.Y(n_1579)
);

BUFx2_ASAP7_75t_L g1580 ( 
.A(n_1533),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1528),
.B(n_1495),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1519),
.B(n_1429),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1552),
.Y(n_1583)
);

AND2x4_ASAP7_75t_L g1584 ( 
.A(n_1559),
.B(n_1546),
.Y(n_1584)
);

AO21x2_ASAP7_75t_L g1585 ( 
.A1(n_1564),
.A2(n_1517),
.B(n_1515),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1552),
.Y(n_1586)
);

NAND3xp33_ASAP7_75t_L g1587 ( 
.A(n_1566),
.B(n_1518),
.C(n_1511),
.Y(n_1587)
);

INVxp67_ASAP7_75t_L g1588 ( 
.A(n_1553),
.Y(n_1588)
);

NOR2xp33_ASAP7_75t_L g1589 ( 
.A(n_1572),
.B(n_1544),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1561),
.B(n_1519),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1553),
.B(n_1532),
.Y(n_1591)
);

OAI22xp5_ASAP7_75t_L g1592 ( 
.A1(n_1567),
.A2(n_1522),
.B1(n_1511),
.B2(n_1518),
.Y(n_1592)
);

BUFx3_ASAP7_75t_L g1593 ( 
.A(n_1549),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1556),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1564),
.Y(n_1595)
);

AOI21xp5_ASAP7_75t_L g1596 ( 
.A1(n_1548),
.A2(n_1543),
.B(n_1522),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_L g1597 ( 
.A(n_1557),
.Y(n_1597)
);

BUFx2_ASAP7_75t_L g1598 ( 
.A(n_1559),
.Y(n_1598)
);

INVx1_ASAP7_75t_SL g1599 ( 
.A(n_1554),
.Y(n_1599)
);

AOI211xp5_ASAP7_75t_L g1600 ( 
.A1(n_1582),
.A2(n_1539),
.B(n_1547),
.C(n_1431),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1571),
.B(n_1533),
.Y(n_1601)
);

OAI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1563),
.A2(n_1539),
.B1(n_1547),
.B2(n_1529),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_SL g1603 ( 
.A1(n_1562),
.A2(n_1543),
.B1(n_1545),
.B2(n_1526),
.Y(n_1603)
);

CKINVDCx8_ASAP7_75t_R g1604 ( 
.A(n_1580),
.Y(n_1604)
);

AND2x4_ASAP7_75t_SL g1605 ( 
.A(n_1573),
.B(n_1524),
.Y(n_1605)
);

HB1xp67_ASAP7_75t_L g1606 ( 
.A(n_1576),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1571),
.B(n_1535),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1554),
.A2(n_1529),
.B1(n_1535),
.B2(n_1455),
.Y(n_1608)
);

AO21x2_ASAP7_75t_L g1609 ( 
.A1(n_1579),
.A2(n_1517),
.B(n_1515),
.Y(n_1609)
);

OAI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1578),
.A2(n_1543),
.B1(n_1521),
.B2(n_1551),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1565),
.B(n_1528),
.Y(n_1611)
);

INVx1_ASAP7_75t_SL g1612 ( 
.A(n_1558),
.Y(n_1612)
);

OAI321xp33_ASAP7_75t_L g1613 ( 
.A1(n_1580),
.A2(n_1530),
.A3(n_1524),
.B1(n_1531),
.B2(n_1546),
.C(n_1512),
.Y(n_1613)
);

OAI22xp5_ASAP7_75t_L g1614 ( 
.A1(n_1558),
.A2(n_1535),
.B1(n_1524),
.B2(n_1416),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1575),
.B(n_1527),
.Y(n_1615)
);

NOR2xp33_ASAP7_75t_L g1616 ( 
.A(n_1560),
.B(n_1545),
.Y(n_1616)
);

BUFx3_ASAP7_75t_L g1617 ( 
.A(n_1577),
.Y(n_1617)
);

BUFx3_ASAP7_75t_L g1618 ( 
.A(n_1577),
.Y(n_1618)
);

AOI22xp33_ASAP7_75t_L g1619 ( 
.A1(n_1562),
.A2(n_1545),
.B1(n_1536),
.B2(n_1526),
.Y(n_1619)
);

NAND4xp25_ASAP7_75t_SL g1620 ( 
.A(n_1574),
.B(n_1450),
.C(n_1509),
.D(n_1430),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1585),
.Y(n_1621)
);

AND2x4_ASAP7_75t_L g1622 ( 
.A(n_1605),
.B(n_1570),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1583),
.Y(n_1623)
);

INVx2_ASAP7_75t_L g1624 ( 
.A(n_1585),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1586),
.Y(n_1625)
);

AO21x2_ASAP7_75t_L g1626 ( 
.A1(n_1610),
.A2(n_1513),
.B(n_1520),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1594),
.Y(n_1627)
);

INVx2_ASAP7_75t_SL g1628 ( 
.A(n_1605),
.Y(n_1628)
);

NOR2x1_ASAP7_75t_L g1629 ( 
.A(n_1610),
.B(n_1620),
.Y(n_1629)
);

BUFx2_ASAP7_75t_L g1630 ( 
.A(n_1617),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1616),
.B(n_1570),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1616),
.B(n_1615),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1611),
.B(n_1579),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1611),
.B(n_1581),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1609),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1597),
.Y(n_1636)
);

OAI21x1_ASAP7_75t_L g1637 ( 
.A1(n_1619),
.A2(n_1541),
.B(n_1537),
.Y(n_1637)
);

INVx2_ASAP7_75t_L g1638 ( 
.A(n_1609),
.Y(n_1638)
);

INVx3_ASAP7_75t_L g1639 ( 
.A(n_1595),
.Y(n_1639)
);

INVx1_ASAP7_75t_SL g1640 ( 
.A(n_1597),
.Y(n_1640)
);

OAI21x1_ASAP7_75t_L g1641 ( 
.A1(n_1596),
.A2(n_1541),
.B(n_1523),
.Y(n_1641)
);

BUFx3_ASAP7_75t_L g1642 ( 
.A(n_1604),
.Y(n_1642)
);

INVxp67_ASAP7_75t_L g1643 ( 
.A(n_1589),
.Y(n_1643)
);

INVx3_ASAP7_75t_L g1644 ( 
.A(n_1584),
.Y(n_1644)
);

NOR2xp33_ASAP7_75t_L g1645 ( 
.A(n_1589),
.B(n_1569),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1642),
.B(n_1628),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1640),
.B(n_1590),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1643),
.B(n_1569),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1623),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1642),
.B(n_1584),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1621),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1621),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1623),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1643),
.B(n_1588),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1642),
.B(n_1584),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1642),
.B(n_1598),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1623),
.Y(n_1657)
);

AND3x2_ASAP7_75t_L g1658 ( 
.A(n_1630),
.B(n_1600),
.C(n_1606),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1642),
.B(n_1565),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1625),
.Y(n_1660)
);

NOR2x1_ASAP7_75t_L g1661 ( 
.A(n_1629),
.B(n_1587),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1640),
.B(n_1606),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1628),
.B(n_1604),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1628),
.B(n_1601),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1628),
.B(n_1607),
.Y(n_1665)
);

NOR3xp33_ASAP7_75t_SL g1666 ( 
.A(n_1632),
.B(n_1613),
.C(n_1602),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1621),
.Y(n_1667)
);

NAND2x1_ASAP7_75t_L g1668 ( 
.A(n_1629),
.B(n_1524),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1625),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1644),
.B(n_1617),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1621),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1644),
.B(n_1618),
.Y(n_1672)
);

INVx2_ASAP7_75t_SL g1673 ( 
.A(n_1630),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_L g1674 ( 
.A(n_1645),
.B(n_1593),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1625),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1645),
.B(n_1599),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1632),
.B(n_1592),
.Y(n_1677)
);

OR2x2_ASAP7_75t_L g1678 ( 
.A(n_1640),
.B(n_1574),
.Y(n_1678)
);

INVx1_ASAP7_75t_SL g1679 ( 
.A(n_1630),
.Y(n_1679)
);

INVxp67_ASAP7_75t_L g1680 ( 
.A(n_1636),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1636),
.B(n_1591),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_L g1682 ( 
.A(n_1632),
.B(n_1550),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1639),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1627),
.Y(n_1684)
);

INVx1_ASAP7_75t_SL g1685 ( 
.A(n_1629),
.Y(n_1685)
);

INVx1_ASAP7_75t_SL g1686 ( 
.A(n_1644),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1626),
.B(n_1612),
.Y(n_1687)
);

HB1xp67_ASAP7_75t_SL g1688 ( 
.A(n_1622),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1624),
.Y(n_1689)
);

OR2x2_ASAP7_75t_L g1690 ( 
.A(n_1626),
.B(n_1631),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1649),
.Y(n_1691)
);

HB1xp67_ASAP7_75t_L g1692 ( 
.A(n_1673),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1663),
.B(n_1622),
.Y(n_1693)
);

OR2x2_ASAP7_75t_L g1694 ( 
.A(n_1654),
.B(n_1631),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1649),
.Y(n_1695)
);

AOI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1661),
.A2(n_1603),
.B1(n_1536),
.B2(n_1626),
.Y(n_1696)
);

NAND2xp33_ASAP7_75t_L g1697 ( 
.A(n_1661),
.B(n_1440),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1663),
.B(n_1644),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1653),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1685),
.B(n_1631),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1653),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1646),
.B(n_1622),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1648),
.B(n_1560),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1677),
.B(n_1550),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1666),
.B(n_1555),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_L g1706 ( 
.A(n_1674),
.B(n_1593),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1646),
.B(n_1622),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1657),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1682),
.B(n_1568),
.Y(n_1709)
);

INVx1_ASAP7_75t_SL g1710 ( 
.A(n_1656),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_L g1711 ( 
.A(n_1676),
.B(n_1490),
.Y(n_1711)
);

INVx2_ASAP7_75t_SL g1712 ( 
.A(n_1673),
.Y(n_1712)
);

AOI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1668),
.A2(n_1536),
.B1(n_1626),
.B2(n_1527),
.Y(n_1713)
);

AND2x2_ASAP7_75t_SL g1714 ( 
.A(n_1656),
.B(n_1521),
.Y(n_1714)
);

INVx1_ASAP7_75t_SL g1715 ( 
.A(n_1679),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1650),
.B(n_1644),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1657),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1660),
.Y(n_1718)
);

AOI21xp5_ASAP7_75t_L g1719 ( 
.A1(n_1668),
.A2(n_1626),
.B(n_1527),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1659),
.B(n_1658),
.Y(n_1720)
);

A2O1A1Ixp33_ASAP7_75t_L g1721 ( 
.A1(n_1690),
.A2(n_1641),
.B(n_1608),
.C(n_1452),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1660),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1650),
.B(n_1655),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1669),
.Y(n_1724)
);

AOI22xp5_ASAP7_75t_L g1725 ( 
.A1(n_1659),
.A2(n_1626),
.B1(n_1527),
.B2(n_1614),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1669),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1675),
.Y(n_1727)
);

BUFx2_ASAP7_75t_L g1728 ( 
.A(n_1692),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1723),
.B(n_1655),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1723),
.B(n_1664),
.Y(n_1730)
);

INVx3_ASAP7_75t_L g1731 ( 
.A(n_1712),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1693),
.B(n_1664),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1698),
.B(n_1665),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1692),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1698),
.B(n_1665),
.Y(n_1735)
);

CKINVDCx16_ASAP7_75t_R g1736 ( 
.A(n_1706),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1700),
.B(n_1680),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1694),
.B(n_1662),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1691),
.Y(n_1739)
);

INVx1_ASAP7_75t_SL g1740 ( 
.A(n_1710),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1712),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1695),
.Y(n_1742)
);

OAI22xp5_ASAP7_75t_L g1743 ( 
.A1(n_1696),
.A2(n_1690),
.B1(n_1687),
.B2(n_1688),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1716),
.B(n_1670),
.Y(n_1744)
);

INVx1_ASAP7_75t_SL g1745 ( 
.A(n_1715),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1699),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1701),
.Y(n_1747)
);

OAI21xp5_ASAP7_75t_SL g1748 ( 
.A1(n_1720),
.A2(n_1687),
.B(n_1662),
.Y(n_1748)
);

CKINVDCx20_ASAP7_75t_R g1749 ( 
.A(n_1706),
.Y(n_1749)
);

OAI21x1_ASAP7_75t_L g1750 ( 
.A1(n_1719),
.A2(n_1672),
.B(n_1670),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1714),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1708),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1714),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1704),
.B(n_1647),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1705),
.B(n_1647),
.Y(n_1755)
);

AOI21xp33_ASAP7_75t_L g1756 ( 
.A1(n_1745),
.A2(n_1697),
.B(n_1713),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1729),
.B(n_1716),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1745),
.B(n_1697),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1740),
.B(n_1711),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_SL g1760 ( 
.A(n_1736),
.B(n_1725),
.Y(n_1760)
);

OR2x2_ASAP7_75t_L g1761 ( 
.A(n_1740),
.B(n_1703),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1728),
.Y(n_1762)
);

OAI21xp33_ASAP7_75t_L g1763 ( 
.A1(n_1755),
.A2(n_1729),
.B(n_1748),
.Y(n_1763)
);

OR2x2_ASAP7_75t_L g1764 ( 
.A(n_1738),
.B(n_1709),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1728),
.Y(n_1765)
);

OR2x2_ASAP7_75t_L g1766 ( 
.A(n_1738),
.B(n_1681),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1734),
.Y(n_1767)
);

AOI21xp5_ASAP7_75t_L g1768 ( 
.A1(n_1743),
.A2(n_1721),
.B(n_1711),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1734),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1739),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1731),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1739),
.Y(n_1772)
);

A2O1A1Ixp33_ASAP7_75t_L g1773 ( 
.A1(n_1748),
.A2(n_1721),
.B(n_1641),
.C(n_1637),
.Y(n_1773)
);

OAI211xp5_ASAP7_75t_L g1774 ( 
.A1(n_1743),
.A2(n_1727),
.B(n_1726),
.C(n_1724),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1730),
.B(n_1702),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1742),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1730),
.B(n_1733),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1777),
.B(n_1736),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1762),
.Y(n_1779)
);

NAND2xp5_ASAP7_75t_L g1780 ( 
.A(n_1777),
.B(n_1733),
.Y(n_1780)
);

NOR2xp33_ASAP7_75t_L g1781 ( 
.A(n_1759),
.B(n_1749),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1765),
.Y(n_1782)
);

OAI221xp5_ASAP7_75t_SL g1783 ( 
.A1(n_1768),
.A2(n_1753),
.B1(n_1751),
.B2(n_1737),
.C(n_1754),
.Y(n_1783)
);

OR2x2_ASAP7_75t_L g1784 ( 
.A(n_1761),
.B(n_1737),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1771),
.Y(n_1785)
);

NOR2xp33_ASAP7_75t_L g1786 ( 
.A(n_1758),
.B(n_1741),
.Y(n_1786)
);

AOI22xp33_ASAP7_75t_SL g1787 ( 
.A1(n_1757),
.A2(n_1753),
.B1(n_1751),
.B2(n_1735),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1763),
.B(n_1735),
.Y(n_1788)
);

AOI22xp33_ASAP7_75t_L g1789 ( 
.A1(n_1756),
.A2(n_1753),
.B1(n_1751),
.B2(n_1731),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1757),
.B(n_1732),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1775),
.B(n_1732),
.Y(n_1791)
);

AOI22xp33_ASAP7_75t_L g1792 ( 
.A1(n_1778),
.A2(n_1760),
.B1(n_1775),
.B2(n_1744),
.Y(n_1792)
);

AOI22xp5_ASAP7_75t_L g1793 ( 
.A1(n_1781),
.A2(n_1760),
.B1(n_1744),
.B2(n_1774),
.Y(n_1793)
);

A2O1A1Ixp33_ASAP7_75t_L g1794 ( 
.A1(n_1783),
.A2(n_1773),
.B(n_1750),
.C(n_1767),
.Y(n_1794)
);

OAI221xp5_ASAP7_75t_L g1795 ( 
.A1(n_1789),
.A2(n_1773),
.B1(n_1766),
.B2(n_1764),
.C(n_1769),
.Y(n_1795)
);

NAND3xp33_ASAP7_75t_L g1796 ( 
.A(n_1789),
.B(n_1741),
.C(n_1771),
.Y(n_1796)
);

AOI221xp5_ASAP7_75t_L g1797 ( 
.A1(n_1786),
.A2(n_1776),
.B1(n_1772),
.B2(n_1770),
.C(n_1741),
.Y(n_1797)
);

OAI211xp5_ASAP7_75t_SL g1798 ( 
.A1(n_1788),
.A2(n_1731),
.B(n_1752),
.C(n_1742),
.Y(n_1798)
);

AOI22xp5_ASAP7_75t_L g1799 ( 
.A1(n_1781),
.A2(n_1731),
.B1(n_1707),
.B2(n_1754),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1786),
.B(n_1746),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1785),
.Y(n_1801)
);

AOI221xp5_ASAP7_75t_L g1802 ( 
.A1(n_1779),
.A2(n_1752),
.B1(n_1747),
.B2(n_1746),
.C(n_1717),
.Y(n_1802)
);

AOI211xp5_ASAP7_75t_L g1803 ( 
.A1(n_1784),
.A2(n_1782),
.B(n_1780),
.C(n_1790),
.Y(n_1803)
);

NAND3xp33_ASAP7_75t_SL g1804 ( 
.A(n_1793),
.B(n_1787),
.C(n_1791),
.Y(n_1804)
);

CKINVDCx5p33_ASAP7_75t_R g1805 ( 
.A(n_1801),
.Y(n_1805)
);

XNOR2xp5_ASAP7_75t_L g1806 ( 
.A(n_1792),
.B(n_1747),
.Y(n_1806)
);

AOI22xp5_ASAP7_75t_L g1807 ( 
.A1(n_1795),
.A2(n_1799),
.B1(n_1798),
.B2(n_1796),
.Y(n_1807)
);

AOI21xp5_ASAP7_75t_L g1808 ( 
.A1(n_1794),
.A2(n_1750),
.B(n_1722),
.Y(n_1808)
);

OAI221xp5_ASAP7_75t_L g1809 ( 
.A1(n_1803),
.A2(n_1718),
.B1(n_1686),
.B2(n_1678),
.C(n_1423),
.Y(n_1809)
);

AOI221xp5_ASAP7_75t_L g1810 ( 
.A1(n_1797),
.A2(n_1635),
.B1(n_1638),
.B2(n_1652),
.C(n_1667),
.Y(n_1810)
);

NOR2xp33_ASAP7_75t_L g1811 ( 
.A(n_1804),
.B(n_1805),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1806),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1809),
.Y(n_1813)
);

CKINVDCx16_ASAP7_75t_R g1814 ( 
.A(n_1807),
.Y(n_1814)
);

OR2x2_ASAP7_75t_L g1815 ( 
.A(n_1808),
.B(n_1800),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1810),
.B(n_1802),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1807),
.B(n_1675),
.Y(n_1817)
);

AOI22x1_ASAP7_75t_L g1818 ( 
.A1(n_1814),
.A2(n_1425),
.B1(n_1651),
.B2(n_1652),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1811),
.B(n_1672),
.Y(n_1819)
);

XNOR2xp5_ASAP7_75t_L g1820 ( 
.A(n_1812),
.B(n_1813),
.Y(n_1820)
);

XNOR2x1_ASAP7_75t_L g1821 ( 
.A(n_1815),
.B(n_1482),
.Y(n_1821)
);

NOR2xp33_ASAP7_75t_SL g1822 ( 
.A(n_1817),
.B(n_1681),
.Y(n_1822)
);

NAND3x1_ASAP7_75t_SL g1823 ( 
.A(n_1816),
.B(n_1634),
.C(n_1633),
.Y(n_1823)
);

NOR2xp33_ASAP7_75t_L g1824 ( 
.A(n_1819),
.B(n_1817),
.Y(n_1824)
);

NOR3xp33_ASAP7_75t_L g1825 ( 
.A(n_1823),
.B(n_1652),
.C(n_1651),
.Y(n_1825)
);

OA21x2_ASAP7_75t_L g1826 ( 
.A1(n_1820),
.A2(n_1684),
.B(n_1667),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1826),
.Y(n_1827)
);

AOI322xp5_ASAP7_75t_L g1828 ( 
.A1(n_1827),
.A2(n_1824),
.A3(n_1822),
.B1(n_1825),
.B2(n_1821),
.C1(n_1818),
.C2(n_1689),
.Y(n_1828)
);

AOI22xp5_ASAP7_75t_L g1829 ( 
.A1(n_1828),
.A2(n_1689),
.B1(n_1667),
.B2(n_1671),
.Y(n_1829)
);

CKINVDCx20_ASAP7_75t_R g1830 ( 
.A(n_1828),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1830),
.B(n_1684),
.Y(n_1831)
);

NOR2x1_ASAP7_75t_L g1832 ( 
.A(n_1829),
.B(n_1651),
.Y(n_1832)
);

AOI22xp5_ASAP7_75t_L g1833 ( 
.A1(n_1831),
.A2(n_1689),
.B1(n_1671),
.B2(n_1635),
.Y(n_1833)
);

BUFx2_ASAP7_75t_L g1834 ( 
.A(n_1832),
.Y(n_1834)
);

INVx4_ASAP7_75t_L g1835 ( 
.A(n_1834),
.Y(n_1835)
);

AOI22xp33_ASAP7_75t_L g1836 ( 
.A1(n_1835),
.A2(n_1833),
.B1(n_1671),
.B2(n_1638),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1836),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1837),
.B(n_1678),
.Y(n_1838)
);

AOI22xp5_ASAP7_75t_L g1839 ( 
.A1(n_1838),
.A2(n_1635),
.B1(n_1638),
.B2(n_1683),
.Y(n_1839)
);

AOI211xp5_ASAP7_75t_L g1840 ( 
.A1(n_1839),
.A2(n_1635),
.B(n_1638),
.C(n_1683),
.Y(n_1840)
);


endmodule