module real_jpeg_30102_n_10 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9, n_10);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_9;

output n_10;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_11;
wire n_131;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_13;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_57;
wire n_43;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_0),
.A2(n_34),
.B1(n_35),
.B2(n_66),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_0),
.Y(n_66)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_1),
.Y(n_62)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_1),
.Y(n_113)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_5),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_5),
.A2(n_20),
.B1(n_41),
.B2(n_42),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_5),
.A2(n_20),
.B1(n_29),
.B2(n_30),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_5),
.A2(n_20),
.B1(n_34),
.B2(n_35),
.Y(n_64)
);

AOI21xp33_ASAP7_75t_SL g74 ( 
.A1(n_5),
.A2(n_26),
.B(n_30),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_5),
.B(n_89),
.Y(n_88)
);

AOI21xp33_ASAP7_75t_L g99 ( 
.A1(n_5),
.A2(n_6),
.B(n_35),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_5),
.B(n_104),
.Y(n_103)
);

O2A1O1Ixp33_ASAP7_75t_L g122 ( 
.A1(n_5),
.A2(n_8),
.B(n_29),
.C(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_6),
.A2(n_34),
.B1(n_35),
.B2(n_37),
.Y(n_33)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

INVx11_ASAP7_75t_SL g36 ( 
.A(n_9),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_92),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_90),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_13),
.Y(n_12)
);

AND2x2_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_79),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_14),
.B(n_79),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_68),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g15 ( 
.A1(n_16),
.A2(n_17),
.B1(n_58),
.B2(n_59),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

AOI211xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_31),
.B(n_44),
.C(n_56),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_18),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_18),
.A2(n_45),
.B1(n_46),
.B2(n_57),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_18),
.A2(n_57),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_23),
.Y(n_18)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_20),
.A2(n_21),
.B(n_27),
.C(n_74),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_20),
.A2(n_37),
.B(n_42),
.C(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_20),
.B(n_33),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_20),
.B(n_113),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_L g123 ( 
.A1(n_20),
.A2(n_41),
.B(n_51),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_21),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_21),
.A2(n_22),
.B1(n_26),
.B2(n_27),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_28),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_28),
.Y(n_24)
);

CKINVDCx14_ASAP7_75t_R g27 ( 
.A(n_26),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_26),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_29),
.A2(n_30),
.B1(n_49),
.B2(n_51),
.Y(n_53)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_31),
.A2(n_55),
.B1(n_60),
.B2(n_67),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_31),
.A2(n_45),
.B1(n_46),
.B2(n_55),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_31),
.A2(n_55),
.B1(n_102),
.B2(n_103),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_31),
.A2(n_55),
.B1(n_98),
.B2(n_116),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_31),
.B(n_75),
.C(n_102),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_31),
.A2(n_55),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_31),
.B(n_131),
.C(n_137),
.Y(n_141)
);

AND2x2_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_43),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_38),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_34),
.B(n_112),
.Y(n_111)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_35),
.B(n_62),
.Y(n_61)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_37),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_41),
.A2(n_42),
.B1(n_49),
.B2(n_51),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_44),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_55),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_45),
.B(n_57),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g128 ( 
.A1(n_45),
.A2(n_55),
.B(n_125),
.C(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_45),
.A2(n_46),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_46),
.B(n_75),
.C(n_87),
.Y(n_86)
);

AND2x2_ASAP7_75t_SL g46 ( 
.A(n_47),
.B(n_54),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_52),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_48),
.B(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_55),
.B(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_60),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_63),
.B2(n_65),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_61),
.B(n_62),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_77),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_71),
.B2(n_78),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_71),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_72),
.A2(n_73),
.B1(n_75),
.B2(n_76),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_75),
.A2(n_76),
.B1(n_101),
.B2(n_105),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_75),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_75),
.B(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_75),
.A2(n_76),
.B1(n_122),
.B2(n_124),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_75),
.A2(n_76),
.B1(n_87),
.B2(n_88),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_75),
.B(n_122),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_76),
.B(n_115),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_84),
.C(n_86),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_80),
.A2(n_81),
.B1(n_143),
.B2(n_145),
.Y(n_142)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_82),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_82),
.A2(n_83),
.B1(n_121),
.B2(n_125),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_84),
.A2(n_85),
.B1(n_86),
.B2(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_86),
.Y(n_144)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_140),
.B(n_146),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_127),
.B(n_139),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_118),
.B(n_126),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_106),
.B(n_117),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_100),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_100),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_98),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_101),
.Y(n_105)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_114),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_110),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_120),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_119),
.B(n_120),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_121),
.Y(n_125)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_122),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_130),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_130),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_135),
.B2(n_136),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_142),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_141),
.B(n_142),
.Y(n_146)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_143),
.Y(n_145)
);


endmodule