module fake_jpeg_5786_n_226 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_226);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_226;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_3),
.B(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_32),
.Y(n_48)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_33),
.A2(n_37),
.B1(n_29),
.B2(n_27),
.Y(n_63)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_20),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_35),
.B(n_39),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_15),
.B(n_0),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_30),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_15),
.B(n_1),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_45),
.Y(n_67)
);

AOI21xp33_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_27),
.B(n_22),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_44),
.B(n_16),
.C(n_28),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_30),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_38),
.B(n_20),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_53),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_51),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_33),
.A2(n_22),
.B1(n_27),
.B2(n_26),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_52),
.A2(n_60),
.B1(n_34),
.B2(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_35),
.B(n_25),
.Y(n_54)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_20),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_58),
.B(n_28),
.Y(n_79)
);

NAND2xp33_ASAP7_75t_SL g59 ( 
.A(n_34),
.B(n_26),
.Y(n_59)
);

OR2x2_ASAP7_75t_SL g73 ( 
.A(n_59),
.B(n_21),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_33),
.A2(n_22),
.B1(n_32),
.B2(n_37),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_64),
.A2(n_76),
.B1(n_50),
.B2(n_62),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_56),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_77),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_44),
.A2(n_31),
.B(n_42),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_66),
.A2(n_48),
.B(n_60),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_48),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_71),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_73),
.B(n_79),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_59),
.A2(n_34),
.B1(n_37),
.B2(n_32),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_75),
.A2(n_43),
.B1(n_49),
.B2(n_54),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_52),
.A2(n_31),
.B1(n_32),
.B2(n_41),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_78),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_80),
.A2(n_58),
.B(n_25),
.Y(n_90)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_67),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_83),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_46),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_91),
.Y(n_105)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_95),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_88),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_66),
.B(n_53),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_64),
.A2(n_57),
.B1(n_61),
.B2(n_50),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_89),
.A2(n_93),
.B1(n_94),
.B2(n_96),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_90),
.A2(n_102),
.B(n_79),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_53),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_64),
.A2(n_57),
.B1(n_55),
.B2(n_29),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_67),
.Y(n_95)
);

OA22x2_ASAP7_75t_L g96 ( 
.A1(n_76),
.A2(n_41),
.B1(n_40),
.B2(n_55),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_96),
.A2(n_98),
.B1(n_29),
.B2(n_68),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_80),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_80),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_45),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_72),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_73),
.A2(n_45),
.B(n_49),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_107),
.Y(n_126)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_101),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g134 ( 
.A1(n_109),
.A2(n_69),
.B(n_86),
.Y(n_134)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_115),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_111),
.A2(n_113),
.B(n_102),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_112),
.A2(n_119),
.B1(n_121),
.B2(n_96),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_100),
.A2(n_73),
.B(n_72),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_65),
.Y(n_114)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_114),
.Y(n_132)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_120),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_118),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_65),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_93),
.A2(n_81),
.B1(n_65),
.B2(n_68),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_99),
.A2(n_68),
.B1(n_78),
.B2(n_77),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_122),
.A2(n_123),
.B1(n_96),
.B2(n_82),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_98),
.A2(n_41),
.B1(n_69),
.B2(n_19),
.Y(n_123)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_105),
.B(n_88),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_134),
.C(n_136),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_128),
.A2(n_133),
.B(n_141),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_129),
.A2(n_104),
.B1(n_51),
.B2(n_24),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_117),
.B(n_95),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_130),
.B(n_131),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_107),
.B(n_84),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_116),
.A2(n_87),
.B1(n_90),
.B2(n_91),
.Y(n_133)
);

NOR3xp33_ASAP7_75t_SL g135 ( 
.A(n_111),
.B(n_47),
.C(n_40),
.Y(n_135)
);

OAI322xp33_ASAP7_75t_L g161 ( 
.A1(n_135),
.A2(n_24),
.A3(n_97),
.B1(n_70),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_105),
.B(n_24),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_112),
.A2(n_21),
.B1(n_19),
.B2(n_16),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_138),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_110),
.A2(n_122),
.B1(n_123),
.B2(n_106),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_140),
.A2(n_119),
.B1(n_104),
.B2(n_17),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_118),
.A2(n_51),
.B(n_70),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_143),
.Y(n_149)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_121),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_128),
.A2(n_113),
.B(n_115),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_144),
.A2(n_137),
.B(n_139),
.Y(n_171)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_127),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_147),
.B(n_148),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_134),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_150),
.B(n_153),
.Y(n_164)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g154 ( 
.A(n_135),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_154),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_155),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_51),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_157),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_141),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_127),
.Y(n_158)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_158),
.Y(n_170)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_126),
.Y(n_160)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_160),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_161),
.A2(n_142),
.B1(n_132),
.B2(n_143),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_162),
.B(n_158),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_146),
.A2(n_157),
.B1(n_152),
.B2(n_140),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_173),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_146),
.A2(n_130),
.B1(n_129),
.B2(n_131),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_165),
.B(n_177),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_150),
.A2(n_145),
.B(n_144),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_166),
.A2(n_171),
.B(n_174),
.Y(n_189)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_149),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_154),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_147),
.A2(n_124),
.B1(n_138),
.B2(n_132),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_1),
.C(n_2),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_145),
.A2(n_125),
.B1(n_136),
.B2(n_70),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_177),
.B(n_156),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_181),
.C(n_183),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_151),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_185),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_172),
.B(n_151),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_148),
.C(n_149),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_184),
.B(n_190),
.C(n_175),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_167),
.B(n_159),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_160),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_186),
.B(n_187),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_171),
.B(n_97),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_188),
.A2(n_164),
.B(n_174),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_2),
.C(n_3),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_178),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_191),
.B(n_197),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_189),
.A2(n_173),
.B1(n_169),
.B2(n_164),
.Y(n_193)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_193),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_195),
.B(n_199),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_190),
.B(n_162),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_R g198 ( 
.A(n_184),
.B(n_168),
.Y(n_198)
);

NOR2xp67_ASAP7_75t_L g209 ( 
.A(n_198),
.B(n_7),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_179),
.B(n_176),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_201),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_180),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_183),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_202),
.A2(n_209),
.B(n_9),
.Y(n_211)
);

NOR2x1_ASAP7_75t_L g204 ( 
.A(n_201),
.B(n_181),
.Y(n_204)
);

OAI211xp5_ASAP7_75t_L g214 ( 
.A1(n_204),
.A2(n_9),
.B(n_11),
.C(n_12),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_195),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_208),
.A2(n_192),
.B1(n_196),
.B2(n_194),
.Y(n_210)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_210),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_211),
.B(n_13),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_206),
.A2(n_194),
.B1(n_10),
.B2(n_11),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_212),
.A2(n_214),
.B1(n_204),
.B2(n_205),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_203),
.B(n_207),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_213),
.B(n_215),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_202),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_217),
.B(n_218),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_212),
.Y(n_221)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_221),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_219),
.B(n_210),
.C(n_14),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_222),
.A2(n_218),
.B(n_14),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_223),
.B(n_220),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_224),
.Y(n_226)
);


endmodule