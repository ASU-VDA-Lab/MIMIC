module fake_jpeg_3617_n_158 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_158);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_158;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_8),
.B(n_25),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_24),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

BUFx16f_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_60),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_0),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_61),
.B(n_63),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_62),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_44),
.B(n_1),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_59),
.A2(n_42),
.B1(n_43),
.B2(n_56),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_65),
.A2(n_68),
.B1(n_69),
.B2(n_70),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_58),
.A2(n_53),
.B1(n_50),
.B2(n_49),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_62),
.A2(n_42),
.B1(n_43),
.B2(n_56),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_62),
.A2(n_42),
.B1(n_43),
.B2(n_51),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_57),
.A2(n_50),
.B1(n_48),
.B2(n_52),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_72),
.A2(n_46),
.B1(n_3),
.B2(n_4),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_55),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_54),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_75),
.B(n_48),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_87),
.Y(n_92)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_74),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_84),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_80),
.B(n_81),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_67),
.B(n_1),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_73),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_83),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_2),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_64),
.Y(n_86)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_86),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_74),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_68),
.A2(n_46),
.B1(n_3),
.B2(n_4),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_88),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_103)
);

AO21x1_ASAP7_75t_L g97 ( 
.A1(n_89),
.A2(n_2),
.B(n_5),
.Y(n_97)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_90),
.B(n_26),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_76),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_93),
.B(n_99),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_87),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_96),
.B(n_105),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_103),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_79),
.A2(n_66),
.B(n_6),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_98),
.B(n_9),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_22),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_23),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_7),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_107),
.Y(n_113)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_100),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_114),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_91),
.A2(n_86),
.B(n_10),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_109),
.A2(n_117),
.B(n_120),
.Y(n_133)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_125),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_101),
.B(n_9),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_116),
.B(n_119),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_98),
.A2(n_29),
.B1(n_38),
.B2(n_12),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_117),
.A2(n_120),
.B1(n_121),
.B2(n_102),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_102),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_118),
.B(n_123),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_92),
.B(n_10),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_92),
.A2(n_30),
.B1(n_15),
.B2(n_20),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_103),
.A2(n_11),
.B1(n_21),
.B2(n_27),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_122),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_99),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_105),
.B(n_11),
.Y(n_125)
);

MAJx2_ASAP7_75t_L g126 ( 
.A(n_111),
.B(n_97),
.C(n_94),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_137),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_127),
.B(n_138),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_115),
.A2(n_31),
.B(n_32),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_133),
.B(n_113),
.Y(n_140)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_134),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_124),
.A2(n_36),
.B(n_39),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_136),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_124),
.B(n_121),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_140),
.B(n_129),
.Y(n_148)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_144),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_146),
.Y(n_150)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_141),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_142),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_147),
.B(n_148),
.C(n_126),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_149),
.B(n_143),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_151),
.B(n_150),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_152),
.B(n_110),
.C(n_142),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_153),
.A2(n_139),
.B1(n_127),
.B2(n_132),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_137),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_135),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_130),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_157),
.B(n_131),
.Y(n_158)
);


endmodule