module fake_jpeg_12324_n_613 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_613);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_613;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_14),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g47 ( 
.A(n_1),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx4f_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx4f_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_9),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_0),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_58),
.Y(n_131)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_59),
.Y(n_141)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_60),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_61),
.Y(n_142)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_62),
.Y(n_152)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_63),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_64),
.Y(n_159)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_65),
.Y(n_161)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_66),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_67),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_36),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g144 ( 
.A(n_68),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_13),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_69),
.B(n_88),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_70),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_16),
.B(n_13),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_71),
.B(n_76),
.Y(n_151)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_72),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_73),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_74),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_75),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_16),
.B(n_13),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_77),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_78),
.Y(n_183)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_79),
.Y(n_160)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_80),
.Y(n_124)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_81),
.Y(n_193)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_82),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx5_ASAP7_75t_L g175 ( 
.A(n_83),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_26),
.B(n_0),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_84),
.B(n_94),
.Y(n_167)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_85),
.Y(n_133)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_86),
.Y(n_185)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_21),
.Y(n_87)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_87),
.Y(n_125)
);

INVx4_ASAP7_75t_SL g88 ( 
.A(n_24),
.Y(n_88)
);

BUFx8_ASAP7_75t_L g89 ( 
.A(n_24),
.Y(n_89)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_89),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_90),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_21),
.Y(n_91)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_91),
.Y(n_154)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_38),
.Y(n_93)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_93),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_26),
.B(n_1),
.Y(n_94)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_32),
.Y(n_95)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_95),
.Y(n_170)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_38),
.Y(n_96)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_96),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_57),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_97),
.A2(n_47),
.B1(n_41),
.B2(n_56),
.Y(n_128)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_17),
.Y(n_98)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_98),
.Y(n_190)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_99),
.Y(n_155)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_19),
.Y(n_100)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_100),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_41),
.B(n_1),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_101),
.B(n_29),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_19),
.Y(n_102)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_102),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_19),
.Y(n_103)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_103),
.Y(n_163)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_30),
.Y(n_104)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_104),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_30),
.Y(n_105)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_105),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_30),
.Y(n_106)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_106),
.Y(n_157)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_34),
.Y(n_107)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_107),
.Y(n_158)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_38),
.Y(n_108)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_108),
.Y(n_164)
);

BUFx12_ASAP7_75t_L g109 ( 
.A(n_24),
.Y(n_109)
);

INVx6_ASAP7_75t_SL g196 ( 
.A(n_109),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_34),
.Y(n_110)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_110),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_34),
.Y(n_111)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_111),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_27),
.B(n_2),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_112),
.B(n_2),
.Y(n_189)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_42),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_113),
.B(n_120),
.Y(n_134)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_42),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_117),
.Y(n_126)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_50),
.Y(n_115)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_115),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_116),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_27),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_118),
.Y(n_199)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_44),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_119),
.B(n_44),
.Y(n_135)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_28),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g121 ( 
.A(n_36),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_121),
.B(n_122),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_49),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_123),
.B(n_135),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_128),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_102),
.A2(n_103),
.B1(n_105),
.B2(n_111),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_132),
.A2(n_90),
.B1(n_77),
.B2(n_75),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_91),
.B(n_55),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_136),
.B(n_169),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_96),
.A2(n_52),
.B1(n_28),
.B2(n_38),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_137),
.A2(n_165),
.B1(n_174),
.B2(n_181),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_117),
.B(n_55),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_139),
.B(n_145),
.Y(n_242)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_106),
.A2(n_52),
.B1(n_28),
.B2(n_54),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_143),
.A2(n_186),
.B1(n_202),
.B2(n_130),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_101),
.B(n_56),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_69),
.B(n_29),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_153),
.B(n_201),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_83),
.B(n_48),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_156),
.B(n_189),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_100),
.A2(n_31),
.B1(n_46),
.B2(n_39),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_109),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_104),
.A2(n_31),
.B1(n_46),
.B2(n_39),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_61),
.B(n_62),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_177),
.B(n_6),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_97),
.A2(n_110),
.B1(n_79),
.B2(n_74),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_178),
.A2(n_198),
.B1(n_12),
.B2(n_202),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_64),
.A2(n_18),
.B1(n_35),
.B2(n_23),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_88),
.B(n_48),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_184),
.B(n_9),
.Y(n_241)
);

OAI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_58),
.A2(n_18),
.B1(n_35),
.B2(n_23),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_116),
.A2(n_54),
.B1(n_43),
.B2(n_37),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_187),
.A2(n_118),
.B1(n_89),
.B2(n_51),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_122),
.B(n_43),
.C(n_37),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_195),
.B(n_167),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_67),
.A2(n_47),
.B1(n_51),
.B2(n_49),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_70),
.B(n_2),
.Y(n_201)
);

OAI22xp33_ASAP7_75t_L g202 ( 
.A1(n_73),
.A2(n_51),
.B1(n_49),
.B2(n_4),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_129),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_204),
.Y(n_281)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_154),
.Y(n_205)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_205),
.Y(n_289)
);

INVx3_ASAP7_75t_SL g207 ( 
.A(n_196),
.Y(n_207)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_207),
.Y(n_300)
);

INVx6_ASAP7_75t_L g208 ( 
.A(n_148),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_208),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_144),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g287 ( 
.A(n_209),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_184),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_210),
.Y(n_298)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_148),
.Y(n_211)
);

INVx5_ASAP7_75t_L g310 ( 
.A(n_211),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_212),
.A2(n_233),
.B1(n_266),
.B2(n_172),
.Y(n_275)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_190),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g331 ( 
.A(n_213),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_214),
.A2(n_265),
.B(n_188),
.Y(n_290)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_158),
.Y(n_215)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_215),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_126),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_216),
.B(n_224),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_170),
.A2(n_49),
.B1(n_51),
.B2(n_4),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_217),
.A2(n_237),
.B1(n_240),
.B2(n_262),
.Y(n_295)
);

OAI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_218),
.A2(n_231),
.B1(n_221),
.B2(n_226),
.Y(n_309)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_200),
.Y(n_220)
);

INVx3_ASAP7_75t_L g279 ( 
.A(n_220),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_221),
.A2(n_142),
.B1(n_193),
.B2(n_161),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_222),
.Y(n_301)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_157),
.Y(n_223)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_223),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_185),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_131),
.Y(n_225)
);

INVx5_ASAP7_75t_L g328 ( 
.A(n_225),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_130),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_226),
.A2(n_268),
.B(n_188),
.Y(n_292)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_160),
.Y(n_227)
);

BUFx2_ASAP7_75t_SL g308 ( 
.A(n_227),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_228),
.B(n_231),
.Y(n_314)
);

BUFx2_ASAP7_75t_SL g229 ( 
.A(n_149),
.Y(n_229)
);

INVx13_ASAP7_75t_L g311 ( 
.A(n_229),
.Y(n_311)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_160),
.Y(n_230)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_230),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_134),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_173),
.Y(n_232)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_232),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_151),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_233)
);

AND2x2_ASAP7_75t_SL g234 ( 
.A(n_124),
.B(n_127),
.Y(n_234)
);

AND2x2_ASAP7_75t_SL g330 ( 
.A(n_234),
.B(n_261),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_131),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_236),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_170),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_141),
.Y(n_238)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_238),
.Y(n_285)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_200),
.Y(n_239)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_239),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_142),
.A2(n_7),
.B1(n_9),
.B2(n_12),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_241),
.B(n_244),
.Y(n_303)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_166),
.Y(n_243)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_243),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_136),
.B(n_9),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_147),
.Y(n_245)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_245),
.Y(n_305)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_168),
.Y(n_246)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_246),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_144),
.Y(n_247)
);

INVx13_ASAP7_75t_L g315 ( 
.A(n_247),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_248),
.A2(n_138),
.B1(n_197),
.B2(n_176),
.Y(n_276)
);

INVx8_ASAP7_75t_L g249 ( 
.A(n_162),
.Y(n_249)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_249),
.Y(n_326)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_175),
.Y(n_250)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_250),
.Y(n_327)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_173),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_251),
.Y(n_278)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_179),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_252),
.B(n_254),
.Y(n_316)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_194),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_253),
.Y(n_312)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_164),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_125),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_255),
.B(n_256),
.Y(n_323)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_125),
.Y(n_256)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_175),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_257),
.B(n_258),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_194),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_134),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_259),
.B(n_260),
.Y(n_291)
);

BUFx8_ASAP7_75t_L g260 ( 
.A(n_152),
.Y(n_260)
);

AND2x2_ASAP7_75t_SL g261 ( 
.A(n_133),
.B(n_155),
.Y(n_261)
);

INVx6_ASAP7_75t_L g262 ( 
.A(n_163),
.Y(n_262)
);

INVx3_ASAP7_75t_SL g263 ( 
.A(n_163),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_263),
.A2(n_271),
.B1(n_272),
.B2(n_273),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_140),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_264),
.B(n_270),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_187),
.A2(n_12),
.B(n_181),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_132),
.A2(n_12),
.B1(n_174),
.B2(n_165),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_182),
.B(n_140),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_267),
.B(n_261),
.Y(n_322)
);

AO22x1_ASAP7_75t_L g268 ( 
.A1(n_143),
.A2(n_186),
.B1(n_193),
.B2(n_137),
.Y(n_268)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_144),
.Y(n_270)
);

INVx11_ASAP7_75t_L g271 ( 
.A(n_159),
.Y(n_271)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_183),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_192),
.Y(n_273)
);

INVx6_ASAP7_75t_L g274 ( 
.A(n_172),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_197),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_275),
.B(n_292),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_276),
.A2(n_283),
.B1(n_309),
.B2(n_261),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_265),
.A2(n_199),
.B1(n_138),
.B2(n_176),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_282),
.A2(n_286),
.B1(n_225),
.B2(n_236),
.Y(n_350)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_284),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_268),
.A2(n_161),
.B1(n_191),
.B2(n_171),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g288 ( 
.A1(n_218),
.A2(n_162),
.B1(n_171),
.B2(n_180),
.Y(n_288)
);

OA22x2_ASAP7_75t_L g349 ( 
.A1(n_288),
.A2(n_294),
.B1(n_319),
.B2(n_324),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_290),
.A2(n_240),
.B(n_260),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_L g294 ( 
.A1(n_210),
.A2(n_180),
.B1(n_191),
.B2(n_150),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_228),
.B(n_150),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_296),
.B(n_297),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_244),
.B(n_146),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_269),
.B(n_146),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_299),
.B(n_313),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_241),
.B(n_234),
.Y(n_313)
);

AOI22xp33_ASAP7_75t_L g319 ( 
.A1(n_267),
.A2(n_219),
.B1(n_206),
.B2(n_214),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_322),
.B(n_303),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_L g324 ( 
.A1(n_206),
.A2(n_258),
.B1(n_274),
.B2(n_208),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_298),
.A2(n_207),
.B1(n_263),
.B2(n_230),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_332),
.Y(n_399)
);

INVx6_ASAP7_75t_L g333 ( 
.A(n_320),
.Y(n_333)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_333),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_334),
.A2(n_335),
.B1(n_339),
.B2(n_364),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_276),
.A2(n_234),
.B1(n_242),
.B2(n_251),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_277),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_336),
.B(n_340),
.Y(n_378)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_331),
.Y(n_338)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_338),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_330),
.A2(n_253),
.B1(n_232),
.B2(n_249),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_316),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_296),
.B(n_235),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_343),
.B(n_347),
.Y(n_387)
);

OAI22xp33_ASAP7_75t_SL g344 ( 
.A1(n_286),
.A2(n_237),
.B1(n_227),
.B2(n_217),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_344),
.A2(n_350),
.B1(n_359),
.B2(n_367),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_314),
.B(n_203),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_345),
.B(n_352),
.C(n_371),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_299),
.B(n_272),
.Y(n_346)
);

INVxp33_ASAP7_75t_L g396 ( 
.A(n_346),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_330),
.B(n_211),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_331),
.Y(n_348)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_348),
.Y(n_380)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_331),
.Y(n_351)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_351),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_313),
.B(n_270),
.C(n_271),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_353),
.B(n_362),
.Y(n_389)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_284),
.Y(n_354)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_354),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_L g355 ( 
.A1(n_298),
.A2(n_262),
.B1(n_239),
.B2(n_257),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_355),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g402 ( 
.A(n_356),
.B(n_369),
.Y(n_402)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_310),
.Y(n_358)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_358),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_275),
.A2(n_220),
.B1(n_250),
.B2(n_247),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_L g360 ( 
.A1(n_283),
.A2(n_209),
.B1(n_260),
.B2(n_306),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g400 ( 
.A(n_360),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_287),
.Y(n_361)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_361),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_323),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_330),
.B(n_297),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_363),
.B(n_365),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_292),
.A2(n_322),
.B1(n_290),
.B2(n_282),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_303),
.B(n_301),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_301),
.B(n_291),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_366),
.B(n_374),
.Y(n_393)
);

OAI22xp33_ASAP7_75t_SL g367 ( 
.A1(n_295),
.A2(n_281),
.B1(n_300),
.B2(n_326),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_281),
.A2(n_278),
.B1(n_312),
.B2(n_326),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_368),
.A2(n_370),
.B1(n_308),
.B2(n_280),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_300),
.B(n_305),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_278),
.A2(n_312),
.B1(n_305),
.B2(n_285),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_285),
.B(n_325),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_327),
.B(n_289),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_372),
.B(n_373),
.Y(n_395)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_321),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_327),
.B(n_289),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_321),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_375),
.B(n_329),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_370),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_377),
.B(n_385),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_364),
.A2(n_334),
.B1(n_354),
.B2(n_337),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_384),
.A2(n_397),
.B1(n_401),
.B2(n_407),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_372),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_357),
.A2(n_310),
.B1(n_320),
.B2(n_317),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g433 ( 
.A1(n_388),
.A2(n_351),
.B1(n_348),
.B2(n_362),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_374),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_392),
.B(n_394),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_369),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_337),
.A2(n_318),
.B1(n_320),
.B2(n_317),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_398),
.B(n_350),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_335),
.A2(n_328),
.B1(n_280),
.B2(n_302),
.Y(n_401)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_404),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_363),
.B(n_304),
.C(n_329),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_405),
.B(n_406),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_341),
.B(n_304),
.C(n_307),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_342),
.A2(n_328),
.B1(n_302),
.B2(n_279),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_368),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_409),
.B(n_410),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_366),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_342),
.B(n_311),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_412),
.B(n_375),
.Y(n_439)
);

OAI32xp33_ASAP7_75t_L g413 ( 
.A1(n_390),
.A2(n_386),
.A3(n_387),
.B1(n_384),
.B2(n_402),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_413),
.B(n_416),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_SL g414 ( 
.A1(n_391),
.A2(n_357),
.B1(n_353),
.B2(n_359),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_414),
.A2(n_427),
.B(n_435),
.Y(n_460)
);

INVxp33_ASAP7_75t_L g415 ( 
.A(n_378),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_415),
.B(n_432),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_389),
.Y(n_416)
);

OAI32xp33_ASAP7_75t_L g417 ( 
.A1(n_390),
.A2(n_341),
.A3(n_356),
.B1(n_347),
.B2(n_365),
.Y(n_417)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_417),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_382),
.A2(n_389),
.B1(n_409),
.B2(n_377),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_418),
.A2(n_433),
.B1(n_385),
.B2(n_392),
.Y(n_464)
);

NAND4xp25_ASAP7_75t_SL g419 ( 
.A(n_378),
.B(n_315),
.C(n_287),
.D(n_361),
.Y(n_419)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_419),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_382),
.A2(n_357),
.B(n_352),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_420),
.A2(n_442),
.B(n_445),
.Y(n_479)
);

CKINVDCx16_ASAP7_75t_R g421 ( 
.A(n_404),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_421),
.B(n_434),
.Y(n_453)
);

MAJx2_ASAP7_75t_L g424 ( 
.A(n_403),
.B(n_345),
.C(n_343),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_424),
.B(n_403),
.C(n_412),
.Y(n_452)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_426),
.Y(n_458)
);

OA21x2_ASAP7_75t_L g427 ( 
.A1(n_391),
.A2(n_339),
.B(n_349),
.Y(n_427)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_380),
.Y(n_430)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_430),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_395),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_410),
.B(n_336),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_388),
.B(n_349),
.Y(n_435)
);

OA22x2_ASAP7_75t_L g436 ( 
.A1(n_382),
.A2(n_349),
.B1(n_340),
.B2(n_338),
.Y(n_436)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_436),
.Y(n_468)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_380),
.Y(n_437)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_437),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_384),
.A2(n_349),
.B1(n_371),
.B2(n_358),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g455 ( 
.A1(n_438),
.A2(n_447),
.B1(n_400),
.B2(n_423),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_SL g473 ( 
.A(n_439),
.B(n_395),
.Y(n_473)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_379),
.Y(n_440)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_440),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_402),
.B(n_373),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_441),
.B(n_443),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_399),
.A2(n_279),
.B(n_293),
.Y(n_442)
);

CKINVDCx16_ASAP7_75t_R g443 ( 
.A(n_393),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_396),
.B(n_287),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_444),
.Y(n_463)
);

A2O1A1Ixp33_ASAP7_75t_SL g445 ( 
.A1(n_388),
.A2(n_315),
.B(n_287),
.C(n_311),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_381),
.Y(n_446)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_446),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_411),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_424),
.B(n_403),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_449),
.B(n_454),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_438),
.A2(n_386),
.B1(n_400),
.B2(n_387),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_451),
.A2(n_455),
.B1(n_427),
.B2(n_435),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_452),
.B(n_476),
.C(n_462),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_428),
.B(n_412),
.Y(n_454)
);

XNOR2x2_ASAP7_75t_L g457 ( 
.A(n_418),
.B(n_393),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g502 ( 
.A(n_457),
.B(n_473),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_428),
.B(n_405),
.Y(n_461)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_461),
.B(n_462),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_439),
.B(n_405),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g481 ( 
.A1(n_464),
.A2(n_478),
.B1(n_468),
.B2(n_458),
.Y(n_481)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_417),
.B(n_406),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_465),
.B(n_471),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_429),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_467),
.B(n_432),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_431),
.B(n_406),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_L g474 ( 
.A1(n_416),
.A2(n_394),
.B(n_398),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g500 ( 
.A1(n_474),
.A2(n_446),
.B(n_430),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_420),
.B(n_381),
.C(n_407),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_443),
.A2(n_383),
.B1(n_401),
.B2(n_379),
.Y(n_477)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_477),
.Y(n_482)
);

OR2x2_ASAP7_75t_L g478 ( 
.A(n_433),
.B(n_401),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_478),
.Y(n_501)
);

INVx13_ASAP7_75t_L g480 ( 
.A(n_450),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_480),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_481),
.A2(n_506),
.B1(n_507),
.B2(n_472),
.Y(n_512)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_483),
.Y(n_526)
);

BUFx24_ASAP7_75t_SL g484 ( 
.A(n_463),
.Y(n_484)
);

BUFx24_ASAP7_75t_SL g513 ( 
.A(n_484),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_475),
.B(n_413),
.Y(n_485)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_485),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_453),
.B(n_421),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_486),
.B(n_493),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_487),
.B(n_458),
.Y(n_523)
);

NAND2x1_ASAP7_75t_SL g490 ( 
.A(n_476),
.B(n_422),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_490),
.A2(n_500),
.B(n_479),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_449),
.B(n_422),
.C(n_414),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_491),
.B(n_508),
.C(n_461),
.Y(n_510)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_448),
.Y(n_492)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_492),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_465),
.B(n_411),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_450),
.B(n_425),
.Y(n_494)
);

CKINVDCx16_ASAP7_75t_R g511 ( 
.A(n_494),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_SL g495 ( 
.A(n_456),
.B(n_437),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_495),
.B(n_498),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_SL g524 ( 
.A1(n_496),
.A2(n_499),
.B1(n_503),
.B2(n_436),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_479),
.A2(n_474),
.B(n_460),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_497),
.A2(n_460),
.B(n_464),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_456),
.B(n_466),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g499 ( 
.A1(n_451),
.A2(n_427),
.B1(n_435),
.B2(n_426),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_468),
.A2(n_436),
.B1(n_397),
.B2(n_423),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_470),
.B(n_447),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_505),
.Y(n_522)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_459),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_459),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_452),
.B(n_436),
.C(n_408),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_510),
.B(n_529),
.Y(n_551)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_512),
.Y(n_540)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_514),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_489),
.B(n_454),
.C(n_471),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_515),
.B(n_521),
.C(n_523),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_SL g535 ( 
.A1(n_516),
.A2(n_497),
.B(n_501),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_489),
.B(n_466),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g544 ( 
.A(n_518),
.B(n_519),
.Y(n_544)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_488),
.B(n_457),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_487),
.B(n_473),
.C(n_470),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_524),
.A2(n_532),
.B1(n_481),
.B2(n_500),
.Y(n_541)
);

XOR2xp5_ASAP7_75t_L g525 ( 
.A(n_488),
.B(n_397),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g546 ( 
.A(n_525),
.B(n_528),
.Y(n_546)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_504),
.B(n_442),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_504),
.B(n_472),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_508),
.B(n_469),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_530),
.B(n_494),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_496),
.A2(n_503),
.B1(n_499),
.B2(n_482),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_SL g533 ( 
.A(n_526),
.B(n_486),
.Y(n_533)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_533),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_527),
.B(n_492),
.Y(n_534)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_534),
.Y(n_565)
);

MAJx2_ASAP7_75t_L g560 ( 
.A(n_535),
.B(n_445),
.C(n_440),
.Y(n_560)
);

CKINVDCx16_ASAP7_75t_R g536 ( 
.A(n_509),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_536),
.B(n_537),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g539 ( 
.A(n_523),
.B(n_491),
.C(n_482),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_539),
.B(n_550),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_L g555 ( 
.A1(n_541),
.A2(n_532),
.B1(n_518),
.B2(n_528),
.Y(n_555)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_531),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_542),
.B(n_548),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_512),
.A2(n_485),
.B1(n_495),
.B2(n_501),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g559 ( 
.A1(n_543),
.A2(n_545),
.B1(n_547),
.B2(n_552),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_SL g545 ( 
.A1(n_516),
.A2(n_490),
.B1(n_505),
.B2(n_506),
.Y(n_545)
);

OAI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_514),
.A2(n_490),
.B1(n_507),
.B2(n_502),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_522),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_521),
.B(n_510),
.C(n_515),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_511),
.A2(n_520),
.B1(n_517),
.B2(n_524),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_550),
.B(n_530),
.C(n_529),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_553),
.B(n_556),
.Y(n_572)
);

XOR2xp5_ASAP7_75t_L g554 ( 
.A(n_546),
.B(n_525),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g575 ( 
.A(n_554),
.B(n_567),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_555),
.A2(n_569),
.B1(n_533),
.B2(n_542),
.Y(n_577)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_551),
.B(n_538),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_SL g557 ( 
.A1(n_547),
.A2(n_519),
.B1(n_502),
.B2(n_469),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_SL g579 ( 
.A1(n_557),
.A2(n_559),
.B1(n_563),
.B2(n_567),
.Y(n_579)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_560),
.Y(n_581)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_551),
.B(n_408),
.Y(n_561)
);

XNOR2xp5_ASAP7_75t_L g580 ( 
.A(n_561),
.B(n_566),
.Y(n_580)
);

AOI21xp5_ASAP7_75t_L g563 ( 
.A1(n_535),
.A2(n_549),
.B(n_540),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g582 ( 
.A1(n_563),
.A2(n_559),
.B1(n_557),
.B2(n_534),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_538),
.B(n_376),
.C(n_445),
.Y(n_566)
);

XOR2x1_ASAP7_75t_L g567 ( 
.A(n_543),
.B(n_480),
.Y(n_567)
);

INVx13_ASAP7_75t_L g569 ( 
.A(n_548),
.Y(n_569)
);

MAJIxp5_ASAP7_75t_L g570 ( 
.A(n_568),
.B(n_556),
.C(n_553),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_570),
.B(n_574),
.Y(n_586)
);

NOR2x1_ASAP7_75t_R g571 ( 
.A(n_565),
.B(n_549),
.Y(n_571)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_571),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_SL g573 ( 
.A1(n_566),
.A2(n_545),
.B1(n_540),
.B2(n_539),
.Y(n_573)
);

XNOR2xp5_ASAP7_75t_L g591 ( 
.A(n_573),
.B(n_579),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g574 ( 
.A(n_561),
.B(n_541),
.C(n_546),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_SL g576 ( 
.A(n_562),
.B(n_513),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_576),
.B(n_578),
.Y(n_590)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_577),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_558),
.B(n_544),
.Y(n_578)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_582),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_SL g583 ( 
.A1(n_581),
.A2(n_564),
.B1(n_560),
.B2(n_569),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g597 ( 
.A1(n_583),
.A2(n_584),
.B1(n_573),
.B2(n_575),
.Y(n_597)
);

INVx11_ASAP7_75t_L g584 ( 
.A(n_571),
.Y(n_584)
);

CKINVDCx20_ASAP7_75t_R g585 ( 
.A(n_570),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_585),
.B(n_592),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_572),
.B(n_554),
.C(n_544),
.Y(n_592)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_590),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_594),
.B(n_595),
.Y(n_603)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_583),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_586),
.B(n_564),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_596),
.B(n_597),
.Y(n_600)
);

OAI21x1_ASAP7_75t_L g598 ( 
.A1(n_584),
.A2(n_578),
.B(n_575),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_598),
.B(n_599),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_587),
.B(n_574),
.Y(n_599)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_593),
.B(n_599),
.C(n_589),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_601),
.B(n_587),
.C(n_588),
.Y(n_604)
);

AOI21xp5_ASAP7_75t_L g607 ( 
.A1(n_604),
.A2(n_605),
.B(n_606),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_603),
.B(n_589),
.C(n_591),
.Y(n_605)
);

AOI21xp33_ASAP7_75t_L g606 ( 
.A1(n_602),
.A2(n_591),
.B(n_592),
.Y(n_606)
);

A2O1A1Ixp33_ASAP7_75t_L g608 ( 
.A1(n_604),
.A2(n_600),
.B(n_580),
.C(n_419),
.Y(n_608)
);

OAI21xp5_ASAP7_75t_L g609 ( 
.A1(n_608),
.A2(n_445),
.B(n_376),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_609),
.Y(n_610)
);

OAI21xp5_ASAP7_75t_SL g611 ( 
.A1(n_610),
.A2(n_607),
.B(n_445),
.Y(n_611)
);

O2A1O1Ixp33_ASAP7_75t_SL g612 ( 
.A1(n_611),
.A2(n_383),
.B(n_333),
.C(n_293),
.Y(n_612)
);

XNOR2xp5_ASAP7_75t_L g613 ( 
.A(n_612),
.B(n_307),
.Y(n_613)
);


endmodule