module fake_ariane_2027_n_106 (n_8, n_3, n_2, n_11, n_7, n_16, n_5, n_14, n_1, n_0, n_12, n_15, n_6, n_13, n_9, n_4, n_10, n_106);

input n_8;
input n_3;
input n_2;
input n_11;
input n_7;
input n_16;
input n_5;
input n_14;
input n_1;
input n_0;
input n_12;
input n_15;
input n_6;
input n_13;
input n_9;
input n_4;
input n_10;

output n_106;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_90;
wire n_38;
wire n_47;
wire n_18;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_34;
wire n_69;
wire n_95;
wire n_92;
wire n_98;
wire n_74;
wire n_33;
wire n_19;
wire n_40;
wire n_53;
wire n_21;
wire n_66;
wire n_71;
wire n_24;
wire n_96;
wire n_49;
wire n_20;
wire n_100;
wire n_17;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_103;
wire n_79;
wire n_26;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_72;
wire n_105;
wire n_44;
wire n_30;
wire n_82;
wire n_31;
wire n_42;
wire n_57;
wire n_70;
wire n_85;
wire n_48;
wire n_94;
wire n_101;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_93;
wire n_23;
wire n_61;
wire n_102;
wire n_22;
wire n_43;
wire n_81;
wire n_87;
wire n_27;
wire n_29;
wire n_41;
wire n_55;
wire n_28;
wire n_80;
wire n_97;
wire n_88;
wire n_68;
wire n_104;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_99;
wire n_35;
wire n_54;
wire n_25;

CKINVDCx14_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx5p33_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVxp33_ASAP7_75t_SL g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx2_ASAP7_75t_SL g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx2_ASAP7_75t_SL g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_22),
.B(n_2),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_18),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_37),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_30),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx4f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_17),
.B1(n_18),
.B2(n_26),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_25),
.Y(n_54)
);

OAI21x1_ASAP7_75t_L g55 ( 
.A1(n_48),
.A2(n_40),
.B(n_44),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_46),
.A2(n_44),
.B(n_40),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_52),
.A2(n_41),
.B1(n_39),
.B2(n_34),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_38),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_50),
.A2(n_36),
.B(n_39),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_50),
.A2(n_48),
.B(n_53),
.Y(n_60)
);

AND2x4_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_58),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_54),
.Y(n_62)
);

AND2x4_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_45),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_60),
.A2(n_51),
.B(n_47),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_43),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_43),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_66),
.Y(n_67)
);

AND2x4_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_23),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_39),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_65),
.Y(n_71)
);

OAI21x1_ASAP7_75t_L g72 ( 
.A1(n_69),
.A2(n_64),
.B(n_62),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_68),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

BUFx8_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_20),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_74),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_76),
.B(n_67),
.Y(n_79)
);

NAND2xp33_ASAP7_75t_R g80 ( 
.A(n_75),
.B(n_63),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_79),
.Y(n_81)
);

AOI222xp33_ASAP7_75t_L g82 ( 
.A1(n_77),
.A2(n_25),
.B1(n_21),
.B2(n_63),
.C1(n_20),
.C2(n_76),
.Y(n_82)
);

NOR3xp33_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_71),
.C(n_61),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_80),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_61),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_84),
.A2(n_27),
.B(n_39),
.C(n_72),
.Y(n_87)
);

AOI211xp5_ASAP7_75t_SL g88 ( 
.A1(n_81),
.A2(n_27),
.B(n_3),
.C(n_6),
.Y(n_88)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

NAND3xp33_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_39),
.C(n_42),
.Y(n_90)
);

NOR3xp33_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_89),
.C(n_87),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

AOI21xp33_ASAP7_75t_SL g93 ( 
.A1(n_89),
.A2(n_2),
.B(n_6),
.Y(n_93)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_84),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_89),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_94),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_92),
.A2(n_85),
.B(n_86),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_95),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_93),
.Y(n_99)
);

NAND3xp33_ASAP7_75t_SL g100 ( 
.A(n_99),
.B(n_91),
.C(n_42),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_101),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_100),
.B(n_42),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_102),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_104),
.Y(n_105)
);

AOI221xp5_ASAP7_75t_L g106 ( 
.A1(n_105),
.A2(n_103),
.B1(n_42),
.B2(n_9),
.C(n_11),
.Y(n_106)
);


endmodule