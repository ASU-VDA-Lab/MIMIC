module fake_netlist_1_3970_n_32 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_32);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_32;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx1_ASAP7_75t_L g12 ( .A(n_1), .Y(n_12) );
BUFx2_ASAP7_75t_L g13 ( .A(n_10), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_8), .Y(n_14) );
CKINVDCx8_ASAP7_75t_R g15 ( .A(n_5), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_7), .Y(n_16) );
OR2x6_ASAP7_75t_L g17 ( .A(n_4), .B(n_1), .Y(n_17) );
NAND2xp5_ASAP7_75t_SL g18 ( .A(n_13), .B(n_0), .Y(n_18) );
NAND2xp5_ASAP7_75t_SL g19 ( .A(n_16), .B(n_0), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
INVx1_ASAP7_75t_L g21 ( .A(n_18), .Y(n_21) );
AND2x4_ASAP7_75t_SL g22 ( .A(n_21), .B(n_17), .Y(n_22) );
OAI21xp5_ASAP7_75t_SL g23 ( .A1(n_22), .A2(n_20), .B(n_12), .Y(n_23) );
NAND2xp5_ASAP7_75t_SL g24 ( .A(n_23), .B(n_14), .Y(n_24) );
NOR2xp33_ASAP7_75t_L g25 ( .A(n_23), .B(n_20), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_25), .Y(n_26) );
AOI22xp5_ASAP7_75t_L g27 ( .A1(n_24), .A2(n_17), .B1(n_14), .B2(n_15), .Y(n_27) );
NAND2xp5_ASAP7_75t_L g28 ( .A(n_26), .B(n_17), .Y(n_28) );
AND4x1_ASAP7_75t_L g29 ( .A(n_27), .B(n_2), .C(n_3), .D(n_4), .Y(n_29) );
AOI22xp5_ASAP7_75t_L g30 ( .A1(n_28), .A2(n_2), .B1(n_3), .B2(n_6), .Y(n_30) );
INVx2_ASAP7_75t_L g31 ( .A(n_30), .Y(n_31) );
AOI22xp33_ASAP7_75t_L g32 ( .A1(n_31), .A2(n_29), .B1(n_9), .B2(n_11), .Y(n_32) );
endmodule