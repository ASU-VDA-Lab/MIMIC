module fake_jpeg_432_n_499 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_499);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_499;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_17),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_17),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_0),
.B(n_10),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_8),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_3),
.Y(n_48)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_16),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_55),
.B(n_87),
.Y(n_181)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_56),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_57),
.Y(n_129)
);

BUFx4f_ASAP7_75t_L g58 ( 
.A(n_25),
.Y(n_58)
);

INVx2_ASAP7_75t_SL g141 ( 
.A(n_58),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_59),
.Y(n_134)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_60),
.Y(n_125)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_61),
.Y(n_197)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_62),
.Y(n_208)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_63),
.Y(n_140)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_64),
.Y(n_187)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_65),
.Y(n_180)
);

BUFx24_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

CKINVDCx6p67_ASAP7_75t_R g123 ( 
.A(n_66),
.Y(n_123)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_67),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_18),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_68),
.B(n_100),
.Y(n_144)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx3_ASAP7_75t_SL g195 ( 
.A(n_69),
.Y(n_195)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_70),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_71),
.Y(n_206)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_72),
.Y(n_163)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_73),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_74),
.Y(n_136)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_75),
.Y(n_174)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_76),
.Y(n_202)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_77),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_16),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_78),
.B(n_83),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_79),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_20),
.A2(n_18),
.B1(n_14),
.B2(n_12),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_80),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_167)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_51),
.Y(n_81)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_81),
.Y(n_190)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_82),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_21),
.B(n_0),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_41),
.Y(n_84)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_84),
.Y(n_184)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_85),
.Y(n_145)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_86),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_0),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_88),
.Y(n_204)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_89),
.Y(n_205)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_90),
.Y(n_156)
);

INVx3_ASAP7_75t_SL g91 ( 
.A(n_29),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_91),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

INVx6_ASAP7_75t_L g199 ( 
.A(n_92),
.Y(n_199)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_19),
.Y(n_93)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_93),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_54),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g160 ( 
.A(n_95),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_20),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_96),
.B(n_97),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_21),
.B(n_1),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_29),
.Y(n_98)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_98),
.Y(n_161)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_31),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g132 ( 
.A(n_99),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_23),
.B(n_1),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_23),
.B(n_1),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_101),
.B(n_114),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_24),
.B(n_1),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_102),
.B(n_95),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_19),
.Y(n_103)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_103),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_44),
.Y(n_104)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_104),
.Y(n_172)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_33),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_105),
.B(n_106),
.Y(n_164)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_33),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_35),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_107),
.Y(n_158)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_19),
.Y(n_108)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_108),
.Y(n_191)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_20),
.Y(n_109)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_109),
.Y(n_207)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_35),
.Y(n_110)
);

BUFx4f_ASAP7_75t_L g151 ( 
.A(n_110),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_44),
.Y(n_111)
);

INVx5_ASAP7_75t_SL g200 ( 
.A(n_111),
.Y(n_200)
);

INVx6_ASAP7_75t_SL g112 ( 
.A(n_49),
.Y(n_112)
);

CKINVDCx12_ASAP7_75t_R g122 ( 
.A(n_112),
.Y(n_122)
);

INVx11_ASAP7_75t_L g113 ( 
.A(n_49),
.Y(n_113)
);

BUFx12_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_45),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_44),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_115),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_44),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_116),
.Y(n_135)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_26),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_117),
.B(n_8),
.Y(n_179)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_52),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_46),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_28),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_119),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_24),
.B(n_9),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_2),
.Y(n_152)
);

BUFx12_ASAP7_75t_L g121 ( 
.A(n_49),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_121),
.B(n_28),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_128),
.Y(n_219)
);

A2O1A1Ixp33_ASAP7_75t_L g130 ( 
.A1(n_55),
.A2(n_27),
.B(n_48),
.C(n_47),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_130),
.B(n_152),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_58),
.A2(n_87),
.B1(n_64),
.B2(n_102),
.Y(n_131)
);

OA22x2_ASAP7_75t_L g279 ( 
.A1(n_131),
.A2(n_146),
.B1(n_150),
.B2(n_154),
.Y(n_279)
);

OR2x4_ASAP7_75t_L g138 ( 
.A(n_78),
.B(n_66),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_138),
.Y(n_226)
);

OAI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_57),
.A2(n_26),
.B1(n_36),
.B2(n_47),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_143),
.A2(n_135),
.B1(n_206),
.B2(n_129),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_67),
.A2(n_26),
.B1(n_36),
.B2(n_27),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_98),
.A2(n_36),
.B1(n_46),
.B2(n_45),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_148),
.A2(n_153),
.B1(n_155),
.B2(n_167),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_91),
.A2(n_48),
.B1(n_43),
.B2(n_30),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_104),
.A2(n_43),
.B1(n_30),
.B2(n_28),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_73),
.A2(n_52),
.B1(n_34),
.B2(n_42),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_79),
.A2(n_52),
.B1(n_34),
.B2(n_42),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_165),
.Y(n_237)
);

OR2x4_ASAP7_75t_L g166 ( 
.A(n_121),
.B(n_42),
.Y(n_166)
);

NAND3xp33_ASAP7_75t_L g248 ( 
.A(n_166),
.B(n_175),
.C(n_183),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_119),
.A2(n_34),
.B1(n_4),
.B2(n_6),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_170),
.A2(n_171),
.B1(n_178),
.B2(n_182),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_111),
.A2(n_2),
.B1(n_4),
.B2(n_6),
.Y(n_171)
);

OA22x2_ASAP7_75t_L g173 ( 
.A1(n_115),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_173),
.B(n_179),
.Y(n_220)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_59),
.B(n_6),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_71),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_176),
.B(n_188),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_74),
.B(n_7),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_177),
.B(n_192),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_90),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_84),
.A2(n_9),
.B1(n_92),
.B2(n_94),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_116),
.A2(n_69),
.B1(n_76),
.B2(n_55),
.Y(n_185)
);

OAI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_185),
.A2(n_154),
.B1(n_155),
.B2(n_203),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_68),
.B(n_55),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_68),
.B(n_55),
.Y(n_192)
);

AND2x2_ASAP7_75t_SL g193 ( 
.A(n_78),
.B(n_68),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_193),
.B(n_194),
.Y(n_234)
);

OA22x2_ASAP7_75t_L g194 ( 
.A1(n_80),
.A2(n_109),
.B1(n_117),
.B2(n_108),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_102),
.B(n_83),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_196),
.B(n_181),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_58),
.A2(n_25),
.B1(n_50),
.B2(n_37),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_203),
.A2(n_166),
.B1(n_123),
.B2(n_141),
.Y(n_222)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_187),
.Y(n_209)
);

BUFx2_ASAP7_75t_L g309 ( 
.A(n_209),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_191),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_210),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_149),
.A2(n_153),
.B1(n_148),
.B2(n_138),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_211),
.A2(n_214),
.B1(n_223),
.B2(n_236),
.Y(n_290)
);

INVx3_ASAP7_75t_SL g213 ( 
.A(n_161),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_213),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_171),
.A2(n_194),
.B1(n_175),
.B2(n_131),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_151),
.Y(n_215)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_215),
.Y(n_283)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_141),
.Y(n_216)
);

BUFx3_ASAP7_75t_L g316 ( 
.A(n_216),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_164),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_217),
.B(n_221),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_193),
.B(n_144),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_218),
.B(n_231),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_123),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_222),
.A2(n_235),
.B1(n_273),
.B2(n_274),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_224),
.B(n_227),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_162),
.B(n_189),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_130),
.B(n_205),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_228),
.B(n_257),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g229 ( 
.A(n_195),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_229),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_140),
.B(n_126),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_230),
.B(n_246),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_132),
.B(n_163),
.C(n_204),
.Y(n_231)
);

INVx5_ASAP7_75t_L g232 ( 
.A(n_123),
.Y(n_232)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_232),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_158),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_233),
.B(n_238),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_151),
.A2(n_169),
.B1(n_168),
.B2(n_124),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_147),
.Y(n_238)
);

AO22x2_ASAP7_75t_SL g239 ( 
.A1(n_143),
.A2(n_194),
.B1(n_173),
.B2(n_125),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_L g292 ( 
.A1(n_239),
.A2(n_211),
.B1(n_219),
.B2(n_257),
.Y(n_292)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_139),
.Y(n_240)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_240),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_147),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_241),
.B(n_244),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_174),
.B(n_201),
.C(n_197),
.Y(n_243)
);

MAJx2_ASAP7_75t_L g297 ( 
.A(n_243),
.B(n_262),
.C(n_280),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_137),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_145),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_245),
.B(n_258),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_196),
.B(n_190),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_139),
.Y(n_247)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_247),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_198),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_249),
.B(n_255),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_251),
.A2(n_253),
.B1(n_261),
.B2(n_221),
.Y(n_308)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_187),
.Y(n_252)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_252),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_L g253 ( 
.A1(n_207),
.A2(n_172),
.B1(n_173),
.B2(n_208),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_159),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_254),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_198),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_186),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_256),
.B(n_260),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_128),
.B(n_158),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_195),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_122),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_259),
.B(n_268),
.Y(n_301)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_157),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_161),
.A2(n_186),
.B1(n_129),
.B2(n_134),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_180),
.B(n_133),
.C(n_156),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_202),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_263),
.B(n_264),
.Y(n_313)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_157),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_180),
.B(n_133),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_265),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_156),
.B(n_136),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_266),
.Y(n_298)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_136),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_267),
.B(n_269),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_202),
.B(n_199),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_184),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_184),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_270),
.B(n_271),
.Y(n_307)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_199),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_134),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_272),
.B(n_275),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g273 ( 
.A1(n_146),
.A2(n_178),
.B1(n_160),
.B2(n_127),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_127),
.A2(n_160),
.B1(n_200),
.B2(n_206),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_200),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_127),
.A2(n_166),
.B1(n_138),
.B2(n_58),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g289 ( 
.A1(n_276),
.A2(n_275),
.B1(n_214),
.B2(n_225),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_160),
.B(n_142),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_277),
.A2(n_258),
.B(n_232),
.Y(n_321)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_142),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_278),
.B(n_281),
.Y(n_325)
);

AND2x2_ASAP7_75t_SL g280 ( 
.A(n_142),
.B(n_138),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_123),
.Y(n_281)
);

FAx1_ASAP7_75t_SL g282 ( 
.A(n_218),
.B(n_226),
.CI(n_250),
.CON(n_282),
.SN(n_282)
);

NOR2xp33_ASAP7_75t_SL g337 ( 
.A(n_282),
.B(n_293),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_289),
.A2(n_311),
.B(n_312),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_290),
.A2(n_295),
.B1(n_312),
.B2(n_326),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_292),
.A2(n_299),
.B1(n_328),
.B2(n_298),
.Y(n_341)
);

NOR2x1_ASAP7_75t_L g293 ( 
.A(n_234),
.B(n_228),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_234),
.A2(n_220),
.B1(n_239),
.B2(n_248),
.Y(n_295)
);

OAI22xp33_ASAP7_75t_L g299 ( 
.A1(n_239),
.A2(n_279),
.B1(n_272),
.B2(n_237),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g334 ( 
.A(n_308),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_SL g311 ( 
.A(n_280),
.B(n_234),
.C(n_226),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_220),
.A2(n_239),
.B1(n_242),
.B2(n_279),
.Y(n_312)
);

A2O1A1Ixp33_ASAP7_75t_L g314 ( 
.A1(n_220),
.A2(n_280),
.B(n_212),
.C(n_231),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_314),
.B(n_240),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_243),
.B(n_249),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_318),
.B(n_319),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_255),
.B(n_262),
.Y(n_319)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_321),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_217),
.B(n_269),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_322),
.B(n_244),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_279),
.A2(n_270),
.B1(n_271),
.B2(n_267),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_279),
.A2(n_256),
.B1(n_266),
.B2(n_209),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_266),
.A2(n_215),
.B1(n_213),
.B2(n_263),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_329),
.A2(n_331),
.B1(n_241),
.B2(n_264),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_213),
.A2(n_238),
.B1(n_252),
.B2(n_229),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_265),
.A2(n_277),
.B(n_245),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_277),
.B(n_265),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_333),
.Y(n_390)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_283),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_305),
.B(n_247),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_338),
.B(n_304),
.C(n_317),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_339),
.B(n_354),
.Y(n_377)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_283),
.Y(n_340)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_340),
.Y(n_399)
);

OAI22xp33_ASAP7_75t_L g389 ( 
.A1(n_341),
.A2(n_316),
.B1(n_330),
.B2(n_359),
.Y(n_389)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_309),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_342),
.B(n_343),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_302),
.B(n_260),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_344),
.B(n_347),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_302),
.B(n_216),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_291),
.B(n_259),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_348),
.Y(n_393)
);

BUFx2_ASAP7_75t_L g385 ( 
.A(n_349),
.Y(n_385)
);

A2O1A1Ixp33_ASAP7_75t_SL g350 ( 
.A1(n_299),
.A2(n_278),
.B(n_319),
.C(n_288),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_350),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_291),
.B(n_306),
.Y(n_351)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_351),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_332),
.Y(n_352)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_352),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_286),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_293),
.B(n_318),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_305),
.B(n_322),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_355),
.B(n_287),
.Y(n_388)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_309),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_306),
.B(n_285),
.Y(n_357)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_357),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_358),
.A2(n_364),
.B(n_287),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_290),
.A2(n_328),
.B1(n_292),
.B2(n_326),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_359),
.A2(n_360),
.B1(n_363),
.B2(n_368),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_295),
.A2(n_314),
.B1(n_308),
.B2(n_298),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_307),
.Y(n_361)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_361),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_313),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_L g381 ( 
.A1(n_362),
.A2(n_366),
.B1(n_284),
.B2(n_310),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_296),
.A2(n_311),
.B1(n_297),
.B2(n_327),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_SL g364 ( 
.A1(n_297),
.A2(n_303),
.B(n_282),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_282),
.A2(n_296),
.B1(n_307),
.B2(n_323),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_365),
.A2(n_300),
.B1(n_320),
.B2(n_310),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_313),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_320),
.Y(n_367)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_367),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_327),
.A2(n_320),
.B1(n_329),
.B2(n_301),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_325),
.B(n_315),
.Y(n_369)
);

NOR3xp33_ASAP7_75t_SL g378 ( 
.A(n_369),
.B(n_370),
.C(n_294),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_304),
.B(n_315),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_371),
.B(n_372),
.C(n_373),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g372 ( 
.A(n_355),
.B(n_321),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_338),
.B(n_313),
.C(n_324),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_354),
.B(n_336),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_SL g420 ( 
.A(n_376),
.B(n_382),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_378),
.B(n_337),
.Y(n_402)
);

NOR3xp33_ASAP7_75t_SL g380 ( 
.A(n_337),
.B(n_324),
.C(n_294),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_380),
.B(n_339),
.Y(n_407)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_381),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_384),
.A2(n_352),
.B(n_347),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_345),
.A2(n_287),
.B1(n_309),
.B2(n_331),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_386),
.A2(n_366),
.B1(n_362),
.B2(n_367),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_388),
.B(n_344),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_389),
.A2(n_391),
.B1(n_334),
.B2(n_349),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_341),
.A2(n_334),
.B1(n_360),
.B2(n_336),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_363),
.B(n_330),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_394),
.B(n_398),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_364),
.B(n_316),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g439 ( 
.A(n_400),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_391),
.A2(n_345),
.B1(n_334),
.B2(n_361),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_401),
.A2(n_416),
.B1(n_382),
.B2(n_396),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_402),
.Y(n_434)
);

AO22x1_ASAP7_75t_L g404 ( 
.A1(n_383),
.A2(n_365),
.B1(n_350),
.B2(n_346),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_404),
.B(n_394),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_379),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_405),
.B(n_407),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_397),
.A2(n_350),
.B(n_346),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_390),
.A2(n_350),
.B(n_368),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_410),
.B(n_418),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_411),
.A2(n_423),
.B1(n_401),
.B2(n_404),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_390),
.B(n_333),
.Y(n_414)
);

CKINVDCx14_ASAP7_75t_R g426 ( 
.A(n_414),
.Y(n_426)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_399),
.Y(n_415)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_415),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_383),
.A2(n_343),
.B1(n_353),
.B2(n_369),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_393),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_417),
.B(n_422),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_376),
.B(n_335),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_375),
.A2(n_340),
.B(n_342),
.Y(n_419)
);

INVx3_ASAP7_75t_SL g421 ( 
.A(n_385),
.Y(n_421)
);

MAJx2_ASAP7_75t_L g422 ( 
.A(n_377),
.B(n_356),
.C(n_372),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g423 ( 
.A1(n_385),
.A2(n_395),
.B1(n_386),
.B2(n_392),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_419),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_424),
.B(n_433),
.Y(n_451)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_427),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_416),
.B(n_377),
.Y(n_428)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_428),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_411),
.B(n_393),
.Y(n_429)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_429),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_409),
.A2(n_398),
.B(n_389),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_430),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g447 ( 
.A1(n_431),
.A2(n_412),
.B1(n_421),
.B2(n_414),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_410),
.B(n_387),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_436),
.B(n_438),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_415),
.B(n_374),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_425),
.B(n_413),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_441),
.B(n_443),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_431),
.A2(n_400),
.B1(n_408),
.B2(n_403),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_442),
.A2(n_445),
.B1(n_447),
.B2(n_430),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_425),
.B(n_406),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_437),
.B(n_406),
.C(n_413),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_444),
.B(n_450),
.C(n_371),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_429),
.A2(n_403),
.B1(n_402),
.B2(n_404),
.Y(n_445)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_435),
.Y(n_448)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_448),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_SL g449 ( 
.A(n_428),
.B(n_422),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_449),
.B(n_433),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_437),
.B(n_373),
.C(n_418),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_438),
.Y(n_452)
);

CKINVDCx16_ASAP7_75t_R g468 ( 
.A(n_452),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_457),
.A2(n_467),
.B1(n_455),
.B2(n_451),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_458),
.B(n_463),
.C(n_441),
.Y(n_472)
);

FAx1_ASAP7_75t_SL g459 ( 
.A(n_444),
.B(n_426),
.CI(n_420),
.CON(n_459),
.SN(n_459)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_459),
.B(n_460),
.Y(n_475)
);

CKINVDCx16_ASAP7_75t_R g460 ( 
.A(n_451),
.Y(n_460)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_448),
.Y(n_462)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_462),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_443),
.B(n_420),
.C(n_436),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_SL g478 ( 
.A(n_464),
.B(n_449),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_440),
.A2(n_439),
.B1(n_434),
.B2(n_424),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_465),
.B(n_442),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_453),
.A2(n_439),
.B1(n_426),
.B2(n_432),
.Y(n_466)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_466),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_440),
.A2(n_427),
.B1(n_439),
.B2(n_423),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_471),
.B(n_478),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_472),
.B(n_461),
.Y(n_482)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_456),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_473),
.B(n_476),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_461),
.B(n_458),
.C(n_463),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_474),
.B(n_472),
.C(n_450),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_465),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_477),
.B(n_466),
.Y(n_485)
);

OAI21x1_ASAP7_75t_L g479 ( 
.A1(n_475),
.A2(n_432),
.B(n_446),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_479),
.B(n_454),
.Y(n_489)
);

CKINVDCx14_ASAP7_75t_R g481 ( 
.A(n_475),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g487 ( 
.A(n_481),
.B(n_482),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_SL g486 ( 
.A(n_484),
.B(n_474),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_485),
.B(n_469),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_SL g491 ( 
.A(n_486),
.B(n_488),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_484),
.B(n_482),
.C(n_476),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_489),
.A2(n_490),
.B1(n_488),
.B2(n_468),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_492),
.B(n_480),
.C(n_483),
.Y(n_495)
);

AOI31xp67_ASAP7_75t_L g493 ( 
.A1(n_487),
.A2(n_460),
.A3(n_470),
.B(n_462),
.Y(n_493)
);

NOR3xp33_ASAP7_75t_L g494 ( 
.A(n_493),
.B(n_469),
.C(n_483),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_L g496 ( 
.A1(n_494),
.A2(n_495),
.B(n_491),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_496),
.B(n_480),
.Y(n_497)
);

MAJx2_ASAP7_75t_L g498 ( 
.A(n_497),
.B(n_471),
.C(n_457),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_498),
.Y(n_499)
);


endmodule