module fake_netlist_1_349_n_41 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_41);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_41;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
INVx1_ASAP7_75t_L g11 ( .A(n_6), .Y(n_11) );
BUFx6f_ASAP7_75t_L g12 ( .A(n_5), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_1), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_4), .Y(n_14) );
CKINVDCx20_ASAP7_75t_R g15 ( .A(n_0), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_10), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_1), .Y(n_17) );
INVx6_ASAP7_75t_L g18 ( .A(n_4), .Y(n_18) );
AND2x4_ASAP7_75t_L g19 ( .A(n_14), .B(n_0), .Y(n_19) );
NAND2xp5_ASAP7_75t_L g20 ( .A(n_16), .B(n_2), .Y(n_20) );
AOI22xp33_ASAP7_75t_L g21 ( .A1(n_18), .A2(n_2), .B1(n_3), .B2(n_5), .Y(n_21) );
INVx6_ASAP7_75t_L g22 ( .A(n_18), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_18), .Y(n_23) );
AND3x1_ASAP7_75t_L g24 ( .A(n_11), .B(n_3), .C(n_6), .Y(n_24) );
INVx2_ASAP7_75t_L g25 ( .A(n_22), .Y(n_25) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_23), .B(n_13), .Y(n_26) );
NAND2xp5_ASAP7_75t_L g27 ( .A(n_23), .B(n_17), .Y(n_27) );
AOI22xp33_ASAP7_75t_L g28 ( .A1(n_19), .A2(n_12), .B1(n_15), .B2(n_9), .Y(n_28) );
INVx2_ASAP7_75t_SL g29 ( .A(n_25), .Y(n_29) );
OR2x2_ASAP7_75t_L g30 ( .A(n_26), .B(n_19), .Y(n_30) );
OAI31xp33_ASAP7_75t_L g31 ( .A1(n_28), .A2(n_19), .A3(n_20), .B(n_21), .Y(n_31) );
AND2x2_ASAP7_75t_L g32 ( .A(n_30), .B(n_15), .Y(n_32) );
OR2x2_ASAP7_75t_L g33 ( .A(n_31), .B(n_27), .Y(n_33) );
INVx2_ASAP7_75t_SL g34 ( .A(n_33), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_32), .Y(n_35) );
AOI21xp5_ASAP7_75t_L g36 ( .A1(n_34), .A2(n_29), .B(n_28), .Y(n_36) );
AOI22xp5_ASAP7_75t_L g37 ( .A1(n_34), .A2(n_24), .B1(n_29), .B2(n_22), .Y(n_37) );
AND3x4_ASAP7_75t_L g38 ( .A(n_37), .B(n_35), .C(n_22), .Y(n_38) );
NAND3xp33_ASAP7_75t_SL g39 ( .A(n_36), .B(n_35), .C(n_22), .Y(n_39) );
NAND3xp33_ASAP7_75t_SL g40 ( .A(n_38), .B(n_12), .C(n_7), .Y(n_40) );
AOI22xp33_ASAP7_75t_L g41 ( .A1(n_40), .A2(n_39), .B1(n_12), .B2(n_8), .Y(n_41) );
endmodule