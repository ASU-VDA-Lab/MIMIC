module real_jpeg_19627_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_340, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_340;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_215;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx13_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_1),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_1),
.A2(n_25),
.B1(n_42),
.B2(n_50),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_1),
.A2(n_25),
.B1(n_29),
.B2(n_30),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_1),
.A2(n_25),
.B1(n_45),
.B2(n_46),
.Y(n_195)
);

OAI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_2),
.A2(n_23),
.B1(n_26),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_33),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_2),
.A2(n_33),
.B1(n_45),
.B2(n_46),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_2),
.A2(n_33),
.B1(n_42),
.B2(n_50),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_3),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_3),
.A2(n_45),
.B1(n_46),
.B2(n_115),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_3),
.A2(n_42),
.B1(n_50),
.B2(n_115),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_3),
.A2(n_23),
.B1(n_26),
.B2(n_115),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_4),
.A2(n_23),
.B1(n_26),
.B2(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_4),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_120),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_4),
.A2(n_42),
.B1(n_50),
.B2(n_120),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_4),
.A2(n_45),
.B1(n_46),
.B2(n_120),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_6),
.A2(n_23),
.B1(n_26),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_6),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_6),
.A2(n_42),
.B1(n_50),
.B2(n_55),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_6),
.A2(n_45),
.B1(n_46),
.B2(n_55),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g270 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_55),
.Y(n_270)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_7),
.Y(n_94)
);

INVx8_ASAP7_75t_L g128 ( 
.A(n_7),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_7),
.A2(n_127),
.B(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_7),
.A2(n_158),
.B1(n_159),
.B2(n_161),
.Y(n_157)
);

BUFx8_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_9),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_9),
.A2(n_23),
.B1(n_26),
.B2(n_113),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_9),
.A2(n_45),
.B1(n_46),
.B2(n_113),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_9),
.A2(n_42),
.B1(n_50),
.B2(n_113),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_10),
.Y(n_118)
);

AOI21xp33_ASAP7_75t_L g166 ( 
.A1(n_10),
.A2(n_14),
.B(n_46),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_10),
.A2(n_42),
.B1(n_50),
.B2(n_118),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_10),
.A2(n_93),
.B1(n_174),
.B2(n_175),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_10),
.B(n_75),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_10),
.B(n_30),
.Y(n_203)
);

AOI21xp33_ASAP7_75t_L g207 ( 
.A1(n_10),
.A2(n_30),
.B(n_203),
.Y(n_207)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_12),
.A2(n_23),
.B1(n_26),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_12),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_12),
.A2(n_45),
.B1(n_46),
.B2(n_57),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_12),
.A2(n_42),
.B1(n_50),
.B2(n_57),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g291 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_57),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_13),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_14),
.A2(n_42),
.B(n_43),
.C(n_44),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_14),
.B(n_42),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_14),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_44)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx11_ASAP7_75t_SL g42 ( 
.A(n_15),
.Y(n_42)
);

MAJx2_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_20),
.C(n_337),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_81),
.B(n_335),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_36),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_20),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_31),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_21),
.A2(n_53),
.B(n_253),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_27),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g299 ( 
.A(n_22),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_22),
.A2(n_27),
.B(n_34),
.Y(n_337)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

O2A1O1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_23),
.A2(n_27),
.B(n_28),
.C(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_28),
.Y(n_35)
);

HAxp5_ASAP7_75t_SL g117 ( 
.A(n_23),
.B(n_118),
.CON(n_117),
.SN(n_117)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_27),
.B(n_32),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_27),
.A2(n_34),
.B1(n_117),
.B2(n_119),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_28),
.B(n_30),
.Y(n_124)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_29),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_29),
.A2(n_35),
.B1(n_117),
.B2(n_124),
.Y(n_123)
);

AOI32xp33_ASAP7_75t_L g202 ( 
.A1(n_29),
.A2(n_42),
.A3(n_65),
.B1(n_203),
.B2(n_204),
.Y(n_202)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_30),
.A2(n_63),
.B(n_64),
.C(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_30),
.B(n_64),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_31),
.A2(n_54),
.B(n_58),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_34),
.Y(n_31)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_34),
.A2(n_78),
.B(n_79),
.Y(n_77)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_37),
.B(n_336),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_73),
.C(n_77),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_38),
.A2(n_39),
.B1(n_331),
.B2(n_333),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_39),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_51),
.C(n_59),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_40),
.A2(n_311),
.B1(n_312),
.B2(n_313),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_40),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_40),
.A2(n_59),
.B1(n_60),
.B2(n_311),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_44),
.B(n_48),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_41),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_41),
.A2(n_48),
.B(n_108),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_41),
.A2(n_44),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_41),
.A2(n_44),
.B1(n_170),
.B2(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_41),
.A2(n_44),
.B1(n_192),
.B2(n_210),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_41),
.A2(n_210),
.B(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_41),
.A2(n_44),
.B1(n_100),
.B2(n_245),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_41),
.A2(n_108),
.B(n_245),
.Y(n_279)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_42),
.A2(n_50),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_44),
.A2(n_100),
.B(n_101),
.Y(n_99)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_44),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_44),
.B(n_118),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_45),
.B(n_181),
.Y(n_180)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_46),
.B(n_94),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_47),
.A2(n_50),
.B(n_118),
.C(n_166),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_49),
.B(n_109),
.Y(n_226)
);

NAND2xp33_ASAP7_75t_SL g204 ( 
.A(n_50),
.B(n_64),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_51),
.A2(n_52),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_56),
.B2(n_58),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_53),
.A2(n_58),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_53),
.A2(n_58),
.B1(n_133),
.B2(n_253),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_53),
.A2(n_80),
.B(n_299),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_56),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_58),
.B(n_118),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_67),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_62),
.A2(n_68),
.B(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_63),
.A2(n_69),
.B1(n_112),
.B2(n_114),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_63),
.A2(n_69),
.B1(n_112),
.B2(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_63),
.A2(n_69),
.B1(n_145),
.B2(n_207),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_63),
.B(n_72),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_63),
.A2(n_67),
.B(n_270),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_63),
.A2(n_69),
.B1(n_270),
.B2(n_291),
.Y(n_290)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_66),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_71),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_68),
.A2(n_75),
.B(n_76),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_68),
.A2(n_76),
.B(n_256),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_68),
.A2(n_256),
.B(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_73),
.A2(n_74),
.B1(n_77),
.B2(n_332),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_77),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_328),
.B(n_334),
.Y(n_81)
);

OAI321xp33_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_304),
.A3(n_323),
.B1(n_326),
.B2(n_327),
.C(n_340),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_283),
.B(n_303),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_85),
.A2(n_261),
.B(n_282),
.Y(n_84)
);

O2A1O1Ixp33_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_150),
.B(n_235),
.C(n_260),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_138),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_87),
.B(n_138),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_121),
.B2(n_137),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_105),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_90),
.B(n_105),
.C(n_137),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_92),
.B1(n_99),
.B2(n_104),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_91),
.B(n_104),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_95),
.B(n_96),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_93),
.A2(n_95),
.B1(n_126),
.B2(n_128),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_93),
.B(n_98),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_93),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_93),
.A2(n_160),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_93),
.A2(n_162),
.B(n_194),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_93),
.A2(n_94),
.B(n_278),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_98),
.Y(n_97)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_94),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_94),
.B(n_118),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_97),
.A2(n_158),
.B(n_195),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_99),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_101),
.B(n_226),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_102),
.B(n_109),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_110),
.C(n_116),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_106),
.A2(n_107),
.B1(n_110),
.B2(n_111),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_114),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_SL g139 ( 
.A(n_116),
.B(n_140),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_119),
.Y(n_132)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_121),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_129),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_122),
.B(n_130),
.C(n_135),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_125),
.Y(n_122)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_123),
.B(n_125),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_134),
.B2(n_135),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_141),
.C(n_143),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_139),
.B(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_141),
.A2(n_142),
.B1(n_143),
.B2(n_232),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_143),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_146),
.C(n_147),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_144),
.B(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_146),
.A2(n_147),
.B1(n_148),
.B2(n_221),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_146),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_149),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_151),
.B(n_234),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_228),
.B(n_233),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_215),
.B(n_227),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_197),
.B(n_214),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_184),
.B(n_196),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_171),
.B(n_183),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_163),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_163),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_167),
.B2(n_168),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_165),
.B(n_167),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_172),
.A2(n_178),
.B(n_182),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_177),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_173),
.B(n_177),
.Y(n_182)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_185),
.B(n_186),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_193),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_191),
.C(n_193),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_194),
.B(n_243),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_195),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_198),
.B(n_199),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_205),
.B1(n_212),
.B2(n_213),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_200),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_201),
.B(n_202),
.Y(n_224)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_205),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_208),
.B1(n_209),
.B2(n_211),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_206),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_208),
.B(n_211),
.C(n_212),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_216),
.B(n_217),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_222),
.B2(n_223),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_218),
.B(n_224),
.C(n_225),
.Y(n_229)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_229),
.B(n_230),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_236),
.B(n_237),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_258),
.B2(n_259),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_241),
.B1(n_246),
.B2(n_247),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_247),
.C(n_259),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_244),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_242),
.B(n_244),
.Y(n_267)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_250),
.B2(n_257),
.Y(n_247)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_248),
.Y(n_257)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_254),
.B2(n_255),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_251),
.B(n_255),
.C(n_257),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_255),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g259 ( 
.A(n_258),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_262),
.B(n_263),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_281),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_274),
.B2(n_275),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_275),
.C(n_281),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_267),
.B(n_271),
.C(n_273),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_269),
.A2(n_271),
.B1(n_272),
.B2(n_273),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_269),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g274 ( 
.A(n_275),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_277),
.B1(n_279),
.B2(n_280),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_276),
.A2(n_277),
.B1(n_298),
.B2(n_300),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_276),
.A2(n_294),
.B(n_298),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_277),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_279),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_279),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_284),
.B(n_285),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_301),
.B2(n_302),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_293),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_288),
.B(n_293),
.C(n_302),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_290),
.B(n_292),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_289),
.B(n_290),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_291),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_306),
.C(n_315),
.Y(n_305)
);

FAx1_ASAP7_75t_SL g325 ( 
.A(n_292),
.B(n_306),
.CI(n_315),
.CON(n_325),
.SN(n_325)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_295),
.B1(n_296),
.B2(n_297),
.Y(n_293)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_298),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_301),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_316),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_305),
.B(n_316),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_308),
.B1(n_309),
.B2(n_310),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_307),
.A2(n_308),
.B1(n_318),
.B2(n_321),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_308),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_308),
.B(n_311),
.C(n_313),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_308),
.B(n_321),
.C(n_322),
.Y(n_329)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_313),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_322),
.Y(n_316)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_318),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_320),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_324),
.B(n_325),
.Y(n_326)
);

BUFx24_ASAP7_75t_SL g338 ( 
.A(n_325),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_329),
.B(n_330),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_331),
.Y(n_333)
);


endmodule