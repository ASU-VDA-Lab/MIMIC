module real_jpeg_32073_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_578;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_412;
wire n_155;
wire n_586;
wire n_405;
wire n_572;
wire n_548;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g135 ( 
.A(n_0),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_0),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_0),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_1),
.A2(n_227),
.B1(n_228),
.B2(n_231),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_1),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_1),
.A2(n_227),
.B1(n_385),
.B2(n_390),
.Y(n_384)
);

AOI22xp33_ASAP7_75t_SL g477 ( 
.A1(n_1),
.A2(n_227),
.B1(n_478),
.B2(n_481),
.Y(n_477)
);

AOI22xp33_ASAP7_75t_SL g517 ( 
.A1(n_1),
.A2(n_227),
.B1(n_518),
.B2(n_524),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_2),
.Y(n_97)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_2),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_3),
.A2(n_104),
.B1(n_105),
.B2(n_111),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_3),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_3),
.A2(n_104),
.B1(n_349),
.B2(n_352),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_SL g456 ( 
.A1(n_3),
.A2(n_104),
.B1(n_246),
.B2(n_457),
.Y(n_456)
);

AOI22xp33_ASAP7_75t_SL g498 ( 
.A1(n_3),
.A2(n_104),
.B1(n_499),
.B2(n_504),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_4),
.Y(n_593)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_5),
.A2(n_148),
.B1(n_151),
.B2(n_152),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_5),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_5),
.A2(n_152),
.B1(n_276),
.B2(n_277),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_6),
.A2(n_81),
.B1(n_86),
.B2(n_87),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_6),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_6),
.A2(n_68),
.B1(n_86),
.B2(n_238),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_6),
.A2(n_86),
.B1(n_370),
.B2(n_372),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_6),
.A2(n_86),
.B1(n_452),
.B2(n_453),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_7),
.B(n_337),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_7),
.Y(n_381)
);

NAND2xp33_ASAP7_75t_SL g422 ( 
.A(n_7),
.B(n_90),
.Y(n_422)
);

OAI32xp33_ASAP7_75t_L g429 ( 
.A1(n_7),
.A2(n_430),
.A3(n_433),
.B1(n_437),
.B2(n_443),
.Y(n_429)
);

OAI32xp33_ASAP7_75t_L g475 ( 
.A1(n_7),
.A2(n_430),
.A3(n_433),
.B1(n_437),
.B2(n_443),
.Y(n_475)
);

AOI22xp33_ASAP7_75t_SL g483 ( 
.A1(n_7),
.A2(n_381),
.B1(n_484),
.B2(n_485),
.Y(n_483)
);

OAI21xp33_ASAP7_75t_L g563 ( 
.A1(n_7),
.A2(n_128),
.B(n_509),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_8),
.A2(n_60),
.B1(n_64),
.B2(n_65),
.Y(n_59)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_8),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_8),
.A2(n_64),
.B1(n_218),
.B2(n_220),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_8),
.A2(n_64),
.B1(n_265),
.B2(n_267),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_8),
.A2(n_64),
.B1(n_413),
.B2(n_417),
.Y(n_412)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_9),
.A2(n_68),
.B1(n_70),
.B2(n_71),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_9),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_9),
.A2(n_70),
.B1(n_181),
.B2(n_186),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_9),
.A2(n_70),
.B1(n_315),
.B2(n_318),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_10),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_10),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_10),
.Y(n_233)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_12),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_12),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_12),
.Y(n_150)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_12),
.Y(n_523)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_13),
.Y(n_159)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_13),
.Y(n_167)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_13),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_SL g19 ( 
.A1(n_14),
.A2(n_20),
.B(n_592),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_14),
.B(n_593),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_15),
.A2(n_137),
.B1(n_140),
.B2(n_141),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_15),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_15),
.A2(n_140),
.B1(n_246),
.B2(n_250),
.Y(n_245)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_16),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_16),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_16),
.Y(n_249)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_17),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_17),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_18),
.A2(n_191),
.B1(n_195),
.B2(n_196),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_18),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_18),
.A2(n_195),
.B1(n_210),
.B2(n_212),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_18),
.A2(n_195),
.B1(n_283),
.B2(n_287),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_297),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_294),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_256),
.Y(n_23)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_24),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_200),
.C(n_242),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

XNOR2x1_ASAP7_75t_L g301 ( 
.A(n_26),
.B(n_302),
.Y(n_301)
);

XNOR2x1_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_125),
.Y(n_26)
);

OAI21x1_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_76),
.B(n_124),
.Y(n_27)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_28),
.Y(n_293)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_30),
.B(n_78),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_59),
.B1(n_66),
.B2(n_67),
.Y(n_30)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_31),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_31),
.A2(n_67),
.B1(n_281),
.B2(n_282),
.Y(n_280)
);

BUFx2_ASAP7_75t_L g383 ( 
.A(n_31),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_31),
.B(n_237),
.Y(n_410)
);

AND2x4_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_46),
.Y(n_31)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_36),
.B1(n_40),
.B2(n_44),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_37),
.Y(n_188)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_38),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g170 ( 
.A(n_39),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_39),
.Y(n_448)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g442 ( 
.A(n_43),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_51),
.B1(n_54),
.B2(n_57),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_49),
.Y(n_392)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_50),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_50),
.Y(n_351)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_57),
.A2(n_92),
.B1(n_95),
.B2(n_98),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx8_ASAP7_75t_L g354 ( 
.A(n_58),
.Y(n_354)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_59),
.Y(n_240)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_62),
.Y(n_65)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_62),
.Y(n_238)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_63),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_63),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_63),
.Y(n_432)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_66),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g281 ( 
.A(n_66),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_66),
.B(n_237),
.Y(n_355)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_75),
.Y(n_330)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_78),
.Y(n_292)
);

NAND2x1_ASAP7_75t_SL g78 ( 
.A(n_79),
.B(n_102),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_79),
.B(n_376),
.Y(n_375)
);

NAND2x1_ASAP7_75t_SL g79 ( 
.A(n_80),
.B(n_90),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_80),
.B(n_114),
.Y(n_262)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_85),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_85),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_85),
.Y(n_269)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_89),
.Y(n_230)
);

AO22x1_ASAP7_75t_L g225 ( 
.A1(n_90),
.A2(n_103),
.B1(n_114),
.B2(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_90),
.B(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_90),
.B(n_226),
.Y(n_346)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_115),
.Y(n_114)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_95),
.Y(n_331)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_97),
.Y(n_344)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_114),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_108),
.Y(n_337)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_110),
.Y(n_380)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_113),
.Y(n_116)
);

OAI21xp33_ASAP7_75t_L g376 ( 
.A1(n_114),
.A2(n_336),
.B(n_377),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_120),
.B2(n_122),
.Y(n_115)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_126),
.B(n_292),
.C(n_293),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_153),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_127),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_136),
.B1(n_145),
.B2(n_147),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_128),
.A2(n_136),
.B1(n_204),
.B2(n_208),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g252 ( 
.A1(n_128),
.A2(n_147),
.B(n_253),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_128),
.A2(n_314),
.B1(n_412),
.B2(n_418),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g497 ( 
.A1(n_128),
.A2(n_498),
.B(n_509),
.Y(n_497)
);

INVx2_ASAP7_75t_SL g128 ( 
.A(n_129),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_129),
.A2(n_209),
.B1(n_313),
.B2(n_322),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_129),
.B(n_451),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_129),
.A2(n_516),
.B1(n_527),
.B2(n_529),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_133),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_131),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_132),
.Y(n_161)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_132),
.Y(n_215)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_132),
.Y(n_321)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_132),
.Y(n_416)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_133),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_135),
.Y(n_146)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_139),
.Y(n_317)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_139),
.Y(n_503)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_144),
.Y(n_526)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_149),
.Y(n_151)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_150),
.Y(n_569)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_153),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_180),
.B1(n_189),
.B2(n_190),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_154),
.A2(n_180),
.B1(n_189),
.B2(n_217),
.Y(n_216)
);

OAI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_154),
.A2(n_189),
.B1(n_190),
.B2(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g273 ( 
.A(n_154),
.Y(n_273)
);

OAI21xp33_ASAP7_75t_SL g455 ( 
.A1(n_154),
.A2(n_456),
.B(n_460),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_154),
.A2(n_189),
.B1(n_456),
.B2(n_477),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g492 ( 
.A1(n_154),
.A2(n_477),
.B1(n_493),
.B2(n_494),
.Y(n_492)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_168),
.Y(n_154)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_155),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_155),
.Y(n_279)
);

OAI22x1_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_160),
.B1(n_162),
.B2(n_165),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_162),
.Y(n_542)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_166),
.Y(n_534)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g550 ( 
.A(n_167),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_171),
.B1(n_175),
.B2(n_177),
.Y(n_168)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_170),
.Y(n_194)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_174),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_177),
.Y(n_371)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_178),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_179),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_179),
.Y(n_219)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx4_ASAP7_75t_L g540 ( 
.A(n_185),
.Y(n_540)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_194),
.Y(n_278)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_199),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_199),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_199),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g547 ( 
.A(n_199),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_200),
.B(n_301),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_224),
.C(n_234),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

XNOR2x1_ASAP7_75t_L g304 ( 
.A(n_202),
.B(n_305),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_216),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_203),
.B(n_216),
.Y(n_365)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_207),
.Y(n_326)
);

INVx2_ASAP7_75t_L g420 ( 
.A(n_207),
.Y(n_420)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_211),
.Y(n_453)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_214),
.Y(n_452)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_217),
.Y(n_374)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_219),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_219),
.Y(n_251)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx3_ASAP7_75t_L g373 ( 
.A(n_222),
.Y(n_373)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XNOR2x1_ASAP7_75t_L g305 ( 
.A(n_225),
.B(n_235),
.Y(n_305)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g335 ( 
.A(n_233),
.Y(n_335)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

OAI22x1_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

OA21x2_ASAP7_75t_L g347 ( 
.A1(n_239),
.A2(n_348),
.B(n_355),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g482 ( 
.A1(n_239),
.A2(n_355),
.B(n_483),
.Y(n_482)
);

HB1xp67_ASAP7_75t_L g409 ( 
.A(n_241),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_241),
.B(n_381),
.Y(n_496)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_242),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_252),
.B2(n_255),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_244),
.B(n_252),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_245),
.Y(n_274)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx4_ASAP7_75t_L g481 ( 
.A(n_248),
.Y(n_481)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_252),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_252),
.A2(n_255),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g449 ( 
.A1(n_253),
.A2(n_412),
.B(n_450),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g561 ( 
.A1(n_253),
.A2(n_450),
.B(n_517),
.Y(n_561)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_256),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_270),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_262),
.B(n_346),
.Y(n_345)
);

BUFx4f_ASAP7_75t_SL g265 ( 
.A(n_266),
.Y(n_265)
);

INVx8_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_291),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_272),
.A2(n_280),
.B(n_290),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_280),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_275),
.B2(n_279),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_273),
.A2(n_279),
.B1(n_369),
.B2(n_374),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_273),
.B(n_553),
.Y(n_552)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_279),
.B(n_369),
.Y(n_460)
);

INVx1_ASAP7_75t_SL g493 ( 
.A(n_279),
.Y(n_493)
);

AOI22x1_ASAP7_75t_L g382 ( 
.A1(n_281),
.A2(n_383),
.B1(n_384),
.B2(n_393),
.Y(n_382)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_289),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

AO21x1_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_356),
.B(n_588),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_303),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g591 ( 
.A(n_300),
.Y(n_591)
);

INVxp33_ASAP7_75t_SL g590 ( 
.A(n_303),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_306),
.C(n_309),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_304),
.B(n_306),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_309),
.B(n_395),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_345),
.C(n_347),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

XNOR2x1_ASAP7_75t_L g362 ( 
.A(n_311),
.B(n_363),
.Y(n_362)
);

NOR2xp67_ASAP7_75t_SL g311 ( 
.A(n_312),
.B(n_327),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_312),
.B(n_327),
.Y(n_404)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

BUFx3_ASAP7_75t_L g417 ( 
.A(n_320),
.Y(n_417)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_322),
.B(n_451),
.Y(n_509)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

AOI32xp33_ASAP7_75t_L g327 ( 
.A1(n_328),
.A2(n_331),
.A3(n_332),
.B1(n_336),
.B2(n_338),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx3_ASAP7_75t_SL g341 ( 
.A(n_330),
.Y(n_341)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx4_ASAP7_75t_SL g334 ( 
.A(n_335),
.Y(n_334)
);

NAND2xp33_ASAP7_75t_SL g338 ( 
.A(n_339),
.B(n_342),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_341),
.Y(n_438)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

XNOR2x1_ASAP7_75t_L g363 ( 
.A(n_345),
.B(n_347),
.Y(n_363)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_348),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx4_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

OAI21x1_ASAP7_75t_L g356 ( 
.A1(n_357),
.A2(n_423),
.B(n_584),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

OAI21xp5_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_394),
.B(n_396),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_360),
.B(n_586),
.C(n_587),
.Y(n_585)
);

MAJx2_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_364),
.C(n_366),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_361),
.A2(n_362),
.B1(n_398),
.B2(n_400),
.Y(n_397)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_364),
.A2(n_365),
.B1(n_367),
.B2(n_399),
.Y(n_398)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g399 ( 
.A(n_367),
.Y(n_399)
);

MAJx2_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_375),
.C(n_382),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_368),
.B(n_382),
.Y(n_403)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_369),
.Y(n_494)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_373),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_375),
.B(n_403),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_381),
.Y(n_377)
);

INVx2_ASAP7_75t_SL g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_381),
.B(n_444),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_381),
.B(n_537),
.Y(n_536)
);

OAI21xp33_ASAP7_75t_SL g553 ( 
.A1(n_381),
.A2(n_536),
.B(n_554),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_SL g560 ( 
.A(n_381),
.B(n_493),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_381),
.B(n_566),
.Y(n_565)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_384),
.Y(n_408)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx3_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_394),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_401),
.Y(n_396)
);

OR2x2_ASAP7_75t_L g587 ( 
.A(n_397),
.B(n_401),
.Y(n_587)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_398),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_404),
.C(n_405),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_402),
.B(n_466),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_404),
.B(n_406),
.Y(n_466)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_411),
.C(n_421),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_407),
.B(n_463),
.Y(n_462)
);

OAI21x1_ASAP7_75t_L g407 ( 
.A1(n_408),
.A2(n_409),
.B(n_410),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_411),
.A2(n_421),
.B1(n_422),
.B2(n_464),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_411),
.Y(n_464)
);

INVx1_ASAP7_75t_SL g413 ( 
.A(n_414),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

BUFx12f_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

OAI21x1_ASAP7_75t_L g424 ( 
.A1(n_425),
.A2(n_467),
.B(n_582),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_465),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_427),
.B(n_583),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_454),
.C(n_461),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_428),
.A2(n_454),
.B1(n_455),
.B2(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_428),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_449),
.Y(n_428)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx4_ASAP7_75t_L g484 ( 
.A(n_431),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_438),
.B(n_439),
.Y(n_437)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

BUFx3_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_446),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_447),
.Y(n_556)
);

INVx5_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_449),
.B(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

INVx2_ASAP7_75t_SL g457 ( 
.A(n_458),
.Y(n_457)
);

INVx4_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_460),
.B(n_552),
.Y(n_551)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_462),
.B(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_465),
.Y(n_583)
);

AOI21x1_ASAP7_75t_L g467 ( 
.A1(n_468),
.A2(n_510),
.B(n_581),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_488),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_473),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_470),
.B(n_473),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_476),
.C(n_482),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_474),
.B(n_490),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_476),
.B(n_482),
.Y(n_490)
);

INVx2_ASAP7_75t_SL g478 ( 
.A(n_479),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_489),
.B(n_491),
.Y(n_488)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_489),
.Y(n_579)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_491),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_492),
.B(n_495),
.C(n_497),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_492),
.B(n_496),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g573 ( 
.A(n_497),
.B(n_574),
.Y(n_573)
);

INVxp67_ASAP7_75t_L g529 ( 
.A(n_498),
.Y(n_529)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_500),
.B(n_533),
.Y(n_532)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx4_ASAP7_75t_L g501 ( 
.A(n_502),
.Y(n_501)
);

INVx4_ASAP7_75t_L g502 ( 
.A(n_503),
.Y(n_502)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_503),
.Y(n_508)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_507),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_508),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_511),
.B(n_577),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_572),
.Y(n_511)
);

OAI21x1_ASAP7_75t_L g512 ( 
.A1(n_513),
.A2(n_557),
.B(n_571),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_515),
.B(n_530),
.Y(n_514)
);

OR2x2_ASAP7_75t_L g571 ( 
.A(n_515),
.B(n_530),
.Y(n_571)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_519),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_520),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_526),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

INVx5_ASAP7_75t_L g566 ( 
.A(n_528),
.Y(n_566)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_531),
.B(n_551),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_531),
.B(n_551),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_532),
.A2(n_535),
.B1(n_541),
.B2(n_543),
.Y(n_531)
);

INVx2_ASAP7_75t_SL g533 ( 
.A(n_534),
.Y(n_533)
);

INVxp67_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_544),
.B(n_548),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

BUFx2_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

BUFx2_ASAP7_75t_L g554 ( 
.A(n_555),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_556),
.Y(n_555)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_558),
.Y(n_557)
);

OAI21xp5_ASAP7_75t_L g558 ( 
.A1(n_559),
.A2(n_562),
.B(n_570),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g559 ( 
.A(n_560),
.B(n_561),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_560),
.B(n_561),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_563),
.B(n_564),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_SL g564 ( 
.A(n_565),
.B(n_567),
.Y(n_564)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_568),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_569),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_573),
.B(n_575),
.Y(n_572)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_573),
.Y(n_580)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_576),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_576),
.A2(n_578),
.B1(n_579),
.B2(n_580),
.Y(n_577)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_585),
.Y(n_584)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_589),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_590),
.B(n_591),
.Y(n_589)
);


endmodule