module fake_jpeg_22687_n_206 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_206);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_206;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_5),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_18),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_34),
.B(n_22),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_35),
.B(n_37),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g38 ( 
.A(n_21),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_41),
.Y(n_50)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_43),
.B(n_37),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_40),
.A2(n_28),
.B1(n_27),
.B2(n_30),
.Y(n_46)
);

OAI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_46),
.A2(n_47),
.B1(n_63),
.B2(n_16),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_40),
.A2(n_27),
.B1(n_30),
.B2(n_31),
.Y(n_47)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_54),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_35),
.B(n_17),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_58),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_24),
.Y(n_56)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_36),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_59),
.B(n_62),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_64),
.Y(n_69)
);

INVx5_ASAP7_75t_SL g62 ( 
.A(n_36),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_43),
.A2(n_17),
.B1(n_19),
.B2(n_26),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_33),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_65),
.B(n_66),
.Y(n_103)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

O2A1O1Ixp33_ASAP7_75t_SL g67 ( 
.A1(n_48),
.A2(n_36),
.B(n_37),
.C(n_42),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_67),
.A2(n_73),
.B1(n_64),
.B2(n_45),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_68),
.A2(n_72),
.B1(n_86),
.B2(n_20),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_55),
.B(n_16),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_81),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_53),
.A2(n_39),
.B1(n_41),
.B2(n_38),
.Y(n_72)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_62),
.A2(n_42),
.B1(n_33),
.B2(n_26),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_74),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_48),
.B(n_33),
.C(n_32),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_75),
.B(n_84),
.C(n_20),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_32),
.Y(n_79)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_54),
.B(n_31),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_58),
.B(n_25),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_29),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_46),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_19),
.Y(n_85)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_49),
.A2(n_29),
.B1(n_25),
.B2(n_22),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_77),
.A2(n_49),
.B1(n_61),
.B2(n_51),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_87),
.A2(n_90),
.B1(n_44),
.B2(n_60),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_65),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_100),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_78),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_91),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_92),
.A2(n_101),
.B1(n_66),
.B2(n_44),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_95),
.B(n_97),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_71),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_52),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_SL g98 ( 
.A(n_67),
.B(n_51),
.C(n_44),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_98),
.A2(n_83),
.B(n_73),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_84),
.A2(n_45),
.B1(n_51),
.B2(n_60),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_15),
.Y(n_104)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_104),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_15),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_106),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_74),
.B(n_13),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_82),
.B(n_44),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_70),
.Y(n_119)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_0),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_102),
.Y(n_129)
);

NAND2xp33_ASAP7_75t_L g111 ( 
.A(n_98),
.B(n_73),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_111),
.B(n_102),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_97),
.A2(n_90),
.B1(n_101),
.B2(n_96),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_112),
.A2(n_113),
.B1(n_126),
.B2(n_93),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_107),
.A2(n_75),
.B1(n_77),
.B2(n_73),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_114),
.A2(n_89),
.B(n_93),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_71),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_116),
.B(n_117),
.C(n_94),
.Y(n_135)
);

A2O1A1O1Ixp25_ASAP7_75t_L g117 ( 
.A1(n_88),
.A2(n_76),
.B(n_83),
.C(n_69),
.D(n_81),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_120),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_123),
.Y(n_138)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_88),
.B(n_76),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_108),
.Y(n_137)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_129),
.B(n_135),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_121),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_131),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_132),
.A2(n_118),
.B(n_116),
.Y(n_153)
);

BUFx4f_ASAP7_75t_SL g133 ( 
.A(n_128),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_133),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_94),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_136),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_137),
.B(n_139),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_1),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_140),
.A2(n_114),
.B(n_123),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_115),
.B(n_99),
.Y(n_142)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_142),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_91),
.Y(n_143)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_143),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_113),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_144),
.A2(n_146),
.B1(n_139),
.B2(n_138),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_12),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_145),
.B(n_147),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_125),
.A2(n_11),
.B1(n_2),
.B2(n_3),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_117),
.B(n_1),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_151),
.B(n_161),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_153),
.B(n_158),
.Y(n_170)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_154),
.B(n_143),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_156),
.A2(n_150),
.B1(n_162),
.B2(n_151),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_142),
.A2(n_109),
.B(n_122),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_144),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_141),
.B(n_110),
.Y(n_158)
);

A2O1A1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_138),
.A2(n_124),
.B(n_122),
.C(n_5),
.Y(n_161)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_163),
.Y(n_177)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_156),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_165),
.B(n_167),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_140),
.Y(n_166)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_166),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_155),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_150),
.A2(n_136),
.B1(n_148),
.B2(n_159),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_168),
.A2(n_152),
.B(n_133),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_148),
.A2(n_146),
.B1(n_135),
.B2(n_134),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_174),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_171),
.B(n_157),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_129),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_153),
.C(n_149),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_140),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_161),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_4),
.Y(n_190)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_176),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_164),
.A2(n_160),
.B(n_133),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_180),
.A2(n_181),
.B1(n_183),
.B2(n_169),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_178),
.A2(n_174),
.B1(n_168),
.B2(n_170),
.Y(n_185)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_185),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_186),
.B(n_190),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_171),
.Y(n_187)
);

OAI221xp5_ASAP7_75t_L g196 ( 
.A1(n_187),
.A2(n_182),
.B1(n_176),
.B2(n_10),
.C(n_7),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_178),
.A2(n_172),
.B1(n_149),
.B2(n_6),
.Y(n_188)
);

NAND4xp25_ASAP7_75t_L g193 ( 
.A(n_188),
.B(n_175),
.C(n_9),
.D(n_10),
.Y(n_193)
);

A2O1A1Ixp33_ASAP7_75t_L g189 ( 
.A1(n_183),
.A2(n_3),
.B(n_4),
.C(n_7),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_189),
.B(n_7),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_184),
.A2(n_180),
.B(n_179),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_191),
.B(n_187),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_196),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_193),
.A2(n_189),
.B(n_185),
.Y(n_197)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_197),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_199),
.A2(n_200),
.B(n_194),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_195),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_198),
.B(n_195),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_202),
.B(n_203),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_201),
.B(n_10),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_205),
.B(n_204),
.Y(n_206)
);


endmodule