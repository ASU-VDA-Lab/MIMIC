module fake_jpeg_3836_n_74 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_74);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_74;

wire n_61;
wire n_45;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_39;
wire n_42;
wire n_49;
wire n_72;
wire n_38;
wire n_56;
wire n_50;
wire n_67;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_69;
wire n_40;
wire n_71;
wire n_48;
wire n_35;
wire n_46;
wire n_44;
wire n_36;
wire n_62;
wire n_37;
wire n_43;
wire n_70;
wire n_66;

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

HB1xp67_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_9),
.B(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_32),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx4f_ASAP7_75t_SL g43 ( 
.A(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_16),
.B(n_18),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

NAND3xp33_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_2),
.C(n_3),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_46),
.B(n_48),
.Y(n_52)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_47),
.A2(n_51),
.B1(n_39),
.B2(n_36),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_40),
.B(n_4),
.Y(n_48)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_49),
.B(n_42),
.Y(n_56)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

HAxp5_ASAP7_75t_SL g51 ( 
.A(n_33),
.B(n_5),
.CON(n_51),
.SN(n_51)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_12),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_14),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_48),
.A2(n_44),
.B1(n_35),
.B2(n_38),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_57),
.A2(n_58),
.B1(n_6),
.B2(n_8),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_L g58 ( 
.A1(n_46),
.A2(n_41),
.B1(n_37),
.B2(n_10),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_19),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_61),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_62),
.B(n_55),
.C(n_52),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_20),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_21),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_67),
.C(n_22),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_65),
.C(n_24),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_69),
.B(n_23),
.C(n_25),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_70),
.B(n_27),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_71),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_29),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_30),
.Y(n_74)
);


endmodule