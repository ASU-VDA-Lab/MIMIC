module fake_jpeg_5727_n_322 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_322);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_322;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx6_ASAP7_75t_SL g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_9),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx3_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_38),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_12),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_39),
.B(n_40),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_41),
.Y(n_102)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_42),
.B(n_46),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_43),
.B(n_52),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx4_ASAP7_75t_SL g87 ( 
.A(n_44),
.Y(n_87)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_16),
.B(n_13),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_54),
.Y(n_83)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_49),
.B(n_51),
.Y(n_97)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_50),
.Y(n_61)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_21),
.B(n_13),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_21),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_57),
.B(n_17),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_20),
.B(n_9),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_58),
.B(n_15),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_26),
.B(n_0),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_59),
.B(n_0),
.Y(n_105)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_60),
.B(n_70),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_50),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_62),
.A2(n_73),
.B1(n_82),
.B2(n_89),
.Y(n_118)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_65),
.Y(n_112)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_48),
.Y(n_66)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_42),
.A2(n_28),
.B1(n_30),
.B2(n_23),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_68),
.A2(n_88),
.B1(n_93),
.B2(n_25),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_40),
.A2(n_30),
.B1(n_28),
.B2(n_35),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_69),
.A2(n_92),
.B1(n_98),
.B2(n_82),
.Y(n_114)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_71),
.Y(n_120)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_72),
.B(n_78),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_49),
.A2(n_28),
.B1(n_26),
.B2(n_29),
.Y(n_73)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_77),
.Y(n_122)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_38),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_79),
.B(n_81),
.Y(n_125)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_80),
.Y(n_137)
);

AO22x1_ASAP7_75t_SL g82 ( 
.A1(n_41),
.A2(n_31),
.B1(n_36),
.B2(n_25),
.Y(n_82)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_85),
.Y(n_115)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

OA22x2_ASAP7_75t_L g89 ( 
.A1(n_44),
.A2(n_45),
.B1(n_17),
.B2(n_34),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_44),
.B(n_16),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_99),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_44),
.A2(n_29),
.B1(n_35),
.B2(n_22),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_64),
.C(n_73),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_45),
.A2(n_22),
.B1(n_15),
.B2(n_17),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_45),
.A2(n_34),
.B1(n_32),
.B2(n_31),
.Y(n_93)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_95),
.Y(n_129)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_40),
.A2(n_37),
.B1(n_36),
.B2(n_31),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_48),
.B(n_34),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_59),
.B(n_8),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_100),
.B(n_104),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_48),
.B(n_36),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_103),
.B(n_106),
.Y(n_126)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_27),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_L g111 ( 
.A1(n_82),
.A2(n_25),
.B1(n_19),
.B2(n_32),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_111),
.A2(n_114),
.B1(n_116),
.B2(n_121),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_119),
.B(n_133),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_61),
.A2(n_19),
.B1(n_27),
.B2(n_11),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_89),
.A2(n_27),
.B1(n_11),
.B2(n_9),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_124),
.B(n_131),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_97),
.B(n_32),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_134),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_128),
.B(n_75),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_89),
.A2(n_27),
.B1(n_32),
.B2(n_3),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_L g132 ( 
.A1(n_62),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_132),
.A2(n_117),
.B1(n_136),
.B2(n_126),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_83),
.B(n_87),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_91),
.B(n_1),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_61),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_135),
.B(n_5),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_123),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_139),
.B(n_142),
.Y(n_178)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

INVx8_ASAP7_75t_L g202 ( 
.A(n_140),
.Y(n_202)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_141),
.A2(n_149),
.B1(n_152),
.B2(n_157),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_143),
.B(n_144),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

OA22x2_ASAP7_75t_L g145 ( 
.A1(n_118),
.A2(n_87),
.B1(n_93),
.B2(n_68),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_145),
.A2(n_107),
.B1(n_76),
.B2(n_102),
.Y(n_174)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_123),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_146),
.B(n_147),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_115),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_127),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_148),
.B(n_161),
.Y(n_188)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_150),
.B(n_151),
.Y(n_207)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_110),
.Y(n_151)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_154),
.A2(n_172),
.B(n_109),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_136),
.B(n_74),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_155),
.B(n_168),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_156),
.Y(n_206)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_110),
.Y(n_157)
);

O2A1O1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_118),
.A2(n_92),
.B(n_102),
.C(n_101),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_158),
.A2(n_109),
.B(n_137),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_79),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_159),
.B(n_78),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_115),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_160),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_113),
.B(n_63),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_119),
.B(n_84),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_162),
.B(n_164),
.Y(n_183)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_125),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_163),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_134),
.B(n_84),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_125),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_165),
.Y(n_187)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_126),
.Y(n_167)
);

INVx2_ASAP7_75t_SL g175 ( 
.A(n_167),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_128),
.B(n_63),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_170),
.B(n_171),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_128),
.B(n_5),
.Y(n_171)
);

AND2x2_ASAP7_75t_SL g172 ( 
.A(n_117),
.B(n_88),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_173),
.A2(n_184),
.B(n_201),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_174),
.A2(n_181),
.B1(n_186),
.B2(n_94),
.Y(n_230)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_148),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_176),
.B(n_177),
.Y(n_209)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_161),
.Y(n_177)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_172),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_182),
.B(n_191),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_170),
.A2(n_133),
.B(n_120),
.Y(n_184)
);

OAI22x1_ASAP7_75t_L g186 ( 
.A1(n_145),
.A2(n_76),
.B1(n_107),
.B2(n_101),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_164),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_190),
.B(n_169),
.C(n_171),
.Y(n_211)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_172),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_168),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_193),
.B(n_194),
.Y(n_229)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_138),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g195 ( 
.A(n_159),
.B(n_137),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_195),
.A2(n_166),
.B(n_112),
.Y(n_217)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_138),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_196),
.B(n_197),
.Y(n_232)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_140),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_158),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_198),
.B(n_199),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_169),
.B(n_120),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_145),
.A2(n_122),
.B(n_112),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_203),
.A2(n_6),
.B(n_7),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_169),
.B(n_122),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_192),
.Y(n_223)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_188),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_210),
.Y(n_235)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_188),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_211),
.B(n_228),
.C(n_192),
.Y(n_246)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_178),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_213),
.B(n_215),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_199),
.A2(n_145),
.B(n_153),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_214),
.A2(n_217),
.B(n_224),
.Y(n_242)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_200),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_189),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_216),
.Y(n_241)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_207),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_220),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_179),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_221),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_207),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_222),
.B(n_223),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_204),
.A2(n_149),
.B(n_143),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_185),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_227),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_194),
.B(n_142),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_183),
.B(n_152),
.C(n_141),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_230),
.A2(n_186),
.B1(n_198),
.B2(n_182),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_184),
.A2(n_150),
.B(n_144),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_231),
.A2(n_191),
.B(n_201),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_185),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_233),
.A2(n_202),
.B1(n_225),
.B2(n_197),
.Y(n_252)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_232),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_248),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_236),
.A2(n_245),
.B1(n_251),
.B2(n_229),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_195),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_239),
.B(n_231),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_211),
.B(n_183),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_243),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_190),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_226),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_214),
.A2(n_193),
.B1(n_180),
.B2(n_176),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_223),
.C(n_212),
.Y(n_259)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_232),
.Y(n_248)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_227),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_254),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_217),
.A2(n_195),
.B1(n_180),
.B2(n_203),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_252),
.A2(n_233),
.B1(n_222),
.B2(n_218),
.Y(n_256)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_228),
.Y(n_253)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_253),
.Y(n_271)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_209),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_256),
.B(n_248),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_257),
.A2(n_268),
.B1(n_230),
.B2(n_242),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_261),
.C(n_262),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_243),
.B(n_219),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_240),
.B(n_229),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_255),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_263),
.B(n_249),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_208),
.C(n_210),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_269),
.C(n_253),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_266),
.A2(n_270),
.B(n_249),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_241),
.B(n_202),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_267),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_245),
.A2(n_174),
.B1(n_181),
.B2(n_226),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_242),
.B(n_224),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_234),
.B(n_196),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_272),
.A2(n_244),
.B(n_239),
.Y(n_286)
);

BUFx12_ASAP7_75t_L g273 ( 
.A(n_260),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_273),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_274),
.B(n_264),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_276),
.A2(n_278),
.B(n_280),
.Y(n_297)
);

NAND3xp33_ASAP7_75t_SL g277 ( 
.A(n_272),
.B(n_254),
.C(n_209),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_281),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_271),
.A2(n_247),
.B1(n_250),
.B2(n_217),
.Y(n_278)
);

BUFx12f_ASAP7_75t_SL g280 ( 
.A(n_269),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_202),
.Y(n_282)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_282),
.Y(n_294)
);

BUFx24_ASAP7_75t_SL g283 ( 
.A(n_262),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_283),
.B(n_258),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_255),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_275),
.C(n_259),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_261),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_298),
.Y(n_302)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_288),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_260),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_289),
.B(n_292),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_279),
.A2(n_206),
.B1(n_241),
.B2(n_177),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_293),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_295),
.B(n_215),
.Y(n_303)
);

NAND3xp33_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_205),
.C(n_173),
.Y(n_296)
);

OAI31xp33_ASAP7_75t_L g299 ( 
.A1(n_296),
.A2(n_239),
.A3(n_238),
.B(n_205),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_299),
.A2(n_304),
.B1(n_307),
.B2(n_301),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_303),
.B(n_175),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_290),
.A2(n_238),
.B1(n_285),
.B2(n_265),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_294),
.B(n_213),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_305),
.A2(n_237),
.B(n_187),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_297),
.A2(n_278),
.B1(n_235),
.B2(n_275),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_302),
.B(n_298),
.C(n_291),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_309),
.C(n_311),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_301),
.A2(n_297),
.B1(n_235),
.B2(n_292),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_312),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_306),
.B(n_289),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_313),
.B(n_300),
.C(n_307),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g318 ( 
.A1(n_315),
.A2(n_308),
.B(n_309),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_316),
.B(n_237),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_317),
.A2(n_318),
.B(n_314),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_311),
.B(n_293),
.Y(n_320)
);

AOI321xp33_ASAP7_75t_L g321 ( 
.A1(n_320),
.A2(n_306),
.A3(n_273),
.B1(n_220),
.B2(n_175),
.C(n_187),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_175),
.Y(n_322)
);


endmodule