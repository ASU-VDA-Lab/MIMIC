module fake_aes_7164_n_729 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_729);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_729;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_638;
wire n_540;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_666;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_581;
wire n_458;
wire n_504;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g81 ( .A(n_69), .Y(n_81) );
INVx2_ASAP7_75t_L g82 ( .A(n_12), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_66), .Y(n_83) );
INVx2_ASAP7_75t_L g84 ( .A(n_40), .Y(n_84) );
BUFx6f_ASAP7_75t_L g85 ( .A(n_68), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_31), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_63), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_59), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_14), .Y(n_89) );
CKINVDCx16_ASAP7_75t_R g90 ( .A(n_23), .Y(n_90) );
INVx2_ASAP7_75t_L g91 ( .A(n_70), .Y(n_91) );
CKINVDCx20_ASAP7_75t_R g92 ( .A(n_28), .Y(n_92) );
CKINVDCx5p33_ASAP7_75t_R g93 ( .A(n_50), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_22), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_21), .Y(n_95) );
BUFx6f_ASAP7_75t_L g96 ( .A(n_18), .Y(n_96) );
BUFx2_ASAP7_75t_L g97 ( .A(n_75), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_56), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_64), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_27), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_58), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_7), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_78), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_4), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_30), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_43), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_18), .Y(n_107) );
BUFx3_ASAP7_75t_L g108 ( .A(n_79), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_46), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_55), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_72), .Y(n_111) );
NOR2xp67_ASAP7_75t_L g112 ( .A(n_57), .B(n_35), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_1), .Y(n_113) );
NOR2xp67_ASAP7_75t_L g114 ( .A(n_53), .B(n_38), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_51), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_60), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_6), .Y(n_117) );
INVx1_ASAP7_75t_SL g118 ( .A(n_67), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_4), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_11), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_39), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_33), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_3), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_74), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_52), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_12), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_13), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_47), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_8), .Y(n_129) );
BUFx2_ASAP7_75t_L g130 ( .A(n_71), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_83), .Y(n_131) );
INVx4_ASAP7_75t_L g132 ( .A(n_97), .Y(n_132) );
AND2x4_ASAP7_75t_L g133 ( .A(n_97), .B(n_0), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g134 ( .A(n_130), .B(n_0), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_83), .Y(n_135) );
INVx3_ASAP7_75t_L g136 ( .A(n_82), .Y(n_136) );
BUFx12f_ASAP7_75t_L g137 ( .A(n_130), .Y(n_137) );
AOI22xp5_ASAP7_75t_L g138 ( .A1(n_90), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_85), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_94), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_84), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_107), .B(n_2), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_84), .Y(n_143) );
AND2x2_ASAP7_75t_SL g144 ( .A(n_94), .B(n_32), .Y(n_144) );
BUFx8_ASAP7_75t_L g145 ( .A(n_98), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_85), .Y(n_146) );
AND2x2_ASAP7_75t_L g147 ( .A(n_82), .B(n_5), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_98), .Y(n_148) );
AND2x4_ASAP7_75t_L g149 ( .A(n_113), .B(n_5), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_128), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_128), .Y(n_151) );
AOI22xp5_ASAP7_75t_L g152 ( .A1(n_107), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_85), .Y(n_153) );
AOI22xp5_ASAP7_75t_L g154 ( .A1(n_120), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_91), .Y(n_155) );
AND2x4_ASAP7_75t_L g156 ( .A(n_113), .B(n_9), .Y(n_156) );
OAI21x1_ASAP7_75t_L g157 ( .A1(n_91), .A2(n_37), .B(n_77), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_85), .B(n_10), .Y(n_158) );
AND2x4_ASAP7_75t_L g159 ( .A(n_126), .B(n_13), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_85), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_81), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_86), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_120), .B(n_14), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_127), .B(n_15), .Y(n_164) );
OAI22xp5_ASAP7_75t_SL g165 ( .A1(n_127), .A2(n_15), .B1(n_16), .B2(n_17), .Y(n_165) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_108), .Y(n_166) );
OAI22x1_ASAP7_75t_R g167 ( .A1(n_92), .A2(n_16), .B1(n_17), .B2(n_19), .Y(n_167) );
AND2x2_ASAP7_75t_L g168 ( .A(n_126), .B(n_129), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_99), .Y(n_169) );
INVx2_ASAP7_75t_SL g170 ( .A(n_108), .Y(n_170) );
AND2x4_ASAP7_75t_L g171 ( .A(n_129), .B(n_19), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_103), .Y(n_172) );
HB1xp67_ASAP7_75t_L g173 ( .A(n_89), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_105), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_99), .Y(n_175) );
INVx4_ASAP7_75t_L g176 ( .A(n_133), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_132), .B(n_124), .Y(n_177) );
AND2x4_ASAP7_75t_L g178 ( .A(n_132), .B(n_123), .Y(n_178) );
BUFx3_ASAP7_75t_L g179 ( .A(n_166), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_149), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_166), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_166), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_166), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_132), .B(n_93), .Y(n_184) );
AOI22xp33_ASAP7_75t_L g185 ( .A1(n_131), .A2(n_102), .B1(n_104), .B2(n_119), .Y(n_185) );
OR2x6_ASAP7_75t_L g186 ( .A(n_137), .B(n_117), .Y(n_186) );
INVx1_ASAP7_75t_L g187 ( .A(n_149), .Y(n_187) );
AOI22xp33_ASAP7_75t_L g188 ( .A1(n_131), .A2(n_96), .B1(n_110), .B2(n_121), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_166), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_161), .B(n_125), .Y(n_190) );
AOI22xp5_ASAP7_75t_L g191 ( .A1(n_133), .A2(n_137), .B1(n_144), .B2(n_156), .Y(n_191) );
OR2x6_ASAP7_75t_L g192 ( .A(n_165), .B(n_96), .Y(n_192) );
AND2x2_ASAP7_75t_L g193 ( .A(n_173), .B(n_125), .Y(n_193) );
INVx3_ASAP7_75t_L g194 ( .A(n_149), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_135), .B(n_124), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_161), .B(n_87), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_156), .Y(n_197) );
OAI221xp5_ASAP7_75t_L g198 ( .A1(n_135), .A2(n_109), .B1(n_115), .B2(n_116), .C(n_87), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_156), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_159), .Y(n_200) );
AND2x4_ASAP7_75t_L g201 ( .A(n_133), .B(n_96), .Y(n_201) );
INVx5_ASAP7_75t_L g202 ( .A(n_159), .Y(n_202) );
OR2x2_ASAP7_75t_L g203 ( .A(n_168), .B(n_96), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_159), .Y(n_204) );
INVx3_ASAP7_75t_L g205 ( .A(n_171), .Y(n_205) );
INVx3_ASAP7_75t_L g206 ( .A(n_171), .Y(n_206) );
BUFx3_ASAP7_75t_L g207 ( .A(n_170), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_168), .B(n_88), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_171), .Y(n_209) );
AOI22xp5_ASAP7_75t_L g210 ( .A1(n_144), .A2(n_88), .B1(n_101), .B2(n_116), .Y(n_210) );
INVx1_ASAP7_75t_SL g211 ( .A(n_142), .Y(n_211) );
BUFx4f_ASAP7_75t_L g212 ( .A(n_144), .Y(n_212) );
AND2x2_ASAP7_75t_L g213 ( .A(n_162), .B(n_93), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_140), .B(n_122), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_162), .B(n_95), .Y(n_215) );
AND2x6_ASAP7_75t_L g216 ( .A(n_147), .B(n_122), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_147), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_139), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_172), .B(n_95), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_140), .Y(n_220) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_148), .A2(n_96), .B1(n_106), .B2(n_100), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_148), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_150), .B(n_106), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_150), .Y(n_224) );
CKINVDCx20_ASAP7_75t_R g225 ( .A(n_145), .Y(n_225) );
AOI22xp33_ASAP7_75t_L g226 ( .A1(n_151), .A2(n_100), .B1(n_118), .B2(n_111), .Y(n_226) );
NAND2xp33_ASAP7_75t_L g227 ( .A(n_151), .B(n_111), .Y(n_227) );
AOI22xp5_ASAP7_75t_L g228 ( .A1(n_145), .A2(n_101), .B1(n_114), .B2(n_112), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_141), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_139), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_172), .B(n_20), .Y(n_231) );
BUFx10_ASAP7_75t_L g232 ( .A(n_134), .Y(n_232) );
OR2x2_ASAP7_75t_L g233 ( .A(n_174), .B(n_24), .Y(n_233) );
BUFx3_ASAP7_75t_L g234 ( .A(n_170), .Y(n_234) );
INVx2_ASAP7_75t_SL g235 ( .A(n_145), .Y(n_235) );
INVx4_ASAP7_75t_L g236 ( .A(n_136), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g237 ( .A(n_174), .B(n_25), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_139), .Y(n_238) );
OR2x2_ASAP7_75t_L g239 ( .A(n_163), .B(n_26), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_141), .B(n_29), .Y(n_240) );
BUFx6f_ASAP7_75t_L g241 ( .A(n_139), .Y(n_241) );
AND2x6_ASAP7_75t_L g242 ( .A(n_143), .B(n_34), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_203), .Y(n_243) );
INVx6_ASAP7_75t_L g244 ( .A(n_236), .Y(n_244) );
OAI221xp5_ASAP7_75t_L g245 ( .A1(n_191), .A2(n_164), .B1(n_138), .B2(n_154), .C(n_152), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_184), .B(n_136), .Y(n_246) );
BUFx6f_ASAP7_75t_L g247 ( .A(n_242), .Y(n_247) );
HB1xp67_ASAP7_75t_L g248 ( .A(n_208), .Y(n_248) );
NAND2x1p5_ASAP7_75t_L g249 ( .A(n_235), .B(n_158), .Y(n_249) );
BUFx8_ASAP7_75t_L g250 ( .A(n_193), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_213), .B(n_136), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_178), .B(n_175), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_212), .A2(n_175), .B1(n_169), .B2(n_143), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_212), .B(n_157), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_201), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_190), .B(n_169), .Y(n_256) );
AND2x6_ASAP7_75t_L g257 ( .A(n_194), .B(n_155), .Y(n_257) );
NAND2xp5_ASAP7_75t_SL g258 ( .A(n_211), .B(n_155), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g259 ( .A(n_178), .B(n_157), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_196), .B(n_160), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_215), .B(n_160), .Y(n_261) );
AOI22xp5_ASAP7_75t_L g262 ( .A1(n_210), .A2(n_160), .B1(n_153), .B2(n_146), .Y(n_262) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_176), .B(n_160), .Y(n_263) );
NOR2x2_ASAP7_75t_L g264 ( .A(n_186), .B(n_167), .Y(n_264) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_176), .B(n_160), .Y(n_265) );
AOI22xp5_ASAP7_75t_L g266 ( .A1(n_227), .A2(n_153), .B1(n_146), .B2(n_139), .Y(n_266) );
OAI22xp5_ASAP7_75t_SL g267 ( .A1(n_192), .A2(n_167), .B1(n_153), .B2(n_146), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_201), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_178), .B(n_153), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_176), .B(n_153), .Y(n_270) );
INVx4_ASAP7_75t_L g271 ( .A(n_236), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_202), .B(n_146), .Y(n_272) );
NOR2xp33_ASAP7_75t_SL g273 ( .A(n_186), .B(n_146), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_219), .B(n_36), .Y(n_274) );
INVx3_ASAP7_75t_L g275 ( .A(n_236), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_216), .B(n_41), .Y(n_276) );
OAI22xp5_ASAP7_75t_SL g277 ( .A1(n_192), .A2(n_42), .B1(n_44), .B2(n_45), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_201), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g279 ( .A1(n_220), .A2(n_48), .B1(n_49), .B2(n_54), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_205), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_186), .B(n_61), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_205), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_216), .B(n_62), .Y(n_283) );
AND2x4_ASAP7_75t_L g284 ( .A(n_217), .B(n_65), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_206), .Y(n_285) );
INVxp67_ASAP7_75t_SL g286 ( .A(n_222), .Y(n_286) );
BUFx8_ASAP7_75t_L g287 ( .A(n_216), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_216), .B(n_80), .Y(n_288) );
AND2x4_ASAP7_75t_L g289 ( .A(n_180), .B(n_73), .Y(n_289) );
OR2x2_ASAP7_75t_L g290 ( .A(n_192), .B(n_76), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_216), .B(n_177), .Y(n_291) );
INVx3_ASAP7_75t_L g292 ( .A(n_207), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_179), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_179), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_177), .B(n_224), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_229), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_187), .B(n_197), .Y(n_297) );
OAI22xp5_ASAP7_75t_L g298 ( .A1(n_199), .A2(n_209), .B1(n_204), .B2(n_200), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_206), .B(n_227), .Y(n_299) );
BUFx4f_ASAP7_75t_SL g300 ( .A(n_225), .Y(n_300) );
INVx2_ASAP7_75t_SL g301 ( .A(n_202), .Y(n_301) );
INVx3_ASAP7_75t_L g302 ( .A(n_207), .Y(n_302) );
INVx3_ASAP7_75t_L g303 ( .A(n_234), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_194), .Y(n_304) );
NAND2xp5_ASAP7_75t_SL g305 ( .A(n_228), .B(n_202), .Y(n_305) );
NAND2xp5_ASAP7_75t_SL g306 ( .A(n_202), .B(n_239), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_234), .B(n_194), .Y(n_307) );
AND2x4_ASAP7_75t_L g308 ( .A(n_185), .B(n_225), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_226), .B(n_233), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_226), .B(n_232), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_185), .B(n_232), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_232), .B(n_198), .Y(n_312) );
NAND2xp5_ASAP7_75t_SL g313 ( .A(n_231), .B(n_237), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_181), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_255), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_268), .Y(n_316) );
BUFx6f_ASAP7_75t_L g317 ( .A(n_271), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_278), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_280), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_304), .Y(n_320) );
OAI22xp5_ASAP7_75t_L g321 ( .A1(n_309), .A2(n_188), .B1(n_221), .B2(n_223), .Y(n_321) );
AOI21x1_ASAP7_75t_L g322 ( .A1(n_254), .A2(n_195), .B(n_223), .Y(n_322) );
AND2x2_ASAP7_75t_L g323 ( .A(n_248), .B(n_214), .Y(n_323) );
A2O1A1Ixp33_ASAP7_75t_L g324 ( .A1(n_259), .A2(n_237), .B(n_231), .C(n_195), .Y(n_324) );
AOI22xp5_ASAP7_75t_L g325 ( .A1(n_310), .A2(n_214), .B1(n_188), .B2(n_221), .Y(n_325) );
NAND2x1p5_ASAP7_75t_L g326 ( .A(n_271), .B(n_240), .Y(n_326) );
NOR2xp33_ASAP7_75t_R g327 ( .A(n_300), .B(n_242), .Y(n_327) );
NOR2xp33_ASAP7_75t_SL g328 ( .A(n_273), .B(n_242), .Y(n_328) );
AOI21xp5_ASAP7_75t_L g329 ( .A1(n_313), .A2(n_240), .B(n_182), .Y(n_329) );
AOI22xp5_ASAP7_75t_L g330 ( .A1(n_245), .A2(n_311), .B1(n_312), .B2(n_267), .Y(n_330) );
INVxp67_ASAP7_75t_L g331 ( .A(n_250), .Y(n_331) );
NOR2xp33_ASAP7_75t_R g332 ( .A(n_300), .B(n_242), .Y(n_332) );
BUFx2_ASAP7_75t_L g333 ( .A(n_287), .Y(n_333) );
O2A1O1Ixp5_ASAP7_75t_L g334 ( .A1(n_254), .A2(n_181), .B(n_182), .C(n_183), .Y(n_334) );
A2O1A1Ixp33_ASAP7_75t_L g335 ( .A1(n_259), .A2(n_183), .B(n_189), .C(n_218), .Y(n_335) );
OA22x2_ASAP7_75t_L g336 ( .A1(n_308), .A2(n_189), .B1(n_242), .B2(n_230), .Y(n_336) );
INVx5_ASAP7_75t_L g337 ( .A(n_257), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_248), .B(n_241), .Y(n_338) );
OR2x2_ASAP7_75t_L g339 ( .A(n_308), .B(n_218), .Y(n_339) );
NAND2xp5_ASAP7_75t_SL g340 ( .A(n_292), .B(n_241), .Y(n_340) );
NOR2xp33_ASAP7_75t_R g341 ( .A(n_250), .B(n_241), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_286), .B(n_230), .Y(n_342) );
OAI21xp5_ASAP7_75t_L g343 ( .A1(n_286), .A2(n_238), .B(n_241), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_243), .B(n_238), .Y(n_344) );
INVxp67_ASAP7_75t_SL g345 ( .A(n_287), .Y(n_345) );
OAI21xp33_ASAP7_75t_L g346 ( .A1(n_297), .A2(n_295), .B(n_246), .Y(n_346) );
AOI21xp5_ASAP7_75t_L g347 ( .A1(n_313), .A2(n_307), .B(n_299), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_298), .B(n_252), .Y(n_348) );
O2A1O1Ixp33_ASAP7_75t_SL g349 ( .A1(n_274), .A2(n_276), .B(n_283), .C(n_288), .Y(n_349) );
INVx3_ASAP7_75t_L g350 ( .A(n_244), .Y(n_350) );
AOI21xp5_ASAP7_75t_L g351 ( .A1(n_306), .A2(n_261), .B(n_260), .Y(n_351) );
AND2x4_ASAP7_75t_L g352 ( .A(n_281), .B(n_284), .Y(n_352) );
AOI21xp5_ASAP7_75t_L g353 ( .A1(n_291), .A2(n_263), .B(n_265), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_282), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_290), .Y(n_355) );
A2O1A1Ixp33_ASAP7_75t_L g356 ( .A1(n_252), .A2(n_246), .B(n_285), .C(n_269), .Y(n_356) );
A2O1A1Ixp33_ASAP7_75t_L g357 ( .A1(n_269), .A2(n_256), .B(n_289), .C(n_284), .Y(n_357) );
OAI22xp5_ASAP7_75t_L g358 ( .A1(n_289), .A2(n_253), .B1(n_244), .B2(n_251), .Y(n_358) );
A2O1A1Ixp33_ASAP7_75t_L g359 ( .A1(n_296), .A2(n_253), .B(n_262), .C(n_303), .Y(n_359) );
O2A1O1Ixp5_ASAP7_75t_L g360 ( .A1(n_305), .A2(n_272), .B(n_270), .C(n_258), .Y(n_360) );
INVxp67_ASAP7_75t_L g361 ( .A(n_257), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_257), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_302), .B(n_257), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_302), .B(n_257), .Y(n_364) );
OR2x2_ASAP7_75t_L g365 ( .A(n_249), .B(n_264), .Y(n_365) );
BUFx8_ASAP7_75t_L g366 ( .A(n_247), .Y(n_366) );
A2O1A1Ixp33_ASAP7_75t_L g367 ( .A1(n_301), .A2(n_275), .B(n_266), .C(n_247), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_244), .Y(n_368) );
INVx2_ASAP7_75t_SL g369 ( .A(n_341), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_320), .Y(n_370) );
AOI22xp5_ASAP7_75t_L g371 ( .A1(n_352), .A2(n_277), .B1(n_249), .B2(n_247), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_330), .B(n_247), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_323), .B(n_293), .Y(n_373) );
AOI22xp5_ASAP7_75t_L g374 ( .A1(n_352), .A2(n_272), .B1(n_294), .B2(n_279), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_339), .Y(n_375) );
AOI21xp5_ASAP7_75t_L g376 ( .A1(n_357), .A2(n_314), .B(n_279), .Y(n_376) );
NOR2xp33_ASAP7_75t_SL g377 ( .A(n_331), .B(n_345), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_355), .B(n_348), .Y(n_378) );
BUFx3_ASAP7_75t_L g379 ( .A(n_366), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g380 ( .A(n_365), .B(n_346), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_315), .A2(n_316), .B1(n_318), .B2(n_336), .Y(n_381) );
NAND2xp5_ASAP7_75t_SL g382 ( .A(n_328), .B(n_358), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_319), .B(n_354), .Y(n_383) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_333), .B(n_356), .Y(n_384) );
AOI21xp5_ASAP7_75t_L g385 ( .A1(n_349), .A2(n_347), .B(n_335), .Y(n_385) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_338), .A2(n_336), .B1(n_325), .B2(n_317), .Y(n_386) );
NOR2x1_ASAP7_75t_R g387 ( .A(n_337), .B(n_317), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_344), .B(n_317), .Y(n_388) );
OAI21xp5_ASAP7_75t_L g389 ( .A1(n_324), .A2(n_351), .B(n_321), .Y(n_389) );
NAND3xp33_ASAP7_75t_L g390 ( .A(n_359), .B(n_367), .C(n_360), .Y(n_390) );
OR2x2_ASAP7_75t_L g391 ( .A(n_342), .B(n_350), .Y(n_391) );
CKINVDCx5p33_ASAP7_75t_R g392 ( .A(n_366), .Y(n_392) );
INVxp67_ASAP7_75t_SL g393 ( .A(n_328), .Y(n_393) );
O2A1O1Ixp33_ASAP7_75t_SL g394 ( .A1(n_329), .A2(n_340), .B(n_362), .C(n_363), .Y(n_394) );
AO21x1_ASAP7_75t_L g395 ( .A1(n_326), .A2(n_322), .B(n_343), .Y(n_395) );
NOR2xp33_ASAP7_75t_SL g396 ( .A(n_337), .B(n_361), .Y(n_396) );
A2O1A1Ixp33_ASAP7_75t_L g397 ( .A1(n_353), .A2(n_343), .B(n_334), .C(n_364), .Y(n_397) );
AO31x2_ASAP7_75t_L g398 ( .A1(n_368), .A2(n_326), .A3(n_337), .B(n_332), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_327), .Y(n_399) );
A2O1A1Ixp33_ASAP7_75t_L g400 ( .A1(n_346), .A2(n_357), .B(n_212), .C(n_330), .Y(n_400) );
AOI22xp5_ASAP7_75t_L g401 ( .A1(n_352), .A2(n_308), .B1(n_212), .B2(n_225), .Y(n_401) );
AOI21xp5_ASAP7_75t_L g402 ( .A1(n_385), .A2(n_382), .B(n_389), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_370), .B(n_388), .Y(n_403) );
OAI21x1_ASAP7_75t_SL g404 ( .A1(n_381), .A2(n_395), .B(n_371), .Y(n_404) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_392), .Y(n_405) );
OAI21x1_ASAP7_75t_SL g406 ( .A1(n_381), .A2(n_372), .B(n_376), .Y(n_406) );
OA21x2_ASAP7_75t_L g407 ( .A1(n_390), .A2(n_382), .B(n_397), .Y(n_407) );
AO21x2_ASAP7_75t_L g408 ( .A1(n_400), .A2(n_397), .B(n_386), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_384), .B(n_378), .Y(n_409) );
BUFx2_ASAP7_75t_L g410 ( .A(n_387), .Y(n_410) );
AOI21xp5_ASAP7_75t_L g411 ( .A1(n_394), .A2(n_393), .B(n_384), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_378), .A2(n_380), .B1(n_401), .B2(n_379), .Y(n_412) );
INVxp67_ASAP7_75t_SL g413 ( .A(n_379), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_383), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_380), .B(n_375), .Y(n_415) );
A2O1A1Ixp33_ASAP7_75t_L g416 ( .A1(n_374), .A2(n_391), .B(n_373), .C(n_399), .Y(n_416) );
OAI21x1_ASAP7_75t_L g417 ( .A1(n_398), .A2(n_396), .B(n_377), .Y(n_417) );
AOI21xp5_ASAP7_75t_L g418 ( .A1(n_369), .A2(n_385), .B(n_357), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_398), .B(n_330), .Y(n_419) );
AOI221xp5_ASAP7_75t_L g420 ( .A1(n_398), .A2(n_245), .B1(n_378), .B2(n_384), .C(n_267), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_398), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_400), .B(n_330), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_370), .B(n_330), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_400), .B(n_330), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_383), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_370), .Y(n_426) );
AND2x4_ASAP7_75t_L g427 ( .A(n_370), .B(n_388), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_383), .Y(n_428) );
INVx3_ASAP7_75t_L g429 ( .A(n_379), .Y(n_429) );
AOI22xp33_ASAP7_75t_SL g430 ( .A1(n_378), .A2(n_267), .B1(n_308), .B2(n_300), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_407), .Y(n_431) );
AND2x4_ASAP7_75t_L g432 ( .A(n_421), .B(n_417), .Y(n_432) );
OA21x2_ASAP7_75t_L g433 ( .A1(n_402), .A2(n_411), .B(n_418), .Y(n_433) );
OR2x6_ASAP7_75t_L g434 ( .A(n_417), .B(n_421), .Y(n_434) );
AND2x4_ASAP7_75t_L g435 ( .A(n_421), .B(n_417), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_426), .Y(n_436) );
OA21x2_ASAP7_75t_L g437 ( .A1(n_402), .A2(n_411), .B(n_418), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_426), .Y(n_438) );
BUFx2_ASAP7_75t_L g439 ( .A(n_419), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_426), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_423), .B(n_414), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_407), .Y(n_442) );
INVx3_ASAP7_75t_L g443 ( .A(n_427), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_407), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_407), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_407), .Y(n_446) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_419), .Y(n_447) );
BUFx2_ASAP7_75t_SL g448 ( .A(n_429), .Y(n_448) );
AOI21x1_ASAP7_75t_L g449 ( .A1(n_422), .A2(n_424), .B(n_404), .Y(n_449) );
BUFx2_ASAP7_75t_SL g450 ( .A(n_429), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_408), .Y(n_451) );
INVxp67_ASAP7_75t_L g452 ( .A(n_414), .Y(n_452) );
AO21x2_ASAP7_75t_L g453 ( .A1(n_406), .A2(n_404), .B(n_422), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_408), .Y(n_454) );
INVx2_ASAP7_75t_SL g455 ( .A(n_427), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_423), .B(n_428), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_408), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_408), .Y(n_458) );
AOI22xp5_ASAP7_75t_L g459 ( .A1(n_409), .A2(n_420), .B1(n_430), .B2(n_412), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_425), .B(n_428), .Y(n_460) );
OA21x2_ASAP7_75t_L g461 ( .A1(n_424), .A2(n_406), .B(n_416), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_425), .B(n_403), .Y(n_462) );
INVx3_ASAP7_75t_L g463 ( .A(n_427), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_403), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_415), .B(n_409), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_431), .B(n_427), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_439), .B(n_415), .Y(n_467) );
INVx2_ASAP7_75t_SL g468 ( .A(n_432), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_431), .B(n_420), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_431), .B(n_429), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_442), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_442), .B(n_429), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_442), .B(n_413), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g474 ( .A1(n_459), .A2(n_456), .B1(n_465), .B2(n_462), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_436), .Y(n_475) );
OAI31xp33_ASAP7_75t_L g476 ( .A1(n_452), .A2(n_405), .A3(n_410), .B(n_460), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_436), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_439), .B(n_410), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_444), .B(n_446), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_438), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_444), .B(n_445), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_444), .B(n_445), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g483 ( .A1(n_459), .A2(n_456), .B1(n_452), .B2(n_460), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_439), .B(n_447), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_445), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_462), .B(n_456), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_438), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_440), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_440), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_446), .B(n_451), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_447), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_446), .Y(n_492) );
AND2x4_ASAP7_75t_L g493 ( .A(n_432), .B(n_435), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_460), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_465), .B(n_441), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_454), .B(n_458), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_454), .B(n_458), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_465), .B(n_441), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_454), .B(n_457), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_449), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_462), .B(n_464), .Y(n_501) );
INVx2_ASAP7_75t_SL g502 ( .A(n_432), .Y(n_502) );
BUFx2_ASAP7_75t_L g503 ( .A(n_434), .Y(n_503) );
BUFx3_ASAP7_75t_L g504 ( .A(n_443), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_457), .B(n_458), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_464), .B(n_463), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_457), .B(n_453), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_433), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_449), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_432), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_433), .Y(n_511) );
INVxp67_ASAP7_75t_SL g512 ( .A(n_432), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_453), .B(n_461), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_475), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_475), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_466), .B(n_453), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_466), .B(n_453), .Y(n_517) );
INVx1_ASAP7_75t_SL g518 ( .A(n_473), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_486), .B(n_463), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_477), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_477), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_480), .Y(n_522) );
OR2x2_ASAP7_75t_L g523 ( .A(n_484), .B(n_453), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_480), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_487), .Y(n_525) );
OR2x2_ASAP7_75t_L g526 ( .A(n_484), .B(n_433), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_491), .B(n_433), .Y(n_527) );
BUFx2_ASAP7_75t_L g528 ( .A(n_512), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_466), .B(n_435), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_486), .B(n_435), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_487), .Y(n_531) );
INVx4_ASAP7_75t_L g532 ( .A(n_473), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_471), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_494), .B(n_463), .Y(n_534) );
INVx1_ASAP7_75t_SL g535 ( .A(n_473), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_469), .B(n_435), .Y(n_536) );
AND2x4_ASAP7_75t_L g537 ( .A(n_493), .B(n_435), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_469), .B(n_461), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_471), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_488), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_488), .Y(n_541) );
AND2x6_ASAP7_75t_SL g542 ( .A(n_495), .B(n_434), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_469), .B(n_461), .Y(n_543) );
INVx2_ASAP7_75t_SL g544 ( .A(n_493), .Y(n_544) );
INVxp67_ASAP7_75t_L g545 ( .A(n_478), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_489), .Y(n_546) );
AND2x4_ASAP7_75t_L g547 ( .A(n_493), .B(n_434), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_493), .B(n_461), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_470), .B(n_461), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_476), .B(n_455), .Y(n_550) );
AND2x2_ASAP7_75t_SL g551 ( .A(n_503), .B(n_461), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_470), .B(n_433), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_470), .B(n_433), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_472), .B(n_437), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_472), .B(n_437), .Y(n_555) );
HB1xp67_ASAP7_75t_L g556 ( .A(n_478), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_489), .Y(n_557) );
INVxp67_ASAP7_75t_L g558 ( .A(n_467), .Y(n_558) );
INVx2_ASAP7_75t_SL g559 ( .A(n_472), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_494), .B(n_437), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_510), .B(n_437), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_506), .Y(n_562) );
HB1xp67_ASAP7_75t_L g563 ( .A(n_491), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_467), .B(n_437), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_506), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_501), .B(n_463), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_501), .B(n_463), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_474), .B(n_443), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_510), .B(n_437), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_513), .B(n_434), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_495), .B(n_443), .Y(n_571) );
OR2x2_ASAP7_75t_L g572 ( .A(n_498), .B(n_434), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_498), .B(n_443), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_563), .Y(n_574) );
NOR2xp67_ASAP7_75t_L g575 ( .A(n_532), .B(n_544), .Y(n_575) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_532), .Y(n_576) );
NOR2xp67_ASAP7_75t_L g577 ( .A(n_532), .B(n_502), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_514), .Y(n_578) );
AND2x2_ASAP7_75t_SL g579 ( .A(n_528), .B(n_503), .Y(n_579) );
INVx2_ASAP7_75t_SL g580 ( .A(n_537), .Y(n_580) );
INVx3_ASAP7_75t_L g581 ( .A(n_542), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_514), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_530), .B(n_513), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_530), .B(n_513), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_558), .B(n_483), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_533), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_536), .B(n_512), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_536), .B(n_468), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_556), .B(n_483), .Y(n_589) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_550), .A2(n_502), .B1(n_468), .B2(n_455), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_516), .B(n_468), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_545), .B(n_476), .Y(n_592) );
BUFx2_ASAP7_75t_L g593 ( .A(n_528), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_515), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_533), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_516), .B(n_502), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_517), .B(n_507), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_518), .B(n_492), .Y(n_598) );
AND2x4_ASAP7_75t_L g599 ( .A(n_544), .B(n_507), .Y(n_599) );
NAND2xp5_ASAP7_75t_SL g600 ( .A(n_535), .B(n_492), .Y(n_600) );
INVx1_ASAP7_75t_SL g601 ( .A(n_572), .Y(n_601) );
AO22x2_ASAP7_75t_L g602 ( .A1(n_562), .A2(n_511), .B1(n_508), .B2(n_509), .Y(n_602) );
AND2x4_ASAP7_75t_L g603 ( .A(n_547), .B(n_507), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_515), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_520), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_517), .B(n_490), .Y(n_606) );
OR2x2_ASAP7_75t_L g607 ( .A(n_519), .B(n_485), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_562), .B(n_481), .Y(n_608) );
AOI21xp33_ASAP7_75t_SL g609 ( .A1(n_551), .A2(n_455), .B(n_434), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_565), .B(n_482), .Y(n_610) );
NAND2x1_ASAP7_75t_L g611 ( .A(n_547), .B(n_434), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_538), .B(n_490), .Y(n_612) );
AOI222xp33_ASAP7_75t_L g613 ( .A1(n_538), .A2(n_496), .B1(n_505), .B2(n_499), .C1(n_497), .C2(n_490), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_565), .B(n_479), .Y(n_614) );
OR2x2_ASAP7_75t_L g615 ( .A(n_564), .B(n_511), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_543), .B(n_479), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_543), .B(n_479), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_520), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_521), .Y(n_619) );
OR2x2_ASAP7_75t_L g620 ( .A(n_572), .B(n_573), .Y(n_620) );
INVxp67_ASAP7_75t_SL g621 ( .A(n_539), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_529), .B(n_482), .Y(n_622) );
NAND2xp67_ASAP7_75t_L g623 ( .A(n_560), .B(n_511), .Y(n_623) );
OR2x2_ASAP7_75t_L g624 ( .A(n_564), .B(n_508), .Y(n_624) );
AND2x4_ASAP7_75t_SL g625 ( .A(n_537), .B(n_482), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_529), .B(n_481), .Y(n_626) );
NAND2xp5_ASAP7_75t_SL g627 ( .A(n_527), .B(n_485), .Y(n_627) );
INVx1_ASAP7_75t_SL g628 ( .A(n_537), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_574), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_625), .B(n_570), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_578), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_625), .B(n_570), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_582), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_583), .B(n_547), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_594), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_613), .B(n_560), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_597), .B(n_527), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_597), .B(n_569), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_608), .B(n_569), .Y(n_639) );
NOR3xp33_ASAP7_75t_L g640 ( .A(n_592), .B(n_568), .C(n_508), .Y(n_640) );
INVx3_ASAP7_75t_L g641 ( .A(n_581), .Y(n_641) );
OAI22xp5_ASAP7_75t_L g642 ( .A1(n_581), .A2(n_559), .B1(n_567), .B2(n_566), .Y(n_642) );
AND2x4_ASAP7_75t_L g643 ( .A(n_575), .B(n_561), .Y(n_643) );
OR2x2_ASAP7_75t_L g644 ( .A(n_615), .B(n_523), .Y(n_644) );
AND2x4_ASAP7_75t_L g645 ( .A(n_577), .B(n_561), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_604), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_583), .B(n_548), .Y(n_647) );
AND2x2_ASAP7_75t_L g648 ( .A(n_584), .B(n_548), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_605), .Y(n_649) );
O2A1O1Ixp33_ASAP7_75t_L g650 ( .A1(n_581), .A2(n_526), .B(n_557), .C(n_546), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_618), .Y(n_651) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_623), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_584), .B(n_559), .Y(n_653) );
OR2x2_ASAP7_75t_L g654 ( .A(n_615), .B(n_624), .Y(n_654) );
OR2x2_ASAP7_75t_L g655 ( .A(n_624), .B(n_523), .Y(n_655) );
OR2x2_ASAP7_75t_L g656 ( .A(n_616), .B(n_526), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_619), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_610), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_614), .B(n_524), .Y(n_659) );
AOI221xp5_ASAP7_75t_L g660 ( .A1(n_585), .A2(n_524), .B1(n_557), .B2(n_546), .C(n_541), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_607), .Y(n_661) );
OR2x2_ASAP7_75t_L g662 ( .A(n_616), .B(n_571), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_606), .B(n_521), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_606), .B(n_531), .Y(n_664) );
NAND2x1p5_ASAP7_75t_L g665 ( .A(n_579), .B(n_504), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_620), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_600), .Y(n_667) );
OAI21xp33_ASAP7_75t_L g668 ( .A1(n_636), .A2(n_576), .B(n_590), .Y(n_668) );
INVx2_ASAP7_75t_L g669 ( .A(n_654), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_636), .B(n_589), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_647), .B(n_617), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_640), .A2(n_551), .B1(n_599), .B2(n_603), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g673 ( .A1(n_666), .A2(n_551), .B1(n_599), .B2(n_603), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_663), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_658), .B(n_612), .Y(n_675) );
OAI21xp5_ASAP7_75t_L g676 ( .A1(n_650), .A2(n_652), .B(n_642), .Y(n_676) );
OAI22xp5_ASAP7_75t_L g677 ( .A1(n_641), .A2(n_579), .B1(n_580), .B2(n_611), .Y(n_677) );
INVxp67_ASAP7_75t_L g678 ( .A(n_629), .Y(n_678) );
OAI221xp5_ASAP7_75t_SL g679 ( .A1(n_641), .A2(n_628), .B1(n_601), .B2(n_580), .C(n_596), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_663), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_664), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_664), .B(n_593), .Y(n_682) );
OAI21xp5_ASAP7_75t_L g683 ( .A1(n_642), .A2(n_609), .B(n_600), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_661), .B(n_612), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_634), .B(n_626), .Y(n_685) );
OR2x2_ASAP7_75t_L g686 ( .A(n_656), .B(n_617), .Y(n_686) );
AOI21xp5_ASAP7_75t_L g687 ( .A1(n_665), .A2(n_627), .B(n_602), .Y(n_687) );
OAI211xp5_ASAP7_75t_L g688 ( .A1(n_660), .A2(n_627), .B(n_591), .C(n_596), .Y(n_688) );
AOI21xp33_ASAP7_75t_L g689 ( .A1(n_667), .A2(n_602), .B(n_531), .Y(n_689) );
AOI21xp33_ASAP7_75t_L g690 ( .A1(n_659), .A2(n_602), .B(n_541), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_645), .A2(n_603), .B1(n_599), .B2(n_591), .Y(n_691) );
NAND3xp33_ASAP7_75t_SL g692 ( .A(n_676), .B(n_665), .C(n_630), .Y(n_692) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_668), .A2(n_645), .B1(n_643), .B2(n_637), .Y(n_693) );
NAND2xp5_ASAP7_75t_SL g694 ( .A(n_687), .B(n_643), .Y(n_694) );
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_670), .A2(n_637), .B1(n_639), .B2(n_659), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_674), .Y(n_696) );
NAND4xp25_ASAP7_75t_SL g697 ( .A(n_672), .B(n_632), .C(n_638), .D(n_653), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_680), .Y(n_698) );
AOI31xp33_ASAP7_75t_L g699 ( .A1(n_683), .A2(n_655), .A3(n_644), .B(n_638), .Y(n_699) );
OAI221xp5_ASAP7_75t_SL g700 ( .A1(n_672), .A2(n_639), .B1(n_662), .B2(n_588), .C(n_587), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g701 ( .A1(n_688), .A2(n_657), .B1(n_651), .B2(n_649), .Y(n_701) );
AOI21xp33_ASAP7_75t_L g702 ( .A1(n_678), .A2(n_631), .B(n_646), .Y(n_702) );
OAI21xp33_ASAP7_75t_L g703 ( .A1(n_679), .A2(n_648), .B(n_635), .Y(n_703) );
AOI22xp5_ASAP7_75t_L g704 ( .A1(n_682), .A2(n_633), .B1(n_588), .B2(n_587), .Y(n_704) );
AOI321xp33_ASAP7_75t_L g705 ( .A1(n_673), .A2(n_554), .A3(n_552), .B1(n_555), .B2(n_553), .C(n_549), .Y(n_705) );
NAND4xp25_ASAP7_75t_L g706 ( .A(n_692), .B(n_673), .C(n_677), .D(n_691), .Y(n_706) );
NAND4xp75_ASAP7_75t_L g707 ( .A(n_694), .B(n_689), .C(n_690), .D(n_682), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_695), .B(n_681), .Y(n_708) );
OAI211xp5_ASAP7_75t_SL g709 ( .A1(n_693), .A2(n_675), .B(n_684), .C(n_669), .Y(n_709) );
AOI21xp5_ASAP7_75t_L g710 ( .A1(n_699), .A2(n_697), .B(n_700), .Y(n_710) );
OAI211xp5_ASAP7_75t_L g711 ( .A1(n_705), .A2(n_669), .B(n_686), .C(n_671), .Y(n_711) );
AOI21xp33_ASAP7_75t_L g712 ( .A1(n_701), .A2(n_522), .B(n_525), .Y(n_712) );
AND2x2_ASAP7_75t_L g713 ( .A(n_704), .B(n_671), .Y(n_713) );
AOI221xp5_ASAP7_75t_L g714 ( .A1(n_710), .A2(n_702), .B1(n_703), .B2(n_698), .C(n_696), .Y(n_714) );
NAND5xp2_ASAP7_75t_L g715 ( .A(n_711), .B(n_555), .C(n_554), .D(n_553), .E(n_552), .Y(n_715) );
AOI211x1_ASAP7_75t_SL g716 ( .A1(n_706), .A2(n_534), .B(n_595), .C(n_586), .Y(n_716) );
AOI21xp5_ASAP7_75t_L g717 ( .A1(n_712), .A2(n_621), .B(n_685), .Y(n_717) );
A2O1A1Ixp33_ASAP7_75t_L g718 ( .A1(n_709), .A2(n_626), .B(n_622), .C(n_598), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_716), .B(n_713), .Y(n_719) );
OR5x1_ASAP7_75t_L g720 ( .A(n_714), .B(n_707), .C(n_708), .D(n_448), .E(n_450), .Y(n_720) );
NAND3xp33_ASAP7_75t_SL g721 ( .A(n_718), .B(n_622), .C(n_522), .Y(n_721) );
AND3x4_ASAP7_75t_L g722 ( .A(n_720), .B(n_715), .C(n_717), .Y(n_722) );
XOR2xp5_ASAP7_75t_L g723 ( .A(n_719), .B(n_448), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_723), .Y(n_724) );
BUFx2_ASAP7_75t_L g725 ( .A(n_724), .Y(n_725) );
AOI21xp33_ASAP7_75t_SL g726 ( .A1(n_725), .A2(n_722), .B(n_721), .Y(n_726) );
NAND3xp33_ASAP7_75t_L g727 ( .A(n_726), .B(n_540), .C(n_525), .Y(n_727) );
AO221x1_ASAP7_75t_L g728 ( .A1(n_727), .A2(n_540), .B1(n_595), .B2(n_586), .C(n_500), .Y(n_728) );
AOI22xp5_ASAP7_75t_L g729 ( .A1(n_728), .A2(n_448), .B1(n_450), .B2(n_549), .Y(n_729) );
endmodule