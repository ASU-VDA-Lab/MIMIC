module fake_jpeg_2258_n_573 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_573);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_573;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_18),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_18),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_17),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_17),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx14_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_3),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_17),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_53),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_29),
.Y(n_54)
);

INVx4_ASAP7_75t_SL g147 ( 
.A(n_54),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_20),
.B(n_16),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_55),
.B(n_57),
.Y(n_114)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_56),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_20),
.B(n_16),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_58),
.Y(n_128)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_59),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_60),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

BUFx8_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx13_ASAP7_75t_L g169 ( 
.A(n_62),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_63),
.Y(n_139)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_64),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_30),
.B(n_15),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_65),
.B(n_68),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_66),
.Y(n_146)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_28),
.Y(n_67)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_67),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_30),
.B(n_15),
.Y(n_68)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_70),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_71),
.Y(n_154)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_72),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_0),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_73),
.B(n_91),
.Y(n_145)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_74),
.Y(n_123)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_76),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_48),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_77),
.B(n_78),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_0),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_79),
.Y(n_166)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_80),
.Y(n_140)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_26),
.Y(n_81)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_81),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_82),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_83),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_35),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_84),
.B(n_87),
.Y(n_161)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_50),
.Y(n_85)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_85),
.Y(n_124)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_86),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_48),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_88),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_49),
.Y(n_89)
);

INVx6_ASAP7_75t_SL g138 ( 
.A(n_89),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_90),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_31),
.B(n_0),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_33),
.Y(n_92)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_92),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_38),
.B(n_1),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_93),
.B(n_100),
.Y(n_158)
);

INVx11_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx5_ASAP7_75t_SL g111 ( 
.A(n_94),
.Y(n_111)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_38),
.Y(n_95)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_95),
.Y(n_151)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_33),
.Y(n_97)
);

INVx8_ASAP7_75t_L g143 ( 
.A(n_97),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_98),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_33),
.Y(n_99)
);

BUFx5_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_42),
.B(n_1),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_101),
.Y(n_155)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_47),
.Y(n_102)
);

INVx3_ASAP7_75t_SL g116 ( 
.A(n_102),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_51),
.B(n_1),
.Y(n_103)
);

AOI21xp33_ASAP7_75t_L g136 ( 
.A1(n_103),
.A2(n_45),
.B(n_42),
.Y(n_136)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_44),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g144 ( 
.A(n_104),
.Y(n_144)
);

INVx4_ASAP7_75t_SL g105 ( 
.A(n_21),
.Y(n_105)
);

INVx3_ASAP7_75t_SL g122 ( 
.A(n_105),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g106 ( 
.A(n_44),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_74),
.A2(n_103),
.B1(n_96),
.B2(n_101),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_108),
.A2(n_167),
.B1(n_46),
.B2(n_25),
.Y(n_216)
);

BUFx12_ASAP7_75t_L g113 ( 
.A(n_62),
.Y(n_113)
);

BUFx10_ASAP7_75t_L g228 ( 
.A(n_113),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_62),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_115),
.B(n_119),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_69),
.Y(n_119)
);

INVx3_ASAP7_75t_SL g126 ( 
.A(n_105),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_126),
.Y(n_180)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_53),
.Y(n_130)
);

INVx4_ASAP7_75t_SL g207 ( 
.A(n_130),
.Y(n_207)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_67),
.Y(n_133)
);

INVx4_ASAP7_75t_SL g215 ( 
.A(n_133),
.Y(n_215)
);

HAxp5_ASAP7_75t_SL g135 ( 
.A(n_81),
.B(n_32),
.CON(n_135),
.SN(n_135)
);

NOR3xp33_ASAP7_75t_L g199 ( 
.A(n_135),
.B(n_148),
.C(n_39),
.Y(n_199)
);

AND2x2_ASAP7_75t_SL g189 ( 
.A(n_136),
.B(n_153),
.Y(n_189)
);

AND2x2_ASAP7_75t_SL g148 ( 
.A(n_56),
.B(n_64),
.Y(n_148)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_70),
.Y(n_152)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_152),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_86),
.B(n_51),
.Y(n_153)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_102),
.Y(n_156)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_156),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_54),
.A2(n_51),
.B1(n_22),
.B2(n_24),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_159),
.A2(n_25),
.B(n_44),
.Y(n_214)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_83),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_160),
.B(n_58),
.Y(n_173)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_60),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_165),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_98),
.A2(n_46),
.B1(n_22),
.B2(n_24),
.Y(n_167)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_170),
.Y(n_171)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_171),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_138),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_172),
.B(n_178),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_173),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_145),
.B(n_45),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_174),
.B(n_232),
.C(n_122),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_149),
.A2(n_79),
.B1(n_61),
.B2(n_63),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_175),
.A2(n_183),
.B1(n_196),
.B2(n_214),
.Y(n_257)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_176),
.Y(n_239)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_157),
.Y(n_177)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_177),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_114),
.B(n_31),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_135),
.A2(n_54),
.B1(n_58),
.B2(n_88),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_181),
.Y(n_274)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_128),
.Y(n_182)
);

BUFx2_ASAP7_75t_L g264 ( 
.A(n_182),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_167),
.A2(n_66),
.B1(n_71),
.B2(n_82),
.Y(n_183)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_110),
.Y(n_184)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_184),
.Y(n_240)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_155),
.Y(n_185)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_185),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_153),
.B(n_90),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g280 ( 
.A(n_186),
.B(n_191),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_114),
.B(n_40),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_187),
.B(n_198),
.Y(n_281)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_140),
.Y(n_188)
);

INVx3_ASAP7_75t_SL g256 ( 
.A(n_188),
.Y(n_256)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_151),
.Y(n_190)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_190),
.Y(n_241)
);

NAND2x2_ASAP7_75t_SL g191 ( 
.A(n_148),
.B(n_32),
.Y(n_191)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_110),
.Y(n_192)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_192),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_122),
.Y(n_193)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_193),
.Y(n_245)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_118),
.Y(n_195)
);

INVx5_ASAP7_75t_L g243 ( 
.A(n_195),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_159),
.A2(n_94),
.B1(n_104),
.B2(n_21),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_147),
.Y(n_197)
);

INVx5_ASAP7_75t_L g272 ( 
.A(n_197),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_161),
.B(n_92),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_199),
.B(n_211),
.Y(n_285)
);

OAI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_149),
.A2(n_22),
.B1(n_24),
.B2(n_21),
.Y(n_200)
);

OA22x2_ASAP7_75t_L g266 ( 
.A1(n_200),
.A2(n_129),
.B1(n_165),
.B2(n_127),
.Y(n_266)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_120),
.Y(n_201)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_201),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_125),
.B(n_37),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_202),
.B(n_204),
.Y(n_238)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_137),
.Y(n_203)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_203),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_158),
.B(n_37),
.Y(n_204)
);

CKINVDCx6p67_ASAP7_75t_R g205 ( 
.A(n_169),
.Y(n_205)
);

INVx13_ASAP7_75t_L g236 ( 
.A(n_205),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_125),
.B(n_39),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_206),
.B(n_210),
.Y(n_246)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_143),
.Y(n_208)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_208),
.Y(n_277)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_131),
.Y(n_209)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_209),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_109),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_161),
.A2(n_40),
.B1(n_41),
.B2(n_46),
.Y(n_211)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_107),
.Y(n_213)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_213),
.Y(n_265)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_216),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_112),
.A2(n_41),
.B1(n_25),
.B2(n_44),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_217),
.A2(n_226),
.B1(n_146),
.B2(n_166),
.Y(n_244)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_143),
.Y(n_219)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_219),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_121),
.B(n_99),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_220),
.B(n_221),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_123),
.B(n_124),
.Y(n_221)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_130),
.Y(n_222)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_222),
.Y(n_269)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_133),
.Y(n_223)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_223),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_109),
.B(n_99),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_224),
.B(n_225),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_162),
.B(n_97),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_118),
.A2(n_166),
.B1(n_154),
.B2(n_146),
.Y(n_226)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_168),
.Y(n_227)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_227),
.Y(n_267)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_163),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_229),
.B(n_231),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_147),
.Y(n_230)
);

BUFx5_ASAP7_75t_L g237 ( 
.A(n_230),
.Y(n_237)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_117),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_142),
.B(n_97),
.Y(n_232)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_150),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_233),
.B(n_180),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_189),
.B(n_191),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_234),
.B(n_260),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_235),
.B(n_34),
.Y(n_331)
);

AO22x1_ASAP7_75t_SL g242 ( 
.A1(n_191),
.A2(n_126),
.B1(n_116),
.B2(n_164),
.Y(n_242)
);

OA21x2_ASAP7_75t_L g315 ( 
.A1(n_242),
.A2(n_113),
.B(n_117),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_244),
.B(n_266),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_189),
.B(n_116),
.C(n_154),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_249),
.B(n_278),
.C(n_286),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_212),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_258),
.B(n_271),
.Y(n_317)
);

OAI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_183),
.A2(n_181),
.B1(n_200),
.B2(n_199),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g321 ( 
.A1(n_259),
.A2(n_34),
.B1(n_33),
.B2(n_5),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_186),
.B(n_129),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_268),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_205),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_194),
.B(n_111),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g301 ( 
.A(n_273),
.B(n_171),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_196),
.A2(n_127),
.B1(n_132),
.B2(n_139),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_276),
.A2(n_180),
.B1(n_193),
.B2(n_179),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_218),
.B(n_111),
.Y(n_278)
);

INVx8_ASAP7_75t_L g282 ( 
.A(n_205),
.Y(n_282)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_282),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_227),
.B(n_132),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_283),
.B(n_287),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_229),
.B(n_139),
.C(n_169),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_179),
.B(n_195),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_263),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_289),
.B(n_293),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_281),
.B(n_177),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_290),
.B(n_292),
.Y(n_353)
);

INVx13_ASAP7_75t_L g291 ( 
.A(n_236),
.Y(n_291)
);

INVx1_ASAP7_75t_SL g359 ( 
.A(n_291),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_262),
.B(n_230),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_262),
.B(n_197),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_294),
.A2(n_306),
.B1(n_321),
.B2(n_337),
.Y(n_350)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_245),
.Y(n_295)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_295),
.Y(n_358)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_275),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_296),
.Y(n_349)
);

AND2x6_ASAP7_75t_L g300 ( 
.A(n_234),
.B(n_228),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_300),
.B(n_327),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_301),
.B(n_310),
.Y(n_354)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_283),
.Y(n_302)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_302),
.Y(n_355)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_245),
.Y(n_303)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_303),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_252),
.A2(n_41),
.B1(n_92),
.B2(n_219),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_305),
.A2(n_315),
.B1(n_320),
.B2(n_319),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_252),
.A2(n_192),
.B1(n_208),
.B2(n_215),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_239),
.Y(n_307)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_307),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_274),
.A2(n_215),
.B(n_207),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_308),
.A2(n_279),
.B(n_272),
.Y(n_381)
);

AO22x2_ASAP7_75t_L g309 ( 
.A1(n_257),
.A2(n_144),
.B1(n_44),
.B2(n_106),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_309),
.B(n_316),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_250),
.B(n_207),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_239),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_311),
.B(n_323),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_251),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_313),
.Y(n_366)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_275),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_314),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_247),
.B(n_1),
.Y(n_316)
);

INVx13_ASAP7_75t_L g318 ( 
.A(n_236),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_318),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_280),
.A2(n_228),
.B(n_134),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g340 ( 
.A1(n_319),
.A2(n_274),
.B(n_272),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_280),
.A2(n_34),
.B1(n_33),
.B2(n_228),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_235),
.B(n_34),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_322),
.B(n_242),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_246),
.B(n_238),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_284),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_324),
.B(n_326),
.Y(n_373)
);

INVx6_ASAP7_75t_SL g325 ( 
.A(n_282),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_325),
.Y(n_363)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_284),
.Y(n_326)
);

INVx5_ASAP7_75t_L g327 ( 
.A(n_243),
.Y(n_327)
);

INVx8_ASAP7_75t_L g328 ( 
.A(n_243),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_328),
.B(n_329),
.Y(n_351)
);

INVx13_ASAP7_75t_L g329 ( 
.A(n_237),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_240),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_330),
.B(n_332),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_331),
.B(n_335),
.C(n_242),
.Y(n_339)
);

NOR2x1_ASAP7_75t_L g332 ( 
.A(n_285),
.B(n_34),
.Y(n_332)
);

INVx2_ASAP7_75t_SL g333 ( 
.A(n_264),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_333),
.B(n_334),
.Y(n_347)
);

AND2x6_ASAP7_75t_L g334 ( 
.A(n_249),
.B(n_2),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_278),
.B(n_2),
.C(n_3),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_287),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_336),
.B(n_253),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_285),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_338),
.B(n_339),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_340),
.Y(n_408)
);

CKINVDCx14_ASAP7_75t_R g418 ( 
.A(n_341),
.Y(n_418)
);

NAND2x1_ASAP7_75t_L g342 ( 
.A(n_308),
.B(n_286),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_L g387 ( 
.A1(n_342),
.A2(n_381),
.B(n_315),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g344 ( 
.A(n_322),
.B(n_331),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_344),
.B(n_370),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_288),
.A2(n_285),
.B1(n_276),
.B2(n_244),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_345),
.A2(n_346),
.B1(n_361),
.B2(n_367),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_288),
.A2(n_266),
.B1(n_260),
.B2(n_255),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_312),
.B(n_255),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_356),
.B(n_360),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_288),
.A2(n_266),
.B1(n_240),
.B2(n_265),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_357),
.A2(n_362),
.B1(n_372),
.B2(n_291),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_312),
.B(n_266),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_336),
.A2(n_261),
.B1(n_277),
.B2(n_270),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_302),
.A2(n_261),
.B1(n_269),
.B2(n_270),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_298),
.A2(n_277),
.B1(n_267),
.B2(n_264),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_298),
.B(n_254),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_299),
.A2(n_267),
.B1(n_248),
.B2(n_256),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_375),
.B(n_376),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_299),
.B(n_241),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_335),
.B(n_237),
.Y(n_377)
);

MAJx2_ASAP7_75t_L g400 ( 
.A(n_377),
.B(n_320),
.C(n_314),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_304),
.B(n_248),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_378),
.B(n_363),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_313),
.B(n_256),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_379),
.B(n_380),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_316),
.B(n_304),
.Y(n_380)
);

CKINVDCx16_ASAP7_75t_R g382 ( 
.A(n_352),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_382),
.B(n_388),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_366),
.B(n_317),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g449 ( 
.A(n_384),
.B(n_385),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_366),
.B(n_279),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_343),
.A2(n_309),
.B1(n_300),
.B2(n_334),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_386),
.B(n_389),
.Y(n_425)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_387),
.A2(n_368),
.B(n_342),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_373),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_343),
.A2(n_309),
.B1(n_294),
.B2(n_306),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_SL g390 ( 
.A(n_354),
.B(n_332),
.Y(n_390)
);

NAND3xp33_ASAP7_75t_L g421 ( 
.A(n_390),
.B(n_391),
.C(n_396),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_353),
.B(n_330),
.Y(n_391)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_394),
.Y(n_419)
);

AND2x6_ASAP7_75t_L g395 ( 
.A(n_348),
.B(n_315),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_395),
.B(n_399),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_364),
.B(n_303),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_365),
.Y(n_397)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_397),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g398 ( 
.A(n_380),
.B(n_325),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_398),
.B(n_406),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_345),
.A2(n_309),
.B1(n_305),
.B2(n_327),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_400),
.B(n_338),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_379),
.B(n_296),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_402),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_360),
.A2(n_328),
.B1(n_297),
.B2(n_333),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_403),
.B(n_407),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_367),
.B(n_297),
.Y(n_404)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_404),
.Y(n_424)
);

BUFx4f_ASAP7_75t_SL g405 ( 
.A(n_359),
.Y(n_405)
);

CKINVDCx16_ASAP7_75t_R g443 ( 
.A(n_405),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_376),
.B(n_333),
.Y(n_406)
);

AND2x6_ASAP7_75t_L g407 ( 
.A(n_347),
.B(n_329),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_378),
.B(n_318),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_409),
.B(n_414),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_410),
.B(n_357),
.Y(n_432)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_365),
.Y(n_411)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_411),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_355),
.B(n_6),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_355),
.B(n_6),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_415),
.B(n_417),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_347),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_416),
.B(n_8),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_358),
.B(n_7),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_401),
.B(n_370),
.C(n_344),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_427),
.B(n_430),
.C(n_436),
.Y(n_462)
);

MAJIxp5_ASAP7_75t_SL g478 ( 
.A(n_428),
.B(n_405),
.C(n_11),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_382),
.B(n_351),
.Y(n_429)
);

CKINVDCx16_ASAP7_75t_R g471 ( 
.A(n_429),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_401),
.B(n_339),
.C(n_377),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_418),
.A2(n_356),
.B1(n_346),
.B2(n_341),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_431),
.A2(n_445),
.B1(n_415),
.B2(n_414),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_432),
.A2(n_399),
.B1(n_389),
.B2(n_383),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g433 ( 
.A1(n_408),
.A2(n_340),
.B(n_381),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g457 ( 
.A(n_433),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_393),
.B(n_342),
.C(n_372),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_437),
.A2(n_439),
.B(n_390),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_392),
.A2(n_361),
.B1(n_374),
.B2(n_350),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_438),
.A2(n_383),
.B1(n_403),
.B2(n_392),
.Y(n_456)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_408),
.A2(n_359),
.B(n_369),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_396),
.B(n_374),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_441),
.B(n_406),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_393),
.B(n_371),
.C(n_349),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_444),
.B(n_400),
.C(n_413),
.Y(n_464)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_397),
.Y(n_447)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_447),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_412),
.B(n_349),
.Y(n_448)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_448),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_394),
.Y(n_450)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_450),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_388),
.B(n_371),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_451),
.B(n_10),
.Y(n_479)
);

INVx2_ASAP7_75t_SL g452 ( 
.A(n_420),
.Y(n_452)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_452),
.Y(n_482)
);

XNOR2x1_ASAP7_75t_L g498 ( 
.A(n_454),
.B(n_461),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_451),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_455),
.B(n_459),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_456),
.A2(n_475),
.B1(n_477),
.B2(n_480),
.Y(n_488)
);

INVx3_ASAP7_75t_L g458 ( 
.A(n_419),
.Y(n_458)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_458),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_448),
.Y(n_459)
);

XNOR2x1_ASAP7_75t_SL g461 ( 
.A(n_428),
.B(n_387),
.Y(n_461)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_463),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_464),
.B(n_465),
.Y(n_481)
);

OA22x2_ASAP7_75t_L g467 ( 
.A1(n_419),
.A2(n_410),
.B1(n_407),
.B2(n_395),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_467),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_449),
.B(n_398),
.Y(n_468)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_468),
.Y(n_486)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_446),
.Y(n_469)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_469),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_426),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_470),
.B(n_474),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_449),
.B(n_412),
.Y(n_472)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_472),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_473),
.A2(n_434),
.B1(n_450),
.B2(n_422),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_423),
.B(n_416),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_431),
.A2(n_386),
.B1(n_413),
.B2(n_411),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_427),
.B(n_400),
.C(n_405),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_476),
.B(n_430),
.C(n_444),
.Y(n_491)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_440),
.A2(n_405),
.B1(n_11),
.B2(n_12),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_SL g503 ( 
.A(n_478),
.B(n_422),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_479),
.B(n_443),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_421),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_476),
.B(n_436),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_489),
.B(n_495),
.Y(n_505)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_490),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_491),
.B(n_502),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_462),
.B(n_437),
.C(n_439),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_492),
.B(n_494),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_462),
.B(n_433),
.C(n_425),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_461),
.B(n_464),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_471),
.B(n_426),
.Y(n_496)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_496),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_457),
.B(n_425),
.C(n_440),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_497),
.B(n_504),
.C(n_424),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_501),
.A2(n_458),
.B1(n_456),
.B2(n_460),
.Y(n_512)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_475),
.B(n_442),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_503),
.B(n_465),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_457),
.B(n_442),
.C(n_447),
.Y(n_504)
);

OR2x2_ASAP7_75t_L g539 ( 
.A(n_508),
.B(n_512),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g509 ( 
.A1(n_484),
.A2(n_460),
.B(n_467),
.Y(n_509)
);

OAI21x1_ASAP7_75t_SL g531 ( 
.A1(n_509),
.A2(n_520),
.B(n_521),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_511),
.B(n_513),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_494),
.B(n_467),
.C(n_452),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g514 ( 
.A1(n_500),
.A2(n_454),
.B(n_467),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_SL g533 ( 
.A1(n_514),
.A2(n_485),
.B(n_498),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_486),
.A2(n_477),
.B1(n_432),
.B2(n_466),
.Y(n_515)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_515),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_499),
.B(n_466),
.Y(n_516)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_516),
.Y(n_527)
);

INVxp67_ASAP7_75t_L g517 ( 
.A(n_482),
.Y(n_517)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_517),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_498),
.A2(n_432),
.B1(n_452),
.B2(n_443),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_518),
.B(n_523),
.Y(n_537)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_504),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_519),
.B(n_481),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_493),
.B(n_453),
.Y(n_520)
);

INVx13_ASAP7_75t_L g521 ( 
.A(n_487),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_488),
.A2(n_438),
.B1(n_453),
.B2(n_469),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_510),
.B(n_489),
.C(n_491),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_524),
.B(n_526),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_SL g528 ( 
.A(n_522),
.B(n_483),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_528),
.B(n_530),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_506),
.B(n_481),
.C(n_492),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_506),
.B(n_497),
.C(n_495),
.Y(n_532)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_532),
.B(n_511),
.C(n_505),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_SL g546 ( 
.A(n_533),
.B(n_536),
.Y(n_546)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_513),
.B(n_502),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_534),
.B(n_523),
.Y(n_543)
);

OAI21xp5_ASAP7_75t_SL g536 ( 
.A1(n_509),
.A2(n_514),
.B(n_518),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g550 ( 
.A1(n_536),
.A2(n_505),
.B(n_434),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_519),
.B(n_435),
.Y(n_538)
);

CKINVDCx16_ASAP7_75t_R g548 ( 
.A(n_538),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_540),
.B(n_543),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_527),
.A2(n_507),
.B1(n_512),
.B2(n_520),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g553 ( 
.A1(n_541),
.A2(n_539),
.B1(n_535),
.B2(n_531),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_529),
.B(n_517),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_544),
.B(n_545),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_L g545 ( 
.A1(n_525),
.A2(n_516),
.B1(n_515),
.B2(n_479),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_L g552 ( 
.A1(n_546),
.A2(n_549),
.B(n_550),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_524),
.B(n_435),
.Y(n_549)
);

AOI21xp5_ASAP7_75t_SL g551 ( 
.A1(n_533),
.A2(n_503),
.B(n_446),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g554 ( 
.A1(n_551),
.A2(n_539),
.B1(n_537),
.B2(n_530),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_553),
.B(n_554),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_542),
.B(n_532),
.C(n_534),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_556),
.B(n_557),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_540),
.B(n_537),
.C(n_420),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_547),
.B(n_478),
.C(n_521),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_SL g561 ( 
.A(n_558),
.B(n_445),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_SL g560 ( 
.A1(n_552),
.A2(n_548),
.B1(n_546),
.B2(n_551),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_560),
.B(n_561),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_562),
.B(n_559),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_L g568 ( 
.A(n_565),
.B(n_566),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_563),
.B(n_556),
.C(n_555),
.Y(n_566)
);

XOR2xp5_ASAP7_75t_L g567 ( 
.A(n_564),
.B(n_557),
.Y(n_567)
);

CKINVDCx14_ASAP7_75t_R g569 ( 
.A(n_567),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_SL g570 ( 
.A1(n_569),
.A2(n_568),
.B(n_563),
.Y(n_570)
);

AOI22xp33_ASAP7_75t_L g571 ( 
.A1(n_570),
.A2(n_558),
.B1(n_13),
.B2(n_14),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g572 ( 
.A(n_571),
.B(n_14),
.Y(n_572)
);

O2A1O1Ixp33_ASAP7_75t_L g573 ( 
.A1(n_572),
.A2(n_12),
.B(n_13),
.C(n_14),
.Y(n_573)
);


endmodule