module fake_jpeg_18591_n_169 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_169);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_169;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_12),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx5p33_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_4),
.B(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_24),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_29),
.B(n_31),
.Y(n_53)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_24),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_26),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_32),
.B(n_33),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_26),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_35),
.B(n_38),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_18),
.B(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_30),
.A2(n_14),
.B1(n_28),
.B2(n_17),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_43),
.A2(n_37),
.B1(n_22),
.B2(n_19),
.Y(n_78)
);

NOR2x1_ASAP7_75t_L g47 ( 
.A(n_29),
.B(n_17),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_15),
.Y(n_71)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_31),
.A2(n_16),
.B(n_22),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_50),
.B(n_41),
.Y(n_77)
);

CKINVDCx12_ASAP7_75t_R g52 ( 
.A(n_41),
.Y(n_52)
);

INVx4_ASAP7_75t_SL g69 ( 
.A(n_52),
.Y(n_69)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_56),
.Y(n_63)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_53),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_59),
.B(n_65),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_50),
.A2(n_14),
.B1(n_32),
.B2(n_33),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_60),
.A2(n_64),
.B1(n_1),
.B2(n_2),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_35),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_61),
.B(n_62),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_44),
.B(n_38),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_42),
.A2(n_37),
.B1(n_34),
.B2(n_40),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_48),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_51),
.B(n_27),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_67),
.B(n_68),
.Y(n_103)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_45),
.B(n_39),
.Y(n_68)
);

INVx3_ASAP7_75t_SL g70 ( 
.A(n_49),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_72),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_71),
.B(n_80),
.Y(n_101)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_74),
.Y(n_92)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

AND2x2_ASAP7_75t_SL g76 ( 
.A(n_45),
.B(n_41),
.Y(n_76)
);

NOR2x1_ASAP7_75t_R g85 ( 
.A(n_76),
.B(n_23),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_77),
.A2(n_78),
.B1(n_81),
.B2(n_79),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_SL g79 ( 
.A1(n_49),
.A2(n_23),
.B(n_13),
.C(n_20),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_79),
.A2(n_25),
.B1(n_21),
.B2(n_4),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_42),
.B(n_19),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_46),
.A2(n_56),
.B1(n_57),
.B2(n_2),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_23),
.Y(n_84)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

AND2x2_ASAP7_75t_SL g120 ( 
.A(n_85),
.B(n_91),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_23),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_86),
.B(n_64),
.Y(n_107)
);

NOR3xp33_ASAP7_75t_SL g90 ( 
.A(n_79),
.B(n_20),
.C(n_25),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_90),
.B(n_93),
.Y(n_115)
);

AND2x4_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_0),
.Y(n_91)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_69),
.Y(n_94)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

NAND2xp33_ASAP7_75t_SL g100 ( 
.A(n_79),
.B(n_1),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_100),
.A2(n_70),
.B(n_63),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_104),
.B(n_74),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_107),
.B(n_93),
.C(n_86),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_76),
.C(n_68),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_110),
.C(n_101),
.Y(n_132)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_76),
.C(n_73),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_99),
.Y(n_111)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_111),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_63),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_112),
.B(n_116),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_113),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_69),
.Y(n_116)
);

INVx3_ASAP7_75t_SL g117 ( 
.A(n_92),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_117),
.B(n_118),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_91),
.B(n_66),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_66),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_119),
.B(n_97),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_121),
.A2(n_91),
.B1(n_100),
.B2(n_95),
.Y(n_124)
);

OAI21xp33_ASAP7_75t_L g145 ( 
.A1(n_124),
.A2(n_126),
.B(n_118),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_129),
.Y(n_143)
);

AND2x4_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_90),
.Y(n_126)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_111),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_106),
.Y(n_130)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_130),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_131),
.B(n_132),
.Y(n_136)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_134),
.Y(n_139)
);

FAx1_ASAP7_75t_SL g135 ( 
.A(n_132),
.B(n_110),
.CI(n_120),
.CON(n_135),
.SN(n_135)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_119),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_138),
.B(n_141),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_140),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_127),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_126),
.A2(n_105),
.B1(n_117),
.B2(n_114),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_142),
.A2(n_114),
.B1(n_128),
.B2(n_105),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_126),
.B(n_108),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_144),
.B(n_120),
.C(n_107),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g146 ( 
.A1(n_145),
.A2(n_122),
.B(n_128),
.Y(n_146)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_146),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_147),
.B(n_151),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_148),
.B(n_149),
.C(n_144),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_136),
.B(n_120),
.C(n_115),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_139),
.A2(n_92),
.B1(n_87),
.B2(n_96),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_137),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_153),
.B(n_138),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_156),
.B(n_157),
.C(n_89),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_149),
.B(n_135),
.C(n_143),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_152),
.B(n_150),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_159),
.B(n_161),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_155),
.A2(n_146),
.B1(n_145),
.B2(n_148),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_160),
.B(n_162),
.Y(n_164)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_154),
.B(n_75),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_163),
.B(n_161),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_164),
.C(n_89),
.Y(n_166)
);

AOI322xp5_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_1),
.A3(n_3),
.B1(n_72),
.B2(n_94),
.C1(n_164),
.C2(n_153),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_167),
.Y(n_168)
);

BUFx24_ASAP7_75t_SL g169 ( 
.A(n_168),
.Y(n_169)
);


endmodule