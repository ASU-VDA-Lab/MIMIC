module real_jpeg_32574_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_332;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_0),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g330 ( 
.A(n_0),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g14 ( 
.A1(n_1),
.A2(n_6),
.B1(n_15),
.B2(n_17),
.Y(n_14)
);

CKINVDCx11_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

OAI22xp33_ASAP7_75t_L g91 ( 
.A1(n_2),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_2),
.Y(n_92)
);

OAI22xp33_ASAP7_75t_L g152 ( 
.A1(n_2),
.A2(n_92),
.B1(n_153),
.B2(n_156),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_2),
.A2(n_92),
.B1(n_212),
.B2(n_217),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_2),
.A2(n_92),
.B1(n_282),
.B2(n_285),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_3),
.Y(n_75)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_3),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_4),
.Y(n_313)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_5),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_5),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_7),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_7),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_8),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_8),
.Y(n_81)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_8),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_8),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_10),
.Y(n_137)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_10),
.Y(n_142)
);

AO22x1_ASAP7_75t_SL g25 ( 
.A1(n_11),
.A2(n_26),
.B1(n_29),
.B2(n_32),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_11),
.Y(n_32)
);

NAND2xp33_ASAP7_75t_SL g124 ( 
.A(n_11),
.B(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_11),
.A2(n_32),
.B1(n_145),
.B2(n_148),
.Y(n_144)
);

AOI22x1_ASAP7_75t_SL g255 ( 
.A1(n_11),
.A2(n_32),
.B1(n_256),
.B2(n_258),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_11),
.B(n_67),
.Y(n_274)
);

OAI32xp33_ASAP7_75t_L g296 ( 
.A1(n_11),
.A2(n_181),
.A3(n_297),
.B1(n_301),
.B2(n_308),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_12),
.A2(n_46),
.B1(n_48),
.B2(n_50),
.Y(n_45)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

AO22x2_ASAP7_75t_L g82 ( 
.A1(n_12),
.A2(n_50),
.B1(n_83),
.B2(n_87),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_12),
.A2(n_50),
.B1(n_119),
.B2(n_250),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_13),
.A2(n_179),
.B1(n_180),
.B2(n_181),
.Y(n_178)
);

INVx2_ASAP7_75t_SL g180 ( 
.A(n_13),
.Y(n_180)
);

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_241),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_239),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_172),
.Y(n_19)
);

NOR2xp67_ASAP7_75t_L g240 ( 
.A(n_20),
.B(n_172),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_111),
.C(n_131),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_21),
.B(n_266),
.Y(n_265)
);

XOR2x2_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_63),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_51),
.B2(n_52),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

MAJx2_ASAP7_75t_L g207 ( 
.A(n_24),
.B(n_51),
.C(n_64),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_33),
.B(n_39),
.Y(n_24)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_25),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_25),
.B(n_278),
.Y(n_277)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_28),
.Y(n_139)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_31),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_32),
.B(n_53),
.Y(n_52)
);

AOI32xp33_ASAP7_75t_L g112 ( 
.A1(n_32),
.A2(n_113),
.A3(n_117),
.B1(n_123),
.B2(n_124),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_32),
.B(n_194),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_32),
.A2(n_193),
.B(n_221),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_32),
.B(n_309),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_R g321 ( 
.A(n_32),
.B(n_134),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_32),
.B(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_33),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_33),
.B(n_45),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_33),
.B(n_281),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

AO21x2_ASAP7_75t_L g128 ( 
.A1(n_34),
.A2(n_129),
.B(n_130),
.Y(n_128)
);

INVx4_ASAP7_75t_SL g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_36),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_38),
.Y(n_182)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_40),
.B(n_280),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_45),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_44),
.Y(n_177)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx2_ASAP7_75t_SL g286 ( 
.A(n_47),
.Y(n_286)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_54),
.B(n_211),
.Y(n_210)
);

NOR2x1p5_ASAP7_75t_L g224 ( 
.A(n_54),
.B(n_225),
.Y(n_224)
);

AO22x2_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_57),
.B1(n_59),
.B2(n_61),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g202 ( 
.A(n_55),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_56),
.Y(n_189)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_56),
.Y(n_231)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_57),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_60),
.Y(n_260)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_90),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AND2x4_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_82),
.Y(n_66)
);

NAND2xp33_ASAP7_75t_SL g235 ( 
.A(n_67),
.B(n_91),
.Y(n_235)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

AO21x2_ASAP7_75t_L g97 ( 
.A1(n_69),
.A2(n_98),
.B(n_105),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_72),
.B1(n_76),
.B2(n_80),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_71),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_71),
.Y(n_162)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_81),
.Y(n_127)
);

NAND2x1_ASAP7_75t_L g234 ( 
.A(n_82),
.B(n_96),
.Y(n_234)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_85),
.Y(n_93)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_85),
.Y(n_257)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_96),
.Y(n_90)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NOR2x1_ASAP7_75t_L g254 ( 
.A(n_97),
.B(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_102),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVxp33_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_108),
.Y(n_105)
);

INVx3_ASAP7_75t_SL g106 ( 
.A(n_107),
.Y(n_106)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_111),
.B(n_131),
.Y(n_266)
);

NOR2x1_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_128),
.Y(n_111)
);

OAI22xp33_ASAP7_75t_L g262 ( 
.A1(n_112),
.A2(n_128),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_112),
.Y(n_263)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_121),
.Y(n_155)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_121),
.Y(n_250)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_122),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_122),
.Y(n_300)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_128),
.Y(n_264)
);

OAI21xp33_ASAP7_75t_L g331 ( 
.A1(n_129),
.A2(n_130),
.B(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_151),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_144),
.Y(n_132)
);

OA21x2_ASAP7_75t_L g237 ( 
.A1(n_133),
.A2(n_144),
.B(n_159),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_133),
.B(n_152),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_133),
.B(n_249),
.Y(n_272)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_134),
.B(n_160),
.Y(n_159)
);

OA22x2_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_138),
.B1(n_140),
.B2(n_143),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_136),
.Y(n_171)
);

INVx4_ASAP7_75t_L g307 ( 
.A(n_136),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_139),
.Y(n_326)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_142),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_144),
.B(n_159),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx5_ASAP7_75t_L g304 ( 
.A(n_146),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_147),
.Y(n_150)
);

INVx2_ASAP7_75t_SL g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_151),
.B(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_159),
.Y(n_151)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_159),
.B(n_249),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_163),
.B1(n_166),
.B2(n_170),
.Y(n_160)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVxp67_ASAP7_75t_SL g170 ( 
.A(n_171),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_208),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_207),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_184),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_178),
.B(n_183),
.Y(n_175)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_182),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_183),
.B(n_332),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_198),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_190),
.B(n_192),
.Y(n_185)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_189),
.Y(n_227)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_195),
.Y(n_200)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_195),
.Y(n_226)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_197),
.Y(n_229)
);

NAND3xp33_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_201),
.C(n_203),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx3_ASAP7_75t_SL g203 ( 
.A(n_204),
.Y(n_203)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_232),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_219),
.Y(n_209)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx6_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_216),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_216),
.Y(n_223)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_224),
.Y(n_219)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_228),
.B2(n_230),
.Y(n_225)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_236),
.B1(n_237),
.B2(n_238),
.Y(n_232)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_233),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_237),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

OAI21x1_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_267),
.B(n_341),
.Y(n_242)
);

NOR2x1_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_265),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_244),
.B(n_265),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_251),
.C(n_261),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_246),
.B(n_252),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_247),
.B(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVxp67_ASAP7_75t_SL g256 ( 
.A(n_257),
.Y(n_256)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_262),
.B(n_288),
.Y(n_287)
);

AOI21x1_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_289),
.B(n_340),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_287),
.Y(n_268)
);

NOR2xp67_ASAP7_75t_SL g340 ( 
.A(n_269),
.B(n_287),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_273),
.C(n_275),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_271),
.A2(n_273),
.B1(n_274),
.B2(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_271),
.Y(n_293)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_292),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_280),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_281),
.B(n_329),
.Y(n_332)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_317),
.B(n_339),
.Y(n_289)
);

NOR2xp67_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_294),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_291),
.B(n_294),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_314),
.Y(n_294)
);

NAND2xp33_ASAP7_75t_SL g336 ( 
.A(n_295),
.B(n_315),
.Y(n_336)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_296),
.B(n_314),
.Y(n_337)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_305),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

AOI21x1_ASAP7_75t_SL g317 ( 
.A1(n_318),
.A2(n_334),
.B(n_338),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_322),
.B(n_333),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_320),
.B(n_321),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_320),
.B(n_321),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_331),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_327),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

BUFx4f_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

NAND3xp33_ASAP7_75t_SL g334 ( 
.A(n_335),
.B(n_336),
.C(n_337),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_335),
.A2(n_336),
.B(n_337),
.Y(n_338)
);


endmodule