module fake_jpeg_6461_n_300 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_3),
.B(n_13),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx11_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_9),
.B(n_4),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_4),
.B(n_11),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx8_ASAP7_75t_SL g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_37),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_46),
.Y(n_56)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_25),
.B(n_0),
.C(n_1),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_22),
.Y(n_55)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

BUFx4f_ASAP7_75t_SL g44 ( 
.A(n_17),
.Y(n_44)
);

INVx4_ASAP7_75t_SL g84 ( 
.A(n_44),
.Y(n_84)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_14),
.B(n_6),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_29),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_28),
.Y(n_61)
);

CKINVDCx12_ASAP7_75t_R g48 ( 
.A(n_44),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_48),
.B(n_59),
.Y(n_119)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_49),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_35),
.A2(n_34),
.B1(n_24),
.B2(n_18),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_50),
.A2(n_51),
.B1(n_63),
.B2(n_70),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_35),
.A2(n_34),
.B1(n_24),
.B2(n_18),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_14),
.Y(n_54)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_54),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_55),
.B(n_61),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_37),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_58),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_39),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_60),
.B(n_65),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_22),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_62),
.B(n_68),
.Y(n_101)
);

OAI21xp33_ASAP7_75t_SL g63 ( 
.A1(n_36),
.A2(n_29),
.B(n_32),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_39),
.A2(n_33),
.B1(n_34),
.B2(n_24),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_64),
.A2(n_26),
.B1(n_30),
.B2(n_28),
.Y(n_107)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_26),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_69),
.Y(n_123)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_32),
.Y(n_71)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_72),
.Y(n_124)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_73),
.A2(n_79),
.B1(n_80),
.B2(n_87),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_75),
.Y(n_117)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_76),
.Y(n_126)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_78),
.B(n_81),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_43),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_23),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_82),
.B(n_83),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_23),
.Y(n_83)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_86),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_45),
.B(n_26),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_88),
.B(n_91),
.Y(n_122)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_89),
.A2(n_94),
.B1(n_97),
.B2(n_31),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_42),
.B(n_23),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_95),
.Y(n_127)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_37),
.B(n_27),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_35),
.A2(n_33),
.B1(n_31),
.B2(n_30),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_46),
.B(n_30),
.Y(n_98)
);

AND2x2_ASAP7_75t_SL g118 ( 
.A(n_98),
.B(n_21),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_104),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_55),
.A2(n_33),
.B1(n_15),
.B2(n_27),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_106),
.A2(n_108),
.B1(n_121),
.B2(n_21),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_107),
.A2(n_15),
.B1(n_74),
.B2(n_96),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_62),
.A2(n_15),
.B1(n_28),
.B2(n_27),
.Y(n_108)
);

AND2x4_ASAP7_75t_L g113 ( 
.A(n_63),
.B(n_19),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_113),
.A2(n_20),
.B(n_19),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_84),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_50),
.A2(n_51),
.B1(n_97),
.B2(n_53),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_125),
.Y(n_128)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_128),
.Y(n_172)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_129),
.B(n_131),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_56),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_130),
.B(n_133),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_113),
.B(n_84),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_113),
.A2(n_74),
.B1(n_76),
.B2(n_70),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_132),
.B(n_137),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_111),
.B(n_78),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_103),
.B(n_73),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_134),
.B(n_135),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_103),
.B(n_125),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_136),
.A2(n_149),
.B1(n_150),
.B2(n_158),
.Y(n_162)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_110),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_109),
.B(n_57),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_138),
.B(n_139),
.Y(n_188)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_110),
.Y(n_140)
);

INVx13_ASAP7_75t_L g184 ( 
.A(n_140),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_141),
.B(n_8),
.Y(n_190)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_123),
.Y(n_142)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_142),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_109),
.B(n_57),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_143),
.B(n_157),
.Y(n_189)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_107),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_144),
.B(n_160),
.Y(n_185)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_123),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_145),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_105),
.B(n_96),
.Y(n_146)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_146),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_113),
.B(n_92),
.Y(n_147)
);

OAI21xp33_ASAP7_75t_SL g167 ( 
.A1(n_147),
.A2(n_151),
.B(n_156),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_113),
.A2(n_102),
.B1(n_99),
.B2(n_101),
.Y(n_149)
);

OA22x2_ASAP7_75t_L g150 ( 
.A1(n_121),
.A2(n_106),
.B1(n_75),
.B2(n_118),
.Y(n_150)
);

NOR3xp33_ASAP7_75t_SL g151 ( 
.A(n_118),
.B(n_59),
.C(n_90),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_115),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_152),
.B(n_161),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_153),
.A2(n_100),
.B(n_112),
.Y(n_171)
);

O2A1O1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_108),
.A2(n_92),
.B(n_90),
.C(n_87),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_154),
.A2(n_114),
.B(n_127),
.Y(n_169)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_117),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_155),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_101),
.B(n_31),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_86),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_102),
.A2(n_52),
.B1(n_67),
.B2(n_20),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_117),
.Y(n_159)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_159),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_112),
.B(n_67),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_115),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_138),
.B(n_122),
.C(n_119),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_173),
.C(n_175),
.Y(n_196)
);

OR2x2_ASAP7_75t_L g168 ( 
.A(n_150),
.B(n_127),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_168),
.B(n_176),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_169),
.A2(n_194),
.B1(n_188),
.B2(n_177),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_171),
.A2(n_147),
.B(n_148),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_86),
.C(n_114),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_133),
.B(n_116),
.C(n_126),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_154),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_150),
.A2(n_0),
.B(n_1),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_177),
.B(n_190),
.Y(n_210)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_130),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_178),
.B(n_179),
.Y(n_220)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_142),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_180),
.B(n_191),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_150),
.A2(n_52),
.B1(n_124),
.B2(n_126),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_187),
.A2(n_148),
.B1(n_144),
.B2(n_131),
.Y(n_200)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_139),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_161),
.B(n_124),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_192),
.B(n_194),
.Y(n_207)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_139),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_158),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_195),
.B(n_156),
.Y(n_209)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_189),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_197),
.B(n_199),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_188),
.B(n_141),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_198),
.B(n_208),
.C(n_216),
.Y(n_226)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_170),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_200),
.A2(n_201),
.B1(n_209),
.B2(n_202),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_201),
.A2(n_171),
.B(n_195),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_173),
.Y(n_202)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_202),
.Y(n_230)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_170),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_204),
.Y(n_235)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_189),
.Y(n_204)
);

MAJx2_ASAP7_75t_L g208 ( 
.A(n_191),
.B(n_153),
.C(n_156),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_209),
.B(n_217),
.Y(n_221)
);

OAI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_176),
.A2(n_151),
.B1(n_147),
.B2(n_145),
.Y(n_211)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_211),
.Y(n_231)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_181),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_214),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_213),
.A2(n_180),
.B1(n_174),
.B2(n_182),
.Y(n_233)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_175),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_183),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_218),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_179),
.B(n_164),
.C(n_178),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_186),
.Y(n_217)
);

OA21x2_ASAP7_75t_L g218 ( 
.A1(n_193),
.A2(n_0),
.B(n_1),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_172),
.B(n_159),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_166),
.Y(n_238)
);

A2O1A1O1Ixp25_ASAP7_75t_L g222 ( 
.A1(n_205),
.A2(n_168),
.B(n_167),
.C(n_169),
.D(n_162),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_210),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_224),
.A2(n_0),
.B(n_1),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_199),
.B(n_185),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_237),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_227),
.A2(n_217),
.B1(n_218),
.B2(n_155),
.Y(n_253)
);

OAI321xp33_ASAP7_75t_L g228 ( 
.A1(n_198),
.A2(n_162),
.A3(n_187),
.B1(n_190),
.B2(n_184),
.C(n_172),
.Y(n_228)
);

AOI221xp5_ASAP7_75t_L g250 ( 
.A1(n_228),
.A2(n_229),
.B1(n_233),
.B2(n_239),
.C(n_221),
.Y(n_250)
);

NAND3xp33_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_184),
.C(n_174),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_196),
.B(n_216),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_226),
.C(n_196),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_203),
.B(n_165),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_238),
.Y(n_248)
);

NAND2x1_ASAP7_75t_SL g239 ( 
.A(n_213),
.B(n_182),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_239),
.A2(n_214),
.B(n_220),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_163),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_240),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_242),
.A2(n_253),
.B(n_254),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_243),
.B(n_252),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_245),
.B(n_247),
.C(n_226),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_204),
.Y(n_246)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_246),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_206),
.C(n_207),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_235),
.B(n_232),
.Y(n_249)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_249),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_250),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_163),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_255),
.Y(n_257)
);

XNOR2x1_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_210),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_237),
.Y(n_255)
);

BUFx12f_ASAP7_75t_L g256 ( 
.A(n_230),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_256),
.B(n_223),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_265),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_242),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_262),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_235),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_241),
.A2(n_224),
.B1(n_227),
.B2(n_231),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_266),
.A2(n_252),
.B1(n_230),
.B2(n_231),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_221),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_232),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_267),
.B(n_253),
.Y(n_269)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_269),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_256),
.Y(n_285)
);

MAJx2_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_245),
.C(n_254),
.Y(n_271)
);

OAI21x1_ASAP7_75t_L g280 ( 
.A1(n_271),
.A2(n_259),
.B(n_261),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_260),
.A2(n_248),
.B1(n_244),
.B2(n_246),
.Y(n_273)
);

AOI322xp5_ASAP7_75t_L g281 ( 
.A1(n_273),
.A2(n_274),
.A3(n_278),
.B1(n_269),
.B2(n_264),
.C1(n_271),
.C2(n_270),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_263),
.A2(n_248),
.B1(n_244),
.B2(n_247),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_276),
.B(n_265),
.C(n_275),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_268),
.B(n_236),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_277),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_263),
.A2(n_222),
.B1(n_228),
.B2(n_256),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_280),
.A2(n_285),
.B(n_8),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_281),
.A2(n_283),
.B1(n_5),
.B2(n_8),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_256),
.C(n_3),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_272),
.A2(n_257),
.B(n_262),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_116),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_286),
.B(n_2),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_283),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_289),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_290),
.C(n_279),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_5),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_291),
.A2(n_292),
.B(n_11),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_293),
.B(n_295),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_287),
.B(n_282),
.C(n_10),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_296),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_298),
.A2(n_294),
.B(n_12),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_297),
.C(n_12),
.Y(n_300)
);


endmodule